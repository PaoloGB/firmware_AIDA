

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UYl0oXbWx07H12+XLY7LSDXLBZxYP6gTZvYTz2TKJK/HlMq0/MaxTmoFA++KzdPqQG+aE6ZPQ+qq
Uf5f81Uxgw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bEg0+1ra2kVZdqsGzhpfcP3LSyFAfoGp5V59eCFSwsKdv16KOkBLDiHpDDmfz4FuBKQxM9vHP9YI
VTTP3KvxWu9q5eBe18cRw11tkuJ61s4QQZID5Pdl7K/z/J91Y+C2pZgC4PyYfdbZV9nqC0rqz34N
t25TMZ4X/3isyExfaM4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uu9uMFaVElOirR8H2+pn9gEMn17E//IYYznJRRoXYZmK9rFyndxvWxzgXxJnpmdqmEWjml6gMm/H
pembPItxQCeo7XrM3lTsic9mzXXAieyH8uZnhARAVJRKdWx7M8NVCShTsM8b9SyZmEbyJbc4S6Ot
QgwnO11NxnwCoi4JadA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mjXvcb09NMDr5cbshxSED/yd+I/z4J19W3+kcWNP/OCSlWn1szLbF7IO8Fo/qEP3dvSJRly/ZKmS
P9xe6HqZi/Hq51kBCz4qioiB1vvTlc/LH1RyHY/WLqF0RFuHmjhEwQpdt4Iq9HALjkDyoFAQOLvh
1tU76/82ig93joc86dKaffZE7U3TM9Jph+IFapSuSYa7IhWH8QczB63lTMnaGHkoVrByWTXAptds
d2R3ikHwtMRxJY499uEXii1jFu5QI26PCikka7w1lgU+SjOvMCKSRdZ1iUl1Jat2MfiNiCqYAMoj
DlISuFAyw9808erW2gozPmJueN0p+foyMN/7mw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c/1c469blILitLPEgX86SdGoVdvoyvD+/mS37IQOELSF9DiZ7DNf22AjlyJ801EIuF2kDm/eFZ7P
QeSl6otd//Msh0knUY7GOjPiKvZrAqibedNiMYmuhgjyAivYhuuHW/qzCXcwxk4zvdSD8qmkBkow
AoGHtgbXvTQrLELWSOJ6kJZrrsBQXOF/LEnLzptFNvsA5mx30A/EhQUwiTWhLRCs0+ZmwoXPja1b
iewVOs+yzFKZxKCXtAslkXwj/v5TAyb7wwAWtv0TZRZmCPLXbG/3htYoj0jStM4a67AxbtJ7ssQM
lCdCllUOr0IzrU5AZgmBqrO+RYeoA12X4rjPaQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hUc2uWOKrgaR6N5dF70TyOCK9ofPYM1/2lX+qEswJVJBduhXVmcxmi0OfBsyfbBOXlaiN9aeep09
buHtyIvGbh36KoOH58SMb+I4sCh75XnlL4Nsd1B7XSIJqyPQs1i+foBbthDqV7JWczDAdgLzhQUT
29R7m/ow9arPbR9LkWhDfFTDRDdhWkgTK/i2hPuXpSuh01iwND2tZY4rwI0aVM/Cdm3eNeMGd3To
gQc1cJ5rut/srYm5QBf8y9aMmvnwM5epeTVH5j/o+D47veCwWGXWno70XbYsJbNWjoWMlR/ARJE6
E+ra4UJgO17qX6pHvFKbOdqIVzF2hfYgExvVuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504800)
`protect data_block
GvopRV4hVhst4X/10vPXB4alpgkR0ai1Bi/ssG/iEieeMNTHQCpoqRGCdTKFUX2/gRJ/mKTHTYW1
c6MASEGsWs7CyZkUdkGxCzMApTk6dWvBGnv67gFpjW9HcZCUbqndAy/44fh9Qc5Cpj9pIc/V0bPQ
wvkqTC/OMney675QL3CuVdaSu110BUbaY8oE7jgMMZhcIJiRZRrwzRRHugROOJcVNGv21PuJjWvR
fqR1jGVo2iFuXPxNff5f7yo9N89CPciXDd6LXQYAySZD3XkV8yPCMPBZgotUP2PIsXcdVO+HY1wb
RYXxDyHlKFtOEG4n3eQHUQ0ZrM3es8t7E6re6aM1zJX/z2BmbwGXFvjGSg10PKDMw+Fvzh1osP+J
4zMFFvMh7xWkqSCFrs9+qHWCcLx6/liOdXsZbnP/D06eEy982ewOebyUEZdnNFqT7I7+E5ZM+EA9
1nA90jWDFs2JjaIDtpPSOtHX++oH1igdQFtJ2TaLMuhfY0KLG8u96BIk8FOv5U0r1zW3T9m4D62h
6oMtR1+rEM7nAiU5vlvXQl34wuJ8Z9KnzzFr3ef1r8BGty//EBSoYFIFqvJ2Z4qQo32I+oSUcK5K
I7OxptTJWpv34wVd94gE53gILeuW9/INWXhctieqHXUOyCEyH5jCjQchUwHUPyIsugJi4dJ4Pq2c
xgVqfG4Mm0hKWJF9fQJoBkNut1wb3eqc9UVAYbG8aF6k9ivcqfLpEOv186M+yuswR0DhS+mOuFFl
wfLUbJmNSpZOFnN5crPExaqRH/Va4x8dMSjFffm3k1sovAxSnis0x7/dfPaPi947fXCpTKlNOxHD
mJc6RJePleD3rG8MKSY+DkpuuJ8j883dBj2tppqGRCf/CgSOAGqrK6mMakrXvonpK2x2f/8hxQUi
q0f4yc10Axy5e7M50Vi63vHj9xRJkdgnyE3pC7in4SMfGou9o+2QLvdwaoe3diDaYhLS+ovzzImf
TL/Zb+RWuV9b64a71V7M0pZao1rVTdYp+ug+AWVrN6834kwKABtwz2EHbG+HKbDsIpGsbfQiKIWP
m9PshbsfHSyPnGxMPupcT2TYVGfdnDIXywmzMGojUg9fgyGz2Ik6rBbBeOPz3pNL9AoSQ3E3Utx8
OaPCn3tdLgtsh2kcgdksTjdzc3MNUQNxoULAWQbQn9Lqs9PJQugFd4w8BCjuVJoI+si/L5dpZHIL
4hWT510uTBu69vKBxwKhpAruJMXg15/N8riOwAx5S+OR+ipZbiqQaMcNouiH3Qit3NNz+ccESCs2
p0ja5IWHu9MQ1VFSldcESgqEb+f/g3wuJR5T0q/5PXGPsCX54bnp6G2h+Ux3OOh3srtsuMrcUV6V
8fIF6ZoNGK5I4Y9Tu8FIOyGT6548WSBqlkVt11X3HJ6sYJk8wPJSkzaKrlKFFT3IlZaWLF1Vkqmt
mBzFyelNItrbXg5NKQgUiPdvJLYDqKNFceftNNeJYiBSau4nXXCNkAZLqTVg9ZC7kBqmjDshY4K+
Co4IRoht/GNN1Km5dAb5YAthdvPW66LybwhI2otPoVqwW0sZr8ZL5ro9DlGVaw7f4b1aCJ0Tl9iV
xdeDUCyGXajPKNKD6o8l92pK7oi/lB3ju4ra/X4QExlWqYoSrL5O4PnOEZaqWsxSZvKCG21Fuf0n
0keV3s/mHZYs6uGjj4qmh+hwcHQa1nZRR5QXwDBoYtHwtbbGZ+H/PUpK9fqvTUDqwX6M5BvrwIIV
Ffx/R5zyXi8hZGUP/pVoMwtldCFcVOkSGGpzcvUI3J1By8NJVmmpQ9Jq89mjnuU7xzee+WVxLiYd
bWzcrreIk3AyyhYPd/mynxuhgIi3X6t7jdQwKOx0QwgzhFwlVVZY3OaEsBn+XhnQl31J3tg/2t4Q
w/1O/q4MRLoNdNFxbk9dWVd1eOc3a6zrrOcN+kQ5A5wadbxmgj/pdeCG+CUSTnOhWdNHx59hpqQY
MxYkzuDeSSJnw2Rwi0RCJ1rTiekxxE4EnBDUtxj9TBWq9v8nMLaR00wN341ZAEuSKNyq+VSXIB95
pdh8z6AWLCgQ34yI8dkg+aqPu+Ny4lHYKgOmwZ1a2dQYD4BPXprjpZR/p0S5PXNb5OaSdkaJrE5Y
eblBoEkvMQ2O42OwsvSJ9hMTz6k8Crje9NjkjfXL2Jt8kM07Sib9FEhSz94ujcWuJAyiFZCes4r9
swJ4vVYmQkbnWQdlAAIxR3iLP9HiK/cybfXWZoSaVSgYqj9jU1Qt5aXE3UBiFNoQuvK6eIcFC/fC
unoYubqapzfkrzX8wJn1Yfz3D8vpQ1WHL4HkVD++OZqLQSr82T0ulo78WiVVQDav6nfL5xXJtMRW
fR9WHE8DNGp1+OBLOGVfXBsUSD+lV3T3O5UrNV4xEQjsbZSiuQ47BXjnLIxGoZFnkfpwvnVwg3TF
ZnUn4ygIj3gbj1FDAlsAMwMajB26bxQDig7gBk0zwX9v841F/UbvX34w/2akqpQt3lmjqImLPK2z
ZIy5ICXkCSxFQO4yAGhV4IToe2JixZ9I2L4ShxUiYk1UU69XNkVCp9/ZNoWQUcox4tN+eISFzIte
USjlxRrFVoKoJ3Gtms81Yul3uisAb0NcMnJWJzD8aCxt8hWA1hc1kNfPZGt6z6S0SGt1rYzPeEqC
8AbvYYhzkESUeSyVH7naAiNvurfZ00a1N7ZsPRGeaDgexpXoFIY55iIFErgzK6otmMslOduQVXmX
c1MpytaiD61ee/OnqtK0mDw/y0SlsuQCfOsBRQ7W29HSh/czNBH2pBDCwc4OxNsAb6lZyMctWNrA
YuQI2n+C3tSO4SAXAK04Sn44jM3MvhV7aJKfVc7NR70NQXYjghlnwv+yoJw0F+C3pPsUrnVSws/2
hHHezQxBk1MJ62Kz6hISnuOKI107p28YosPnOvmkjOwB/9SNY0gD8mbzhehO1+WGUWnz4vP+zhW5
hnMd/qMIi6Wo7w4YElHOinH6od7eHmeT6ZsSSGzHNai/hkyh0vxlrncuc1vDCtpWxoKy6Lz4OyiN
XVocy/zVhl24rZUxLe86eUZUXVVwsBgHGLub3GVbV2Dbr3coc+O7diuUC9Fic2ghSnjeESVJxadK
F2xZmxMyBZAn3aLjLroiX2RgKmUqY/9lvwWX09EaZIcDX/ZCOIJRJ1Xbz2rrBhQnRlXfbSyHHqpU
BUy0zOxl90hmgp8p4jbo4ExnYEI0XaA+4h1KgPORY8Auz3TBinnFVnVCAZvZRT3TeMZuqbfakQ1m
O2lmCXwCg2zx1fgvoSVuP03DRxI15LguqUfqLy52MJJvLY5JO3Xt2vPj6HG3hTUgyyfVSxSQ99vJ
3cEFU1HQVEIZ8nCoEk6PgP2QEGTXFTcpK8ATGp/rxCZL6qUmt8buFZqyTbHm7Dl/hJYbnV9aFBWS
rYeQBUNEvuu9k9kfFvljaM3MSYTwBVQlK6HcEU+N5gNQpQdFnp5gdYtiAjPtCekPTS+m7dxu3gk4
bEuzuhoAeow0KYZH6PadDu6jGtHyDfxqdggiQyUFbzmXCopcQsZWBOOnDDLRsh4fu0zBHKfqV89X
uU+r+wbT0+4AxWHgN6raiWHU0MzITfHAfwYAFSyHq7E3DFZBKZgxlmz/xmj/4YCWzXv6a9TVQoLl
8zcz4hZlispQIvPF466jO2VSBkiw57OopgyzU51ltXeEvyXO9yx/z2G07d7bP2cvGpQFh77/nRFs
uUhZCiepHYXl9h31PpUQGgoceIYiFM89oryR4yCbUCMopuWc4CkLm1yND/2A64bGGtQLuaFKqqEO
26yI+BhOlnoHquHSmklVyyLHfmkGceEA1BAXQ7lhsMtE5QEGTlSFONVjyDkLGArW98qlWJOgz5bw
XkfallGN+OPVD9Q3/qwYk/v3lkbCHlK4BjgMx8BZHEU3Qy/J+U/lmjwUcuuKHei9/WudiAnePCGS
IrHPlRd1yWuhjLVxQ4djtSUxBXH/5gNCijgsy33irF6A7JgW5ins9IxdE8yvP3tr1Wz6b/iVPSKl
HLXEW548Y9vqQiRd0i6BUcOfuJWirf7C/roBDvQAlGpSL7KJ9leSbeilBtHPd//8YBsuHI+m7jCl
sGnIJUv7XgX15WZYRobqpcHgimUacyZtsp20OSVzkBQClbayDDKNBd7Ce0x2m06yaxJLsSB1JaDq
wPw2WxAS/8neSfBtGCPDYWY0kaVP5/QVnl5DmEZIFYEP1ULJ/ZYm9W5+qJuX5KXTXUVU9dej+CiW
ehHwMhiC+VxoQ5hL+zAq6bOd7VqvrYsLnlRdzZwMvzP02qBNaJCf/vWj+/nbDGDJBsLh2aDUn5b6
+JSNixoLgJE1QaV/2MdrjuIRGcpOXwgjp8Xm5Gmo595BufCEkeawv/vKGUlvpYbzpxbYud8yK6rD
f80ChMW5FZrSELe1G5Lds2DfKlEGGVcP4MJL/JBFIGoIqi7M/iL/GlnSiUf9rr5I6lYYHj+2IoLu
zdB8OHMLrUSOdCKDGZW9Bvg1WwsFcw9J0PqMV1OaY5OhZdGbyPxrno3cuwvC0BsGZWkDCJiBmOAI
vEpHQLK0r4p0fFg9DV/rw23F2TSs7SzS0x5cCBIJCxrUB2JizpZVrgm1ijYqHrKkHnaePOP0RE9D
uN6zjYbc2zImM/03vYuAzb4SRZa3w3yUjEgmJeStLeALApGVw7tv4IwmQ6JBiaDs6uIu+R+GDRVe
HeE514nksiG1sJeYSbbk3IUY6GOH+S96OMLIyjgldVwwqYtpQ4o/Y8kmV9n8REsAATmCSMt/mLkl
UGCQjvRSw7ZhISrL6cSygZdPDMzEcY7j+/9EBI8C5GaZUeaBFMF2n65t/Y7OjnMhcqjHsbdX5bkh
yfHq1L92LasHCk17J+TMruYeDJsPewz051JA4INQIOpiI0vphRn2MxhZuwd6NmpuQJ7XFOHXrVJj
+CJts8N4w7goKPAX8l96QYMwkYJC/si1XDB2jK7tiGbN9yWfDAz8lIMgIOKTRE/J3C6qxy52VK3K
2DkUiKByOen+XRKn0UDlioHh6Yi5nzBaaEq2sWxpcy27QVCzwZb0XLGbSAlk4H0rJQvDAZ+xjF/z
0xgGmvu0G6WTpu/vwIoC4txyxbC5bi/wsNKZ1gWVBAYGUiG8Zic5kh5jLXI/ZHmGa00SuG6fDKA1
i/wsFUAsICzFudbZpdH40c7ifn91kirDnucrEhleMYfB09p5CK9LMlYUN25sBmqqXdZfTN+WsrwZ
qiMNPigZSuGWMezZiU8Zm3x27B5AkAVJFY4g4CKJbC3yy6ukXXRMUti+/zwYVSypPnCJirH8HOST
9bXfoz4maMxKHyiAqZ+TJu+mVq1AaAHY+YlPe3ZK0EH9Hp6yKIbeZNHBJpJScNNMCh5dDz1OtKxy
3V7qvc6zF9VOLjqXovh3u0Sudk1VbfVBvA24pvZNHv0lhIIBUn3efNCHNT3Jd7eGz9fR3BJxhnTd
TiBXatt7f1xTbdr0CNIFQQyXPHhpIfpEceYOkMgLG/i3SF0d2RR3c/dM3cf/tFPE+oqH+lPFsZbL
Q2VWwzwYpM5HwoPtuuxv0lB1gcJdXxSjIKfCs1fbp5xMm7g8xaAps41VInY4IAv4F6DcGTvJDSr9
/pw4VkS2CSdKoJgrMPDrw7s/Nl6ruiixoUAB6Vw6pxsCaQamVOQgV893EM2FYqraaekX7NwgQ25H
DP+wHHmzjPvyWTnTBr2qoNWAzJ+yQyORPGq/0E98cFFwPYHs7+QcM7g0rcfJCA9vRpQloVtGvBqQ
qQ+IzSaWwWiFnELvVJIjO4F0IWfGWY9wBMkhft4rHft70SporkYlbQb37+G0ms70hadMSRTSiAuh
v2NDmd5rlFN3T8sdjd2i7LsFWq/xti9tHLT5zCkDwJuF/+AyaG01sxo7eLJ3eL+t5MJGS9TnzSey
7P4egn9ToUKLV5KUH7WDSnmDrrI7Kca4b3jhPVEoTMEuiPy5AD+qJaOjl8bwQl85Rk73h+5F5+cq
Zg3vALB9BxzKRA0o5B0gadv63NS+XLlw4/4Ez2IcwlO/KSedRVHVkiNUgM43ihpEvm/USFVSlj38
ajzAtaVILkkclQWuINSS9V6FQKEbH4MFqWt+JNIdDuiv4oYyBRDre69rY07cilmrbVs8btcbldv0
jVNUeR1P+BQxGiSHL9PXrzbccGxYz4UTV9xTY6POwpHbp11xSikwByBccthj53ZxFoiPMfYhBEMt
3bTu4LVEXzMV7ma/LyKf/GYKzJnEm28JSja+KVsUvmbq2+d0wia6p1Lz6YKI0gVKFYUd3+Vtwp3X
vjJXng4uGouIDoKsp3QG0mFda35V3UePiGD0E867pw0707K3cuZFhiZ8eRcKac1c5wG4pvWj280h
aiyPwZaZ+Ct+XUwsuS570+dFC2QaDQupjCbApKR28Bjehvppa4flsfTaJP1FFoYMi1UqgjnHw2gI
/BFxII9JvLeFH1hpSVr1t8yWrP2MpL8HglE0mRrOEEFGlFdCD5f3R0BDHOZ61nn7FjJc/2WVP+ZJ
Lsps9o91MQOaiF5tFPL6tRZN9P0G0uZtAhdCY1FSKyoYIxdaH0GjfxLTM9ZjEOPPfBnKI9S28Df2
0gCOWPtLZjFixU87/g9nEO8/WNPal1o3aLSx/3hcSXCCJRm6zfmZyLJQ/GGvwIqNHZAIpTHt3SZB
1g7t4ZLOEuqxAMj+xKavwPUHeWrCAcLsKKXhOQJr62QG5pp9uSx2REhFqcRQ6jxJwkKpCuoYxY1y
q9QpxbhDlog+K92nbPmPnXHPOzYVlobfQliqanluvA5pc1DIM416vCgwj4fGUfs0iNWi5w24+65Y
5QB1LEFYdnVnm5J49PStD8smVQd8QQANEODEB9CHN1QxFmJeV7Y1SKjfmsdWbnIt+jEP0XrooxHV
vGzvhbLV/cXEaqDq9KQsFTXVzNjl0jn5/4iFe+y38h+i/WB5zIb+hmIEJpnS4O2ZorH30F+a+ycA
5DVZ8V6w193+9ahi0Rhn41LSZufO6PEnd3tCgBWDhyYqyjd/RIKcaxINYJ4M5EZcrpHU6+OgRIF2
RlYe2BZZ25y+zFHDEDRa1tayOZoFN4dSbrVZ/bzUXsnV0XLZTHReIQOb+pQkPDy1Pbqf9OzVl98i
cXDA0jzPbWDhK21Jl/zxL71ey3nfkRbdRM2XjaVdUjCnCwWuvyDelW3s4NAAPFV91wqGEeOaIGOd
Y8/twlEdqm/igWenWPyVZTT8BMms3AKa44Osf+VtHpNEccSw67gc+rG9ZDKmJuo19yQkzRL7Bicy
L6pE6IdtyM9FKTBU4kXwfNeF4SwUe10b/bL0HVY6Nd3v5EPDJiHCRaS0jQGXSMYxDO8hGixMcYDe
W63C786QqVILzD5NSXMfRqLbAmulsVNF4FMw3v26ASZ57NLcaVoR0JV27qY+/I5Eb3/FCKvfLFHe
c2sVhtVsUSoCCzrSgBj15N7ZKU3J4X6HR84s1Sra8J0BrsJ1D0fEdtPY7G/tiQSIdsi6DAPlDgWz
lHdgOy8uFJRzTREXJYp7Dnhx6if08efACf8yB+RMGgF/o6+QlsOlQRDVy0ESt2aH2/shb+IIvAvR
9PO1AUDWEEawIf+TVjCRIfjpb39YRixkdJVuiDY2OqcJSxUXyZs4G2IhFxGVCAvHKFXy6a/oJ5Cj
WJ8QmHnO6XuYxAIvEOP9pKq0knQjKINGqVQag5TxgBWQhvNnRn/9sHC0yKuBPLKZVCUH/fl/ho3v
xajYI9koea6Per4YbalQ5qDCvVZ1dYWXlwFVwr8m7UMsBpZ3AGcV2lUhSG8MGP8nYAT7FW7kRHl+
U9Frj/APy6p9sGGrzFsym14t26/brK4/bpeIq17sp/BSSFie5pH4ufzlP/JdyDTYtFImzz3gxX9G
rIFivqMU0J8FzpBBaHY53fooNW8n73mNwLwhL2Lem2Z1LxWgWEtYCDd2f2sx37aFLbS2EtxsYOBC
nbPqRxMiQ1c5CfJ3w4q/GvMPzrlubuGiWvS3zfeadT6JPY3pgIhBvbdO1Tu1c+G1X5iZ25Wz86gZ
sRyMywhS5Y3vZRtIe/CniPV/V0+LRjoKos7KpsDLOYY8zCgDNrDycqzhCZ3w0tw3UqkPRgLCOq26
dfDSKnkIgMPbSpQcNlrkDx/3m5yxUwP95+73NpkXuTY1+RDLA4oiKUuGRr2AeXXhFRrpJlML+Rfx
lpCyhNVuErFt3AVaw4DoumcgMR8aeRJX6/ukgh4KN/A3erUpzRteRq3yUMN0+NTRrnpTyXJrkhMl
0kKKYNSeR8mxc5gEnRYaDmUYhDm3pXsHovLy8zWmAzRe29Eotr7x0rJT+PoPKsqeskKuTeGPPLSu
ki4ZTmYV6oFxSGGS50cQLROJl2JAxvQ4ce4864La44YYluhj9/v7BimQQYsj3nNCc/tj0yZSp2As
HmqpKC+7oxtGFVUqTsqA401nJSndvosjL3OvwPz5f4K0L0pt8GMad97LldMKBdvHKfvHRk6lKWIJ
8oLxikoPjgyGbeTAUGvV9l7U+pst0yxVubc/cBtmpb5H+/dJoUDy/Um3/ujltCxswYjlQMHO9xw8
hhGVhi3CyuPJyYS+hyr8MZW8vv7CpJ2ofHAgJHj2sE+rHbYk/GWtTqNFyjMG64udc+m3/SJ4MLiT
Aww1ivgwDwmkqhS7DfBzi+hoRALhQscFLKYVUn+Mj+3Me50ZnXjnshD9vbck29sxUN7epBLbdFN1
TOHAKwg4Q49FS1Jy/C9a4vpDqVh2UdB2JOAoJikrKQiGoBSc4fIbHZK1q+pP3vmKEwppVLy/dnqt
6hpVHjz+W90wObsOaopuly4pW36aj+WOFX77jMYtF2TgRnO/Zqebz08ZhUxHyaWPgNOYMqv8a0UP
59U3K7GjRywRm4cMILzroOfV2yrdWUY/vUzsocPiUJsNTNM476OjfZEstejOF4XNZuFbhgeHVPsB
/CAE7Eqq54PhH7xWo+HwXSq9jy2K3cJwL4nnF+iQbAAgJXLaU3B+YKHACuaG7N5+HNESjEba08GJ
tMyf/5gEAYfxy7rq3+H61vpm2GVGTydzUN7sF93xwLXX2xTt5QT6pdB4dlVjOkINd0dMxNYaHPl8
RgJUlvVNVd5mT4kgzK5OqmgeQjoNdoAetcjQJODSfRwqGwdwe4C4UGczE4g8HpxsUjV9MnJxZNla
aUUz0Z1z7R7cciqa58wLEtKpqCl6gvb9LgzkA0HupfZjkCOi36LAm9baZ9hxYsTUpNL/tVgOqFXR
p2hrYLHBVbFcU+G1YkZnPVpLqW+MpQ1nfZEX4bOBv+JF026krPB9x0bJYi2Y9lRurcQDW1xoAaPc
6fxBvoq0UDRgHqYcYi7YKLhsH08m15UFX1K3ZUQsIMIrkw4OLQy3j7GRJJwOuO3t09DyVvHD6m75
RYLMPHHGGSLrrUXKA4kTe5jJrhXYbLLAjDV6nijLbQJO5FTVxYtFJx0294VO6dQMuPVO2webQxoT
omSfwif9wRDKhNd3Vlj5W2N4Fuy59Lu3oWlKI3Ox3RZC9/FRdIUXho+Q8450zJIyBqsGE1UTHGkR
uz+7vGk299+iw/kgF52mKoi5hZz7pBQlGZQ1vffl7oOZ2qBvKcE9XxuSd4g4xTsYPgQ3XAadoUKT
is75HOLEEcBiw5TNWZGNoyYszGa/jgiymwubIQhpNeCEij9SqYPJOQtDRosnDWPKhnBmzwzi/3mY
ZXvw+b9JTgEHoZFL+aEq35avD2ybDxVytA0mBNlOmcvvMXspKetsc8T8bGSXxIyfbiC8begdYobK
AjaUsJp2hqnO2mzXzBdYfUNKJMCTjEMWHQ5ww949baITLZxZgoo8ODWiHg6/DHgUIMriBzBpLlwq
RtByQuqDIVLflJQzeW0J5Ig4LO+TcQ6L7xVX1jGgC92egBZmah/uy7bFmy5FmZl95JEiZm/GMoIB
xRv0eiuyJvttNjrFJNFVXT/9uvRU+gVu4JcPj45wUqZ1UI64bGag2dSQtG+gRCfeg9tXUN7J8s/K
Xe7vimLzQHIThB8KQYTU/6TB7b3YfUso1f+e2idS0Sq2UHqvedfDgwak0D6T+dNmYt+S3kAz6O0g
rthfmlEJDsk45alM4S1+dJXe9wKpPjZtkDT/8dUrUyI/s2zX1aRzRSFAUHJCN55uPpfemVw9BvjZ
b0Kjgg0cbv5bj2AunusoOKHOmUJDbXlVAQO8x7cxxRu+QVfXN3F7F5aUG49XUeDPqAlY708FShy3
dRqBN9VPSEj7NvS7Iz8eJk16aI+eH5yZ213r5VC01e7lm6ic1bhZdBZ+9oXGoijHivPBt936927n
3rZTCE4zNFucKCvZ9TAWMCTLqlpoPdx2GslYqFP5BvS8c9tsuHN3W+QXJAU6ukgPl0Lfy1h+k5WL
sQjJ82LOCo55kXN4RKXnz/r5rI71WcyaYjEyjYCtCGV/91TEId8x/XOkzFfCmxw3JAls9b3yc+Rk
hLQANKX3hbHGd7drIPSiP4hY/o4psw3UT3uItm5mQL2jx1FtuWpMi1b1I8WW7jOkc3oyI5m2u1yT
i0B3L92OfuBOpxeUSQOv9jQCr5MQctS5khrFqZRcjAhPgil/K9sLrUJo+D2oljBlNFzzaHoLQMxc
t1bKjgo9n5fCxEOCHkPpWLEv9aB+iYaEzMtbX51xj6W+YRUKOfR8mE7tzCNyemxII0s4QSB8lwdy
zVKjsRAnK/QsmYtnQPeE/1V7tBB7BWmAtqT0VS2j5w9R6mVs/8DA+QRJvtXG4RTfRmi3lu1Nc6iD
hZ62MXX3kh9kLm+KCQw8tzn6fVvjgnll9tPc3+g1IApmVpYdKGmY4meHn1NscfBIF4Rw+kXUPxsn
EW8z2/7P91Y/ys3MRhSTmKLqMqBZ08dWZ3zsdYJt/TQ4ITbYlxG+WWlPFo0x0X0w3CSLK8albV8V
/FOTuNpegNy1lRUzf+U3SbTzEZKloLgKxyf8B+0/OBVbOMyPwwmnr94uNABQylNWdI5QhTKQZVqA
OyUxAhgniPfd7qw7jklSnsKSlmVe5SOeqr/LhZSgQpZJOv/S0Y8OdKy3C/x1c0jh/XGqWxofZvu4
ZoTSTNDWxpbFMWrUdqkQJjkNFAQAMoaiNExfIqRWcTIzajXwm4HMeKZ32XnZVIRrdh2PnXIZ6z++
ncqbAXrGraPCPgmEXcc/lW+nhQXCmUT3FhmpVMCR+zn3OSB5cACHn6Gx+L04T1QBCcZ+Ag7aIBwt
lgxhN7qr7IZYt9jXNsiVRteAQ+UvEUOvPvvO1LT+p++BpGvByM+p5daWW5MSG0Mjkl1YzSOG89uG
0B3VGU5I5MbbkLVM1JAxzvA3ptunYoGKWO4wQOFndqCQq/+VKo5zT6gRMupIjPcOM4BAx9IW1nEl
SuMdgkWlPEeQJwsa1NOm1+RojPGq7qvwsmD06cAdcDKOQUBwXNidwUdSpOuI9ZFDDq5fq1hhEuo8
1k4RBhfrWHZZA5RvR9aM9fQ1u3GWul4zW3kT+PowXJf9jlhwgvlWhJ2Ujc5DALJBTTWxCErscX95
L6rYTA4tI/bBye7RGHfX1EllY1aoe2WrMvX9mDny1BY5WAXjsOGN2LMtE9YYMSnFudIcVskKV3JD
b5qlKwAL+kMSFXDOtADic63anv01tDkhyP61RcH0rzvOYOwg9zyiz/IbAsndnvfEsU6LJEyu00Au
vWYCwoikJdWFgFXxpEUh7I5Fvqyig8hKj6zyupqGvj4RlVVcT1LHJQfPj3KYJ1bCB5z55KuV/SPJ
slbWxxa638TGqwLX3LMEQ8WZerDyNpaugGyybF5PfTpNlEOAjsoKLtFAXnaVImhWUnYTN00D0OBP
7aW7cCHGg65cQLpux/KOF1nYtfLGye10KhT1Mgn/8cIcWoBUbPB24IM0scvNQ48cag03jp0Ji9e+
txn16gmpSre11HkIhtbh8mswqeNB46dL4kvqPmozcPOuWwfbh0S+JFRzcQmflj0ZsyM2scb5wVk/
xuKDCOPwq4zbfeCSbSEdaQKXvsNl16G3sedZsdOlrMGM9IIZtno7f+/J9bS1i+7qNTCCuBBhNT3M
KkCDJsTo4N3lhssIhV9E7sWDHJN8GqAR5Jo4Xle7laNXwllBxtYErtDhOdu2yzvtAbk1zv8JMJFP
HM4501PDOzMt80r3wVbLpOxWAxy3LafQSKzXX18VHHKn7KHWW6av2zg17rCdbGQ+xrHbXWVaJLuy
ir3JMr37DIYg0N1kvHL7VJB3rkEVgEoHlNO5g0uhY14crp158rJiOCrdp4Qiw38hrXYC+dJj2/UX
K5R8SlOpoHz6wK/vZonTSfHcX+yh7PtMaVi1u9Fka8nQWwtsJK2ADxhm6InaGEoTsk2YtuJyV7NF
ygKi1VIYd0t8pwh7s5cT02sT5HwVmXirBr3AFpx16xAgZiP7jbRgce3PFUV12fcePlcBmsH81eSj
jnWOkJDPACQvTDFv1iS9fdDpTbwIdz8Uhx7pv4brPSPMmJ75HHxuCxDqUD4DBXdwHf+1hhLae7CG
HWm3d3TB8CFXD52t1EWwudkayrDQrIILKv4enGlMt+z98a3I+RbNKKOMc7pOoi9sDW4o8p/PwRJV
qo2PYURGbdZTxrL6WTo+g4zXlABR3gbb55TjanvkXA8iEKQUd9MDHeprioog6RZLk9CTVexTG76L
6PVxauFkqfVMIojNMQlVmTi0jbeKWs3xAglPX6SzQ2YgCcfTzJS90Id/tbhGFS/wEKAM8Y0+uAgM
tIF1ChnTxedzPSxBs3SAiLJAWLXjA6zfxVj7Wz1l8RZvyaYFO+52VeZBGOlcOZIlLDgAPAuMRhja
AP3W2kMPOo6IOT/oYmxMMJjh8rNRVyRjo2Okchoux/IvaoL9xFPSHbxSGAX/AWC7tzn8jULuJsjg
BJjFcWUOGWO8FVkOWgLb7oP3XSvGMPG55GWYNOjdCmIavTQNkx9BGiadnhVU9p2baxweSFGUYQ9s
5GjAozgRCdLHRDiMajmdsGD4PGZf4c/3ZbWjU8wGH0xoCsJ9UgGLPkfide+KpKROHju9I6+JaRgN
KNktBmxH6d03yi7Y1pQo1XvqL7rgOR+mHO4HcHnFnI+96HAfwFxkR8eWJcA+ZbbkWXOkxFC+Gfg0
JvGqnLqdtOG8UbYZJYiV1OhFTPibOqHfjFZRcDuPA7k+ZIO0SEIz08O/AtGT1SpMJkKZrOS28G+H
YROCs5GUP8xV9ci28GNKAKK1ZdewunoYc57YOuJyHCXKbctX22ujJ9te8Tzsh3AYrt2TG7UXuHF1
sVkOl0KYIv8hWkLnFZVhptQDUAgls+gHTQzRsZW/EjTK+cGMAuRy6iNVMIdDZYcZqnVvfPxihxXk
ktgXLdc3eaxFVK/X7PhGGZU6RnUicHAJcDeQjt89cH4ZAcO9jxC4TI2U2Mxv0itKMCW65LMuuJEg
iq9LTWoGujZ7EsiylVJL5GAMFJw4bvgsR1yIMblq0NpdTenMXIjPjORF4tYV8WWQQDezhtPL6QfK
X3d46F1XNkJIe0l+yP/iWaQAWLCJhyZAJ3DU+dMJ8+P8ZCFOjb41gmBi1HCpOUb0kXgketM5+ZYM
F1DZt1ihQaCze70rdG8yd68vVHRlZJgqyBfREq52jJ24yBPkZbjvnwpesoVLDTgdMlIM6YGhxgU+
hoi66OoaE9yiwu5Ly046oz/Gq507rLPzldSThCiaYghZcNuKENdQHpCzz6MpEqYCdjkItu/VvXdJ
+cCQY7CQb6qCtV6bziQEOTIOa3EcO0w2xHzYwUjyjd/ZooqPQGutwxrk2LvJh/OQHIyxeXPbBW3S
aCTZJvW04RCVpD5oGm4e1qSJtfi+T40DP612q2tQt0HoYlVweDv9RzjvRVv2AieMnfMNKjoW1HQV
rjtcyponQbyMjDsuA//iYfCvJc+vtXX9+OWdvEk9NdS5R8QEUygjx26gCY2lsHsIU+mjGOPYh7C8
Q22T/lQyRiFSjLNsNdZFrtpocpO8M/8CrrHdPHL5SHpyddZpJXSTh0tGd2xG6pOAx8j5cfnUsyXo
3O7aJvDJw8fA6XT1SYIqdivz2M1hqY1LBdcEKvb8GODBMX1WT+yUSHQP2EDkHK7sQatl5fMpZwv3
AEZ+s41Fe0UkNh4UZ9G7wGhoUj4ILSSB/VPiXF3xs+UnR7QmkqZFQeYAgtfFnKnT8rRL1c8z4wZH
6yi2xHuITqollbHc35ZNuW1gdTKdVlxpiSgthwkcgSpUD6RvjLKKJ1BM6I3bPMiODlBPTBRwfpl4
6mdu3rQL/ERRd5EpCVuG/K8vuHo+P2eA5tDWQz6CW5/+/CZejmqp20VwJCMS9TiIvdl1HuN0jALa
IpnFhPGbuFqBBp+q/O5/Ycw1PvObOiWqbqcUhkazt6zij6zlzsB+roG8jPqAH5LsSHB7sPtA/l8T
EdUeGyXeAbE47/N61hWuTq1YoCQCSdZ/HUDrDbeM2SrebUJSnpEfGZFrVlOiq3yuOxHV2JBoCeyY
7XjFKsEEG7/05JYCrk8lhsu8+qhMffuaHeTm4DQSC5FTeEfxyWXI2EFJXAH329tcT48USN6whxvO
9/XonxWZBj11tXePLfKs9c/ZcTPuKt9YMpg/jgGFrMLoPzqHJhpzxXD2vccT38aC2BzDDwtYGtm4
Zz2WAjUrG122izuG7rCNcZ4zZ2OnhQuY1LhWFzbXZLmONBtsICkmsLMSgz+PtCzTMCfk+qXyOrQC
kAbfgQsl2VeOG2lFtTLSNNQ6//xACPNhxPqlur8z1BAIwMI2LwBJ75TADlef/ZSpPn3Nl3P9ciKr
AGISqvfBVXaXt1EA8vC4QrXuDS6upfM04sxToSKrOJEmmBwmRQVQm8CEUqqnqNYDX9VqIaIKlZFl
yBbfGfAuLdygOVzMtoSxwg158AqBos8So/vQk45y6dJvvfrnHKRDw0BXcPiKV7jObj0bp/q6Ei9Y
watJYZBeeJ77UrdnRTdavUJx5cZY4zviRTIt+7N5yrhhgzMfYIxcqF6JufPBtq2+OyqcJd8Xmgok
aMNQ4DAFqYG5dPNCULWslL/pZQXXqPOG/RfSnrtXrBsxRZ0N/BG7WdGZj7HCW8O2TtoPT8P63hNg
DcCrzYW1k3tjmWaZ+dDf0IozG8mlgiTkwhsSMFnmFfospdUHxJPR2zOXLsreYHzmlqsxK2wAl8zx
f40LphEYUaNuP9cD0zFWzx5wjjKpEqgguUXhtGOZwli9apQJpqXHH6opJLoHRm2d3dBZ1zzZw7qb
Uq9MVEK74XZ+s3rqO9Z0LI/65m7Sm3HwKlw91v8AP9yv92SxYsy6lm6vc6UJ+Qe56OZXTdGezYfW
0aaiN4fm+tU5jQPq9NpZpGMKqC/OCGLeDQ2GTv09Pn3hNXIq2ecqLUz/t2HzE13VuyHt0+wmaEb/
alRIqfmrh4ux/03NkUjOkza3ZyRG5xYADlwawYHMo8wIOVYMDreqibYoeUWp4/jB7nLaNeZFsBp5
D0PVGYpWTyILc2xq/83pGtuR8aZhcviyI5W7nfu+3xaxZqU2o5XwfxLZMPLeVp9YwzKfbjgaF2XX
yqu83BDglOy8oGU4tec2EO3XLMFppSTYDUkbYtc/PqSmyK5SNpGjGWx4TzSgaqxNIsPguVV2EJgh
h43faFIjOLOTMM5BjVYwIR0MoYbuch2ZN5jWjPGJaOqnmdJzKBm+Oan1UVOwJPzrBCTsSmWzPf7f
yP7/SGWgbgx3RAGRKLhBly96APpNL/gIWtYFGeG1ddO0vN5C7vl/sqT3XpBf3ktl+SIz8sx1XU3u
xVd+32cvVoB1K4WWIPfCPY6IX2qfmmq4FtB3lVhihLGPlsBjacn7NxGZD4EvNeGgwKisCi1Q4DBp
Mty2VW9stWX/f9UiYvVSu521t30lQ0AG8WBZ7lkBJX3BYYkMP+xjpFSeGQ4DGHKnQ/kuCkFYFKo5
uz7jFrXU4XNI8rL2y84Y7+4DDGLgjPtpcev63D8HKH7+pbsXPtYJvOHkot/eHGsHFeIDozvEyIEV
2xzgb3i02S9gvD7oaBPscWXdeqHVGWXfQO3r2vHWN+/qvl+2BkzDgA7yRhaFbc57WkgITJMwAQM7
WDj/1nGJ1FMeY0m27lUwJtlHO4cDJWAKNzsdND7EGMMACti9ZsnDAGhMmo3VHlKQ6/vo1wS85yVR
7Qh+UfcwlDQoOqvEGfr5vSlpTzzmJ9RKbgXmYdw/MixxXAUl0qqebYbAxozBBzbhW02AP4nPmMKE
bmD/b0xfOTswFjTGdTKAOnm/NSMTZU2LbruHRej5HzGo5YcjHMoSiA6iIY2b+5sYGgnPz1WoUsw9
c/GnQoX7RZl4cVmrYTcjRVg81IS2wN+jTaQeMY0f5+y2rCNdGIoXTMfF4S6Kt0l96Xvq09Ns0H3M
bpEUxzuhWUry9eND2xbkdRK4reyIYSHM/M28guNmlItjxtqzLDraeKlQq2FmrxzERjXusVjmD95t
3bFlbveqEYcZQPMo8s4leTpW47p8flaYhttmtB4ppG0PTGtOezBBDSrpwjfAG6JGgPwTkax2PfIf
Y+ArsR+4k02HJQw6WHrXYD7knJkNJdcMfKdyb8EDkDPpOmKAet+b5dGydbAoep5utYZXc24dgSXA
LoADQ5q7YHTHiHf4WQ1UaYxqRM+GwTh/IBLBIgdUD2n9hoUFDVidpp10rBfxYW0XfzNgEbJtKaBx
+7TuGAB8YgPZoTnCSOOIY/otvMiNGgYPn3HeHNY17ZlS+AN31x32vv9PHhD/3z5LohgyM6HtBnaD
dO1GC1FePpHaJ10++KliMocSdmUogVNwVmmnaFn04jX918utwrdmcNPasb+FF+oEn6ls1JhFuYTr
uJa8EpUXdoVznnqbxUH/dHT2BK83P47O7+e96rU9W4fHaRJDtvx6Cvo/70fm2/CMCT9Oib74DRJB
4kxy06wFxhuoAM8baRopl2CoQrO1/GvV8yatuuRxvdfwXnMHJwfTNvyFBeLHsIscaFpNPoBMclUJ
vSisy7LnEjXqzwpqUFrsxy+bilF96oT0kvxzSUh4DZp6v34U239MjXIaOY4KLgAyJR+RxoSnvGrh
UqMB8+yo0tTdhV2J7gWvLPAwInsbHkWPA0EkAvNmhydxKRdhuYF2A54ow3LkD+9Gi8xej0sYWjOE
dJo7idTRNbj/2utUyIHIzO9nsaMWQGKZuAknyLU23OyR++W/EH3XDDBwYgF2/AN9qzJzxIKcM8nd
+jI21gZo5OgNwLff6T5CgIUY0XPA1IOpwRdhGxSTOGL1QQUEkrKKoekTzeV2df9xEHj7kG/YMUqx
MiwlcaRZAkyuHtZx7WtYoanPsckR/MHWRFGUxaJk+cHj9NZ156LHsrkxts3VvjfECNuUtQ8dxJ6r
kKMBjyFRlcAZ/vbM0n1+Un8COuOm5yc4fPgfsmK1zbBbU6VsxdOwyLcYP7RZDDMHGTegGNGp8iY+
kcQEVMerp/OUZXpPBvbvEiCpI8ltgZNWpRsLuuSxY4Eg/gejsPDT1qWj1SUqYdSBg4baNc7L8sgH
4qJg8xQU5IGhcZW552t2+mXAYWBJY2TFH9gzjsgEvcTOvwIblaWn/1QPo7L+r3dcRxNTuVleKdHf
3X8/UA4A0vQRiq/Z8DR7/FMRDUe09UoS+YAmY54RMSyz01VdS4jUrnkBKtKEmFuR8JMOi659GhW7
Fkm1sjGHABmbrvNljzPY4ASHozr0E1YuHMNPSmBjR65M/PNrHqspB0aI9FrOmLzZas7ZIC19//C1
Gu2cdUGd341H/Ck0d6RszoCJdrdbWW6Ej0OYwM/tyzQ/ZRGAhb7x/pp2IR6KmlDOocU/zZcoM1Ak
uY5xp55/k2AI+L2P+BUd1bqPW+kMKESOp96i3kyHJcednSgyqODz5mnjAjHW+vpxVclXX3b8txdh
rdNKb+clr/1il4R/C+9codpz1eJcEqEl/LzsfnVTPbwQYf36UppH72ah4Y3RkiD9NH4CkagT2ArZ
YpRUAiU7g+Lrp22JGKhx2Y0kk/BcbWILD8p3tTv59fZV8u/gxfo2ANXFppAnpBXDeIF1dExEYzMf
QRt0roWJ/hLoTEW0pn0MKFKG+TOhcf+l5AdTVpd+Z7L2IQfi8noCKTWZkp46krVVpFg/L/Mfbbn3
4m1hErkweJIahKr5XptKJ6Zff6fEgsdN+Gw4+s2MO3+p+bubQbIFunmYyIAVVMxSnb+cwOuhugtR
Z9i9XNrF66r0hjV3Px3Wc2KtEp9Mao8J+Y6VnRls/rPo8OqMjkuKG7XQ2BBOqyL15Y9w4ord4Flv
r+75snh9ZwTLfWkqq3ISHAF/wuJqzoQeEggzmDcmgu4UbPrCeoEeoKwo/+EtW6bclWVBlz3lA3lU
LJQYRbRc2epMR/OVJ/P66mR/sNH5vjUwyc3EY0PqXtaz1EZce3KPIWAWcRItdFaHOvhXFG5ucqid
MupVvXFGVmyg4708gIwNmjcjJk/m1FEJ6DAUpScsSNu6Z6ESAI26VBnNU3t92by+dK5e4AZEvhlA
yvZkA3McSM2pcdL5/pAdB0f5QfzjCoFrT6+aQka0sIlZFU+1nW47q6G3nxZIgEcvnjAepCm4Z7hm
uAelShcMaAc35PlXVjIyyQq7tNBYgKQlBI7wFhwSnR6Eemj/yAjy808WiS1UKjN+XjN/38FV4r8P
iYdEE0WAD4idWjzJVWk2BhA+yro2chKlj7a/TJP8/rgeTvQ3jDhKhoqnjiGpRilgn1MTFE0FvB2e
YQXOTlAg4M9CmEoE5xMNJHkC3G0fSJrKblYaX4Vljylu/oDzyZFxlZ1KBsD5FdEYP+bje6e4cho/
1U3C5XytMMoqyj9mqtrwUe5d6auH1lmjKYk3SmVLgKQBmqsYa3kuilbW1TB/J5qhze99VFngzpc2
42vsA0GV+vyvodo5yqs3Jyhc8SzoeH6Ty54ciUt3fZJ4DVAm0wpvC/hVHPeAi1o5BMd/6XtePDWL
Hc1yiZBi+UJRVpmEfg3QdAKNnwcreEoJLSeym+AjLxzGA572fuJTNXk1lNgHO08YgTewT0uGaPcE
fLUtjXyeRb32KZIo9tYWNP+nsDdCHqqQml3F90Mkg3D6g05M54bgmTu9YtMsjlllGF2fPavjxrrv
e3UFeFlb9WaA5hCELjZDFIBYitFVdC7Eypyq7i7PBzFrQ+At6RCTr47G3MGsJuBL7Qjj5qrEr0rQ
3ZpvmA2aatCn+VLx4mK3QLXLrtl2tOr5+dgxlrFmQN82/KTLw6iS+Ibml2iPMf7ewAAnXmpTDx18
6Pp2K5SHCnV7f1kvdIodp9iamOEJ/lDuz/eIh/p9snBCuTXp+3SfFPUiE2m0uJ45w8DkZbfWlhLK
CIhm6r9wNuoshzin1QOPkD7HQkDGVmopbk/IDU6P43Je/7E3dpYOoUngJtGakIfOchd8udiY/6y+
E3NQHgShBZa/5M2iDNRRy6HAjMNuvo3FYr1RLsU3CKqtch9H19bsYtFIQibaX062eUnGrDTN/0qE
PcFZqPK2WiCyPcAfRS/Thjv1tIzLAR96vmQDdwMF88+mKYWkIJDT19TRtB81RETpbsFH6/Cco1kp
mvw4cxe6diGcWJQ+B7niMTBMv8mnq7SINDcGkkhpdJuf1cZz+Fo8QUiXayr5VrWUX0gNIWQA9h10
rmm209Mmo9oupLMJgw/gK4q10DVFB8oUC8anhUBtmokzCBQLc66RO80r4BXoKvYHmVt4tHpsBVdM
Z0OlomhW8hlAOsPCswbPNa4bsXoiKaimotCNsZ782BXJklBi5gF9jEznwu2ZmeJkMSJthX0vebBG
ivEr1jPzn8S5V9eSOnR1Mp0D3Jgav77xYQa6ZATE+G9/p0+shkZKEmvnZJCpYl40fcxHh+5v1zSz
kyTVpRDNfNAxY8BdN/82qpXjODoab4CNnzWUx8eSw6avQetZ7zVpFTSkvkgucTRuii664XKHnNBC
SMui8Z7mMlYVVLskurnhFGB+p/s0aWInsGJp0Zi3V1fCkisjD98t/aA+MtIijzQQqRYjsv0YV3NP
IVT5MIO5v8qxtmPE/DwCvZaGrSvcVSnFqADPQMIcVKUxzlmB2JRPRvkUxZ9pWVWYI496eBXmcWan
BFbRLPFqvilwGjNuQxlmwMAP7FmF0ETZYzgcJr1sOYmcwXDNnkOS4vzRZ82OAuFQ5rTt3ArJQs2S
Y/3LZJAdbyPEAmc8CucSr9bvseca/eNKaP96kCXUVq9BzDQO3gbBPQlVsRg5siH4ImeuAN01jaXb
Xygg5AYLMM641dEV7YKYGdoocTZr42xi1z07FkmVgRMQWzgox9XwT6whZ4/mgfQ6SSlNxE2TN6+K
F6m+EXxBsDxQk+yMqAAAzyg74lLZgkruKb/mvLbfoR1k+leW4i+W7u1P5bkNcQjXg2j7hdIJi+3k
hKnYLEOLr1I20JhQLT54vy6b/HVn+ldqRM0rpyoJsXSJTTYBEEhkrF/s3xH5y6gANqk/KD5jf7+J
ZLGJZRyymhU/GDg14dYH1PqIKO6IK7IE1GeLVWY7nLsGpQNp3+cuHg7q56GOPBfvuEBNS1N6JtQy
Q4PHwE4YcXG25nuG2/slRI7SGM6NLmW7x5U/jyubndnwHtzfI6GhIrXkJRroxVhjiT3sG+15ryhO
5M7cMFAUKV0iAGtsiVUmziLm8y99Nmk9lBuipqKwERKxsQnzCLiA/EA8IvR6BZKC+KQM0Z3+dyEk
VdzBR7444tPtFp/J8Fl4J6DsxcZm7JrDsahuzjKddkytbi7n+KEhOEyypMdxNeycBcSgUxW6UL8V
xELZVbDsD916rX2eF4MjCCq377/mDGDRDI9qI2baO1eaOJ2W+niQDHs4NGjli7thZMieKzCjx5uI
2KWcZIYGFyApnfZcGzI8jjJgkb3dLDjMtowBbeoqTDb+hnQlRw1I1vJJmBGilyzhcGjWi5/06Ub0
F3Tq4Tb390MZT/G1jop+Fiu5wFk3ZHvxBsxO6nqGgvf4HO7N0mAIgngbNSe9FCBO8I7suP/Yf5hw
JryjGGQGoH2ruhOG1VO77UUCa+X1H6n8T6DkG6rBoacydy4xzRnwLN6vjjLTxQaRkUeEmiF/9Ns4
tW12gR3if9X55LnhqJDc3WHZ62K87kl3D/zn1CAz+vJNL1642oaMlWnjMYRk8kcuKTxND9vdasvT
gQEwBvI81/Va5ohm2kWIXee8oIpyRhECrOlGqCyzsgwrXsMIGMHJCiClKBoCRCFQIVKg+LD4/+Zb
XPxlQVcS7OuHS5TbEZ+xssFjZiEJkJmtxQ6MZFQh7pbM76bWWzs5Z2Sy+4qZ84/dVHxxPk7/xeyN
OLxVarI4UlgBK5N6CfHl9J4zZUmxKdCCJgdOLnC4H4X9fiEQ70+YAa46aVpxeNfPwJ9hlIDp/Mvd
Orx0FPiYeV1MW9X1qKaFip3fpTw3AuJHAIVElc0TPbEXL+3zC4l+yWhCWsIT/jjX0Poggblo1AHr
N/JQorbDbDsMjui1auOGGvvKs56+6xNb4d8qY7dAerkkcS1jk7lKTPnJ5QuUsuwdGLLnj9v1C0qs
+BmzbD4VZr5HzmKlbhHMRNyacmU6owN9/CVGD89VEqtAvqWq8LD/LBfmECBOsAFlqV2s33qdJyjB
WD8qlmNU/Dd2MvfBq0IXDvLXWFTdpfNzrnZI8ziFuMR9kajQnWmrnD+UeKGSpbLdWBA7mpI9h5V1
O4d3I//ujbUTodk3RuZqGuFnZNqZcvsIs5mQBMNYFKL9QzJPsjJUKvOwOFLNK/o4woHq3jTtAhyP
r00/MnBgejOd7dNgWgfGsVFDG6rTIKD8LQeYYX2GWeoGz4yBNceiszLtdJwrNjnZIQiMCZJGs0Xy
cs3UcIZ1sAKTOIYbVY2E0cDdVDJWA9k0JGX1a3AsyvcPxLIK14HSPxWP/uFt34u0VzxMvgplZeCS
AOK0zf3gHKCNvkR/F5m6t3Nmx5ILtCRKPl9DfpobMedkQlIQOPxQRSwQzKroAztEWU2E34Yr51Q6
KJN9EVxjHfPFd+Hzb1IUgc3tywgMkNhB5J8xheqYQG3uZXDI/ezh4ekxBd3Tc3UbwY2eEuUvDUD6
8T1lXotSvcJmmVIAfPcz+fkEdZkturN0VI1d72506PxFPIc6AT0IgIUtCbGJ9d8GA2M519QeSo71
xfR6MAqaj+KDvnO2rk9dt7nw/tr73BqWUEoar8AV5iKZGXkiXV9lmZ9mKH+2ZdpIyrjm1TjNgP0P
1cTNPq6od1xYkXg8dyURWSPUjJgiaDsRE8YnEmYV4c1iD1XvzCl/AK4GttFNjPUgxFYbo7NsZnzV
h7v/jQsHHxrA1+L9wDKhurXgvMhju58tDFd9jt3FnIT1j2b+tOUXHdnimOG141EzafcYYQ2jdOtC
CpI3jFMSYTDUa+oCOBpOVP6CeGWyiwuygH3p8OS7pZIeayvRdUKbFyyWLWRsBLYTOtah2Dd4y6zA
DKBpP+seYambSoCU0nuhj68CuaAw/Hap43wUi1h5NFhEvBdhSd7+jrQ1JLP05iy4ZDOh02RFLKqN
V9zuVT8zVLmI/RZkX76cDcI5nXQyw/f6M77/6EOQRol19MZs6eoKEiA46tQhOinBKCNxFubIKUx1
qTd+d+ATWwr5dxxaQ6Q+gk+Mmma+odXa12MjILzSIWLBRqAtYpHDkjKhlwtDvnHfk0AwfEcJXUty
Wk0/HY2xQQ+407CPijjTnz5hlJkyo/zn0H07lwKKKbv56JfW1bZwabU0yX9b6Sr5T+M/lqlzIprF
BVXGM0CRcKOOZMElbmNTY5LJYituGfRjjER5p9GPIDaior8moYSv1yH37oKpEWwZ01D7/PYQSM6h
eAYWyNY62M+RWCSKL/TyBBdNB9454i3qhbE/gSYvoXhUyeusj5YNv3oSJhb7MQzDxtJUvta2+5K/
zYZkZ4+nPoc+o2JiBrc/JRnrn9XAAORQyczdunn6y59+v+Nkat+eoHKS72hh1lFazQswCt1DBcxY
ecDUjsKcOI+0ctYPnBEzfjvS+uwiPyE28NUujI8xBkA9Wl3/hka35iHxSL3R3B9+ralPGjRKhasO
3QtVcHbVWJbfBWALLI5wvKzjR4Oa6+/WSAt9dmd5Wky0OzvqssQzL8ZOUyzZf/DpQL5Ad6/8MW9n
VoGMxkft8T1pEMDq+dhuUc3wmrCsH/4a0y/ZtHAlaWFEMiwc71uPBYzbhZOyxy9H0rrgTFtVyMsa
o/U6WWJtkkDNLa2Ew1LvhMjom+IpgdRHnTu66wgU5UStX97LKdmL/Dgw2WP9P43pyl0g+t91iFCT
rn1yIXUaGxP9aR/NUX/HQkg4cKdCN9YR5U1I88Ekkwid1ElXyUkGGwtEZ3qJWt6SZ3a1+dGWBgvy
db9CleSyQrwI0o1LuW6uFlzmgMVa/0PNDS7qeourInb++19kXhzXIRAAfj7aw/hJy3o5mVYRUhjV
GyZhzHzW1B1catLAcVusu1+UaDZC654rc/uB5ruQmAYoqUyEQWi9/eIkBQRciU7w6fW7EEWsZai5
5UdjGoXi6TX0IBRmnFEc5q/olfi7Unv5M1A4wpTn6sm1o4fF7rNnVmT37g8ag8mbW4J4SkxIgRPz
u1wWORgh09M8Lr9raRWOBZ7iEgwWc0S+ZvZsbwh3GROTG0fzeddYRoq+DOeB1F6yi7XDh9y7fGwj
mgqv6FP73+GmsRBRTFkATouXT9HsFum+tpGamJ7nHF9b15HIV5OVpbW5ElVb0pdIzGRH0OqbpBqY
KBHIDYrLp3ODoRiDXb7f+gMPpmHUhgSsvjof57ThKFOx9Woxz4HxpbC0rnTtrtTftnQ6wYRetNyP
DFJr8MF6cSFjVthMe4encTNtn3Nwpde2TmO7D84dBSi8aCnGS7yStnDqd/gGh0uKESiVtl507eGI
Wh8vbvV4SsHKN2BK8CZv6a9C2hR17j3wJ3b2p5wLIRLWHWrMdRKGQVmZsv1iX8K6MiqK0dnify1I
swuZ6h9RCwMZh4MclQ0Ooxy+DIajXXExB5zVeHUz1SwxieRZ2X0TXoJgiLqazXNjWcYCHhhSAD9K
3YspVuZXKezb1dZ36u+iWCAGSd2uMw39I87vrvcB6xWKrbYdCJkS9YIzLFyM57Xl1JrupcqsEXbV
AgOVsKSHyVPGsEwpgHl1Iw0jQnvc/sDjxn7eyTFMRFeXYtJd8A7pUDiv+Ij9yZj8KBoGwXrEIg5u
Deb7JWOOfDTBUcQ9EkGELWhV02JwjfdIr8ae9KmLTQjZY/w/SnLbwiw1qcYvR1YvkwXyNP+tgSLH
8H9anYu8484run26G+3e51mqm/j7LsRVrhRbPWFou8jL+IZTrKyaZdRTv6vOZuqHQbrvU90MJiee
hCTfZkZrNHAfDICkDz3WEJFl86eZ9OfTHTamj8d/UrU3EkIvml+VSwdos+CtUynVZo7oHiVXBIOL
Q6fBp1T9aOKucGcYUliHciI8RAAOOSLtzCRZkC2h42iNPHe/wMyBZFactbj0ZI9QrnDHhbmi1zqI
5VIHHUdOER+0pHcsBQQFGY+vI+T+TRNUtDAcTO+wLNookMgmgRnnV2rvCCUBMAUE7mak8lk5/dwK
z4uIuIXeJUyJO1UPo6sGHw4Q22W6pI3w1mNgDqvVCdkN4qy2eygPDN781qeNElQwVJqhvm/GQGME
U+kGP76BeEr9zS8j8ef2hTYGTQH/5h66S0dHwr6gyh8aK0WLo3pB3rhn+fVasN6Xc5UOx1e1pHIv
eYLkfBliqCEUX/APECp2zqSkcTLwTzhwrvuzRe0nVYLu3Mj4w8G+BhyU1WgR7RCHnvq4+hxvghrn
RluxDYbghSggxIgL2pEfI86UPznOzqxUZ48HGH+M8lCL3FkvQbmLCoCzs6GYvwGQljYDjJrS7CVV
oWaQ6uiPQZU/Kvn17XwBNd4Cp9kDFh36as8Gy8FBPmbfulpoyJdbxE3q1wxu4SAqafBTwac1Pubq
Rs0x37AnloaG4aVnRRfVbzrCryNvkg1ScqgjTvlkXCcBTAztSiYQV+t2iRLwp2rXgVNSFjr03aBz
NrqCtp6Lg5M4b1xBxRACsVTQGT56jYkHcPKqlgZFzCYCRdC8etU981MpYXWMtrse7xRX1OT1B7t/
abuiBjtaYbcEthCNLlZ55dVcm4yPviY/HSlwMPUcYSTXN3pUqvalpHUkzbtnE2WZ2WczsmKmE643
DwlZrbdtNrN4q1hqvz+4r6Q42clbfgsz9N2D+EeKjcWH9h4iHAfJqQWxHHCA2zsj+8O5IjRW1ayg
8nYl4PUGlT8y2Hy1cnQdYFUjki//AiAGWa+zvio7F+ZWgyLYBqnrttVMlaRoYtWkn+fmpT3HRG5s
JDNZonLtyhUFweuUU2GuPogHhXDECRuSIy8Y1V2TbJUcWMBjpMMcYGfUwjYzM7j64/Ng/bDDPsxo
bv807p0WXfgGcM+SPodGk7t5aHOJtIlWMT1+5qz2wQT4S0AeqLV9kMuaxoemBSjBbsaNlnUi0D15
54C9G5W9GRSnj7YeBcGUd51dMwgFboIr3iIIPvFQIJxkR/irhfKRLuVDBpafUvtr80s9TKLUCp8o
2NhK/8B5QnbObEBw53joTsqShfDM8M8hq1vRTx3n11btWdl+dwpLEo1SAfeFSC3FPHArempgvSTP
/PbH0TwEkBOgulM2OqKCiSzQXx9I3uDGKqguoN06Y9FpFCprOEFZ+LtnTuiex9DVnEjl/rbnS/p1
ldv9GLGtRhWxA28MU5gAh6prc7yiBh1UlZ048a8e0Y8kdsSJrz5LkbfbFzmmNdkb2GKhlNVKRjwc
fI78zK0YNMqWzBJxOQgTvYJEzJx2Ckr8AHtVmQ6HpS///SbqczsCCFfpGjKyE5mR3d5+/5fZBoN6
zw+V8BlCRFtmn4yZWo0e8VSTJfVV/wHjtdMr9lCcqJAoCizwIOrPMsOh4uW44SgfFUPMDZbg/7n/
VYKyrLmcp2KarQvPestpjioZIgoFDRBh4bzfc4VwP+nWKk50fERlQac68b0BvmCdwXpUbBnSFRaH
F1yc6POo1eG0FvvQ10fYPipPq7Emd4efdWHEjhAe/08t72yQoLBOqyd+mn/PV2ZL2DqDckb+2nzI
Dk5RS2Iug1cB/XsevHIejsTy4l03w1hKNigJryZIDfg8RTUe0jMuPeHwPPJCC6Qsj9vDYwrsfEiS
HH/iwHlXaqsWXd/Gs83YS7Js2Y0HYHyB263vuTeUbZtA4mVMtM5SPrl7VR3iDMIPumlsZQ4BM3ei
mNJqf3pjdhg64VG5zUhoUOG+oIUGiaJENsicStajW/3l/fnPHWV/i5HgR52PbScczipyqw+Rf2EJ
QSJsAhMggRE5RgY+JNco8nYWoVGSsH2J/eemk8OXrCB1OtwErdGXPeyds3armkSFjPBcT7bYn2Wx
T/aMr5LI7xyB0oIU/c2QNQK9lToE/FKEN+stPlk9K64G3IU8Jnv2yeKAe64wrfAQhti20/AYGiqZ
FriNgFiI/EyWv7zN3fVJfg7aLselKhBbhTyCSLMrp5RNnv7WhgYV/0jHsYhKuxM/eyqatc/IMPOp
YFZvSBjBa1jLIzluoD7ug42tkpSUWzOCLy9JaoaR61NzCunH2tneEA7bPfmbnhucutGLVTocWDDJ
8RkYnqZAec3VtdcjXaGNqJGpV2NW3Jq7DDa2l3Nh4bZrd1nFS+2NgOpBE+lW4oOqxzBDjoxNbyTH
UlcfOr6RLkyLEJpwZu/jjlk6eCNhtQq5jQRiY/xW8xE16+gBn8Ab73S/1pzAZzwpxmgMyzSVqnh6
UXDGeLJZETUTFrGMcJTl+0/b2+VOGKuvTqYHek/84Stk7BxnZo0VJDwabvtE1Oy0hX/2+r4VAw2w
cc1lw8pPSyCFetEPmBmAotaxsq3S8Ci4UemXw2D3iWRlwddJYtPIA1fv9735+FFBGGuoxEPj4p2e
GT6NX7ksrVZtU60c76MJMW2+fF/B505NS/rsmSPE/kHVMx7SzwiSd3lvrHVISz/kxenySC8TW/Wq
4uil8sgfHlvWr66Dm79hbeBfRVZcGeR6lABtZkH+jlajbR96HUGx/uH8YTvMIN5bkodPBGjoCIDC
kuyJGz9UnZP3+2VuGnCKCjhFhCfpce72mcXTzuBrPBvni0lt/TCSvb/O/RP1hu5J4T8SXM0jVUUv
fkVzz+JkUi9Obuk4caVsrdJJTCi9BbGuAh/ZXMUYKuNgqtLQkSbdAjLUi65tusFeO7G4rS452gnT
8IdHm6QcHjMYBC0IDyqvBTh27RWyXhs/xLbtEdoxGgogAnDp3u/AjoygUXbICmFcKBEa/mFNACd+
RekFBbiRmTY4fAXeX23XocFLiLBDnNPxXh57wETR35FXmWL2mO4tleYxLCYA5+9sImlWh/dV1KMF
P/S8LkKTsmtKiHGXXouNP0R2u93fxrHsKEib28CretWiV1VILXq6t3opBZHecAGxUZRL8urmPMq+
cdJC4mCv7Vz1l7W6VmlD6SV5e2BnQG0UEyGJdh+g8KX2BC/KQs+aaodskh2idd6Fr4Dj8JQIONG6
DM6jgVqsTRsmhKHcJEg4PIMra/vel30ZZCd+kHy3rmSHHhwW5vTC0cV+ymLQX+bAhbXmmC5rRrrk
PeRpbofSm9h3yyiETQqntVXfBS6ZxN22VLjTHvw2lwJogt3Fs1SdVgvJr6VQMplsVS9cNqL4IEXz
ZIdyru+NQyVnHsI8bS94vhiwq5JrUiZqCfnGa3gTj3M81m6U2qu0ymBHFJGbh7UhssOqIA9AYiBp
siorV/Ux8KbIsWAxmNsCDWlJmx99NWVRKWEG2vW67m5rZ8Nz7FEvIM6LETzFLb+A33BnNhCWrGNt
lF36E+TRsV9BXetp1uSVy9vhvN7JIYi/jNHmSNACMgyB13nh8plyZhA3wNSoilHLS+sG4cHDDBqc
7b+bk8dQTRm/UeVuCWClN9BIG9+vXIzRFpKK0DAVVX8HWy2arXEZNH/aRRlDMmaKEmHJTgKR5jAo
OZubUxITRVNm1fM6/urBwCPYWAikyQA5kfLDD7l221qvVsK/QGKWKiuje0rMTDSuJC5kWubmPb0X
mlfH5Xe8RFGmuSneHtEbv4tCRlAW87fTsyoxIRLbvxgRuN8JwmD+MizdlIDQMloHWSCeggx/m84a
Ln5Z/UIWudma8rXZ/ln5SjkSN+LwgXnKlt+M+pHmR7zxwo3hLGpYX7hvWSJIo7Hh7J2Cad8MRYUW
GvfqJAujYuoXWeEl2un2hhNWtrM3bI/UKgegKBS9Gqajzpv7U/bQE77et+xVtwvf0wCDVyGufV8V
Umr/uWncc26PBvjul22TTAD2sVOrLym5p3i+mMiNeo5eQfm2r1lKDm1qw7eWcUUcLP4vnKYtba8q
VAEsHxNCn4ibNtZTgwHEiRtL/5ElHrTJdVB6cZ63mZ/t3V+YfkRn2X4vZL6zErzob5+SwiQD4ikz
BbZk5u8i4dl/0Zt09oHVmnFmZ/9PKGFydWrKXcWpdsmxCe6pfJWS6kYjGT7jDjyAj6hP9DM9KqEs
4wtyscWvJFI0LSqYr/uXpcozMxFZCQxo7dF2lsP/c0y1vkbabFr8/h2wt9UgLjjRJLFWU6epNO4D
bE6TyG8qg0N05VQv5BW//LtRyZxVB4+KVqYZwLvcVynejt+eR1cVP/c6EssFr2grA/uuLSin/kPR
EPz4NgfSEmOyXhxnu+0PI78+LK90/Ct7GtmyFIwNK27U5jLtjbH+uF5e+VS0caONvj6wvjfz3io3
Tc4UjS51GhJIb7Xg6TY+E1923coQvxTcYKfpjnqSpCFiSo48FQHjhR7HBYcCyLq0I+SDF8j1iUUV
Qs8Jh0IHEUTLiE0uvSH58u2Im1ahVNiYb/OCeyRJiXfopitIfz1NSGbEi1rW22tVT9XIYqdNgXMU
yKrHKIKzGPJLuEAg/+/X3lz31E3uoxncC6/DwA8wjfDy8bE+Ta014LkX5+pG2TXtSRAZPqUzKFod
N+bvYmNuZ+mwBSvqk+M0P7qecOMqgPm6q+F5qDC/d/quN27kNR6hSUDSVQwyM2LoMcvqmQg+HpGi
qlSOatZ9IuZqrzWsbjfv2gqs1oK43RpKk2S0AcPdqLTF1gCSph+33FJttDrkymNdQtTgyGHhtCAB
tUJKeRsT48oAz7fQXF+kDz+uUsq76902ULDS1IzWdroKSm+DF4OKVK2EO74iFgN2aLVXGqyUAvvC
kuOq+pHF+S7t0e3OWmPMvTP0NCrD4iPMjIhiN3HVL6Wjnlq/2YZpKoiNKpF9NWd2OtqQ2PDySXh4
+ABVZBNh+KXyCABndBNqO6kE1dvXjV585XcgfOUqPyj8EYSw7MaTjct7MZiRPV94cy68fiEt1hwO
QSRa4pQAdRFq2UUnp193rsu1Uaq+dru99cjUyoVlZQs99JvU/MPnogp17S7JCLw1Sjl6e8xyXkP8
Nc6wPzDJ6LvS1ac9yiB+sFUlVV//tUVnPOlDcePUhHq1LQtnFERM6bhNJEEwRuEFK0aNKVuLsfD3
virxjntMYdspHP7Hd8ZG6ZeG3as+0B36KJzb3DsNUgQmnWd0xYk3M/0xLNsYpli4J6RaZRyIHWy3
zZrw9dXbkhBlwn5vWjbe46PTOIxjGIV6yH9UbsdbSTuwnkpJosafdyfo1IH6bketLVAwBWydOUM/
+0pP/E4tmXyxCDSCABhcgf+xtEfM8DjIR1sjPPyD23OxmModsXdYqhNLH3Sb/2doHO2/jofV45J0
9YSLUA+4FWm0cX1hjEgeea93iBMed0Lq59NwypxIRWVA1zv2vWQhtIghqa3144XRoWXtiirKYEEL
vnSOpAE6u0/r4tSi03UR9zniEaUpckM2TmPzv2eoGdpDCqnFp4s/Tz33f85huIlsOeGD8rIGtXoC
o5f3pi3d84ZyBTQZZCioU9E8WxxyagBPph+VXJgN9S5pKOWakikXIA5clJ0qE+Qky5eMn2jUFsni
mHxArzMBb2O9Vz8Z8QVyp8R3lVFZVLvzz2YlkUaPg/Ap6FQpWJ9Ay7AOYqrRIQit0FZ4Josp7sgf
+pgBh44VS2kMyW/nvdsWF3+ZULrSF9R/969M5Qoz5m+br77VKIR/IFBqEjcgpa39Q5VG7djudO1y
K2xkujF7YidLKmSLwsv9vT8+SBLqB2DEpsh4hewitCkby4jaIb2Z/13cDFZIi8QgEOhZmdNvotHU
ATF4BGsKfFtnqMRVrcrxMCaaUF9SNAM1Oqxi7UYUyomY1KZqselqp/g67kq+eXBAyaaBcacTR3LQ
oIzZMtmrW9KhIeYu0y85CIx0iAp5HKOZ6JfF9lJZ/ue9vB7RUwHdgSiC0nUwhg+07ebe5QDxWEJ2
rZWxyc+VdnQ1bw4qCvSYZm1XVgPZEdMcioPfcU6T4xrk328UKXKHPqyZpUcEfris+usUssvl87bk
1tD007U6bs8UhBISqPqkn64Zak50N/Nx85DIAWZMNkvMDgrdiK1whFaTK72ypPZaaeIXqir7PSAZ
p597yR3PLoCTNSnky0HviDoZqKpnqrew8fwyeFZYzX1Xzju6PiC6ZNCmIsCNo9Bzn6Kv0gbA+7te
QFBzxIYzlTCIArw1t6EVFHK+jw82LdKPOQqN81VeP4rhFMhb7DSX5mB0fLSA+dZZsR+eK7S1UJnr
6SWrVlTtcqovxALR3ndyf7fTFAEBLwLnMJJnIBi1r88HniR1nYluY0+wfjLWMDUWlaaZYKjz3eYn
eB4+LIOLqcP3EyS/RZhHLUHH/LFM6MlFklu0yO7N9rF0KfOrr87PkJeudkFlw2U36Z85k/Lh4zGk
+yzoul3KnsDTmgVOIv99Y+5mXxTMcKBNiCRBKX++fT/mXgn8A8gmJTROIheySsq5tI8vmWahL+vK
zvJNroAVaQKhU4qUSvmMPn9pgCxvlst44lIULvdhr2V8GmSbDsf1ThNsoW4t+g3/U7/sSBEW2DEv
KsnRfgE4V9UM10VT62vZxPQzZ9DjEXLjE06DRHEPuAGN5xB4iVv8HjFInKdtIx5jbxdQ5r8BnTNb
VP8hRejYz1kfyhmtF46UTL6ChkTkklCA0CX11dDBE6Of5LW5EnDo/b4/B5iboqa/2ZECZIiGS4Zk
fOaosvFM1ZgsmNeE/MUwl8Ti0M6TygvBfw4u/Yh3CapnaIb6gu4lzlDk1YfSRXs7eyPGd4l+OV+8
cgoxA5rVDYwHXTOcDDYJdEgPijzCYI/xv0QkVw0lRgnfTsmEbQP8FICzijE6fmoxQnqeWPLKYGqx
w81XJed6l1X0EoL4bZ9dnIuXKYe85WdnzhS1y0lTtDxgfo4jDsSdBPn7R07VwiXfRx5s8BBhoGrX
0QUgF06V/fFTmStMH3G4oLCOZuDTxHiebn1Jt8n08hNr8iFHr03nf+0+Gl2DKfIXBVCpOzY+DolE
zJMlZ6z/aPwIBDge24tgGkWIsjZMYfnYTHpHGA1XAMcTf3bxAWi09WJ37TQVLfkNEY/SthPX8fSd
Om8fW+tjUzl42eTiF9NeZRro7BsyZYAxFY6V99hRSt/J2temvsuEZ2pFEquzU8HMrEiEvcR/SD5v
o7t/G+DHH8+ur7G+ZRVP0KZw2mdMYyUi/3flonbgVf4o4PgYH5LG9pE5u7l6n9BDriTaTU5UhjjZ
EGjIKTtxpqoRL9xEusyrcFSCNcbLU0lko07k+pPFoNZFZ3VWq5vptTVVsB9aCUgEPY3ohdxQ/44E
41sxDo2oRV6e4/yiwvOLKJt1ko/JnI8fIulY2vy2TwSFCB+B7HLGbZRFihHuiwtrCBJNor4/4U7W
EOo3qbmEmAmMjKFbNf7HxSFiRvxldz+kJXSjeh6vLeMKzfzK232Yr9b2Qx6iq95lynHik26lEBWt
pvnTTxzHU08965Nqy8J2sM3XnpCztdGVXVchJyVHqP4bIjoZpxl78LRf1zqrXzZYUGFDxDcqYiSS
D8FFW2hQZ9aBIckx9nIZwSKdujipvShvbj46H8KoEARjKnr6DIw8Je8rLzq/KXFNXmjavVMvDe+V
NiQKZsQjM7Pcj3yPi4qYXdwwt7e7+apaei4V9i20uqfmz7ysF6Ha/Wj7MiQ29mChqYxLIsslIFxu
Grg/UEjNr5aYF+VfnJ3xxVA1KVjpIiWyuIJmNzrxT+84/6jyM37YmQZBGJkp7zICLzTzwRgIYefD
EXk5DJmvpdJaXRLulrmNindD6Yq8Gme+pg60yANr7sn00GltGMBuqOHCnKinr6lE9CfUjtNtthtU
VtKTx4E88r7iMAz1fY3bX2/LsObX8TIdWk8OHOJHHDYVZV9Cp3/LlT1RvleEThbEH+/oLhqz9NVi
ae3IA7UoJRM1/odWYItY/Zd0nj211nw8J1cdVu/dZCOm6vEWvKo2GHj+Ljh3M0RMb1hpySrG1/Xv
Bi3q21JYiFG8RkGwc4ik/ZU77Yoig1wTaoJftXxkHYNzFZf4eM4rLBkRPJKNofqDPtuA5rnlQwDq
q6U8OAH89D6Z2xn8coXO0hvT8hzAwzwceO9+w2BXT4ZUKvyJ10Or3y3Fpav5V9HYSlSmRzFSm1dJ
csNxkPPW1oRMbq7HwcRiFr3l2TattTj9J53i8yjHO7YBEfEJw2nPc06rIx1C2XCBp0YCCp3fciVD
qKeNrMJ1Ca+AK8HBa3TbX6C/eiD1Ortzhd5nNed8fdXD1GJBVMUPk+luy2jD2IB0pyCaoozAU7gN
6s5KhbwZ28RB/865jE5r2+kyIs/HjcsHhnonFVtasXKUQzm695vB/CdSTUgsPcvegZ0/HWk1gPTY
d/dldS3uqI3f3yZxvPyDbf9LZJ7EdFhJH6yjnXgOrpo4YT0siLEzU+WT+UU6jU1LjhuhBOi65chz
EYJHD+f8lKga2iDFwo3YtNWcCCoBUypKt6nOHyr7YisxLxI4V7pcSBQMrJRUtq42vcnXWrcD6s7w
hjc1UR3LdWEva5+9xLK6VSHD9topewPCjLH1li9eZOHpg5QTL/ZwvBu9PopFChyTO95DnH19O9y6
orT7MygTp1g/OF3SjQX3AkrnsRhwucVcumwvbo6tPK3hfSIOx/BiM1l9ByqKA6QpNrHB+5NEUH5m
aZ+oZPLnVWCeyaRkF12kVAYq+YLyHqCBxI1bNU09w1pKwKA/8AoQtvovh9pkVpEnvEx5Tf9InxWY
jpmwzTq2z+K5V7Zl3ULNYor8sBXHI9rNpE3COPhHKfbRjhf8WkdPJ0698aD7ibN9rEVjji2FRTVo
zcR/WdGwL843EDCQflsLOifQ2wCruu2ct5tLPcc3TgSe55VSPGeqW59eEmz1NdTzuMlHpj9a6Bkn
FP17es0yc8E++zi93FXjArwhYlIj/MvfSktGaG+RP/JWW7h9TO52eoUJIZ7X1rT7VfXvSedtqQH8
z8S9Ya/5N2WCXDjtKpn5KLzGaxGOImrm5xnG/YKSwG2+12S94RcjezRAGy50g7UzFgYvXivZ9lhH
KtapvUOvI+R+KcQea/sxVvkDNAj+d9cU9G3T6LLusZJsoEHlT2QAMt2w9anVRa5y+AibSB8rOthh
L76ybTH1RL+0uEetiq5K3ui9gADjnviw4CFuIu73Gr/6M3p2+gpOvlsGwlzoYvTXo43zTPX77wPQ
8bCTBxUyoTe5Gj5TVBFi438omVfBTt113xG0bwLs7xvayikP1MLGU/JzbT6hv9OmhB5s5RaZIqFE
7ImzrwrsYoxphnnI3NwJW87c8gAWEJNUPgOTFzJWDTW8C8+Z9ZzqFvQbfBltHJ5bAA+gsfJ5jwFb
8lIjAamYV2xU8Rv5W5moQT/ou1oIV+sh50/ZHULb2zRLEWMm4c92PfcQGGiR9SysdWgH92jRRavF
Nr1tmxkV31m0TvAVYtOpDFuXy6xPEqlE0Kc4E8v4/gghmEjlU7sUIx64klTL3bBuwncZc4nnJDHK
3Cjx18qJNMGgx9yZnG+bQAvX+dB/IVlA6Q6g4Ugi04gmTBmDteAk+hoZOPIIf/tEpyXYanAjattI
S3R4IyFkNjy6focorJ4Uo3Yb7QC8XQ+vnJNg9DhRMIhvZ7dWUxTNdABMYkGNa80gGHwipZGBd6u0
TMAV+5ibq8lbU9X9qCZUo6142wBPr+xv6YI5SRVu4ZJ6e3QEVBu0GWtM8re5Y1Xp5etyTb3qdcYx
BmqPkYk0mwtOJES9o1YbRbw6t5mOzu8CP6NXcl2eGwtqMvdmCEJSTSz86I4R3sqNC1k96Ev4nkyB
mt4P/2gpms24pZhKfrLYYJjTQI77Y6ivQCBBa9BVwVrXvqk3ah3poGrRn1fXx225JQECTr8ccV+v
kYKHD0bxLOQkt1lv3wIqLcx+EwoBI4DUnyFltjh9pUfNy69Z7f0k33iov9k+QIGWhlD0bDCtO282
UyR3SodHuma/mvpbsM4Mc98qrHWHu5e6r7aoYvCQRCAMwU5LRC/5IsDD3tYyIFG7Eg3rMu3lE5mo
TpfNUvXoCWnEoIXzniWR/gcLBMOxpmcIL/ICnR+mvtuY/0jKWSX7v4SClnGN6WEmHkDMohhFqHyD
9rKn0dB3+X4ZdkSitVWZq8sA6mUqGCNPYBrEuE+q4hsikkY0fD4/vdFguFzyTKmg5HbnA2DVY1WT
ivE5hZwy2ZKAvC0Dlxu+eWHp7lwv01uFLUtrZ6pfrvmYmJQ+HPM+s8Lxa2Q8yHc19Edm/qfqZbs2
QtZce1FE0+0poOkiiMCFTbVfacNqNSWXZanWKNFl4GD7LgLNrVSIaB0rJIl/O1aojwrnNSTynB6P
oYKA6fYAL/3u1LL3hpGOwh7o3+8GcZ/507HSfhzpMZdy1+unGgDMC7932GHaW0J6m+Hfd04TbEzQ
YgmyXe+nzunYwfYEk0CJJ/hYB2mfxRPwWcpXJ8hDOKFdNjF23FTS73w+17To4wwmMkBUAoZCPmwk
zQ3O3YqUFLxN/LgQ4fnyJjgCEh6vhTB9iqFouV6/CfXvwkc8rSozSPheC96bIdED5rGUI0ScUQCM
HF3geFDvHLUxwSQ+32glMsf+23BmiRP54aNITR6eQ9DngnL3bKrw5w+OO2crzd32E5qtjXXQxWw7
C6KlhdDN850uS4uAeMNince8a5zHMC+8t7rPB4F4N30092haR32G2Cg8Em4gM1OAnn0oqk+6TODi
taJN+j5X9Dtmg3EhfftjmcJsk8S/5oeBCSfiMXIr8nodTiBmULphz8TmrszY+dRnrUwx/r/npYhN
PQyhGjFkUoqyAIGO7ywdtsPMBokeJDMj3xh5fxtTqdkZrF5HjBTaneA3xRbxS+t+wM1nnBQZcnu3
T/P+O6aG9sfa3y4CRzmRYo3XfJgL6b5dom+Nw8hIedXCjXGBXIG7XwDrk2BkdnwtlOSxnPzQyoue
LJaxHIcNdcuO2F0Lg9Y7gxlGK5R84qY0hB/ZIPj7vqRmW1g92GJzrLHMcQyvz0N/SjDB5a++Trrv
TidqCPktctm75unzDFT4T7YVUE8lSvhcDPXlz+faleUtqVxZ6n7cijvcVibAlUtc6iZ/GMt4o4Xt
7PJr0+6W4VbADiOvvYZ15OhyAhDPClLgNG0nkPsd72CEqIr2PQvZ9xlYED2XpWGhGP44EK5Ozvcm
rL5HoCEOJdtHAB9IYH29t6viYMpbriFkjwCEFT09UakcNW0AjWui0SQpyCpudUIvNY69wAm4CRXp
kIFSjVIgKynmaEytgSUxXeZ048BwnDtX4ooCJYufkj8xvpg6VxlDSV49ORusqPnmIEPPHPLuy70/
nMvGqAMnCUlbhym7kkkv6dqRfqcsoA69TPAD5FRBXnDawA0gcENKxWmdpE1Nk0AV6qgUnTEPEPq5
X/IbhZHRsAKHcxxUl9dtqBrFCzI9TT95PeojHbdL9k9nA0VLUzo7pIOkLtzO3+Al4Bl9Ws8BN0Mg
P/ABqiAVAuTTYuKU7H3dphlGXyQbax8jY1MrDwtcRaYwSLTotKlmP/IRLJFFaO/UQG7N8/iDwzzh
gzttYcCXu2J/bJVQDH/zBQdGCJYV6aF993fTiZllZB7+UOlEI6yCRwoS1/oFuKzlcKzxi3jbJGEg
g5X7qb8vvgOjezPSCwlnL87Z9sA+FNX/tNdbxTq9F4cg3AuNO1anV6Iskyo8a/7xXatm25uTbQ2v
y1RFiDtmUyqakyL5ZRTW+FJs8U0L6xgmNn1dKdXI1KmooCeHVtss2LFwYBtigH3Ixk/hNZfMSHvd
pO9s4CZUDSHsvMYTnMbdVXRP7sPFYjqkikfPm8f2W3kA4QKbbtazQqT119Y50Sl2UBwNnJo6YANX
5Hi1L7nvnU9Yl6hl5zbLy6KtxH8YZQWC8JsJtbaQ3I+lVh9R4NsfGqHu8C9njPyY/bFeuXAp8s02
3ne5jtGt+J3m67vzbdA3gD7fK+Hx4ejSqLmUsqcPMskyKG0SxuyPog9X9iLqs6wAtc2ugR9fR7gP
mI8AOKg0HZHdTHh+HjeDz8Kt/TjU0WnvRD1die8cK7PMK2TP58StAIhSZco+JGXDGK6jCkLcWUQ5
nSb6n8OoFSCj635rCVxG1Si6iL5UEGdwryKkJMFY66hAbpl6b1vyWMKRX94wgzUwGzTzhiiMG4Pw
B1Nh5VGSaLfeHWL5gHay7dmugUxm8MGQ3FS54ISPyrV1f7TPWggQbiMWQJdVqKWPWlL1gQo/5gWw
p1Y73AiIhe+9Kchm9AvXyb/VJfL3TcG8Tqay247OdaCkYXnia7SxTMmOFjGJdzw9XAQFEHDUVGY+
a96bf2pPeW3+LcgE2ER+QR+vp+vymWBT9R6Cayv9AQMATRkaNWiKKVes0ZtRGQQ+wXnKwXDk/GZS
uBh/AL4DohKgcJrRRgUMVXkwmDsVnx9jas5TW3fvE+AME7DdX0PYN9fgpN7Xhx4yXHLXKYB3GENc
7+vWDiUJJ9ryoQR6G9lPEw9Lf+vaOvrfDK0HHkB6NMjymNIK0oLRCb+bnhpTSX0bSvWTkY+HQPay
OU5krUTaomoh2fRFDgsWXCxfCsd6u8YA1U3DDBy1duY+MV0EzA6Xz3cjF2yP5m6Dxg9qRvUxFeTC
moKy+8Z/Wvcu+TjW+5bXSnO3wnw61IfG6SFWcdYBf72iOP+4GCEIAzHz5sSJ7Mna5yoP+2fjQO9l
VZM2Pd9GXhXzTXcttp1PyV8ImGqe3GyrM038cqZj77+LkFl3hyWpU0xhpGC8v14Q0rJeWrVJV0Zp
iCEmc6mOeKvg7ilH0+jlGtH5RdUJTfZvfbYeqFSza+MpsUyXUR1P5bgUmYhuyonBt3TIaIQCkLuZ
Tzmovyuvex+na1aMdRKHAjyQUyO3BtzqwCVdhbichYsHEtsyTLvSim329AXwR4I6UmKZqbu2b5XP
NfdQar/euZAIRGJVC4Me6C3xtmWpMTrsKNRB+mSfYnV95opqz0m62SzWy0O3Tg5BxRv9t8I8hmG8
mdKxuxJBtM1GmLreTLqu0lk47ZL9XWh7shprg1OO+aov6oFcLdVO/MeJ0YJr/bCPr9hpiGpZeG6P
qtp/ZAFd+Y2ua0mV3puRcxxiJtr0qz8Sq6nAS+xDySUP8yv/dcD+0EbvPAN5Kt35g9BL2rhpcsyl
dH1MlgBH1jNFevgv3us1P85f1Um/WxW4rqfQCP2/XvLLY+20Y7sLD/Hc4HOWSNl4rzZSbQcu4Iq1
BI8bVZ09YK572nhSqJk8S+3sBe6wIpJBViH0N1RCEPq4msnLXXCXPK4mTTmcVUL2sYq7+GMyshVf
Qd/732aqsCcXodlRzyazJLNRcISCuRoSEyOMidsATRZNToMlQ7CMsXJUrEvxpy498WPNAwz7hqSL
yc6WGxsdlDn2R5oDY5Z3FeXxdmM8Ufm6SSOcYkIg5jRiHj6lmigMAHLpC3iUmpFe77rpON/lp2O6
bKht6vb7LA2Hb484z5jO7rD82UenNh/Om9tdEpIUjXJ6WY+J8tOJtdgTmYstDlvnxDxa6hcsGE7u
iLGJXN1UMf3bO99rMEefN66YnEA9qGLI/J5vS5R6uMqb2ebMb0cRBVGkM1POIInXhr8Ki7SW/TbU
efvRwaBxSl3pZTNhUG7wglc/TKkWkcK2QfuKEebyotjb8CL+0WU1q+zpcNhkJ3++N/HoT/rBzDRQ
xDH6mcVbriGZtB+w06SbJYsQ+kZNGd+8vv8U7xwvRzOhOoEXVv38ANf5pn4vZ1diaKyOx2dT8HpS
z+F3ytN2yaRkF7bzauPefeg+dN4lNRMKFf3352JlCOHO56sSQLuYb+IeDcWMhR6zZPNOJxeAm9Gx
yHQ6GOlGGrFTHU+hxTPX88faRbnXdlG82MPxSGnlO/k4ybpoRyZ5ie3Jo8X+Y7IanoJetkG6qprq
YMGa0TDDXLVJ8q2GS+Hjcql9xQVa61kTpjMNRwIFgexTQgd4lj65XCRaHo6bGtl+UX7AgDyfFRrW
XH1+xhH8LGavwRL++IiBkMC40VoLGJjuD3EXtmPVTACKRuJr3pIMzbROxhgzzYQFCAc3PwpnwOSK
y+WqlLzdydyq/JruS1NvS1mYBd9Fgn74F5gA4gK/ZTYYdpHah+8Y9VUrfgmwhSmiSMH2HSYsdiTC
kBXzy/DxkPISyJvf3KHiZDIcgtC8ftNdOVb7UawabVvtYdqKG74SZzJudaOsOV30gCmOEVjfW10Q
ELsmHjsNHKD+dMbMXR4S1hVvAk88jX7Y/x3ryW5SrXSPiKWK5+5TZX/W0bU4BvNG2llN4MKeKbgc
MVCc+p8OwJbOFnjifoVrchas4fyX3KSwKQnTEkxmZ/KYzvRQ8XkOokzMCsgrkQF571OkItZDntxe
bVMMwSMSPlsN2m2ogtchS08gSVeQirKQ5v5LLdjoxRnwjhS1gfN//aTicbloP/QxcfDfhMtFkC79
UbCb0M0EaJml66ftEOUbhh21uR+cQ5yvdIFcjyhQ6glRO5ZauULH+vSTtD7ElRpYyEULyGk69kHk
WAZK9qc4qty6qZuRBEHsCRxJtzmqFk/Cju9M8Ncp9UvZGw2fHkoqBXudG+CpuAqG6uZ3EUSwE49P
ojGCkVqvIQPIdIAji/hH8JIoXsb74fTCJUp0Z7vPpiO+ING2AbQPIGEdTR/8b7MjBpV4KhjzqDRl
Gj4ynBYInatQvYv05u7g8tjziZ7CXP3dNa8VPFW2WL+DFNL0p7U134weY4SBGYIl3opmqKmRlKJK
0KzapdL4NDb8yJLw9myKIJl62R/cjW9NVNX5e2qtn09xTFG3fqR6skju5oAA8kgUOKkt8zkJF8PT
RbiC0Mal7NnOHwsePSzYUqxCJUxbgush+0tptuGG6EkQcl4gAQBd0flPg4N8hjovRgLAx1lw2+kP
ggqA5E/XZXfOZfq8I45XjF0Eqjlj2CtnXLU3b0S83HCg2ksnKINkjM3hl6SNzwquRgrQU7zfrpKs
yT5ODskTLXkyZX9Ny2zbpM8VjeesbFT9vGn2Z9nbfTC04PBdtOzg/VNJo84/km4vYzywh5VLzC0y
kI5N8rkYNuJuhXKT16RVSTlRwC8nsCpIrqr7IcMwiG6pYArBRcf93u3SAL28XOle55CP0IfpeMU5
sWjeAbTxUcJXKOP7pUMQmN0JtUoM5GUWMnzJXFYzg9LnosNUpHHT1+8KMhM6ALKpHag/RsLSj7kl
YlAve5ef6joIHEcrhi8jsJkMj8sabh7TKwckcNkEcBLz7ygIQ4rcYzUQaVPj9HFoTbWlpHyiWKkq
+m5J9bdvd5fA8lHva+ppBbl/YcKNWCbwuW8O9c9/dzXi+VjQD9Tdq6y44oAWAIffa5+j1cwgo/9c
JGTkQ6EZ6x49HLh2+7aEQgsSM9MZrzxdPy06LRZK84yXG/u3t4LowA8Cie3xyOf2pXQhTFq6Za+Y
jRwHCUz94pzzt61ZxYJzspEjQFSMFR6Qi4PkGIuYcsuX+aoU8N4Rglil7LHy4jYKRhWBV8sRb3Hk
8L4rba9jw4dIY6QkEyV0jjyQ9hM/7iN68U4mKsbEyMVhGb6xPRjLr3DW7tYeaDWOwtsnYz/7SJeK
5W9akFAT+He+lVPEwi7f+/s/fsOxGdpYH6gKPEkQoaDdPF91XuDevXt9v6jdpgN7Dz1ZfsKmIZzr
jyRJCoiBR7trOh324Z0BR/TGEAZ6vhIer6iAqxT7tK80KyEH4RsqcPqkLZgnQcMkVqDlYQhLOi6K
XZrBz8ycFwfeNsRKCplBVbu/yLAN3MImITPd/9OfrH13u75LopTv4s9GU+IgRaOzChbq4tzuKAUt
G+mIr0DQGm5z/EjVGvZQ6qxNz3xRpxJmi5nfzEJJ4YTHRZE8w1pSbyeUC3I68QSMtAnNqMDEJnpx
CF1FJ9JLADXc7g+WGEmIErSWtf5UNWQjeKMxnIM2Rsz409aXS3h5VuW62soTe+ynGgqbXShB0fW1
gGWS841+HXjrmAfHz0w+qTUfk8vzFhFhgYzgbbakV+stZikyC8zamiJzWu/nVfLeQ5PZmvHV2n8+
xl9DtENfZXGaYLaCkYtmlOokVbF3ZI6THzJUseGO1JP3rkOy0/sIbwZU1n3VBt2oiMW0FyRG3Z6O
xWdJuk7N5Lnko53C5ncUn2rJD7jlS/EBVTcD7h/yq7kZA0MT23agFPr9dmxNOB7L57mQ0HuYURFg
a6TJ0ClVcKLN3uPKqK6tlXPWgi14pGY0Q38cNURM/STKcxsRDDNjVdF2Loq7dyzZjhlVgbNXWxv8
6hJOYL0JZaZc368NkUDyGjioCcQa8nbQ1++24AdIRau38a/kBMdvoBVsSvlex2qORpS5+Cf7Sz4Q
BN0eUq+JKD1TbAplMNVJ5VWGRHsAtNH4fJxyy1Dz9ek4Gq/wBLrr9fAaKI3CMT/7r3zuB4PWTlmV
GgJwCr8XHRAoZRHsj2PzzD1s/JCkwqE/RECwQsqvYrxZDoCGd3TOkeRub0MtaeKFGpGkq8dyNZ1E
I08KXnl/h8TzvV0PbCZkpr90mjhbOq3VHFNg9RH2t3LSm7Gl+J0VUQN80opFaXGI4sslVFM9LiT0
IeDDX2n7YK36LtbTtkhrsohevADG7A40I6Q6IOobtf/JqWJ6594xvMqQp9nEEQKdxw/+XkcXR5mh
Dx02VwGk6Lw2G3cHBAgv6DsmWM2aqD6pdb+UwxsgHaNn26kdZzfC9y8gXdf96ecum6qmHUARcPC+
HUiHg5HKtc95yv4LoZKGMHuhmIJieA/a0cTkpaPxdqqngqPFH2Rii8TBxFEm/kQ3ECWZQTKWrMB5
YEzuDsI8dVF/zekVo20HQKMsb32l9C5bpe7w4JL7rUMgv86qaLYaxtHcSo4pA/noOiO8xQPaZANf
QVEtZspxErmmQvrFErkRA6aJe6Fa4tKGAVdBlWoU/0mvt+qbBHIuXNb9LR3jMV7dn/kMK2OQKhtO
Uha8LxWG/nzgMAwCoDA0/iBVNMgTWxl845G8FajWQ3XpAt9EtY9AwuzUltpkJA9dGPwKiFN2zxqS
eBm2e91dn9MTLQ+4ymgKQP/IXCgiU1LtbB1kbiiANYwXK9MhQFntAtJuLQSo9sCi76pj5RBZsw3Z
laaFWpxPbo/fBvR2QWeuCMkK/6I/c4YTwEGhYCcjVhftkijaPdu9HS7JxVFOubhtaHVIH98ZXDYr
uU1ncKHCxudubSPzQzwSGLnU2nfbeDynVF7UBEK+92/NXnGgPGnvCmN0nQmXnHzc24ErAqMzssAt
O+FTcgXwcAznUhy5VentYnm9kGVUmg0fR1eDQt8it96KQYrf/oWgWR/sgrvLN06JBrLORheXNTgr
X9fP3HPO58uvJIHnGA/frYVC3IIsXFWQdeTiulfdQGubjBQRw4tIEXonjexoCbx/sqrF1bP+LEGB
dgaqDHalZHBId77MchdrDoquhZvg0Y++5qjj8em1qEnatH9CKromTd24KMVtTGBytS7mco9HfXm8
YxcUQYGAFWhKOWtZcuBsU09DPE/v7n5B1ESbQVS/gYgsyLDuy14GBpYJtdHAm0XR/3opa09THng3
p8ATkOjErvxCiNSSOBWVh9pE2Lu9XJbqwhhlahzXrHiU2H/C68YaArBTNLijd6Nb5y6OieW15mEa
4AOeqihdLvSORrldkf7pXTbgOjhQLdZTzxgb0eoxRRtG3cGSfuDmJZf/cDsTQC5uyeVMfl9dTViz
7BwkANYeuDxjWBo7pGUEPWoOE3Ksuo3gkgIp2kkNPUsCHTm+7a7t/eL0etD6bphs7v6i4fK+jN46
expoKWjIffPdazo9sZuksdIv1V0uBq8ErnEVNyqyvdzSOCCOHxfVpMwq6mASojnvwSpsmhjfzKVJ
CnUOZ04h1BDXI7WGsrb9IOZCOn3GJMqMTLodWTddPu9aKNZVkLvUtATAEXtPWx/wCiHlnB0/jgea
FWpLVO3l1peyU6YEfiwhQqOxF2A86Y7q5Yoq/GM4Sals5DpieViVJ6CE5sCCaiKi9uWwioTUU1my
ny/dHoGu7qRfBtOM5u9TyTM+QIBJwa4T19cn70DBpfdl1o6WDYo7c/QmlYyfjve0twMmEYGApShg
1jzKh5//Q5r8OykIy5U8vw7C2Iv/vYEmN2kgAjLRewDlUbzh+MDu21EXcKNgf5xEpUa6HPyererj
3Pp2K1f56fimt8ca4/F4YYcmAwqA0GyBNeG4RqsLNLE1xhq1RLwfNOn8Ti6S2FKvEDMigc/fx4hZ
KkxXlUsnvSclzvOrLxpxIPE+H9BmqGXqzYoVTBlTNYcqdhi6Dn0KZ6bbrLvFVhpsb533B8caKvtg
HGU27sGfddgMrACI4mkFEzMtZBP3tpLie5i4jT2lW0r5WYKCsVF3d1KCNcEvkK709Bp06TMcukGg
wcj/uHDZhHw8QHsxGFBgS0bjDC3CiwfyFpJ02P5rnYALohTbq8uLPdeCNa1tJdA8YZE2TtZXMwXw
SMi4qTVLF4WuqI+SdJVN6fhBNpYW9J1xPpbivUAQCGCQ5T84Vz8Hi0j/wq8/ZI6bZMKXPzoAgIbs
gLoaImdDZpQkW/qWDEd8erPrIsv7U2PueANOZp1vMSrYEstJ9a+kVO/m97ZhUQBCSk3mJCY8mFhp
4ofMw6Xuhl6THy2zU6go5PkgdWADWPT4YKwwMNAK8pqIue17vDXgFcTP8cJvQNKcAvc0GrdLPlEk
AgJ3VJY4loXHyytNp4I9JlGHCfpNc6Eus57+twtZlxCYRw0Z7Le9TkMtif5rGn1K9Xapt5577zaD
CfOmJClTNsBrFdPb8kwarwnShvU0og7ZmUdgAAKoZGQj6Sd073mjYiYqbijAsyA/0vZUyckfAgEg
xyB2DLW0T4bwuJ2tSuyLSmDMw5U/FB/+acWalrO6o1lPBVZNJmteszVDf3tGCRawv0DXavSwcq3r
v10oO3xiOnBwzQ+W54xBZ2Sz/qrLsTVqNDFbrJ9TrJYIS+8oFDTGt6IfQ/2x2rnVzVpGSNI4ydG4
81YIVT3aI++jmX9oUUPhNOmhVm8YJxoYstFPC4eO+0kWl6rQlkKUFRXy6yO8sm84oenwmXI7SAkH
IsDZCOW7+r6+D8attNJNmSyTZynn+IF7cnrQ+HMJJVRXpzjSDxFwyVyt3TeFJSIyqnO4I00rxOLN
lOP5unLn+q1WVgajJZToeof4H43hDT6BmlK+dre5oM9mn9O66MDZawOV/HNz93c/LILAbN/vbfVU
nmJ+vaG2HbMDaPe46+SmRUEKssjrwmuwrakik+L0IpaRWaPXY0t2/rAn6p38OzrRWDa2hQ6OstXv
036yLXgmQzPH+hu192RKysJdDPl97uiqE0qzBr2NTE5Jg942AslgABeKN0FnkkeY/p+G9TIP6b+5
YMZP3uHqaw3ek5Lt/gWF5u3G8k+2DoTdTlJi95cJxGag0crO6e14XkR97jTlmQfk5yYVAJYvPw2d
MkavlZrksJY3ugHrjpWZCq2OIzS2/B47VSoI5fuFOufTipERrGgrjo1JXvkZo97JqGtHQaaHzTIC
JtbQbynycHKhVV5YR6HbnBr9NzO0QLbCPryowXbWVUMWQWWDD9sGkRUOqjnKzvc/7V71tJ3eMZbO
/v9l4fVaeQrfNeXqfS3YCBWVXDokkmTSp+PWFhe81DNVTLEKd+k6Djh6hJUVLcl3mUOZHq9sKIwX
zhp6iUen87Ks62tNUee9rAfjBNZUWRhXlwHstiyCnfPx6UN7jZllMApCG6JFtYlke80WXPyfR3aE
xsxgmEbHxQqpOAVpPrcKnQoL09CSDEIeTvXnAbbsrP2Ba3xmPRmemJXvFOwmQXhqQR3TE06lip32
nnNNhTBTpWBYnmI9MDLLAkIJVbEGWtK/YNmTELklEkx7t5TruapEcoH7d6RUc0xWwW3xqZDoeSb6
5PWrpo981FPDMjiVA/3QxkQOw2ArxNQ8WFD6/mOqnkqHmQPMVMHJ/oed2L2rscZ15nd8Hvcj7iFk
yOvUAMdHZ+v8n9Fs5j7f2uTA+UukkANegFwF3LoAsWwBWm0f8tS8eE/u5ZaqrcoT5a2OhvDMv6yH
IXYxuTDX9o6tWKp10+V/GQci9zM8IGb3H1fe6iacGneJF/f2scvMqMODpg1AUBimtQDjJDwK2eDy
X11aEhmgHH9sMsUHtRjKiQPriBWI42jWvJXOhmb884TIWPb1Go4jaeb2R0ulFwteovpIuMeuT10n
vjWBUqgrlawt17W20jotlyfMP4+A3pJNNnqoWBjDJ8vNkE3f+AeltRNntFORT81RzxFyGz2Eh+DO
cF3zvYo2qzpmR+KTuTQLNMMkOAPex4x2XXcy6HhvWZT3NMHJLndYlLoQUt2mMlnhjqdxThxu0QYN
RI/S49w3rIEoDUgHmn7neDBvGPk1Vdwr888Qqkz+z0rUVtvMZrC+4ukVKeRSPsXa0aWO1VpSXCdy
j9advCXoiF7Oj25aKIFUXaiQF4Bgcv+ea0WhuPQsobpB3otkb4MtcbA9WQakpZmQqchWYdYj9nI8
SfXQb6KRc1chNyaaTEHzElaOdZZbW0o7+Y5+WSTOricrpEALkgUOT0m4S4tqGWNBLDMVabnwu+u+
piXMpXJzpVrvhJ2DZh+/Xkt0N34RfA8pNZVEk1otwVpQemFHXwUXfkq74Bcqjj+XmBUaWSfAlUEd
tGJ5XFr2IjtHOQWTQ7RSsiO6ymgi2MgLs/g6cZSLNEU95zEW2uefNbuFzc0ig1t5DKW7rC8JJ+Ju
zD1539D0DkJe919khkJqnRhM/cbzjFFK90DG4XJDDQe2lrLDdv94yZ3fxKkRA20OJhDvfxPINxZA
2X0C5ZDAS3Ff93Z3LJYz+ZsuwVicsTcYrV7z+BptGkpRMhz4/jP2dVTt6hgf8yvrOrxKe0Olcar3
nqpC2RWVnSjf0gYjEZBmqci7QUGOGsaEe/BARXOpkfNp8/wP0bzQKJW2UHIi6GpMoQ6EObD5+ChT
zs28KVj5JTHqxuv0uM48iTxwhFb5s5TJ6QvjyO1rinGXIWw3B3HSEVzsmcsXhdAfOEpfhMyP3iI1
us7Bk5tSEbGL0W7MMhrEyZAZXhfqbmArU4/1+9NEJRsubBLRe32UyLrIb1kzE1bfFb9zPjc57F75
/eg3j/NZ03jeuIR2QjzvqKfJchpAIJHctXaQDOXDZq4oLzHUkyAIH60Nt8c0funbBaEM4cLDvpJY
hM++8/E2v0EfvcJT3xAmo3nUItxnGZrt/677IcyVnjT+ywzjk6Mi/nRreuyjCc07FdFjRaj2c2ve
GfjJdMGAuOjLlceVmB5r2wcEpcSGFBSYkHvvnQX5WUVv+opuvEmfjstXCmIsR+4SLuQ+y3JKPzft
IeK1qIpFphx+jFZqMHGhTpr2NYyDWlRTe07vM+kuzBtCNzdhZhwvCwZ1DNdF5zwyYordgdCz6SSy
1plLWJwZTh9JOGNpYBp2RRK9fIhx9uDfEQxlzu3JuFP9ZuBCShBCcATWY1SFj0LR0NO4vf9m0Tbw
cHvYoQ0ips7lgPgvRWUu1f5gXpmmXutXHIkpcDt7tqJ/lYq2E2HBeqzDk7cG45f24BvGL5rDjjue
JBu9fgyy4YQYHHYZPCPNGNcg2/eSVsoxC7tWvM/4M7Q8fJGQ6+Ab7mbtMwePjvc2H23RmlfZ4Cgv
P/x6MyC7pI9hPfdnRqXoEv4Ui/xM6vFY/4kzcPPrKaJp4kkJfDfsqUz9kVJweIQD1g3OfVWvJwU0
ZIaHm2afO+OCQz0zwVVcfuCpav6ll6mlBo8PMpXtjduIjnUbW/94fDU/1u5j4j6Rmkscxp3ebfMp
zFZqALm7gzXphuvCzYYH2d0tBg8uvPAOXP286bQUbJ2e1lalzu9eImZMaJc6j2dZyxjP3ybsSF3m
VnHIzZyTxc3fudA6UyzJxIJF2av/jE7EQHnGcgpoldaV5QBgPG89iuqhWJO8NjdWWtONgh1eF/Ad
+mer6i63Duz4nGpbFY3EwBy5wLznFOcuAMdgvT6Av3Obtn1gtRnmsD75BvCTOxBROLgJBsTdwnte
J1eVlCHpADwAuArW2MYvXAEAGW9u8EvsGHcooFHiBS4wtQ4FXMdCX6/f9uUaC6WPy5GoyghOTmHC
fud3V/gtWfCWbLjVQdbyvHTAOceSwGQ94lxGylLgyYpMewdMEJptzbaz/mBqR0/YaAwcv02lqdZY
1+QftmsNOofR3tdE6wrsW4JU6+HkTGyclruyUkOgtHTvFh5yK696STEU5W7jpvoXEopMja7XY+Ej
abqwgAu4hpTk1B7gOnxg68Izlh1yX6XCW0x1U6K+/q5WId7QxjRdJ4W0e8NHXSd0EYd6fypb7PaF
oubuvQ+7uq2wIQJT35lKjpqhgNAw71uL3v2fgjgG0Z09ZDKs8tM+GQb80tNqGv5sJNCnl99MoFxw
HGzbg00W6A0MFEipLSJoncAp6iU3/iKwltJ54j1onKSUnuwfVPi12Srk8gpB2SqvNnA5Mbk+Bv6y
X1lGKqdYS8VtpVcFQHwXZAzQI1hkQU7O4B2YnBF/vdBSOtphyJ8tI/gUFQYnrl+LEp7/oCa2g40W
9PYSyA5fWDwfGLaJf/B4PMmp9xrGecZg3PDOQBcrsBdVFFnsN4121Zu4RqPbpugfjNbqroOEuZHf
gjGCZcWE6Zf6FG7kopCH/H6EG1e0+PZADTETb2Ob4EhFjwrmAQtcg9Vna8qirtmFyzR0ZQYaTlfq
etQenbJjBHhb4zjbWEVNdnqPVbld/YV+BM3zawBT+Rg+H4/SKGIJ5EhjXLVBHxB6Q25Nbi+iQ8l3
vdFJXEgExR3QuMp4U3L1DOShttvi7wOnnQm3XbcZQV4Zak81dcS7AwrtN2n2xtdDX+UWEtEPsOkW
suBn9d17DWNcuFy3DgUtYQrXsuFXoSNtuEczSpfj72y3MrL5pOMWyT+9G5DjvnyCFpl7aNOWK+Ch
QILxxZxH98SX+O2FTyvmFSsE5lf1poc2Osslxw8lndEFGF75xGd0FRgNSRr05/fokqcQDN19So/x
DrAh1kWitoI4hyZZDP6mFSLNm+FtzIuM8gq+BqI8C2Jh2BNzE+H45LQ53gd0zvz66AGNJtW96REF
6rYJb6AOxOuUBSZz/gd/KdEsiGJrg2j2EA+lkSnp3R/GkAHQWkPol4zNwP4oxbjr7BPZpOOs49Oq
ol06vTJbo4S7kArTHYoldtRbXkcccDZTnqgF1wbDFOLJquEe+12JQ1GjdQVixvU01YI7rVi4PZoV
YvnHNWgr6djtAmZvG8yUpxIxbEcwzWhULea5cg0PErE7rk/dFlXKM56RJpRs410CYj89HjqxnECK
OxGyhoFIxbXi0NbUdpxtVD3Q0rFKCWS+H49fpqkt3fHFtaR1RKm2Dl5IwB99L3H2pvYfnB4Ph7I+
bXnvKx0+qJhETbSc9Rp2aOMN1zELtOg7FkLiqvIO6Go7JzcZvtUlRhPAJi2IvVFNvlgaJvl54OSm
hx1/ieD7SDY7grNR46sGNXJHEa/xibpSDhbVQMlZEwUiprZTh0Pe18f36nR5GEaMhrZE6bjrI5UF
pfIcfjPhH6j1/i5AFZEiN3b9gbeVYKc1c1uV6s5GmLMO0Ffq7IhVKxzoL1GHZOIzxbSu4n8zvaG4
Y7AfLoqorep2Y498nehK33K98xjhLykomYZDkr9+HDMClc5SbI55mb21qDP5et3c8u4gdsJaMp11
fztVCYljrYt2knAV/EQGQwlZGJjF4rpAi0rkKRIylChDd307ylF+VJFn+JbdY1Ws7kEgS9YWWKG6
gnrqVKJFnoSO8YEdKAUneTa/afDSdiV3lM5TligBRiYH4meYwQQ3Bo/tq03s5uMXkMFc2ETC/y0i
PKmE5+MdJjd8OClOEcZGqUoMD08nHQEm9ug2PAbhqN6TKiWlH/OLZ8w+CZVI8HK3CCvnO5pUjK7r
tJ1dv40xt0sVdqMVaJvI6szKpMwmfDwVQAqkAkiL3RyQy6MLG5Tujy145CjcBrF2dXKshwdgiJ7m
hY5dJhX9Dw+43HhliNVvIVi30XTlwr8oSw/4mrTthl/tYwnmU9UCKQ9B185CxIO6VfNvQulF9i0v
eshxeVR32kyjJwH0lGDFA3gJoIUwZIT1W58HMaOZDIC8l4F4N17hgXknZL2x/sC+bCeV1M4ENaD5
DWMf06NjqYQhb2c5FhuX60rl6YiBEmGPoZpKEjl4xJWhclFw76Z9R05VXBGJB3r3qn8xUh8Xtz/7
M0rBPDqz/3bvjaG/fu8vAnCusNsxVpsWSMB+efj0osPqWD2nLpxqgY9s5tA98SAgFtxbETvk6B0k
vR1j+s1ftSE4nRPcb9l+/kT1EKBK2c12X3bUUzFmFH6gBFpBiK56ThmNNQgwnRLLHIdAgeD25shd
12b9bQ1Z9FYG0us3Jo4iCkz+s0be9mTKghOszNHwEJ3LI6V00mhc/lBUzCSPMdQRmqwG0E51kdC5
eDbmUqL187wPcV7ISvhC7RpxfpBdVKTb+TRkNBQadVOnFtfMxdOjb2QJ7paTjqPaBttqGM4DGOSb
CET7fEtT2wDyP+OI/arHH8oTQ89izYvoRLDYsD1brvy/F9m+0PgmawGgWDkTpROCYYnZUela/Ude
ZR224vGZkIwfa0pNJ3e1ZDPAnam2FNXBdtKXjepr2OEnyERlDNqdnIAaW6o0qQWj+xTfMx2afaM8
FajU8e8Q8STWrU2LW+dJJND4VxgNvbjIfuiW0UG+N/Wz80GICfzx8xhcjQLDG17MkpkP3+HwBOgf
ilwRPRVujmuskerZzL+6L19Gzpsas/ykdYAjRRBUKZQKbPCPPTNdaJOJdGNzW5LlxVespfkBe+oQ
jwt9KlNbpJvnL7c8EJYt5zbJrSiC8r68McEXguAmAHBjOMr33CH/pzCGdZ7vh1YarQPaR4eNsPNC
68tFIF3Uqijf7chA0Q91/eS7py0HAv2p8M9L4qk56MvEIdYP0kYOLufbwIGhU7bWX4DJ8y9izC5w
/K0gRKRMNqVPct1UwJhkirFM9Bc0abJScoBHU1fHQWidA1GCFHf/zh3ZBg5bQIBehI6PehqlQnqW
oivYne5LC95zHygpJ8LFn57qR8O7vcJ02hGtCKsS3mZmommjkM92mxqfxjNs05RZV7C7E6uCzVHi
UGyCkHFjJFrWoSaspIodgmwtBZRwGDOCQeGdGB4WeQlcf+dluECAGqtO61UWiSAnqf9HA6q/ukQ8
fR6fShRAcJD2y8bAY86/9DJYzLsnVDRZ0yb6jtis8w0oQGrhqBvUrIU67G8auzWP4WBos1oS2a1+
WXOw3dAOc3hUS2KejKXDgd2dGnAG8sLU/zFdVMMpk47Y4i60jSYXDPny9hgd3R8Yv+F8uFnELFPc
uYi6PilUpBZjNWSJ6t0ju5HTUQfa3qIfhvgx4eSGRPxZJ09wbkCyp7vwYhEGE1m03xUAcgdYrCCL
KjsV7eLyrGVEgRzlUksFa63e6k4v1xbyzIa4+mX3W3fEhrRATbvVBSrxeD9MLgybExQR9iyliapL
J3pgr++HNbK+UvVFGyERlXXm4Y0llQ2Y/x9YJ37/VS6aP81rIXBTbA/lYGOi/mQMSznLTnZyPJtO
4/4izx2Zc3pdfMSqm2iJn43W4Pk7VYfWxMJYz4NX8dUieb3Tu+FotqxnhqKTkGDxY3Lbjry0txqH
o3G3u3tqqC5wJ0GP/g98hiIJHeBUw+UfuNjOAuvCS7TGrUag8qbr9vpY/rMSPjPIhowY83L6nmrH
sQMoVWPOO5slceaZlt3PdOG9SaCOg0BfgWHR7UIgkfEb3Mw00LK83dzcYAGXogwLSgT9who57ElN
R1THCDHHDP8B0nLN9LKjaTVS4Qw2J4ovewyxWWaco64IZ4ur2NL7wgYqIbJBPprTbCy8EoMr+RZK
4lJr+PKqtixv2cPgLDneGqM47/CM0FGwVg1t31nEFr//oqAuL2aW8wKRuuhSoWwwkY/0V9erbMFX
FQgBBbvLpYiJ7+9/DAAJIjbrgR6uVl7sFrW9FHVnvhplZpYzjC+H99WJzQAP1s+t3O1saDtiO+It
dfvdkyFKSbjyDNhhTSH1UtyeHlVVEIcs0Qq63t5y4uxcxvDcs3f9Dk69CJK8HPwoXmx22vsOltUx
tZoLPijmDSfDlkJZBxZS+dUdo0b1dS58a+pzIw+CGubWMkNd/QXuosatefcCwD3AQtetxvZYmt8D
xSY1juDCs1jvggthgKbuFl+QSXYLIDn7IQnfjcITsREIJM7A8WTbt9Atvx1RB/DwxiuauwlXqKoL
JBoKda2QTk7cvd4w04/DbIESXXnSJhaEbZYZQ68E1kYRcodLACcvj9CZXedDbBcvZn1yBGIKnbyd
L1ALFTcT9b6NsAji0/l3+ATSj0Mx/n8k1sCqyDVJ9GJDROrTnZ8cd+9W0S2RZzTOA8C/7zE9mDl5
yG+qBE7fOgEzRltM72pmZ7PwaEL1yTyKdgKlbecjPXffJV0WHUqlWfuUfE6gnjqnbexQ8wtIJefn
hXGv6JXg7Ww1fGC7MnjAWxVonFHxwZ8lRvccRee1y+oqAxbhOS7skVZkuFOXJR3BVdmR5YG5uIwt
m/oH1es7mJjy6uMzxM725hfCCNj09VSc66WRwKgnOYHy+z5KUuG/AUgu39U5OXJKeyJXloiN3TqN
a7metKTCFWs/Oc/1jQWBD4JUQAtYiVsBX1WLG8ifGTG9sHOY3Kn7ZGrN+i+qERDDQ4K3rJboK+6Y
p27fPsJCSoXBlDt0oBx1voonRdlHcdwF3+5jhiIvKJr1Kd1DpBrSUvchvCFS56AktlGAYvsGG4om
uIyNaYpEzzihjUh0Ra6rxcFaq8qp0pNB7BTiUueEFpd99jtS3cfwYGtXmw6uDAeXXkJ7bh/usf4M
HhyQZRQ0WDxt8lZM9+1wlZgv/3NYOtV8H19hhGI79fm+AkhUiwwOwPEoJBlXz0JZpdS1ZKDz8qx/
wIwI2+3FMNoEhNka2hkR9GhAEm8G387IQQ1KqkojueDaUsnnX2WZUs56+yh2l0zpmEMqrZ6i5Clm
KYMrsm17A8xQdSu1cJtlr99A9g6bpj8K/4UEYxvxjbhDWIhUguarT7G7YCOtlXO1RrgqySAF0a7G
/2FCBDPZelXLpi1+ZrlBAKjg+QM+ewv3QPcegrpSb/m3LyePugx40Y54LfVmFw44ASyI7IH+AW7I
4TrgcIPJoIz1vcy74NT5HzpS/q3UmV+YaDDpK3n+qZIkpLCAE8KVv0SL49b9X+CBnrSdhxx6Ws5R
r7DNHvQ8Ts2vtg2ci7perQbp5ZdNtSc0b5Z5StoyeJ/SXbT64Yv9BOH5WsXXUZwPCOXXVit3MiH7
EqqUi1mYt1B+aUaKck6vtuXSUun3WcyCmCH0xEtnBTQaQ+5O+HEIN0ouhGbLYGY5JGTy5h9tYWu6
nhOL4HWTZvIqqdzM471jSsA8XUi5bpR2JlY2j4+e8I2fsubiy9leaHRbqx2bLPS8U4BWwr8H81Hu
f7lWNdlAdCcTGGKZev6ArItts/qURLLwThchJzRyd4Ayu0ubFh5tF3koiyxUzmKut+Xh13byDwXb
WVgxnFXACzvyYlObq8dbkc4lf7QzZqvb9gjnu9PSbbWhumtN5AOLt1kiEpTRQZZupjcisPoxBrxq
WqSUXBlF/3Kf4ngMrN/ZcGuBsvqzucOboem8EHtWDiF0+YMHoRx8GrPLOADKCrO5TRSHx5lOEx32
jiwJUm6MSRqydfLYayUzH2TtM6WpTfjE1Dvrp3fGVj9XRTzhVaL8sGM9J9fsJKeBFKsIz+5WmWtL
Rw+JcFJrHLKpLGX6t+pX2zQjIMrnVdbIBLV56CkZ3O73nQJLIQpo5WQUmbT73d0aKCESaJvfhyru
9Tt7kYT9UmuGK9MvowBOZUCeMUBZH1JJP138jVDUSCuoPWJApUjsngmlPv9+amaxgqQbdq2tfpmO
xyADOUtKKQysmJD1g0hMIuYSZsfokDNVlXpjyPkZy3DvK1Tl7JI2KBJwnqIBeGRJmWpE6SRNOknq
HdtDah4DaMxMHIULEG/cdMWHCngrbm2iddFySdqV2g9n2F7pR3gAAe6quXMrI11moN10ePUnpiJX
lU+8GxK1nCZe+YNkA19PRfB1LaDFg8LdfKENukPxAVoUDOXtcZTo7UCWHTwQQYcRmE3LzegGjo/3
zeXmnR31pvnQ4P5shmKEyInZcqXqYGoCBu5DWPfU1/cZ3Kmc0HYlPCeTzHrca4zHlUBhEK8rzYwo
o0g+xmnZaMWLym8XnH21bWud6UZtaoJZD7JZjgD9X/SFyGX+Q+QS3DDNIyw5fkZTpgYSaQolQoAU
QFjNOosJIZJuKNiaoNA63Tcrgmg8OMcM9Qi+Ri7evpXGoHdDJra+OK1nc9/ylyCWcbPNfuJb42ue
h7tHdvdKJH6AtTPBJiSK3vV59dtx8AbEEnv95iDnDWXCh7kzVzl3TecCaAsqQiWH8gFaWMJOvQGH
kaAb9oxiRM7g2k0LTFvhvBzNlBEXe933GgAzUoROqQXzHDS2t0IemP7/+4oCf0JlUpAtuCkFaaw5
P7cIO5cwy11zLCy1ij9qZZ0592jpqnwLLaA5v/0BLfeTTCoxJBs+vP4/Lf01aKFzHvskLLRriiv+
vN84hnRf4T7JJb/SnJtzlBt91i6ATxW4i++FMIKtIRHplWFDbhftw42NTLBHtg1e+hSfPTP3+m3c
Y/JNoEkVYo0+ZavKkjSKEZcdQWyKamNWGjEyiCtMBYkw2nYXVpJ+3HzgpXuOO3+UIs4UH4VknDG7
NNAKVjJf4gN0Z5HzlG08ivmsmmQR5kmqWin1Z1fUj5eoJTp2DyG0vXS+61QwCD6g4z3HZK4BtSHT
IcD/J5EIikXYnV4Ib2EmaPi/2hxOutDeXLskGcWmvWMNjEwbd276EMDyFg80b5S9WQbYFksbX0iw
piISjFK/fKkuuCDhB7TcpdQPdFpT9z4MmGbIXcQJ+SvBxq2zLsJKFOGOnVfUOhf0+SI+k3v/2jFh
ocBZ1921bBWP73RDUWZIc2chG3eF5pufUuklqLsBHIpUlaBLebDmxG9oUqdETxno45P/H8H0iVoh
UqnPnd/lZ24hHgCjvQduRFknNIV189jSQMNP8LojhNAcyRy16g7ZwxY0vRn4WHYYSXr04IlWVrnK
CBkPXYGxzFyaFWqlEu0ct7T8+y2LZQeOFzpJcRiPyOnZHPYdXYp3iTdY4QrjLYc+6o2iNunND535
p6Dc4jQgP9dDcwRbvfqUNFE13q8g+LM+s4IPOpjZMOAWwJ64Ad2sycPtRfTcS312NYnGYEMTLfo0
Fj9H5CZ+QyrmYskMwD14XnMRkL+d1SZYiprHFcdMIupUtfppTZaT0ZjB/IXHuOXKVRPqj9V/l161
LIab7uWwRgdt2rrW1GofILLfpUEnAYcsmbRYSn4A+5jzWoD6oq45T7rUhklWzi8ZSMwHlYp2aqnZ
2QpIZuDLYmlISp2fqQBM+Ev4yzzfZtcLls/C3aC+DCkdu8WbBSlSkvvGH7ln6OqNrn8C8Gb5heX4
kW+HHJTcMuM3XTqU8nH2TxrvqykWAdSsF+snB8/2UV2dUZIdwkKlNBkympCZi5hJlrNKQfDzzYdw
4UR00XD1SQQhDN4vPhPXhkfsPHsOjIJO4vDwlEb7QSaWOfRsHZZ5zgL57VZNSe5TAaFCXo5QO1MW
u/b1fK2LYePYty1dCeBo/nUIVRlDHnHYmf+1IO9Wt+QQb4UXKAtKRIepRnFr0bDTNs0uSOmPJ46Z
qtPl7zOJ+49Ok08GhjnxiwwSGuebnTFOoen9A9nk7ikSJpqihyScqVfUcLIcIedJNBJrs4FIsiiN
apI+X6UQ7AimW2hg+mKEhBOK2OGtqtk+9iFCRi1Od9PbRKrTQDeHCPB0EbmwF1fBxTtt1HuSTmb5
OqeMzw343LtOBPQHXgNzquqAJCabzZa7ifwKs4QUDpUWlFFjDsqDtQmnBt8kcBx2JkiPaj4GTnVF
KcsSBYHBFOlMJPtqxuLBvUWmA/fROeap7Xd1ByH4QaK5If9zIR6bSJfGkbNEb4mAmbo992xkizTG
8Yc7lmUh1vfefvl4Z1B71rwJP6tbGZ00t3jOHbsKGBDcn46i4bO3NVODgzUXTJvtZA7E36yRv6vL
BUfmKJgZ6LYwuVSkW+vui092yWHoIWePEhNpl8hAkp9zH0VHTogkbUpKfUEaHSEJv9haEE4oncZn
MuQURXH6amNLfKIdw5hTEkZwOTojxl9c2NuJ/Ho16t/wzTLq2+sWXQO3gUuyTp2ZtA8cLZeJjSlG
4VsknpMaHqiu/FkuA5D0ewGX8I7/LdK6GYJJkK+8du4lzFCsmBDbFEf5Eu9BIUZl2oASZD43oBrz
EdHNMa4hrkoq1mOnQvvyX/OL8JlB3R8MrWrZsG2eRv82ltzymylvuzwL636p5xh9zTzAK+toeyPj
xIAkYkkocxjjSj9YWcnD3JdGOHvMPmYrDpDX/sUu+fPOkh/XcmVRJpKQ4F0BpcZtnaJ2jrjhOkq6
p7ZXeW28Phj4nosMuy0W0NaC1piX2PVxOe0AT5jZETlhea3K8VXoEDFxeCDX1zIap5o2Q1BXL/va
xM+KUSVszFFdj/QfndV2XTWkn65lvO94hYzZDWJKbuMAnTYiAvWGYp4L/xKsDb7K1xJ4h691PCoF
j6DN2sw9D4ViT0ZVJIauZKpsojnwlIiDxzrDHvqvvvWS6VRYU1urlRxNOq+aS7vtQBXQrIwiMnzg
A8eJ4PbpBoRL+W+sSeeVqlZ3U2OtOBhNiU0htlNf8T8XJeZeifSB9m8o4ENOINbQhb1OO14b7F/i
1h8E58SWsLFVJQ2PLhZbYLQFKDFUnufj0+5quKJ4G7V90EJgBHPxIXGVMejQIuu33JQYQn+pcbTw
2uYzHLopScP6r9ju+0rFbpiCXmU9VXUXdbXPWmLOk0reB+kGmEZHRQDzcIF4sRQ99aagdtSSG1KD
js91nnf88bQYv0LKQh8ElJeshZ/eQ1tH6o3TK49zvBL304DCH2frF0zX6UdHKr3YYoVeqIcFC1dO
ECiveF3VqiuO2K1qb1Yvn/zROk2N+EQzk8Yn3sFcarjNUp9q39ZHe8L8F8poo/Bu4qk3jH4A6xAG
+tn/T8pbCxuWP2AybrjnKRO3sDoO5q2oPfAdEGunYcx+L0k8cGsLdl4n04FZiT7zOiGqpVALxEIs
YipHxdjndS0lod1vJXxcFSoReYtyaAYia8qr+RsQ16IOcHOOAUyey83rNOtGml3CnewL8oTM0FL1
vTae31eLzwF4H0p7+yNjK92jNoW6r4QIa/isjD2HsUzfDsdu5AjPDLTVglHUuL/eKLsVnIhlF4Q4
4Vc4xbMNhufX9JXlk5A4yw1RbkBREIgQYaX5QR7i3xxo6AvQX6wZ2CIN+0NGBJAy/ifvDO39ubld
zK6QSCPB7CrsmRTPH8vJ6d+GXbrH6GQROkcNH3vtFarYVixg/XpeD9qtAqsPL/YsBNO5Sr3O4FxH
UVPu3RP99lm+hw6Q0bHuM3Mo0kb8b8DmEM4gWwBOaZc4po2Z6CILBE1PDyFPUXZShvPxAvBkHPVv
z6gocFwtEJ/+PrLY+I9axKYkAUCTioiLd3V2rvyr+kJorMx9McFszYaTQBbqA22moeNeNyLcTh13
V5Fk4cJGTo+Z7Tvu/glzlxcMf9bfJRehgVrM3+AnHC/o5VGQF0uQ3FJ6CVfkFoURuKMBHsVLuIG5
LKN3PZkJWA7jSd0v03I/T1oaSQbe0x4Dw3MMUv2TycuJxMVd+yWlvVKIRrafanRvV0d99ln7v314
EVq8o7ArWAxsnudi8gH4ZswpmU5pkJsBT+ENYZxJx96oIz05zl9dmr+PgGgqpIqs1psXaWxhPneo
7VM8eV7p7rOVfogTnDb0vxGQ4XHiJcEVHK/jGqH4GGq5Sh0Wqrr891cdBzE597PZvsq6kCiaWcJI
DSNbeb0Or8FE5Fk7k+hVX4v5qs8eOsNnbiV9At7NVPZARZ757UTUVcLmHD8h2XphI9De7hYXkyOT
g/r4h2N5nBguDWdLFTeXkiy2qxyHQbPYokR/VPqUKnUo6oSefuD8MhEw9FOnFle/uuBqH+olvUR9
M3PYQTfLC+bcMd0KVP7UYv9jb+82W3jcJuKc61IrlwPlY4MQDGe6FeRivtZVjRaBreK4zB658jlY
pfElCwvIOt8u+ZX/PROH5QaRlSCZKc4Y5J9zjw/OW1Zu+h9+skTzNdJgYobpY4rqDdWxCThoQp3l
n5squEr+mM0NOLgn9M7zAu2P1BPplO08SGXOQWbCUXGEbLmKr4MbaOtMRWKQ30nI5jX1KizjJLs3
uZEByTsTdicCcc1BaPnBJ+hj542QtUaYf7q6/AOf9yRYYWVn0ddcvoaHGhBajAYNExG36xjBFTQr
bszVERK0Ug/aevxk5CIVSNwdbZGK1dYvLzNKsGqwhTQ75474r232TB42b9mbvVHVjEltZdzAUSVz
txX15IXdfz9U528rj5xllCHs0M/ho+GA+S6eZrYssjN36CvDZXnmGCLPXpDnhTmfWaGZygK/J5Ju
qnYhhjcBXNWj3bJY1uqCE9vnKc381jNIeJS1rtRCny2v4kXJpT9huglllXxkRBzBPk8kK3i4TyHw
gwbFSNHHSdu7fSTtw4eeDpbk89/2I/GXlQWNaO/YEc7hsMQ7LoRzSw0qdOjPhUpD+KiNHfNEHS5l
ovm9xktot/DfdAtyVpDh48I+mQ7ADmEbp8jpHTAlyVzn2TKqUy8cgW5mZVnM5JHwlDB311PwgOP/
yakt3JrBG7XFbyXWMZDA3T/LSrJ3UcKVgIkLipZ1E6p8URHJpKIXzDsUt3dRctjR1mmsTjg0Kvz4
jR/JAVUKGD5YYabE9DBTSWmKw4cXaLLvmFohJsZ7mmIPBkPIgHez2amDEYHuaO7z8a7kHSaXCjFe
wwubscR8MKgXbGpd9VAwygMx7qg7a1Vh+xHvfskC5n4rR6rz+PBRRTHhoI1857Akhr3jYfZmtEuF
w2v2e/SiYvxeqzJ8Y565t0qwvyU9AYhm1f3WZFOf47rZEevfD01/7pYeaDPpNzTFGxy+MVVQql94
GNL0Z2DfXa9QpD7OTVigu5+k9JHQd6LYdw04p67Wt/XeeU/ivbOqHLUGqLJsjLsgZlMPqrG0V73U
YwUHMVVJTkND+U2KEGoAQS/gBzS34FZonXd7Qdh6S94z3uKFOCDweHdh7gGsW/mdqKgiYq4Jx6Rr
mkelT8qsL9KZzjadiyHM5LL02xqjCvnFd12G+TLbPYgxDlkJI4u+iiOv+guvc8ymSHMfYTgkTmeU
1Oy5zVULK3ayLO2T+YDJExRZbmWtbml7/i3HwM1AzCrDN42e6iflKpXWqLq0S2s2x6UUdCQcxBmy
tSHJ5saEApYelegEgDOmmhAHbzHwiA5uzH0KHHCd/al4/pb7R2lW5B+kINpqubbNQ7X9asrv04Bc
qvu9q9kDU1elwlf1Yb3HLRoqyrzZbMBf/I6Iy/6uV2s1DofKmvcqkHZ5ooVlAxu8VNHPz+z2g99b
W7+hR7SeWmyu7Evo/hvzfMgxhJpp+MM/6vgT3OA6S6yUNGsBpa7q6G9COZLQ0FkdFW6k6H7Xw26c
G7m/Br0O6cEuIs2fbeIipypp0F39/mf6WpH1SJBjgaipAEBTxOVy9b5SPElOsw6KpcU36TXdp7tP
R4+Svy5HFKVMaWFjI//Vjb4MXiAKKBjB4QLCETzVdGgZrt81tToxOCpVmimca4QS6n3NRwpbQU92
KoNS3f80LgpD/3mQXysukmnDrI7GBvclvoXyYOnP5X/aqfj8VuKNPism2AZC2UwW6ZZo3rxLGdaO
Rr72tvGOOOqR5X+OVCEarniBd5lbkssDLFfOxk6PGcHbED8WVuiMGelnTZUp+O46r5/iDicBWJbs
bz4GcAIHyj5lO3B6dYnSZY2mS4qQHeQa7GnTonrvscLqGmf2xZGDC7sDE0zO81jFgQK4ND3i8Qsh
ZkQehcyngNYXnA5OXjAyI5qgcRhX2KgM05bD9s7Ts4+bgMjc5pYPNzI+qZ042GpfxvkRV6wn1tyc
IdMFzqdjhI06HNpRfj+CJQU+boQmZG6WQ/AsLxQWYLx8OUzl5FfYIbuHzGxz69uzv4kthA2EKO/m
PVXAFrtXADL+sjeLgUbLSFvnfdzGVHW+AQgDxmtYbfWC3ebiD5DZTqN4t76SzxvhB6lq4PhwxbrA
q1V2t7MIePYXYTqZ6aNuOVvXY4P2FqCxK63CI46svIA6We9a6jAB5GNiM1q0s2LSuuSyynxiBW3d
Ke+TFzsQveBUj6zNg4AJJi2Rv6R9K4bZfSMvSvELCCeosyHH13KPQJugjoo3VZaMgQKe8/QPz0bJ
bAPI2S1hzRX/tCauN040ru4Sn9+AmQC8gfqFCUZDrtrURYgFUU/a5d+1EK3oABYB3MOema8D81h7
OZo/8ZxwSEWXpoSbIGPcCoPxfZI0HNRi5QoBctKftqCkAxGaOlmwAXAYWZ78Wci/sNMmaKv7Q3Zj
PbDJBNKPeupVS7lOqaCPljmqlkr1qLuSyXlPDlMrX81+8+vE4tQN7B68k6WMvc+QLUpL1NYlwlY0
/OYmmD/rN1ypeA5rb/6W1sdIVXBWkJLFz3POcRPfQBjr0B1CVV/hpm/IboxwlWKeZv/Xz/U7nUn7
hXtNTA6K55SxnpVGnNdscTJMqL6Z8ZkyNcC+VKLv194rEmlrBAWFdmMZ8B0ppPoBIY0QO3vUFnFi
R4EHCi9/I6ywaDW98+FGLt7xb2Cf9lQQ9KCYHwYN/i3IQQyrqsFrAplG2AuwLY4fiekQMSzBIAmQ
J8gi45WRRJsslBFeuc2iwbfVhq5ph6Uc7eI2cwEcui+HJfV74i6VtO6o7Xm0dXWUl3uo6D1gE4eo
08WJpteSUbk2WgLCX/YZe2YXXKQIT58UPX/9ZRfq/Z2L/nDyJghTlyAETdw2GxoaStgWjCFIaDxi
zp3in5+j+LC2l6LoB1J7bmbejVhhqmrTld1199u3m1RwYJGWV6KzdWgIjgL+HZqL2D85BrYMzdaH
V6kJOjLWAfNVhGUuPnhOriVwW5lDk0Vo1wbYPmEiodWGmVriuiqF7yxOhToDqOT+uzdJvIjzgWaq
BY2xKbyQB+dLK/u9Uu878TBDuuxcHrSFsggo+n0zWFEPdy5dw+LMn3cxraPwmDU69KohEoT3FUcj
H9W2Nzq/NXw2yqa0b8ak84srMcpD7LLN9NQ401P+A8Ix/Mb8rIvJl1+aCfqc216VAfu/qPSINH4U
u+sWx8UaYb6L4zQ2FcnY7n/6LIXdZAb4Ifwgf13BveZ/9KF8mIm1yQsniTum8awedlFkgOXxonr+
msxcqLXdBrN7CoCP7z1nJ6PBCMdrPHjsWx2HJSpmsxL+mPe94HAEhx+5RNa2Irjhf7T3koE5fo9J
7Vw6L7fjkfkA/a8U/i/x+JGdnvE1gCuMZmUWRniXjIJRBi5hDmL2tVglaWGps3i4fDvntb98w4ZS
WJc7pEJvWk7uiHvWzszgWmWGHbEWUoZO+NukmRKXbaJ9b/DklcpfpSnQnWKr1cq1BWPg52grW2KS
5dSGK6mE/nHnfj1FNeVAR47apJY8pdrXdpxpAb6nokvM7/FFHC52XH/xkeyjNgyt4otBymPOS4SK
bgj59XspgH/GSFhms/4KS8C2i7072iteJZV1eW05ImurTH1TrQ+2KnsSik6ttA8COzj/oWp+96sk
hhWcB1IatWTX4wLK2D2+3/o3213W24/yOGFlxu4etecSdo7jUzROcSuh/LP5KRJfUe8VlE4Wd8MS
Ge2scQ2ne0LxwKGcWMoGLp9N7eNBAfV7gkt9h1r7YyVWFbvKzKK5Ru4mO0Q8XqsJzpRg8IfVgEnu
VYWMT3IWQLV6/EG2LIi/+QGswj3IndrExoodkPzusK1UvRoYJAn6xCGPjS8gznGBP2m09rhJKG+/
t0D6UlcCZX/VVRsAlDjmVQrCp19TIPGU46DV7++uGxYDK6mB3sN5BT5pM2IbvFNsYb4bi83JXlil
5lY+eBPs+leAzv8kzhJU70aFeh8oRnePBSjmyCfhKD9EqVl8l5ML5uISKunpvxq2tWJztxMcjCn1
ScOo8LAvj/haJ0ekHhxyyK71eDp8o+6xmIf1uBHZ3PKhyUMnEOb9E02IXyv5o5frUUmgEzAqa/i8
AJW+GZHZYDdHFEpR+T1hC+OSxPFSIomoK+dsZOLosDQLvYoq7OdbfCseSGIdzopa1oYiHJv4CohR
m6ajQ1n7wWSPe5De91D0wpM3so7JHRovfkdm2UvRmyovZU6PoiIcGh+nnZLXz15zex4lQMAqeN7U
rRgqx7OvM8xziFkZGITpgXIftvK+xZZqpQrPzOBSxuQY5RKmRgWdCBWxxFlq1tY3tj3WyL8WxvkZ
yH0uSbblxPqA990qlH9MreXFLp+w9tuxio+4PyFSMnuCQylEvdRy3VDqtQkoVqq/S/M570gFd3Ev
uU1VVUp2rDD43+UF8pn31PMEz4jWkcdJQ/35kwq/pqTjIwBSThQZK3IESxD5ZxImh5+orJa0RQcD
3I8bRo4XLOw9HH07smQJt+dC6E9mT4LbewOKwWL3ymNcQqE2c+0dMVESB8xeqQdFc7jY4QxYluCQ
iN3jG1g4zzgDaBswTJGu1Sj6s8A/DZ0H31S7M0VVKOekNy74ohSoR31cj3S/K5hUOm2LkrzJ4x6J
0vcUjZcM6F/yH4sDDIY5pNviEaCtr1RVpF4yA/uQrihCpB/gUpdjF+xZpMDPMjZvvID2gT1ExFrL
gTwcBXVHOhyLzk+Mfe9WovrD+0Huc+2qtBY3uQKuNNrLknlkDSl66Mxw5XurnGctRsXNLXR63cKA
+0BN2mmNeGNZ4FPZnb1DhAVy/xwuN9t6k2Y02xgilr4KYDL1TE1BNl1e/eoXWCFaDXG4M7dW9/zH
UcsoJtRUbJpGojK9yzl0UKDxTbiBWjuGxmvRKd2Kd7o16C57vdL6njLdvd8Q4TyvkHgPUu8ILft9
2sX5/QKrSYOM6cU4Eu8pctWPveiaQRR68HU/78M0LPLtGnN0/FFmFPxYUhu6/uvDymFofdTLB0tN
X4sYkgbHsUGBRonHpoMFZYmar3KuXSVaDMmvBnXDQviLK8mjds8rp+cRFsku6y1ZUrD9T0JtrfKb
FrFqbJnMC96KM3fi4qKcFK5pchN7qKImhgZlRaVF8zxaWAO/cZmejdRfvFXe8mtHls0Ri0sVDJ0B
7aJHGzoGUYtNZFIem1/z9zdASo9gANV4jCFs5GgsByjp5NT0kgaB9lc7mNNq8SfmEE0W01xGQn0H
xywip7QkktX2G8v+RQyjUWsVkSkHKls8QyZFisAVgOdDUPIK1HbOS0LGzjNd2miVag7whIAMddgm
63ZdkXrve46uuRs/LLsMjUMuv1aKbhz2voWkW56lzxUxfxi5Ey/FXYR57j6qbUJnrWethJEH2sPh
PloaYa+peJr2aZRV7HbgTgp9FzcAu7KafNAi7SIIg/NOmNSgCr7Dg4VMFV4/1A0lOqylNpBxoSBu
/SevogQkdl+PfcjbM66LDLz0BAXwirXaGLEA83Y9QmKikTE1W5I33LKQu7dWDOW3FhP44zUCUJD6
XJhSvJQdRq/NyP8Ew6vi2av2rG/iAs9j5cjHmXeIys+vl3Fwm1ztcV6sE55CBaSZ8gdXv0717pXy
Gkrjsqg6N0YGSozHQM3aFAvTN0nlt0GGtUmtM39gUHAOL0UhEZhnPus9dmTE1Uc92V3VJS9GtD+s
jyuM05xyM+ktPZaxRgV2gAoxTfnmwlkoi6QOuTD7nKqFB5BmmY0+vhspDR4b8dik3Xz/5Ym0APhS
oMP8dZxkFUow7BWiIqtwzzFwyAFiJlHF16H1EIK0aCeE1ouoXbBRUXKONLx6Ml/IvvDeruCeBp60
HoZaQphT4dGUV7DLr7AcD0TKjXjU6vhssuKkF5Dp7/YyfJVfsdPPpt3xThPwqk2rTFnEqaznFMmY
0uj8LhKBTSU61OveO8ZePLLIjydArP/gw4XMVcXU0JVGDGuaAkK0IU4RGAiTxxPELw2ssFvFhI8M
25toPdwehoD1P3NFjLGwdjwGMJHwsGxyvWPhor2rTnfCVLOlRon/hfSgS488pienHRqjHFmOp25B
6AQZOqfZelTxBt2crdtVmg3z7zuVKZUTN3xZOejeapBD0DeHXLMQKVv+6LEGfAqi/4VhdHB6r28s
dpstzRRNUGYK14OESIFkdmMrPPU9s6y8Odq92/UINS8Zjco7FsqJmlADrJT2K+8iOhqMUQFnFvhw
2wxvZSw3c+qU8uGm1MIk5S+cTdyYaz8Y9N/oPPmiVK6kCa5UGO56Mjd9tkuRin7BRNOjqPg8nNJH
t+mYCt4T1P+Yl8IhUiwka5U4BbZBDjHE8DUlgjbnuuMllkl7MCIVyEGRTfRNkbEHocwVEkYd0RQf
HsNrN33tYrC2eTr1q+AYIcX03uVPG5yaxryZWd0qad5SErSgF4Qps8EgQlKch6ajc6bJ9eo/woY5
HiqoPnolM9cudrPrlqawvjPsYmZ/y9AFrRrxktqZ7aAYnrUGFRfqnhKZelSUOlpQFGaddvt7C/Pc
s09ZMruB/gLXpsUeScSj9/oqte7sQEEBJPXgRZN1HRZOGw0Q2545/t4f59oSMZfFndN1DOaBylak
G99hiJdkxPrNGTGWDM00ofM0DMdDUhZpTp7/56C8CmMRBpB3YWgtw/R0ORi6xESgzVjIAQ3T7hR2
xNCDPTi2ZJb1TugN1iMeRGEFJHqyHgcMEFcfcLWHPSqJwL4+cMiCwD9xfxRzlzJSi01MvWB1GyTD
WERUUR5L5BfkjVP2DBlC9p5Rfutx//OJsPPx5eSCBLIf/vAB15LpXuzd38ujfFlgweFWs8zpqCr1
am2sYzaWDFzalGqiFnHOKTzmPu37d0jgRYuHGucMTLyemHpowU7RmFL+xhWbaZB951M6GZGRn+d0
ueFJYYL9Ay62EHf9bXcND/Zx/IuzMNWlx+Atlja7oSibh+NTnXsg53dgZ+2tiD46RbG9cIovnVOF
au/DIFVnqB2oKLLXQvK8TxD7tvuA0aJy5Hf5UBXqk2ddeG9YSsxBBDl+lTnhb/NpofUiI4dl8/oA
YMUuTLTx7aI5eE58WftqhXXgy5+6rgtQIjyQVQrjHrhRcIg/IdvFRghiUSlmUp1BlVjTOvUd5DYD
+BbbQNqFZhYRTGn1v//B1C3NkSHh+ffvEjfzfzLc4gYH5HLAxW8ioRVgBP4Gcfa6HR3qIko4RV2j
tD8L4/1TcZI+7wu0aXGmmNOmKE5P28oU5h/+X10fhp3IDnt5MQBHOtTBlj95J/IssOztEvsXH8VB
ZyYdWwUlLw4x+8szMOfMp8TScGI2+pqIzdKMepugRU8F0pd/P/yQmPiGAUP6Dxg2Fq7rJUvu9302
e4yabWv+upl5rGNjT3l0KT7SEqB0SBeAz0I+0K4St/1yJoFrE0RdjLplsYd32Sp4vkhA4REatGbw
e2uDDydBTg1KOUh5UP8kmPJIdm+fVJPSW22bGimFK7rx5eSVDeRUmAIykbcDZWTd2C23yqGhvp5f
zDUCUXlhFdwXg2f25BEzEz405hHXF7Cv0+iYLGNE7EzR6fTpqgKKzcR9xnsgkv5QKTJHv/zJlnES
N+yDoN7XMINXaJIep5jrogGcRek32bwwRbwl/W25sQF4fVWowRdhjpaMCxqu+rYTiUrshNvV4pVL
N82r0LOiLFvl6apsJPSm+Nkq4fCEYlWHAxkA7Mb3OyUl2o2irR1WF4O95zcaVld51HvAN0+x97wr
0HcH3eEPHF6+RkhPiIXTvm8WGA5SNepNZincOEjZKn3s5dpCZHotU4C4KWH5okZOZ7jv8qgD0z/l
K0Yfsn65nJg5ytLJEAWuNtGnGn3L7vN8VKhxNK6B54ADG0COhBWK/fnaDSwz5LpcHhrPPvQ3jq/X
T2HGSGcw4Je3KTySTG+j36QN7J7fG9N/zsPkj95c0Wo3cZTKTwmiImAe6zDzmFUbmxKFlMRRmXnM
gHIIBUOTsjk3+h07sAOegwElsUkLxFDGpPstBTt+0JPWr9ebJlqwnPu/tGmAmpxARTL3eJX7nCsQ
EGJ/nj6h+jj2W4emC/C5sQ+VJn9foE7qGQ/7yPJ+b1o047aCTyDfiHI/WOYb14hMBufSfakYEHOw
1waPqFvmTZIO/HViozyPRdO33D0OLr7sKl8azjOVXysnVk3oS1QTmU+9J2PpMTkgnt1id4CpfmJb
+xUjLZTI7kiUU/+POS5tEHl8g8Na6p4wDDByK8qhlsb2h/tmnfZxhtdIs5lv0UGJDhMpMXYJou9M
Kzp0vGRNyLY1ag8CNOt20OLOAX7397l2AxYtxflCp+pQf/zQ/7pmnF33N1jhAOn1vKA+8Jfuq1mS
aO8Axav4OmLwpSemDyhzCC8H80Jmj5f4DQ2c9Zu5JLbNdJRJIYsxVK0oDpNC9Nug7dE1BASQOiao
YNp1qbmA2HfFoOOd/OGlg5WhFXwix5oFyRVtxyXlqJHZj7lAJXHMQnKRQ9Uej4SKF62SGyv7JMGC
kBWoAujirYmaH71F+GkLol2GIUkkXyGRce7xlrXs0qYcF9maG+Mdde+mvTTC5OO6qBeApK7yG5gv
YFojX4inC8Q5LU0fLGweYhyocuqiEoRyib2Ugi2q6FJrxJDg4LBmcPtI7VCF/iR58MGrIJ7SYsef
MDLKBl1hmTK32AT0V5B7V05xUfyPWX20Xqp+xfPBC3IPZMksPngmqJReGObbN9koEDumR/pGqDhB
V55vggQwZgzWiuBbDQzUDH6BaAUec1YQwfbnw0u2XXRopD7PanW4Gq/cqK955uNEOxcW1CP5z2Zi
nNEVLdIMNm+m6MocQvlMIeRGLL+xPAGYgEYRtl2P0DLoLyTCdEDeO2buBsDAE+f9BWUbQiybT9Cl
2Jiw/90nqtZgaawo0jVK/IrtOvNOt6g5VEUAVPqj4nxR916TZ1PlgzRijX/hi2B9qQ3ECNiiDnIl
ug4bJP6deLymLrD971T+fY3bxPABsp7Q8PNZL207mIyqd+CFajsM27QEdrhCx5YwnpTFZViKxjic
Rpt9mPKA7AmPTA+Kx2aGCyuuN15NSt2/vVWrNBjSdM90vP5zducS1iS2DNvl8YlaaOVGk2P59fzL
dZ47OEEeaBGg5dN/FPjPlqsH/7m61cI+cGCb3RqbGQC22XndjeyNk9+SKwVhiPwhNDDUNeQP9+EJ
v2isxkhD5ZVGxCGMa0PvVGm7tgY06p17+AKAQsLokg9ajstWnJceM5dtS+wQEvB6qYnuGGRksfiH
iSXkakhr3jnU8LZjd01l2839M8J1xqr9CVsgD6O6lcFQgdpX51AeuC9qPL8iNumsS140Ud8LDbtv
Myuxk3mfH1GT2vQj75y9rwo0s+3t2QygEuPAgx/71eMG4olpxwbqLtDKv3CFio8oSV/4hZnHBXS8
OT6EUB0LLz2qpjJNVRGNMiIyK7X78uDheGKrseRYxgUWCUGmE6/IiTNl46XzWXWber8W+0IXDLgJ
K8uro5amt+O8pfJOCjYe/jGI+60ybDxtwXGAAZS+f2tTPsEwxfqDNYPRQdDJlq5LKOP7/vF7/GtW
IHwyzqiltOtrR01zgTqnqNBhm7yvhnyTyu6CVXOMkJ7NMeAANOANuUfKZdei82n2t5JCyyRK3Cak
r0vh6P+qv7v6joV7IWftsXRI8nTbmu7u/dCdYkhF4b849E1Mg/Dxahz4dFgZm/dLci3dkC+Wvoux
b/pGjIMSLo8xLkvb7HhGP7tlB4Svj+VvhqbhW4b0K3P/QFhtsL15Y/QKfulkJRZbCwimn3WjGu5l
jQ3YjuZ9jpFZiDjAfmNkxGy5xSsJCNf2DcHME622uAIDpeYWj8rWAUJWV1L89NvUCOtRQF+VwrLm
rDAS6mhGCgUDftPBWWfX+4y+RrO+Ofx1Qx5gedUiVYx6B7lBQHfT6cDyc36fU741tewNLyLkl7uo
cf0hmP/BPMu06JEJtrnfF+VxkY5qsTnGviG+M/taNfPgIWCCyWD0HD1qeA6QIqOz9ybW7HLPfYOT
oZKYHZX92xS3ZzMTzjyevnjkK8TmI76SCIKpApBCHtOnSh59cvgrjr9zU6VB8JwPYOVrLM+riDn3
8DQ/gisnEFE9KfzKCXoPUsBXu583Mv3jfWr7vXmMt8HzDdwgwTLIHraag/EYOf82Hy0BwClFsXg8
RhOH8GeVA7qumj5JKqQd9jVJxlRZfVSt56L6cGn4p9HPCL2TJpbZErtneT0AnEwQvKiQnmszNdQw
YWiyq21HVcktfGdxyFqmFftWe9oh29O+fXO7+zWQpe9oV4Pp1/ZbAdBc1CtHpg1lpa5K47WQgdUe
ArTC2xMXA6KQcjynwA2yRjqniOjpNUsEsDSp6jJ804leyvpAoEx+ZOcaxusnMyNpiIuyKw2YUuek
spv9GO5Le6wQ/XfB3HV4GIKHM+crOCgfSsnuYJi/QS4yA7iZS8S5B/qK8HGmPF4dhhaowc2DfsqV
WjKqd9xT2VjQcuNlEp9AzFvp6zj0f8XsSSqFIHVGRIASxZKhnYPD7nlUOhyh/xYOTwc16z2m7JW7
IQk6AeZRwdMp8CnTBF9V9rvKqQD6Px7eBki8MA31DXJomB/IvZexZ+xe9pCIbtvoIn9x7y6vhrxK
8bEM35+aQnjJMNXD/LOljBtfSz9fDnslRiLXiAJpST3PoYx4HuxYMxPKg2QhKvKaaTZuwf1xTwZA
c43mzOhHJ4BmlEgyzBPKJfG0DwwfFI+1iWkjrWWHFBFIllCRfn//FQrwVeXtwu5Mzo9SgA4LhsqP
qRty2TYAm9rxbtVmCdZg+gKZm4XGCKbaFksQoYFkHDAtmuZjisbTDAKwBFWyz8cODK1fhAeHw669
CTDGKrKKg91BnzJa3D8oxOwQ5DFgltNmFWo6N1Kx6+x+LYmtGe5iKeaL4IYCy2B5RkM/dEcgG0Rf
tuizFNRUXY7VAQQUC/LO0i3SuZNw2EDe7DVUlcGsy0OTuAiq8JyjVQ1DR/edPkEev+9xStbvYDLI
LsaB1e5PzLQQiKUfVifKofsSO2zKf4Z8LuU3cBsx9HIRMPBaCNwiApw64XFFp6H3EwP87nFaSU/i
ZJmw8wZ/oP0VCgXcHNC5GI4vyj//TPY3nDTWxzf3G4pwMhev75s6hGI5prJjQ3w8iyR+GoRnNWKl
oURUsQJllPTjOnowNCm4l+R6D8tiA6io9dQO9F220nbTC88xL9+oVGC+Yd8F3F5ejS4BwYGnYd8q
kemo9+4N3Rt6fNDDPUQ1yFWt2ENuE7i03OGG9A6hLP+FEOWzglSosCosdz+Apr+na572nboa115W
vTpUmSCn3dG4LKd+1ZszHG6SfMWQ0dXsceJhluIzAEwMHjoa5vxHLel2T4iGIwAA2CeYcAT0fl/0
GpiA7ZSIod6U9ZfJsTDhQDc4Mp1+jchmFMj3HNQ4XacvqB3NwlGfWlolrlp4xKyQ7manj3SQ4zJA
uJSmZjotak6eHEIqmMjrNRqd0xXowgVJfC+oRNU7631d+Kka1j99lUj6WkBRECtbsYx9o5FGMGRE
8iAvYM6t3PKtw0y8QMlEFrHAjYGDA/KOSUso57I21z1Nfiq7ekVfBda3nX8eANMRY5R1ujA6yWhE
RsXhJn4hxfgYCGlfxkSpM30Df3ha4pnaMjdz0oWT+TooTyNzXFlVZwUh1fYdko/XaaJ0z9aqNRit
rFTRFfjFroFthvf5iU+zPirckU/pc7AmoaZCBE3isPZecw2H4vTZjs6ASRgpKcOnSsnydmlLt0S4
dF2KvJfK8iQejqeL+56A24Xta0yYXEqUp+5Ces+pXkdURrfV7U72wsM1fvWqq/42ft0elSIGtvAQ
PcvP2HlpwzaOqm2ivLy+Kue7LQUSus325whAfqIEQUtqEF/h1UfClRegpkmN74dzbtEzeosAyJpG
wsbMBdgxa8kDzaT6QARuqVruWPvc0lnm3UCuGXvc2R9bRXYPenO2qc1DAjcqkXs9OGPraDis+ppb
bag+/B1uflRP9peVxii+5IJ5+eUSj5qWtowhoC1OHJO8wBeh0maTxzWxSdQhm2QHg8cLELNRokLn
tfjYiAGyK0N3+T+Kc1xDuvIOmrnVoHchcIS+BCpVOJ2XMSpGW6kvcsIMw00CG2H0bIL/wB/ml28B
yhAvaM+twjnl/BzFMz+/y+DYgx6qNLhi9z0tDLFrGhOr2fD8y2cPrJYUcPwIEEXlopH/ciCWbqc6
zpPt+lnbYOEAmIKEgcH+htJ14i0EFQrvMa3NZN76Qn/qN1u2VA7djP8D7a/JIjDMPTlaL66JKiUI
SrJ/jrBo6Vm0u/0MWgmc5JmvO5Me1vOVV+0XM9sGNQK+vhhX563db9N90b3nQgoqnp4U33YuGGn3
S5NYfb5hH5DGO3GHE8UtgxjxmA1QDn2ck3yMMRqJlQzQX+bfDEXppvC3tA8BOn3kCUGUneCqFC7k
JvHFlD7kJ69+4mlJgbRSJRjtBy/0GyTuu2bRQQWEk0BFhNUevtK6B++EV3qXYz/QvJfYV/6gqfQg
tRmqpoTdQ2NmtCIT9cSpFg04jO0sJnTIgTXpdzRqyYcUma9w6AxKPoMJy5iQ/bWZGTouEd/Az5Jl
u31fws3CkXJu05r1gz1ZdBIthzsGzYNjeHniUZyzPw5o2SGgj3tLypkQqsnD8a6bzBeU1CEpScbT
ziNCS2imBc725ZHvGbGiRwhsHKcOAONok85auc0W2n7XNOsL3hI2qYh7xOzSs6Z48ammpnhoewbO
0didnbDzM8p+jShdmDTu9Gub4VhqPwbWbXYFqSnsKuUyUf19NJgdB1UDkZ9S38Tj0DVSEG6854U/
ZY7Yf8QANmKUKeMktx/wbSvpN1Giuzaq7n8fJws0vUGMV+pV2mYYkK1L2Ni5YK5LBoFepGcuIpZ7
PeFXaakW39uXxKvEWvyR5ZZSCUcVNdH6zyTiVG/SYjF0xrLeWAHKLMIF8x4bvoHPsGmZttLRt3OO
OGMSlA3VgcwcY16UzkMdkigQdI8jHRaC3TlOhcPDzLaKCyJv1ddI9BbLAkLt9shKnwh3324RpgZm
23apmnuhE2xfyqa89ENpuiG/76Mj01XmsKAMvuZyo7Hb/irhppamBb/XM4plAP2LItDBapi++Md3
Qt+Wjdpj6JwxRB6UF2BNkLuBMuANEGbpPSPfslyWgIsbiH5e2n3wRrbuegY2lWSsqRBY7nTaSyzm
LE6+JOoNCf1OvGb7pCC3JZNVprE3GPIDroXc5/e9YqVoz87H+3lBxf8WvHD6O4657ctlqdLqVhsL
cp3mFdAuXLjKNclDzMcWefdiKh/BHt2Q6Vft5HNm0ZaY9SGmW0JWrADLELb2UFoRressYYKOzgza
JjMmWATfM8K9eXL1+k5whWQToaJemoRGwmLR4MVo2wzDMP5BwFnuffPgmQh/VyNCK93x0BFXlamL
+IK+4fAlZR8dSI1w7LHErFFWzOcWw4hQdeDMYecOAKfXVksjJDWIR7CToqbXIvpeaOTG9Or5SJb4
05/kiA6hdgHftw57XgN/HLWNfHpvH7NSNL9oFMH1XFoGterimOZ6pKuiTis8VYuoHd0eezNtn5H+
0uBO5SrJ2igU7FxG0cMtlhikj0D3wOUMAXkD6/Og7l8ugOQH9j51Gkn0kxj0TvL2ES9xPxU6u0Fw
3eWh+ODUZFWOL6L/mMM180Pk7u51XqqaKh5vPRBDZfZ1OyVRht4TdS4nBBdb2SkfbYYOtlkirgWR
oa/SB58e8JwArOXsgliaV0/27PazyY82bTAehrt535ZmLURViW6LfgLAByZ/zSo265eJvnGR/xns
w/tu6/de9QfFjvq6txtCzsqqFamgrj5V3Aa4q4BYAfwXMbAuUen1G1A2wKsL5yNrBq4D9/RhoWBu
zrbRabz7PN/qcYIoDO28MlC252yyIKvOl1xmvdAzqWpxFKdC8bcHorTKgJAve00HyRXP7OuKV662
eCGijVXpGg7GF7RXusTaXX8SuOza6yfawtPaAZh884S6Z2x/RfKLEkkv85kEqyz5t7cAlTaJmsKo
x12JsAuSXjiG2Ln7bb7DzKVJ3dTk75dF+RMAfTreLM1CqEI5krElzKWeTQziV7pIK2zdCOInuRjd
5X/9JYEGw+3zY1WcNJD3m+XwVsby67MJeXPD3dk1pNwxfA2DDZ1/d3htgbkpWF2e8F8gZLT0K4nr
OhyyjAoCldO1wq5eea/EZdr1Ep8grjGUm2R8Ul/J/C8jaTQEwpKCiWVbzRubeoWVGR6fEtgbjFQd
eXHQSoehtOhTE36OJnC2jeznKPEq33lXfWgHNItBHHIBSsvKrqw0K6ih/3kwQWQmngnhe3gxOPpH
2d9kb/e7zyWYbL9iKmKxLq9IcEAdmQIPePhQjBApswYRJHtRV/1MU5o9492tNOifbHST3snesVHa
kpvmt6oJv3Q7WdQlw63ZI+zi0xDJf/qL3Z5fItcTeYs3iRP6AB4lcUMxouQQizfNDrNWfPchbeHl
F9nNRiFUTvQUjy2UKu94jJ8IpBTGxgSlkSd1b667kVnoz55JHYt0XoUu9nKnOZ8FNX/inxvuuZVU
/vmU60cYygMRqtyUYxXO/bxadYNS/0IQGDjdgDO6A4WvRQNAwahvjS3qIiV2zsAsxdEuOd5MwajI
U+fBYo/KRkmVB0jUFy3uoeeChoHJ6Nyly559nYE1vhn1My3n/S6YFa8hxnAQMamTGJMIL2xfj41l
NFeOoKDXBpq7vKVnB3oEO3doef4LskpAn8Cx7mTb7py29xjHQMsA349ok4Hw7TyupccE6ZqBhmXD
5GOMqz/yzZ2IIsoajOiadlYXD4nrOxETU6M5VzZkFgUPImBh98GKdlRKK/TnyYXzx7uZ2fl6t2jc
5M7gq0S8tH34Z/nRec4KIxFojhUVRm9TLk0vIiMFqpxTrUi4BIX8Id6XETM5k0ImLYN103gmZiKe
pplrTYfJwu8QoV2Nzfh7Xs19fVDzlrnOXJd8cupxy6/l4MYZqZMiJ7mmaeKLs+JXa3l0b4AM1rW0
p7RdTgI1smNdcqrGV+9+stACnhpWyYON/bzadeBnnADyBUufXjkyBqXqOwHzYQ+F0SlWUhw+DrRc
VzMaU5oVGWYbAiiOwDfujg0/bXYhRHpoilK0whm1AhRG8W4uYDAy/vhv2TvF/QCX70BMtAoc7RgF
Qz1eX7fO5FR467zrLRdSZT4qGsIRnK5iJBVWIeFYiu/7A+oQelsSGmYBN/Mc4/xY9R3Rz1ZpCrQQ
0R2lUfWNlR03C8X+kLZ78hSHHtskgmz366JyZ/khRfluskK+eqy08+Os1xSv+XLUu2n1pGo/bOAc
S6wg9BJljA/VGJPNRPHbYcAgjQxQ9gkpQ3xPOnWz5BvUVxJrLi132ETfj/rxbPAkcKaT0yyPDjuz
Zbri+uoUpwwrycxtnv36tL+Q/OywM5KsZowPMZdWSyzMYTlpusTJ1WE+fVm0c5ZHzM9JkOF22B3T
Ve/ztyoObugraVvktR2mMIAizGD06P2oPu64rF25/YMWnHnYJA/Yr/Zlt75Lnu/OJlkNA2naawFp
2Mot+tUBOl5/DUJM8jNXrsCeS5dwy5Vpv8kgYGO2HEp6ks8MkKiqZ2DmR2mII7rIbYT37LuRtvbL
1pgfIC6SW+vSmTveelsg5qJuqjASlgwDpTmwwQXV4mwirZhwnG7gJBZubVx3RB36+mxHhNOKiCOk
74KZiVCAIW525WBIvaCtHFd+5jgg9bcuJDHknqDxHRFH4jqK/0UGvXsOccVnTxlVKsvhB8v1wcYW
rSqV6JuQPd+Zlb1VX5rGRSlRbLVkRh3Xh5nqu5GoB3DjuS9dqRrO7Pc6Q1akdTU0xOCvcLvgEHyz
uNQBbMKRmXn84IAZJmox4143Wk/r3i/WYU377P68l1M83HEE0U6S+btPubpDnBwA8BPIWGwA4OOP
IGjKFRKiyCIaJC1wqUFVtqp/Q0RgwHtdM5Jrw4xMjeGPwng+kor7LQ/9wb5imzT/k+ixdj6hEpKc
y+A8+o6Wlz5mgXUwTdMDY3LMfVaAJiS337P2OkSLI0JMdPNX5rl8DBvyV8ISlVhsRSeB/HbUao+A
r2sEXkXqRy45qNfSOC/o+RUn7ZfNvjpVmP40Ww/M9+OxO0DWiShstMSTFo7rvktNkqXfQ8GhhDex
NWWUgyi9XmOQdgeQhFnSqvr6dGPXlo6MfjLutxJ/TCwbUKI+iX2Gqe0ShPUS40Xi7cQ3IvD8oloS
P22DT9GtARj7jfRZ5ASMDQjFgf4hMZw7AUAC/+vqkNBlQ/1z0OfHliGDxMsIIy+fl5wI8wzWGiPO
m9rjiAL+tNOQLrX+N//7P67eLMnvjxuPIhbhWlLJDt/AoY5/Ftpbw2DCMsuumbAnKfInVoqYe3z4
Bb90IiquEcSQlATa1JBUL6gBbSmRiPPFKcNuhweCG7Ny5NwhIjd6jbSw4ZOkvFnhD9swKbTS37W5
likDUYiqtVXFaO/UcR6Duwf63U1J5pH1B200HpYrhPFVtEY7RcgRoLX5gez36uh6wQk+6dKLaR3o
4DVKyPmBxVVps22JmHTV/empcWcRRoIwKEoWb3HVsScHTrBBiu5kDAQyDfzPBDcwdXm1IEfctsGq
QzRuQu8YNHs2oCoWFi0ghaxz+DBsetoOJV4l/ZovqdIaHGIBhDaB9rUeWbhMFLICR9DT0+gDPyvs
oUqnUDbY9CZZ+xE/AQaPhoNe/LLAbzIc9HEniTTGjiJPYgolwbPPowvFbPsyRtwkD9oD1jXMsNKv
TixqWc81jIqPZs9RIXrsH2uDjQuXEWJpsiOlsbRsaiZK9uFKIGunVvq7ufPMwdUfmTAGckr5ZVQQ
ojaRdAfwe2BwDAOIsyeobuAZOeUEdTt5uxrFPXDhSe0Ffc0oQXJsWjDbN15JeugaUaucrGieuRoM
2sLquXnT6/tUR9Wvop/gW0MUOrYxXlXyQwKbb0R/NlmMXDB3bA7URDMGuOEiHqMlsERmuCa22BsN
UEnz1f4QQkpsDET/5qeCDZ42/bI5PNlDDCs1vbqd6Y8o7wYdXuCcj+L9nmxihyrCvWzKJTd2ZzZv
nmElrktqGUrKVNYXeVCOOUNU0RoIwH+ODlnzC+4hJJxJhTVtF3Rc8VCGSX7+zfp5GKbLTBiACLgG
1mPLkNFE5kSky6M3+nqp0R5go6cIvWAuPms+gJdXeeSlQ7/msMF4tLatvcnC8J93wCQIrNNoBJ4a
LnFDg38YlgCIrGmje/WQr5AWZzFaTQfUBENGzQu0/iTlU6c2LzU/Vr3szC7IyJd5nRZz1IXcX+aX
8Mvfey5fsN60d82voU8za/EEopGRYyq8HcVHiPitZtohEr4cWKuWdsCw+6ZnK+G+j0I9xd/KdTN3
crvX/w7eV9Bx5sr7u04qM4BqzB2bs5sBBZTGB3tzUg6WGpZTd3sBAjVMvmNYK2U3KVKutIRfi/mu
RvPkAc/ZRl3RNAXEFep6wnGQtwPRXp8b35YoVdqoeCvnAfEP5AYwqimLuFBu7EGzE7bSwo0AHWOW
QhJ5F1ApV+Vpf35j1GqcpDYIDxT95atWI5JlV0l0rakdCDs8dFbYmzNOmPOY5BbnrW53sfoIiTLS
mgiQiwzATm0z7phB+q+6ZmA/L99OtBX4ZOeR7KhM7uM23zl0aZSDp/gw41DP3lWc8ImdqsQuuBcr
LcZ6yFF/WTHrNE9QwxojpFgqmY5MluvFZ83oEffO7vbTI4q28NXZ3E3gorbXAhJPPafofkk5bBR+
BsEAsB6P0TfFdVTCVM1Uq2jBl575pjsAfmpXcS6HlKptLUI+xsanx/DxFkXvdWVxuUUkxEXXvHrz
IJfXE3EcpWHQRatGbbi8KhJ99E9iZssPFKE7AlcWYeItB2EZ5nMtkN6FsugYrOpP0e3YbuM/JNTz
UCnUz3hW4AeCl6yI07vzwscr/hcvXrfIa8M0/AlVbgOUXho7itFLmPS+Hog9egOT6ry56D6/U7D4
mQpwYf+L/MqrkHBEycnxMf6tuy7KmqGylprwzDsPMrJlp3gQ8q5JkyWui6XwoBTLoUCW/NpXiKW1
jpYrcKwwATBRZObMSXap9uVih92Wd2BJLLEqkFascaoCGOagzcjjTWR2G0txBHO9erkKuzyYN7D8
kTA6YI2SpC+M/d3urPUEBbnaBBJQY8OUCJQmgPlFvae8k0C/mks+tgpkrGCEm3hmTdbYb3dnIRtb
d0QRf6Xyb3ZSAIG+3gjFDQeMlE+xdpX4uFcSzYZOg3gkF4NLx0DZ0PBGCJxnzNFy4M9R7eN1Ste6
Z/H1E95sgyvpPOgVkMa1oW4p2CPxQPG8ORnxXt2Wo/TdRssflOgLYHu/5ptVgu9480Q7bNJ4HDE3
FeawJihyA4F2f/pKOcxol7AZarTVe0QGgizCoOxd1l8SSGmAK2Xxn7K4Vla/lc5kZAiIAKwUSFhO
yM6KmuY+ngJ62SeX1rpLCGIFU7PxYB2tsReo3Dbcghfyg8mJbivlfWcTYvP6jmpJYyUjPl+WZ44r
+wK3kmVSAEBgmMT/LApU54pAWcJL1u6/eOvq6Fqy/KFuPuE1FfTtUbdhY8shQS/1uMibn47un2LN
+hLClDuPPJp5yX7Xj33KiBUwBu9tovNozIKvZ+qJm9WjCJxK9a2FFIPGdIZoNEiy5lrGyo3RmN8Z
k/BOT5LSbxNEme3mIPlZKuy0Ix5qbKvlfxyQb58E3cLS34tE530WS0C7ApxN00ffv90uNp5Lgcpb
CBlPM9mmKA+2weCIYOZGcshu5pBL//gVml2snzWP6RQzwXfW9u3FR1vSRjzcYDPRjrXk+aJV+QLO
V70TRkDsyatqGqGz54GCCLvO2MjQ4vFtcH5zpy5E1xjh5ZVVf6MTca4QAqB0CbXc81tUlJufI0lO
qgSwrx9CjVMjhQr4DmnOjp1wzSmqYpL8lqmU2QdMFWNvdaDktNcOyKeFw9KCw+wZXxds3VwQMoYa
DNRed65iKS9OZdTG+plrtpFFUyXH4HrTVgxpvv24nKfXUaEyIx01KVajmJi1H6X0xkSB+Hamjt09
qWGtdcVmWVs2dwo8+39YyyJUxAHCgPFXqR+iZuDnswBmTCptX20Ok23fooO68nGNyuK2nAYCWHgu
v8U0RfvjBY+gfPi1zUciQ71De603Az4YEfWwNO3pelRRw3+P6bfSoFlZ3vg1So9m7kXiPTGQyFg1
HVgLEPqdLMrUA5uBoJXmR7aRhovyb91TIrlQ9Ocn7bEu4yytjwrCxo4hO23hAvqzk1OP8UIU5AiN
zQ5wCHLBACUIs97hTWeJ5vhaIRyZfryGK1jTaKO88tyeiAuICK0BBOhJ3KougoWXk87iIVzWnW6r
OhRt5U8Fs6g3HOudJJTf+s+y/jaUXs9St3CMhl95gFT/NF390oFtjm3k80KGvHxsla+/i7eRG9Ux
yZeDONELdxXBBH96EJ6R+VikaVA37pHU3tGMIPeq0cb7/WZTT9H1Dc6WAjmibv1HVNEXLBdZz6t8
ZZzY3rHotBQOglajmoQ6xILTRASjMZe0mv1tqGKLl3innhe+mp3+pngmIGVwAwrMFslBODuCNroq
nQjxEXUJyxOKTAnf82EsP+NkX5K9yaoMiAUFpph8s+xwbcX8W216XMPMYjidMR2R4z+xK2g90sa6
rA1WajUr7ew/HLG9wo+vVq+opzPbCYUO+/6q6criWq0v0L8fb+Q22xnKnv/6tqwkD+5QRUomvodF
2Lp6xsNbGXidY/7uSO6kIPYkk8eUvHRfSnpc0pQKTvPX6GjfFQXcaNumJKNvRXKmu/03Vwg7P+jG
WAx5zPk+bqNtrHIrIKCYhWkJpy4XVAui+p/mC6MzQPnSu4a8JyKt+jjQgs0v72yg7ax/+NJwT2/H
FcIvtkDR+nCkYXK7ED+H9szgVsZaIAb0mj8Wx/kHNrDiqOJ3unCLrNgj/Bkqop8AyFYjd704fUef
z2f6TNBWePBSXoDeLrz5y1yWsQRfRp+MZ1WwY5gXSgPmQmn+5jwFmDqPrqrBtj6q60zq722HYI6N
97hVzSOS5rvUXdP2ZZOP3iW2O2B9+UuOT/Y8IxuQlZDzRRmWj6sqhKvWXDPWAoCPs6YAIJwkMgSn
B0VvFeonawH0+wYbYfU1kD0acDFWaVI6ohpcZKFjZTckee7KHajJFyGqY2uddC9bXgYLW8vHH29+
alekIoDN2M3hRH9/xiMZDO0u/5+rnYsYHXKtQEjZeJWmMhozOiKEkmy2BsLtE9wVTSJLSsbXMb40
ku5Rg32wsiceNPn2+PvR7PrBJlMCZIhcXorYFJH/fcpZ8go+ypVC+1IWxhfYSoIlwMfIsNd8oxZv
RTSH4TOLz36iK9+XUqzN5yDtDjsMlyUq1HB2PcLcRT1vhM/XilO+WcEIZ8fvSSXrqe06hSiMUl2Z
UNCRV0LAUZOSZTxZr4nfWL18fA91wgLo7SApbEmqr3/MYr32w2cq/pJACUL0m7cOyZS9XzBMZ88y
VIUKOC5JPldg2hxjkMmRapAZc2YhkPshxPe/Iu6HJ/eGzafG40Qc+oTwT9APiPAkqI9ly3E/CqVi
E5nm7+o3BCZOrg8TqqTpzYz+bO6qqeVJXTK6UTGcNbbVhajQzic77j0lsI0niBxP75RQvuzPc7kE
DiR5+5kzBVQjT2XGN9O32RAyjoEKIecglvN7DBx09fz3LXI1MbEkZwUU+aaKKHF2Zksfbnpx8nqA
+K8nu6khkKENTi4JZ9BrySGFzB7lKwmA3RXPKjfUTZU+PVOGu2ebXjhoSkRmRfsayevYje7u4jQ3
0U62wBrWtsR06iSOCy8Nm+q750BsfQiFYvlsrl8Rv0HEK7CG8ssE4heRaEh/Baz60bZFSw0wbAoG
J8XQb9GBOL1RuDof7UYv4Opg0ERKZrSjDa/5LQZ3XxCKjyfDNmy7U6WxLXo6BgDwahdZLkGPW38n
VsHR5Rq6ScVQegH05yhObByoYkIFeeV91YKsM170i9S2RxEQUtMb0LzPHfqLHUr1bWvAGeQO/YuS
f4NwZU4tfPMeJnSfCu1Bvfjj0ib3m/hMD7cg30M8qPXdX8XqZruEwOegnQsMF6nn7oZxIT+jH25D
ne+C7rvTsuTmLU/NZOgG+t/+EmY3Wce1sJDF+pCJs/+6lECkg7aMV5TikaSOKIRCO7UuINtTKyjG
hJgFX41Xw2ati1NHiewUjaR09JJ+flTKQ8hSb48zhi4X7HlpNAQ28iHt+aRwx8Gjd+ogx0l15ute
Dv6hEewNfYSUamZUSaKB6sEQE4pBAdNQkunAnI3ZXW7l6n+aCyIBsFePvntb3DsD7cQkYRXWLBBQ
OCMSSS0AnOfY5Xs5EqEI+OP64krZLjUniAfg9YpuCBCRn7Mze59QPk5yHwx6fF4c0HigB5b6lX8e
Pl4BGinaOJhs63bI5Mlnpw10UnKaN0CkMRij6NvR3+qojeuUr+t9O/AHIR8iKrS9rceRpgUNuC+h
nQu2dabn/v2VKODwvj3BV1nm3rodRyTkaL2/g8TxOFENnNIRCC7Ew8H9iiELN30ZRISaClRWdbiE
u6fzxAQKUF0FpHJL9Q+0xKtHqh31uMZTs/LY1QsIsMKcfDPRuDshWX2YiTrk1YD43+KhFVFOBlsT
nSruLiZkjbNAanz7Vb0seaNnJjW1MruxbkeYWjgTpwy3lTmWrcnwhE7mYywZ5DK+ZerhNadvK6SQ
YhztCNmxnPvmpCIf8jBVD2SlMmF3jorEomgB6XmBesdepQ6cHCTW8U/tqkPqQHArM4z2Tiu163VU
AMWzVqBXANKZzP9bLYd9g9CUvpSh10SsrXrZNKQ9U+JwcIrAsUoEJTnHiFZR+oLOD4bF4t2oYktM
aFdMG/+I2xe5LDGXTLZUnoXYC8C34yIL7GklK/0K9gclwLa42zvVqSScchdN76SkSR/VJ+CwHhx3
7tPK/9pmVRK1R34QZBardzcKw0FMtbjf+GRA0/saxWUE2h4cbZRhfpNn2XVm6u2pZF94OD12fHLo
VQTZKoJkLgH2fj/LnCyxBSsPCbm1yw8rUpCdp0gmu2fieejinWr6XUQ+yHwbRW8SAZ1WDXdw1D3H
9MCDKkTyw9RlW4nX4d4lICVpeExuKDjUuufEXS+vtmq1og24op7AjFEZGov37mJbQOLWp76Xdqcb
Y31QJIEEZ4VrKrQBLfBjvBf6Wese1JrK14Dt6st7eAec1jzVPnbDYYM3ZTLsCsWEnrBrVk/4AYL/
qwRGQr2FgELCQ2HqVgZtNNDo4pKX+TlgSY38NDkAB8IXpqnakqariIfoiQWGM7oYN2Ly2TcjDygF
mOHd1uyxHtLAkA5ZhI7xr/405j+xSHUSlh5v733N1DbmjU53ykn6Ag1UZ+hdKAMlZ/0sWMH4Suv1
TW6F5cyXPzpwq8tkkQtAKFGNclnK9+Kjk0ytZMqOUKXmDPClFs6Wk/3Te1FeGB8HmWGBhXcXybtd
q+QNkkxNITqfwjNfEXWcZ4DiqZ/5OTWRAE9ZC7GIM0UeiElalcbf29MG0NwfUUsqThnvP+iqE9xn
m3xPPt4A8Jm3hcFYamlZeKtRTDcj/HV4dLHVllET7wFT7lMub1lJxugcVkB189+rI6fDXnGpCyMY
qo9VissaaoaIQ4nqBYud/EAruOJYo9ZN8rZ804SLQazRSb59YTTnZgl1ne8wGDu0nKRg2EA/4X6X
jmivW4b/1JaCWOevK7OtJkhjcNq2U0SWjCdOatHXTHDUTtqOMWs2NDKqGR5XOQ7LMHWr/2Lpm4MQ
cg4ZleCJ8V3Als+Xas1r1ARzYo6dTcKXcMY5G7ooblIPfLsNY61fsJX2+GY5uZMkymdEIV5vyfbu
Zlq6lWpAlVvDXKchDOBbMUu047sjdqjNHmUDcuGuc5g/TGo3R0bfFhf7DgMaKr6U+0jZCDoHTmg1
AgguuaDbgaAfnsrb9PgcspECwz5rK88SYTxBPhVgooTC8YP9hXonROaaBELiIKQyY2nY22h2lART
c5PPBZ6pMAWy5nKLMZM8hj+DEXnmY2dSemMeo9Ndbcr1PP+ho6AMrfHIrRXbq9cNpdgWEu+cfpQp
hc51rQzndy8T3IXkG8ETPHkT/YpUncWJod3qNXpFItV4meDdWEYLxQwY6m6ar+PNNWRecezrVQ9i
LcrcV5gJzp7Af4lbHqJTxKVqrrUvgmEyN2bT/i2jvWA+6F6sejAOmndiXi+oeBz7snTX2XImb0Mw
35/gzEPbZREpkdonUFc61R0j05635SHyP1ZakUpFM5m6uAVyIgaZkRQsr6IMe7veKF7gMsxtsO7K
44wjjeVytJwEhnNGkGItASQdUwU90ZeNGFA6lSvCQ9zQbmtOeg8HTIJoNW+FV1V57MUPBmVOn2vX
Dlx8WWXkIElxUECBMFXHoeyyVqDc4Ko52HP6nQANiv6bdRlDqWuewCkuKzkEAX56A+uryAznMoFp
zK5jYyo1+nAIS2OVrOMWSR10XXGG1OnAwmKS1MwkNZAr6j9obnxCM4Rbml2djvJgF5v8GqGgoYCC
hWdQOIYZm4V51b6Wzl3B5skIAaCTRBGl45IbVePr7SgE0tGs8gHxIKOvgPtWSLv0I50Gp5tyQR2M
wpJDr+GBDVMSZ4zTHENx3fdMdnH0JGjZlXRyUwWzwjHfQF7gsNQgYM2vXuAnwVTtCema6vhJcdIu
WGkT0ejhwVKV9ikSuEJmc4mxIvA0nvewamDaXtbUpES7S3ni1UDpObrS6X4GiVpw6tZeWanYepK7
prqFLoNyvOqijUlJgwQU8WQSXiz61/qhipQJc4gofBNW8Wvktf21pP25owpB1hKI2JUCj0x5kyz/
oujO8FR7bxNKh3jgN79gJ+syE8cIocrMHdefdGZqNCILBIqq1m260wi1unogWKD+qF6XzParMuLP
ROqsLPqXFdAUkQsOZIGXzur9nva6zQzZu8Aal8/XZiK/Llrzwq5FyOso8UtWzQ1HXQJd54FpnPgE
ZgOHvYJbxBAHQnsE3cAcvsV/vBRCokN6zd/XmXVycL774Gyp9RM7ROFXsYewVjKFjFJ7U/dEvKHy
3RgJ9eX2kSlvTYJtHQOJ3GLdXOtwuxhqOgMFulCgAs4xAxWOxxJK1nzhdyBnwmgZppLYW3lUCl7z
VYx5cd/js9g4g7AEfWwmgvuVr8GIQ2mRlYUO3dgOH6ed5D2LwZRr9dxUp89H2g33GK6BWU8+3THj
Qdk9Cq7EONlF7R9fkf3gQlI2OXFepqEQB4kZn8nev9/6Y9aOxw14zU6y+mcj0o1vPUIFcrlJDWra
5wGN/EhO6mlvaB0c4zrZ8+BiiZ4wQdpSBgAI2wsj/RkGXrMiRCJ7EsRMaRQJ1IgJohqs7mfgKun/
3UWG6e5Xq917IIhPfFVsbkwWhB87F09NiPoBkReU3R49YPe+rkdjBYVf36SG48SDVDvgk8rEb6Z8
VKCBgMCh1IofQtYM3nBve7ZbH/4gnpIcO/RywS3RUBBIutxvEv8NLt2wPkHiwCGMLWv/cbbNkHgt
C48pwARbavowzGOM2Er0gxoYKHwiOopy81cLoHxxZJF6avLQ4OZD8d9SiQLGYRvrHPqIjAkES1J7
EsWGhdrj1ZojbJ/PgplSmQiFbnqw2d9eS/1A0jDdAKK70dDfFtqLmHVlPUwPHzYP7q3UnLNE8nEs
AgKAyLIpj7cTckwGAbh1LYACflk2VqW9uRZssMmAqomfy4oKr/CvEllme7cBzcFzMzCpqbsUjpjs
cL5NNN8JE8IVXm28k/jZ7FAyw49uB5mxKryNfNwzjSTw1SD4foL2fOHyeQGkcpEIqujiXJhILqMz
6AoVfSJfYhuidtL0p8OGQ0MswqVuJejJUDd/SdePaQFbeWGKY+4IpcD8LdKxiDuyptA9H45Dwqvq
+rcuku4nIqXqT373DliypKcw8P6gmAtaKumdfq9yEeeQgd5Ksc6MeMBinumY47+zE7UdilfMargL
Lb+lCTRMrV7mzgTBNfwaB4TcMxbHA7tHoerV3KmZA3AzEZHPB1liLTmzx3192MdkY+nplEsGH1UL
8z96MMuprNO1k0rqVqYQC4tBR6+qMcFB4eQZkXsrHMt2fpmvkInl7jgkk0YvXMSSwcWPo9FgG+N7
BqFF0ahTJy28GPIH7e4nzOwZqimBU4UHru7Oaz3uT6ESY512qtbADkplN18QWwPkSnMEnP6ScRkZ
ACPq5plaDdawAI0oglvILAlGfQAJdFMnIUIyHFo2i05kwfba4RXukCSpSwCsPhEr79MBLGVymTxl
+P0WKi9mSGPWLXIhOU0MhfdsQwdRXxIxsPgvpGoBXhgJqwUOQBIL8tYpBcwCPr6s4v/VLgGzAiH8
T2LsYudiK+tqbcL5seKQfLYj+Qr3gfs0jbMDqQPwlxE2gt7RHMbHrcJ/UWQVTt5/vPRWMMJb+JFG
+hxHGEeABD9vzOnASzUtbb32EdiR8Zb/fm8cGKNpUIPZ/+zxlJS/4iGSt2Ea3RpgOz3DxCKcYaKC
bZkjGrsZiv3qd53GruaYvlcXV+M+HhxcDb0qBtdAqu7Ji2UtvfZ+N83/rxPjUnhM1b8dIIb7LUqj
tCP+dxzrTipnEmWTMIGfwvlDhVml77+sF5rn0vDp1PF5d5UeH82qv9UiaDVNccA4rponXkwwyj+6
l/HOZSp1vYU+fjnTQW1eAiiYz4PYZYlxO+Yjpc0EmghBTQuwQtQcdSpRrBLtuezQU+rMJcJ2dn+9
BzEYGwSIkKskkSp1A8otm93bMqz/ViE8na4l4a2YBdlViJXVmR54FIlRIkfWLVsFM1AtxUqFgD6g
GfLEbHd8e81LT/AiV2dUKDQODhTr/LY1y2uk5BEkReQr3ORVBjeRXQbkcU/vnwkCxl/epxmiuUVA
4IshqLSIsQr1VKsoofgiEGiVIPLjot47+lT7XwUYFNo/TYlPTdzwhDFqXRCOZLajT+ZPdP9o57bM
tj3B3SQG2u1wRiHIB/fEAO8TO53wYTKvDiV6UahMOCr02cEUtk7BKIU0MDEzpN8Tsi1BpMq195S/
xi5TH3u7cAZeaD1p41TuhvewaGpmKZBACEYzk2YMpp0rpPd+FKmlw0e/6YBQK19WW9NY6NI7DjG7
+5nV3xjYbFXVbjqNf0tNI3qZvBWOGsTzMJEofjqhQPtiVymcA8H6cA/YC4s/sMT5NXH+Ntu2fTYw
pB7JnLGqA8CItkkrmEoWp9ix2IUadJYdnhI9OYB4GVkzdyUQQtiuDEH2xliET18EKQij9kQ82Ku+
ZPDFgN6ZE79aevCS/VeRtzxxdnjFUEB0RK5ZSaViYJo02OMejCCdf7Qg3kRjV9hKmEY1j3rIxamQ
HCHIvmQw9VCh56mnYjSBr4IXB+xYtl+lJ+t/iOQRRv8zeEZQG7Ljr23S/AVKs2czNz/4AO++ZX1e
44leRA8wNjivfnOlx7mpjmsvBtk7fv/uJ1SnoKa/AQi47MQY2Ljek3+K+UcQOjR4tL2/51S5/+IC
dqEfsOKHNql2a5gsc+jiksxr2R9EvnjXyfZgwrttkiypW3mm8es/1YJ+f0oyhBdJPM6RfMtqVDJb
56gImMp8LuyvS5el7HD84ru+MRW17sZMaP20WKAyU8VW2d/277Bd8oicjsURGvzBz7DRc4MkI3MU
bo2cQI4Qbn/N8ncunT1/QtF7vraFMxgaMDTen6yw2sK9qEugdu5kqns/CGA6/yz9BMxFQWF3Gbr9
14MDWQ3gwAUd8+7gTlBZRba9LnrjjjcXI5Ug/qUro2tt5Owjqf/1N5WCxT9RPpKEUXp/DM6y5ueG
4MVEAxoE0zm72Z6CpN5ndZsgB0GmHXnhnk20N3YMENw4xXSyEVgWwXMVbS236gradxRFyA1U8jf5
6CdoLLD7U7MGfHeikscATEI26Yy+rfIskKlT6r11at3+Yon9sTzWE7QYVL5IXjjqjQXqOB3AR04k
JhH5tplSsp6+hqjXZA2jK4IL3Ip1n97RV379SpC1T1nWI13PpTUXMzmTHstpAVz6VdnIKT1uWiQM
9zERPaUiht1MvlXWm3HLG3WdQtZKA2z9/WhvsUUaOUEAfg45ulOck2F4SMZShfORhIGvjku06R5P
FiMqtRjRCo0aASyOGyEGRq/T/teFOlV0suaHMtU4Tb/DN9Q4HVIeON26G0W4o0nn+JZttDz6jHiV
xxpoeNpenwZxymPNuhIyglR+EoCGHnSZy7/3w9FsQjadT/TyLeI9jG3qsPgk6DCk3Qc06qpQ4VAC
kqElTDj3jcuaMUbF/Gyw+gSC7cgXfA0LDnn6OB8gCSyo1xueNNG8GXA0gDbmX0DFMiMFof9Kyq6X
xZm5ft6GVcFousaagUO2UyMr/I1eFcJrJDqXfuLSQXPrA9TT/HLt0+tGTkwX579FKAtXs8cxmVlJ
r1OtibQxrXjQFZki0DXWpCHxS4ic78+jU6I2CoDxmcaPqFuiiJHOdnupaVKLgcqYDWCRRUZ3urLs
GwiRQ4Mdr7HBrzw+OMFnEHF9qi5cVduE0/yqxtR/Xxi96eo6yxxTmZS7PEVTVgMLf2+GG1NrY+w6
+hE66wtzvqhDqZGi+pKSD9tla4QCkM51RKq9g74onsZQzVXmqd3W+dCj0HiLlJuXYM4GcCE+C2qu
iWPNL/2MIN886s1/66kHoUUtgxKDpYcxbL/T+u0Zbqa7a4cf2ZMWjZags18OY7ot5YSLpFzrrP3x
/m632uLFHar9imCoUtEFJnAWR7HzoK0CI5ffef8Vb7uGZ6LCYeddYJ6MruXKMwg9SeR8hWcZxhhw
345yJavnZ2gH2ePILzJ2YW67Zw+v0UEA38zZPJfCRCkJcTtkf6h/9zEW0/agju9eA2AvSSXM0oTS
Fv1i6lIdqGWQjrS18YK0om/Zo7xVnrI8ZvsLweEbxFLVz4NRKk35EszWASV7jKMIDx4paV2c0iBh
GNDBFjRyhFzgzKrZleYPfJgAgWDehObwR4NLhMyIeTwgOqGKyYoD7kHod8+qtkPVAu9L06kt8Vq6
iFXjtaO9FofDFgljZDInyZVWymTi/5+qk3loOsBs0t6oho0UTFSpYx1jI2HN9IBU/N6JDz21XaXF
wl7df8PVu+UBTpJYbw2jfV/b+/xOwVYuntgWMlVnQu/8lCbwObCVq+xfubhCKA4UvdxFSnadhDsG
Vq3VMkbPKRkmOPrBIFr93nvfy+VuAnub3XRlyWfdIQM1S/1gcZTQgMhoM0JgPj7fq2/6sVCWWZlf
lzoqOr8MbyZq9jsn4B6L1qTY4Fh60Ei8d0xejpWEqlliHyeRvAgDk2hKYuwhNEq6EO+fNyas3xd1
PfFpFsyt6DQCkBPXUx+KREFec2K1hw13bDQCHzGAk6jTG+qg6uL27ZWd3Ujzrr5uKT1rb6fc3kfJ
hFx/5t6dwnlUro1L8oj5B/J/YXv6P3qCgyY+DQB+Yx0NV2V/Ja9t3wZpjXaiVWu4WicslvIQB6pK
T+uI44Iowy2LVlM0LZsMgZk0Y9BfWFzHhKvjh2Y4qaDEYhPUqe6qxQamP7gCxxip6AaQpyr7NFB3
mM6K/o5pMVvjtahsZVvjm5kXYHWqcvvw1e8r4GY7zg4F6yOyHnYOFQtooYR1dEcG+tgX+pHapeQ9
AXmhlg5134BJEm0UVAfj1dj1pjtvsDRRZncw7y2JAOWu7TRwvDBh8Hxdg/apu3wlY/vBj9IMSLK+
cURjYkP2L2R8QWpNZAkaY5+VPLuP3wEyk0Q2MG1gMr37SNHHUZI9nR1VU/omSPyjTtBn2duH1Aty
LFzoD5C/5XIAbBob6Y7+TJYR+O+hduN/MRqW1QRaEtnTmyc9VU0cQgC5+MToAY1kjkJTpd9oxeEW
3+LwqehCBwaFcB9P8WIPx6kf2EKwLHaOQ/UicNMtoUHmq/rhQVxiyyRtAR0sP9DVwaitVNW+hu8E
gPcQzDfuZIfg67Vrm3NeEta0yaznISxomEGm7p3YUW6OMpzyMR8Jnc8nJVz/EdRhJUFLGoq/hkGl
FeEXcp03ef+PDSH/xMtGPKKrwuGvReHJ9mIUleN1RFJ05UgWs7Lvtxl+ixrDMzrutl76lOymRoJM
sF6cff8RqJkBdGQcYdr3pWdnhKeWMdXHFHVMpIsK0WTcloORrAwe/nF2ietbdvi3WshFyeKfC6A2
FV4j1OW2mFMrofl2sXW+9Q7mNizJppcwQCbTKSE6X3DyFI9jZXA3lNc9uqSof7VpVwU3dpaXH5eE
27XpxYCGzKFYsGFDwcrhU/ZwnJM7kjVlM3CxKMgXwp6sh9V9DM+33qqPhlWEd1jzpqY1rjtb1AH2
u6Chf7tHPfhtme0G1vTnJtYDTf4xtq6krmH2YElIH5aFxYxIhh62vfdCmez60Sypd0X9OxFbe57X
ez55Bc7LNdfpg+V2Qf1jlHkRyIpECmkV5/JGqnLOqEzJR+XjQRRynS0zW6l9ni7RMu1jNjWNiLAt
JG9/HaYGrfeW+T3y0xPXaR+KgJEeBxORsr44Bh0nyg+a/Zx6dPdruDG/W9Ec+4+C46ekBSDS7JtD
ZYE+uYSvu3EFGKi6wRYCrhSs/u4BcZGqdoDXWr7oVTnv40JZTktf+ysdboGiVtQWFguMorOg4p2e
AT2JclGvkBJ8u+8t45Kwg/dDT9HAG0IwrAAYt5qCQnA5Hw4ro++UICG5yLJtjBxeELiuo8UCdKpU
xEOCGeecR8sfjuc7Jt48tq5w/NUUlxhB60nY49bR7eI1azD06SKNrTi2tMplpHd4/d2J4sL/0iSl
cv+lHUP/+37Mvf45K2bWT+OHHO2HcSM3hSiMzbr6HpAValpIpg9E/+uopSIUjoox5O1Yuz+AktIB
xAhM3drUPaTQziz3G3O90H7tqOEi/ucA7uIwOgeKniCrkWypyaOysBOJyxl5M7IOkp11kuL94VHv
zxNyRvfx0vykTmSsLUjaNzQGmEiTFizNLK0wRSUBJzmNpRo1TtRWMiw+10+F/3l9plCvMHtgFVxK
IZZKySxjs2ss92zlitFpfqX2LqOixO0NgUu0fbJNRvHTLlqaCRlZVLF9pWTYjTA9y69jYpIcb5v/
pNZ6D77IyFeaY7tqLEFHIilEor7z7fEg1RBfLRT4S9pp9l1eoe2dRvjOgn1q0+3xxtjf5IG/EWJY
wSsWEwzddV4v1bP8T2+DOclHExfCrm+ZDVXYKAs9EcCUlo1sINizoIjjtRyuMD9d9NtzZgWUyzsR
pGPNUFllNazDav6j6VOlfP5qXpPNqv7Do+uFfuYTU1UpUY80Xb2ee9olOKLDWxetTgNANewk4wlL
s24s02qbX1Kdh+dvHZsyMqUYVMJjxKJbegnh8yHyawQwFMmObfgzCNVNGFSFEsv1DfuFKMsqfm6W
ZPjIdneTeVumMtL7dJnPbZi6okHMEAHEUYYrTTSjljr0yUD4LnqESKjFmnbMOnaLINboeehZGt6x
WjDqcxdA18d19hSd75O+PLSIwEWirhvhG2ZfTcSAbgc1MXb7Zl0HymsP8g1R2oK4085b6Wq5wnJF
MROufA3movtohId2WlACiOYQOQrqre9ELmSGDaiWAVXCrTL1lLGxUB7pvr9WPo65SOwbqJTtXPpF
P6c9F1FPb6LH5fZoYUSF/Z8WP/cnG8nW5/ttcYvsxqaQS1LMLgI5S94NlKNJCgRvjB4Mw4fs918o
F0KF/doe7dpItSR+O3s6yYaf+KDgM7+qONmMK6+ohE2YOmzdecGIQ0TtwPqn0BDDjt2DgCWVyqAN
XQ+AHRq2BYV3ZiZoYplWN2jg6aRSrQv0NU4q8W3oFLEDc0QP4z8KE5QS9siHe7D/dPv3vP7q48pi
ELAADgQHxfr4CqWSakAahvcs2qKSr1j3ONAFcN1EErTEsAQYdV0/YK6oO2lII9mVv8bxqTfmKCjU
eAv+UMPSUONjCiL7CmjvLkx5S5SqhKSuq1kuJZnPK5W1DQxd6pOTejVF0EIWga+l4bKPf5tAmYYf
GhS7yhFd4jjV8geQEw64vRN5JeNnVQjm7Vahg/BdXQs2KOKxnqoq5S8pbkt3c6Ewut8TbTi8APO+
SQ4IaFsKWXDzj6iuehpIekZtEU7zy6U2p57JTZHhGhvZBG6Ugk1mv+FqPS8ltEtWszXPM7EhK6uW
0FlcjQ2RGScTGstsIUL1NbMVP7WvGlpE0DsNqqyKczOAm/WWbHMoIWnXsFnEdpzcEeDK8CuilTnL
pGnLBzAT5/N86PiAMrVRVjmFO4wgbHdt8qZYDUlOj94mOF/BvW4ATMbuUCrD4ZhREOKV8suPx0Iu
LbFWGN1m5Zz6e97lr6GweVQsv9U7oxrkWHD0lMjRxxWWSC8ZqYEcAu7coIB29xJrMMYsOnC5I54w
fdpyrm0ZzhzGVGAdVEp6rCjC94zvRjDH+EaIhdnEnlNCe8ABzl0dYIQZoCpJc+rJl6tlSIQH1oAJ
0Wb29/Lrvc683ll/18/xhq2cp/zb+CuRbYfcQr3NULZIa0KjITxhgMOFXP+m6Ja2elBZpqCq6pUI
Up27z082Fs+NRTvYjAJ8rJBvCm5YNh3D0rwasMCigfTJUdgPyrv/AMVma2tOc6MGIqo5kyQi2Ksv
MFgOusvW6Bk/3VBfX4R7woJoNbWMc2BZr9+vY28ZZveKAyIVhKsU03ye9wucRX+mKHDNRdKt8Vfo
VrlsYI2+p6PDckeBgKOguQrbi2TilICrPcrZWk29FjjlesU+v4fpkGHjLv+0oED4bmNvM5cn9Ckw
z2Yn7mh3alYBly9BM3+0yUxqHOwhf1C474MZG5j42RAzvkA+u02baUeJ1RAyiKsPdh7pIEZ2o4Lz
O4SLb/q6EP3+u3KPCgJu0c1NLMTHMu2WH46KOshLYBw0riHNApabka4L6R7dHWcYT66c7pOsnnxP
xfX+ewpFcF6WCUA+t0T9sg5rA698pUOeGfkIzn1O7bQkHl7Zs1tNf1tPD88L2p6d3WqUzQJ3vWWB
WXhmSq6Z73mKy9IRmHfJs3oXIAfz1kEC3s7NO+kjhamK/ugTbFmnVvbDmPKIpkF+r/M1P20H2TTO
KR4DlW8Qy/HmZq5vpDar0yD0LTCz5f+XhbFdu8m372mFpO9Uj3qXBAjmNxqcox+dSoWzlOE1O57G
oiTC4JwVWaiNXR7UK8RrUb9tpvet02mzdYJB6t3Yna59b3m2M/DuRH+dKPL7O55KfgsY6DAu6pfZ
tWa5iGGHJ8RKwZhSv4/kBenahC5MfntOrel0TCAyrdGcU1vmILee/hpu9jPpSzAPYhU8cpYoDGyz
ER6kH9z1gi/E7TTkJsOeQDAYZF/sQOICnLmc2z9Sq2qpWHQYf6lJGovCDldCZpTdwdxaX4g9Q6UH
7jeeYTPtFPGC+VPrcVLO43m9cTspX/QJknVnZ4/we2uxNAZPclaS9HIsKKCLAfxukunIJwUZ3wRz
Qseb6wldh7bipLwstL9PrT6/jrucALNACdXUQBOEGtrpCZ3+ZhLl2sOtk4+EuwBZIRa45Euy3lqq
vVIYpYUEjQKYHROdeZITaelevKyeDFUMizOB7Q4R9TlpkSgTsyJbCpuEfI7eJ08eBW7779ecHaTj
Lp+M+/p/dP3SoFs/x+D7fFEPZ9Z/AfyhJnfsSc43qrGPvtFOp8EIXjlG0Nz7NeEii0kDmOX6Ky8b
YopKgk3KF1/OZG8jWtmG+d7iBr5TdntRqdJChnSz+Z5f4nnm6iMHoeyiAGZabbBiFhGao/fCtThk
80XNoBIAAD0kOHa17EHW0W9naiWqs3jEETtEU9r91De7+tJpQ36wbTF9n4bHpgcEs60FS4NBKTf+
qrc+CHIwvZ0mOjNROgDfKbFmX48k/dxWIth3TyR0QRd9LIxE02QDPMDMQeuxnlUxYfYAuEJu0po+
ONr+1CLmK7OXBsEFYMggGnnxcC7gmHP6hWs4xHLqTOa41JdWCugFDzN5CCc8IQIU1JCfKI2k+8Xd
tahc5ppPrdiLJ5cjUCKhMopzrHrRQ2RdQ0hGuIHosYzjWJ50/9e/v0NN+oEkbSTDF7bsw3lq1KDB
hKJyEYREt0zX/OsNwkdHhArZaxrgcL8BoWLHY9CvVDK7ARwkZWc3j+MVaP38gjvBQb95yCkSDrct
SO0Jxj7wZ58dTaCe048WL43ks1rQMADDSQPLzWb3NQ2nNkFVbbL8WeB3KxGuaAiaghv3geKPLEaJ
XnjDf3WhdFYmqnNc7vebcrG1WPuHmDovkF1K/DI50lvFb8fHs9aB7ruhgmDrau8NyJ3hG/gwCmvg
8eGrH2p35VNEzTfPq3hT3ZOH+1qGN7oRabo+ALGqMrza71GQXDK6zLK7GgzSrJFGI4nhMuEhHg1B
ugyeke+iAghAgShHHEvqcDUyDsNROVKuWhMSc03c6own34LYeskGltEgblJUlLYPwqPXDpOyXKht
iGC6K8q4xA3wO7Mqkj5X7W8HFDy9HonFL9t8bDZftO2rXUcPIuc6LTYwLS0rLzUfdiQqJkJm0zBZ
4g5BdSClBGplGHBkEBD9p6wpoHOZTqStky7Wg6J5F3d0xwyVDT4SO4IbnGsZs2WhaFRs8TfJXVE9
TJ5rJHIdGW3fmQHaIyVBn+0PL+uqm/hJYZnWskBR+uDxF5iLyeZEkT3FHh2tGFXYZWRrkexO+e+o
N7Yse7RRkLK+HV1qhLWnLg+JIcl1glwCqDNb8KNnnqOt4Lpm3gZaAPXcSuaK/Gmf86NKz6/xBnn4
iefpTiU2wiZsh46io+yVB+rBVw1I+y3JCo/yaUdlWDZFs9dQ+k46UISiCrXs89khMRF4Id5+8UL2
v4JVBrCwolITHE5Q6xsX76FD1v8dat+mWj+u2MhsXa+aYvgK3fPr3ALlQcKv/2AU8Gw6/toq7lGX
wKY95P0jjidzwaGK/XArleeOHP10z6b3/sA2rqyKwRdaY0lj2skSzjmAiCB2IeQ3TYXZ5PR8Ljtf
848gwP8hnE5V/Fbt8835LlSawgfoCb9V9NpWm8Y5krrJDxWBHxCIvx2D4Pmn8T9HS29tspMIzJ64
lRoIbBDLQ/68umaE4vc5uvnSJhhhKxGkNs4LpwS45E1spubeYy7eIY6Azm2on3DYjjGINAeUSUqr
Qv2SXUALQbQBFbqC0Aott4AIDOJzF8qyKpYjnOQs9y2tJSSw2hHaiLkQFYh/gqZuetOH8An9PRYf
F4/ASpq2DvGSfu03wQloRzxeqkeaO1VzBdN1vgFfHr54qVND8AqqSC53bohZSsOG4IlTpddI5PbY
FTqIX8/Rto/ksVClcnwjgaFzSWQRM+Sk+HwQ9/3yit1RkSz24IGNWDPnVp9ud6GoVA/3TZBm492o
sFBnyjhgPbY1JbXfYqD0rz8OgZTKIF9ne6/dSDm6julgn+pdTWZVolcJHjewNmQeROwq5L2MNQJ1
UG5tpje4SO0G2XPB9XRvogZuYyVQemlqqoU768B8LMfkrvDCmjjQ1VSq7mtgfxSmR9ZxoqDzhHrN
m0fd60vQEyBjNCK37B8tGIzr0448iCr0cWotu3lffvE8ngtwzqDrT2bmRl7jeDWutbPTc2eaBF8G
nK/T6uEDGg3nCxIkIyEOphq/lsaSlvcvGy0ChVycKaI90uiGK3znEP4jdFeKrhoZIxcE7t4RpC6k
5Br45BZrVMLv+iTVLPxyXwxh+ZBeTh0VKMEFB0LK+3W2c51K9Z7xPSIqUTVFngjzUC7QxWCALK+m
dESchM5pneX993ER+4qhFKoQ1EmUbzp1EAMcpKger3W59vQEOYPa1EkIevuHFmrSkH7teWMVhRmN
wuDMzx9+Ys/WsdWo2xI9y8vSPXy3hW/8LX5DAfy0FtzXmIrR6XLeJyJBzylpDDD/GiuZO07uyO3n
np2MR6vvdzdTGOvqOIL0XALnU9MsE5cBU2mCGKLhO9hYnYI7URGS4uKXqVu5gXzysmDvCK6bbIsC
aZ4eVE2j2ce96qTAxuhL0y+Q+PX80P+Je+dVlDuOzEcH435cL9JOxCSb2UBZfzRnr0q1cIwxOmVL
dROY3BmE3pR83DZtP2PAIghRIl/1I4kF2DcqmjEW0Da3X1w8mz4QRJPxNPmC1VuCtmlJDbadp7T0
ERbAdkSMAVwjFGvVzRZzJjTasM8f5RCiqi8EOs7RzJhCiv8dDYtO3vP0rfHzuI+mZpg0lpPHtN4e
MaSChegXIjulb/lOL0so6qJmaL8J/eYy5SyPqEp2Tm0YsCXWWFLQ9AY026tkCvU9r9wkj8ejfPGH
ndJhy35kJWyTO45Q2PQMdHiy/UyNnTiE7/TySPAcBXopNkZBxBO2KCGxZeg0WG3Xo4clhpn65II7
nqvuYvudFRmGO4e7780QQ5ne5L5xr+e8YhbPQk7ylw8djonj3VWW3c9pFJxZ3wXbx6JQMskkDDLb
gwu/nvnN3JZ1HLFOx693uyx9susPCzagzpSGsP8504sBHqDdpa36vtQFVvFpAMoCE/vSla3YMneh
Li0hkYn5/y93s6T3rGfWlyLHXF2u0Ilr7uSxv/2jk1rmLSZbujDpAGqI7A1PkI8fEVJpjO/nR1k+
wmc4VucKeYJVwtGa04uixYsrdxqIkQpp6O6q75jISJOAIagEFxqoBNKefK88viiO/qwCWGiL0zTt
DPX7mJXkhesfyRe3PkJdBFwWegJmhDYP4CsEzGObIPbFuSKWB78Hvcuz1+24e683tKZcUGZ4CKlQ
J6KX1NhCV17XsrWK0B8Cj6f2pNmDcIZBiJmEpA9rc0sUMUPHEY2hIfw/68VaKADLCN2vY0t+pH1S
45JoiZhMDdgn20UBeecoSUQ7sEjPz4FesPUCiZW7i0ixegOq39NGTcmPn4gFXWTq3crovZbxEZ+7
N6sGcrgJdyzVXBBMQ7W0es9EvaVpV1E6pcgSEaTuBZBES+jpmpo3OOT1WARrxixJRLZiDrTlYPPS
pGm9T6G6S0m6+ZVSBs99HCDgjGquN9ZPzfb8x/yIMRsfCyDOuQtMAkPxBYtCeB7WMUOBQ+F4YUdf
jt9e6ZFlyCOyGUTZfKab9dwZvLa7+5/Apc/ghFelCRZyqOVn8aS8lJzEpANF4TaSz11jnJu/0KMC
7rcUKvZgL3jntiRr7LcsDR0+ke0yI1V5pTcs4YhMBCqafbaHRtV2S4n1u5o8ktL+hKJLXJqggdIw
gSMVdt98gKo6Dxk5X0L9LvO2zbOaGX0SQupv2rrrerFFWLWw4ReJBIEtO2IPRCpSRvqmWubZIWgJ
WJS5sMGqRNrDVRZq0gsd5+oXuBUK7itBkND+DU1gZkdngJ1ivrPinLYbEvhcgaQdjfn/oIlqH1rS
w0gqGq/yFg5Y6uA2SJXaJwF+OD6Qgl0d3fXCJxC9D3lzpoT9zpxUgmFPxCwPsDvwYB8vi3YZ3fiF
8bOYOJILRjMlCMBFjH0W5HiRI1rhHocOBnTmLtSkBOUQ4bTp9pUTZe585pv9yAOB5DQE9wHhIMco
obLGVUSrVPi8V/fLlOExwRJfF45nx7X0a9s3+jLH4uBNsotZN/i04OyhzRxA3/3OEs8MXpCoyL+j
O0Fn38W+znRQZ5i0qoCfIgVNo6RS4XPd0RXNSGidouhijJkIrN9djENYa5mWea8B3Cgl6aYc3PIR
HpzYwLE35OKIII83CTSRwZPM1MXpfpaKz3zTEWtX1TaoTjh86z32Rd0t5vJyRBzfYH9+6QHkfAQ7
0flSl/qp5RdrOjLAxVfCRCy0VQZBhkpxpkWuSUju4WEBwB6qP3a8vn8OYp0hWXp9Zp1P85jWWLs8
uX8SN88E+IgBnyon81utYHj4mIuESr+BbIrh3uSSt/qbESZfLSRXElqEbeuJyDIXvvx9FPywY6nd
CqZGIzVj3l1YNUAY5crNo7zN8Ekjb++kVsx7fWmCFE4SgNdgPVM7zZoME2OChBrlcF7Wi9IZ4nvd
b3bYhW9i65WjSwl3fiosuICJgUgFRbwFIfeDp5tdyF80DXMZIs6KmcTZYKM/YzgvWtvih3w802SE
bHLNthhWmiBeswha/7MjkKMhwwo7yoCMuOjYEC3DEMvgIyvB5Zi0nR/PECkZC4EsB/lFi54uUF/G
z5c7MiNmYdYQoSrG3C5SI6jj3Rnu80HQPnf2W9fyhNZyw4yTcNOao6GGyEfi+ikdNGWAzp7o/yTW
CYNFEBko3zJr/y/OAmO4IZCITRcGLJXbEB9WLybusf7fMjU33FaFcyBGaif/Y6xoLe0yDc9Ft0j2
P3SOQSP2AvK25FNDyFoCfYNinrf1RbZRsDRgR9uoFioSPMIWfBjMec6oQEtl0VrSnEa60L44ahR3
RpIvxRRryJL50wEhjBkJQg5U/tfh1SGdbgtjTowcYtp2WkYvh65iTTo4QVbvJ/f/o9bNlQ9DqmyE
qlbNt9XOTj+5/cJk4OPquhhICe7bRs5nMy7twWMNzsD9LPaI5AxZuTl4yH81nDfYiWLkePvSdxbw
wX32TK3/Knq+XkLofsVLnUmolZ4oCZ+/mJSWziSi58iUccbT/Q20JTyfUGK2bgGE3lzMLrOpiKXy
ur1tRVCipRM6H5TEaWKnaIPPXnClW1w6y7PN51u0r4tLckrsxQoakTMrJhHCIrbV0iShEIwvhVkR
sIF8ryrsR3gpCAEzrJnIfP0KJzGVExTW7SG8Zn8kXeoy3lY+Lm9+QbSA0KLQocbA4QFOKfm5tJ/d
llDCxl8gWEt5JVeuJ92u2Jjq1IpKPHhWlvkNQZlZLhYYOu96sIID8Jvr27uAcyhaDcQqbGOqRBS4
fLOxeKnvo/o46w6lrNJDOsy1EBO07XODkA3C32krCp14w4JBMi6CUA3OX/PBRU2OzuPB1KpTdhOI
K7XIc5CLKurnLOT6yZNkrFQTfwWdfEQ95EBYjaJwU9WEWWbkwn06gCuAnlR3nc/WP+GxVeqReddM
KKbR/bPbJMPiOyznBDeaHAK+lE7Cyv2sbHg81CbiUtogYbfSV4lx5auwG8Q7KnmKPFnf+7S/PxdZ
5L3uKb9AZubmxGJwqeRtmwWPMgaWNP5K64Fm4c6iOweHjE3e+Q4/1kQdR6LppDNsA7NbqyfwCjrl
iFN96MaxHDamz8mD1K1Q+vzTK8VmAP0knJzH3bL4W0bcvRiVYoATflL/CGGVVIEN5cVOp1hznw3U
45f0AZaHcSoV07kITKTd/ZVRzLaTejiOdtgFxVgIcsoBnt8v8vsQXLTh9a3ZQigXb/1t3bl2KtWg
a3P75cPCcR59sgNjdfEME8xCoGWv6a6qLrFX5N/untTk60TkZs9S5L9LHBQlnQHKD9F42eJtmYqJ
VHz4X3WURBUBRiNIrcnXOv7zyFds4tCr6w+Nr7kH3cxO5WPBBV36xZtHbl02j83soGMWhV9/ADE0
BVxbk8OSkLU9imLZH3yGvlpI0mrF7mipQcvwvBlFvHVIrFk3fdJKoSgMpRzEHdM17JLyo2OptXbY
6DG+gKw3BeojdClvsuQTzVJ/zFCfjl+k9O7nJvlO4hgVS4izpiCQbM7PYfMufcN0bQ5IkQtdbL71
8BMNlcNjqLNizSyCqXZW8J26nq4b5hY9jPqXzRbg9lnLH4Y74YmV1L4zc8hO/VWhQkYioeOPQcX3
34lcKeqJl70DtH7R96znJ3hFDrSmvobiQUDV2Q0qrP7lXNVjTP2gsC/n1TKbbcNKKdK+nO/pDhjH
sGf9T9tiPOdfAiQt2KMGtHr0/lWlABtbiI/l6wpkL9xXRRBkUJnxua0qnP7qZv/B4ZJpuv3NX/nn
Xv92C5ePRBfiNQLIs7xfoOEoOO/wc3WYheY7eNRONpWtpF2bMdVYdbIj2yVLnO9Tb4fDcK0V2XYn
2VE8skVqeN4xXI+FYBnJ9QjxvhulmenWkAejxYrxO1Z5+J/MZGQwvRnln8jpE7HLN20mwyEUuAbC
7d6CGJjg1Ov4AqIo5NavNAicu1Y2N3hgTJWEnBJr3ULHbkfiCNEfs3JVPDbitd7mMQMk+/ST7qMy
mNMhh5HQTqZE6612FaSN+EzlRLPLxnfMltvcv+KS0BkjjoRJxQHVHkwP7Zrqy4gWaT3M9FbuF2r+
c4gLUqbOPR7euQnPGBL4DNhiPi642JVNhfo17rG8orczFJonkPZHP/XkYmDchEBFeotNZBYy+EIt
UNOPiTvmFpOxTyR+bSDp6Hto4nzCAKlljXgFyfVF6Mv7kCyOd4w0ol6eOZE7lPH7PFnFfsDRJCox
7FoEro8/eQEz/FjaMu7UM8IWLSqJsiiUSa7EZ6Rtf94qDqKIJni3F19unxrJpMxWntD6CflvFiql
wEkc8pSooJ+XZ9+UzpsQxVY/QNpf2NjNZMeJZmuTWDNJufLeWWI4MscE9YaN8DD8U8USZQo3S0yX
aMldDG2/pYTprvIFI1qI35NUDKgqe0BFuuR7I3LBjnRuuO6caJoM7XsUgPvunZmFQM0mB0Zq8bsv
4RfmdJYRYto4Sd6sVXKqvUwaXozollx2hIbzFYcpROez1vCyl5370B8yzpqU9uB7F/zunbX5dsQ1
nX5/XWykElBi1v7p7jtBEXPjaVeeIt0Tcvj831z1NLAAlVwgwe63VH5JM2PfjXkI8egCpmm9OxO1
r1i44z0zFzj3x6S8QnLkbj3Ys6Tib+etYtYr1MQcaiIxlZNMLuXEfrG6VVuPMdsymOwKjxuaVczT
Ls+kPIxVDJ40w9BuzlKvxzVNvciBafeDOaWjbdMtLtcuR+5DHyrOExvBVpMkeQQrCcekTxJUxiSk
JBhYf57kHh/vjdwx4N6WAigXXoLwh43nm6Bzjft/h35nwSWVpTcRAOxfRlZu1yojvosDHpd6xG1W
jaCPBitV8+p0dRRzIZVaK/Sw3QQtEUU30C7Zyw2ddl6E+w1qF8iVe3pWeowRUPeRFZb9x6/yyd9+
XIaUZMBZgusypeADv9PlWQFKvy53ksazxIkVN5kYwFxGVadPkVwWFfaETqOBNsuFdr5LIaVmCipj
kpQ0K968aPqwl8lQ5q5RmnwxfN7yqx7W815vUpsFNVgccbFPh5UTvV6d17e9Gon/E3lBL6VrIQQB
f1cia7ElswxjOZj3IKE3KLB0h9+y/CaV69opzUunZ2BDrE1ToRdj8rskag1QkUCr0KpGPHJTjGMC
On7uWbjOvyA2OfJfztiysYNfeopzJq+nwSe27CIdEChcV81+E+7AKBcwkQOw6iwS4Y1kujBLT5l+
PnPGVqahU64veeqZLoHntWbSCD7NK6ILoWFu48Ig1JJz7pUJ1QI3DK5J2cnPL8wsqcrwMj3BVZQ7
4RHG6T+jbo5iChZ4CmyBqzKYcLE7njDtJDyPNG4iKM+XO6kpIWjmAYBfxOoyb/jSfplm9GJuAmxY
wU5BTi0Pn9hqucpvcR7jO6omtbeT/fVchOcvnD2l71HCazou7LTrRQOa7XUpS5sAZN/M+G7xjVrp
fNWLkGIMUeIoFU/fOH2c7ZVgcT6wtsEM9zbSVZGH4d4aFP/X/c4DP7bkHTxbe/HlActkwISu3du0
U+c3eGNMj8d737gFDgz66bu90ylgSe+9a04sjxaXxT1XwJiuXepnwi/y4U81BUYugrTk+/yWdP1g
KpHmFqOOduga9NL2mSN5ckUV/vBr4SDkuGQnDicdA9IdWJqkBD9MMWY26Pgg7AqXrGzm+Rsohqsh
lbBpLLfrKzz5MxXXz1iWvDqqLrUhBojiHKTdCkjlPxNIO1DF9W4rT4uhXN3YnKCmy7dog6cpl97w
/KlctTJ7Z87nPGgxMjGyLD+Q+fbVpRXqWh9I1BOS03SwqR6FaqGlrCGMUu05amOz7DU86SiF9Bwf
AK8tngkxHF0ikMRNV1ElnFEjFpBhkxsGiid17IqRfQyQI9GpOtUf6Dy7nnFKlQ4TEK+FpWwTUCyh
IuvFd1DbMGv44HE0o8t8h6TxzLwynNkVrAJVgqNI2LizT//XkTf7a2iS3rHNKKEnV1MdaWTXe8Hg
xbLw1lGO7M6UUr+J9NTTaMjtq/p+8YbaFRfnQCRdGKL++yfKhhQHmhEIXgMMJcGIgsacoj8jT6yC
EZLOAyfZWRNJVB0ocezgBbqUhFStBlDeL4WP6cqliFHjhiW0nWvv3SiJQQzi/B20aamEt+O/kxuq
MCR8EOuF5LalcccJ5yo/vu9mfUA9Rj5TveOq9TZBH7W5KBQprKjg89FmqOvlEigYbhA0Y1vbG3ID
g2axxEXtU4ipHdf2vTWcE4KO+Pw3CrghRxf5ejbjM+sMFZPBDqdK/gQy215y/7HiqHRW8Zy0RJZX
ouloDYQuykiqGCAHwA8VEJ/nwfz+Uizi7W5nW3KVDDaBYpBvZZlvK3DTeNwxUMHi0vnrxcQ0+JCJ
G+A4IavwSLlEp4mO2lqcDh5NYINPh2PcKjqPtz0hUaEkDZMMfM8tzuZo8LRkyiRPs4sZectHsjwO
I3CXS0rOd3lZ6ogITORLz6FEMK206i8wCLkFyCAl653aCfuqTRezrAacpai4rbWqyg9r62DhRAqP
bpH7QLVCqCv3jYU4pbseW8gbKvsU1jhR1FFLJVfXx5XKeo0NpdGaB3CaHu32mnl9nbsj0jCnXfKi
zf15z8pW5s0iZTVhcnp1wVwJ+1YvTOijT1hlFYUkhiwxJB7q30LskXWgqickBPRsDVS5NOb3qils
JrRArMgYNnIOatAQ619PMXuHznusZjcUBA8UZoJ6dB7+06U7HLyS4LQeUTM8fgHtKaxW2YWptTYO
wltTsp9DB2rVPtsfV8P4yoHTtQt/2SYNU05Ybir3ibDlE7SlNtllM97Hj6MWaITpvbEnrTsn+xJO
4UFhsXnv6dklG84eRfd4icBi7pEoge2MNRJYEzjec4hxTil02e0AbNZJLH3ykDZYyafXO/xh0VkD
I/ZOxDabTr3o5J3DsUudwXfPlNb2mCsXxFjowj069FqgZRmKkuZYM4bKvDpFv2O/X04pH0LTwfZD
ghI7Ju/rBJ39c8EWj0UufxVQO/+a66C2OwHK4kwslpkhuh9+nln0uevvuagtm6GKmrQVR+1gzUk/
zOEBsOwgo0exKIT+UfJkku8HlJikcV6pCObLqg5rrH6jE4vy9QhNIqP1onXkK286qiPOCXxodoZV
m2NxeHbpoNia3TaDtwYY9yA4L0iFpJGhsM0Zt67qJpQDUv5PUm4BE4JKTp6YSq5GV/wYwXt1OsiH
jvWzvv3sJqoQ0FIqUq5QvlmrSDVYaU9KjQjVes7vVCMPI3sgADaVH7dy0bPyVfp0QqjLIyG8GzNT
TktrWfb4z+QGyG8WnN5SnOqXSbMaV5klNnwAS5gVNrz6qKDcY8xOWfcqyKJrGUi08yx4wtZMKobm
VzF7P11kMijbCYuU/lC4EHL4dlhii0gTj54ncOgC1+5DZOQ/XvDm2Wofoi4QZyneNwjWZ6A4MrAU
p+q+OlXU0GVnCtspLp+0xIuSiOCF4y6hdNnR9mmuIEdQZExyiiWbaXbua+4SqZ+jDc3mzR0qM5V4
4HzhPqgtGOE6Uuh49TiaWTgL21c7+EkMEcphVoFguMfsQ4pCjjgMpX6xY9LoEYLX6sx2gRyhW10B
O40j9u5W6fJty5k5aDGB6t1y8beSLGuG538yYxI4L9489M4fjGI3xRuP1g3v1H1/kdovSDUH13qi
V3gp+gi1hEBBUun/fzrow7Ukp14gR1xIM6+hcBxQHJt2bCkBB+71yB9fM0NYJ7ViVHe4aRLft5sK
HbQr+5kOi6xdnBR0JZ9fZMtVPuvyioJ+pdhY7xIjsmIFh247a5gSKY5AWoSpdzhxaimqKLBB24/n
OZe3Ggps0Gxb+qHM0H1LKrNWv5nySaapI3DoC1mqiOU89YcMBh9uBHiZAyIoYTXv9i5QU8xyC3jE
FG0XhfiZIYSUC2doLtWF+Wtek2CHwl2+rZmfHKQHyTiz2Hwdf7/amOIjqW26H8Yg29zX+/pxVBdZ
sC5K1dMFVRU+qzdNXUsLSHiaLbDiWu+Gs3a/FGJRVpckqvnKlJJBxsAa2bRy7ytfI+UnOiZ0TNf+
kerVOP51P3Qokd2W70NiSMdrB7+zyD9/NzYJAxplk/kJhopaBzUNoJNZOMVtXtxTrpAiB1R9BJ8s
aGcOAEV2X9qmRkJIomxH0tm5dY+DYqfD1VKq9Hnw4Hlzd9zUXXP0+cY4ZtVIB/DRgK9jNUDVnUFd
DMO9hqGE7h+qcFHXDRtCmN1eJR3YlapEkh7s6Dqy3LDkiakcNhDJ40BhzkR2H7yWoFHJTRI4GBcd
xvHg+7LWJcFRSVr8K14zbCZbzw4XB+FVtcBLDnasC1heGri4X0rwINh9nGN55OKxCPFGWZTZEp48
1XEYNLVyRba7JqM8cTubGAEFSksObtGZFzJljzRWcSAeNQ7mJCGCfcQ3s2j9gf4ifAmQ0MRCAi61
PTB+6+kD+T4Ro1Cvv7WS4EhhyXQUl9ohXCvTFBTVsYkowN8tJBRLARptsUSqzdRI2YPI9Y6RwtH6
5Y3/Pm6mHZ8UPeMwC66i+B33W/joReiq6SDfgJ+oQviNSWLKBJXB+HMygAGWpnFyatCEyWclRXA7
gyOq47SrxyhmG1V/IEwowduReNKSwoxBmfiteFU//rvSIx7A9KAF5z8Ay40TwHaSxIzfxOMp3fhF
+r0Pz/tG+wthHptWLM5MlP2if5RcGUD0tZK9hKYy1ntfRBdZz3ZUxjkzBQ+E4ZT+1EM3D/rzcMmI
s14Fwo9dVUu7Z4GqDp3ZQUbNjegtUHtY1tY4kY9S3AHbTvOG7EuiIZgCQZUjq8gXISTl9CEtoAW4
K46ME5OYptSvIbNlNuQ+5j+WotC8gr/rxr05WyGGNY2n2pHTzbdBllcLznZtKHhMhJ8D3wVQp0of
dd7SPXewVfXyrUWgEwq4e4ibyUhoAp4cllDVTUCuY/qzakwJc6AImpP2ySC1fdsHGeOrL3LhunnL
6rNRQbwh6rp5jnJpqUWtE9ZJbDxS+5RsA8xteqCHqvqgCQ3LFfbIs9Sg6JrYMT5UQ7/sFO48YeU2
W5jNrUsWMMpBhxoONRDnqsfGUeaAbTDyZJZC5RxwX07JQ3OAlsYaydjvUyA3u+mlLrRQGJxJmTFs
YdKjzzFXyfMoseiZNubVsnfAXDXGF9AqMw6EmwHtmov40fXDhd09Qu6SNkcUKdoaZiNP7fPxHHAG
aA2bc2JJBAp6xduw+GsIi4TQj8h+3mxWntH1KTJat5z29VH/BmWJa26lMA9B8pTOqLDZMhV7qo7j
8pTj8f3VnCkcegpWMeEY2iJYJXV6f9z2a9bKqByHXcetmmRgotb0g+F1dYsnaGjr+IAEUdldD1gm
ujxnzXbAN0GEtkpfVVXEM31FbSGV1hEUltU4I7rGE9C0c0dNswEBxu3vkQpOOGWz6mE+tzyctMWR
fke3Uap2K1nVO9/QHGeT7pbVol0hW3k9hNgq2w+BHbNBeBLIspWjwiKy7Aaw2jnuyLb9kr9I9rfG
3NW/OgXbauAgRtXINVXNQKJAOjjHCl1b0qsAxv6VQre+9jz5nkNI6+OxIzRYnFoyyg6c5BferN5X
0UySPQTPv5/hWVxM77EyU3jtARx2VSn23vmsMpOcBqLfDqlINCBKtL0ZV/uku9vZiWY7e7vWkgc6
Mt3Tq0Ef3LnLl3kPXs/YwrX3jhxQmRsNluNxhNGHQPH9aKDZ/MITPFHfHWt2Kaeinzj/ZIgx4l+I
cVh83aSUQobScvZtgPJZoIFgPX6rLa2dFhDaPOw1vWthUtqzEgDOiPbUXo7BvZGsLYPvR5WzwMry
INSVaenEXCc6QbxzruNTefFCq0miz5CRGwUBAMsjgXOu/fMuAYzpc2maxbu57cEYH7z6qU5O35p0
WBhZ6rUkNaVPr7MA3mka6kDSAy88emjmm5SZ/C5aGarbOMDZilgjmh53EpAT8LysXLuoppGJcnaD
Kow8GAEakDhDMq85ib52lqvuK2OwIZ3psAmwWy4zF6lY0NoFsu1VARhpS5Gdpb2/MOIrK8e0l0nR
fTaktsfqxe7Ac3oHK9rN+pRQ1jn6+5zWhXWQelLhYdCBataB/YR4zTN3cRPVvTgqaIRgkzEKcrmu
mrQs4XuqcQvMF1k5IQaJ4EdIXKE1A1s0LPcScydpUeZFgPG14BhMgrOJOJlSWcFaAgLt2KD1xJ7D
8fbusgbH+Pqsn8OXLhjBLgUNjXd0Rbdt8HmXwDW2yCVo6Tvvz2nciK7JBbLF7iidLAvZEfu4cQsv
iMiFmeMP6v7vUzvApdB2vtrFqS/Fd3/vQcCLyNQBBe5hm3lvTzEKgnP+maKZDW7efNjcB+uPXrre
afTsluDtWWKPcHr/P2kk8g/MV8Ro2SPmE376Q7md14If0HzUVAuIfqX3glmCSLpo0BZhydeEbPXp
t3uv+MbMMopX048xOt51dgrb9OdC3SEjK51AjaM3b5x6RrF3nUIvwosTzb+wyhoYTtUu4vhJofEy
Q6JPY3Isa/o8uRFd8XXdUDO3H+X1DALBZfF39qmde04gt+l3t+whe0v88MrT8gUjzvAGi4swt2XQ
k2PNfXR6JD0J2kVxl7fAtnxbDWnFfFazoF7rvcL8rrLLy7fh0DXSV/i28zev/RYcw3EN7hR8rQRV
Sw/I0RKCsA+eraFRy3g6OXC2XReTmEv08hPuFpwwZrZCGc/6VTWaiXFjGP6KU0/sFkAB0vyOO3ku
n0kHZIblKulw4Qe5GvvFtMCELwstggjG/t1kiyXGUPlIrOd806a+oQ9QungqdKDx5oc8ux7Fm0ze
LtpDsC1xjrQ2qTw3cmyCgF+6UhVCptBTuhAJLJXDwARa+5Fmlt7VyPGckAqvtLeVkaVI8rijugdA
OC1an/r6lsrTJmWEA5A8eTzR9F6kOA/0svxxhlXGCqP+QW+6JL4xaz1drlaZda5sPaAfmldhIlEA
jrd4CEtKaBArc6ktCP1y7gTyEdOc6U4z/7ID1iaSfM2MVUCzJfzcQvmF23zIkW8JhDxEc/S0RHmP
x5b6jSToSWQdxhedahA/WN/nhxyoDQiFjjb8ih6wgT5TjggnnmKbqioYwUFffVmuUmZyJ95YqQ6N
KgsMEQxlXJGc5NeAneP6twJSVMe/fKg73kyEOAZK0fVACc0p0Eag0y78LJ/7sGS0lJzJMtiCWfec
GM607oE5HAfyhoR6msN894qQQ02LCAd8vWWJC1haSxK2R5sB/da5sl8oAbdngVeZQ8ekP41Uj/oK
gTZlHM1amP52CG3nONDw8Wk1/ibHjxg85gnyipcCTrApUdt3mDPMa/kzTVcVgZSHkV0m2jSh8A/E
NjOqXyxNaj8IIxz+RTyFyEgv0quUFnNRQYXkIGWPmE+qnOA94Yi8B8t6fTaI6VrHjLQIAXsSMqZ+
AZn0rn96WxnE62+N5qmZzTU68GNru8TYJiy9ms1CLmUPifK6X3JEIdeF/2FOfm7AFdQZY5T5mrK0
VsWOorFsny/D0vM93muznzuv5hhZKmBcZA3h9QHFrjsmFjHmIhLfvhYFJ6OkagUNvJ0qzUq5Atxd
bdOBQ4rHKCB7lE6ft0kH9wvJiY/iD4pKq5W1HEMwKsT15064p4F6VgjGAuCXVwTrrKzlGXxpmvpU
+kFc4K+9hLcPnoq7DDg58UzpTQGx2rFuWqcs0S7POP9fEZcpgl918Peb/HFimvzkUjvPPAHWrBRH
8Jx/A8mp1W9UBJGxb3jHtEufgeweBRZBECCiF/mi3UAKP+6a6YPn8XWi9SLZp2S/ifE5ivDvlf+a
dP967Z3vXC3NnsHxnUArrrl67/YLnMgWgILFescsxir/3oD2lg4FfMaAnHcGBCGJZWrVhKCU99++
X0qulWcto3dle7FEQiUbsTsMOLov5NGBttI8SvDpWNxfv195zXq60UnY/jBGrK/8f6QDOlzM+f6D
i241kWcCibFS2o65k6WHylt77pjrKxD+JVjHlwanZYi2Q+k286mMCKn5X7SfV/wVven8w+b+tDgD
69v6SzXdN+/n3oCEgdNgp307DsE3tY5xI2aSVpwT3DfTfnL5xA0FvR8JhhffuLq2ZJ4mNwRnRgsN
Z4MYI2C3ttIhRJWryfDt3X7zoF7tZUCfJgz+wi2shmUoiFJZCe8SdQZxe1X/DiqKRn2I6L17WGcp
wPfIuvuoQfbA0x1u5OeSUvMD5qylXPia9RTiJyCdNgd9XyfICcl/YdDzzfxU5zmrDZazmSkx/Wnl
P+7rJwqnsfp0xR4hLICP1ALcK0GpMH+tg6LL/HPPfHTY0OQ0OdKESHdXfnpMj9f+z1brUCz/4fwd
EAkVeCupNUhNCbVf3RFOl/try3yppx5yvjCcAXoZ4dGY0NZrBnh4pSdCdmd+dlvwtB8zMza0Czom
6E2p8jbz0jkKyeQK7lvm8qBNqjRMe4SfjlPmaRIEogLQA4XD5VeYpwflHNk1as5ECaUtVG3PqvnR
YJhS2TgRYxBeaZhcHxFeq3ee9+W0OYWIR486eHzsErv2UjMlILenMGeEU7OdgSVs19YPSKK6oI7w
Ny3+nT+79Ywo8vW8tbeThxzaK/5M3XcjeYgbkcYYwJPterthhVnDgbEgY9CADMUJqxu9Z9agTCAQ
5h1wYOmo+HfRhqfjcXscIBPSKLA5KpVMHtLNmC38nybJckijDvuRCE/H7p5aSmtJQk3vX5v9SfkD
hT72D47TZWPYHuwsuKMCDFGRTzL3i95978AAmSoKkpoDipfyVmepA+R7Q+2i0eA5Fuu05vGnpQw2
H3pAsSjQUxB+E/shgGttJWQW3aFVNilXQivqkK92ORZqabqY3tp/MPQZOAma6R50waXzP5JqTXyB
Y2eGjSFHJsAi/hIEo0mmlB/2I2jY3tdHfBVsvFz0RMbIfSsbVkjTYB3ddheAsms7zQ4o7G93Scgo
8lzHDB8PORVc09dQl9a1+1GX9WookYj/3LWNO7GqKmVDkRAEFQXZnSoSEFR/fbBLpWLeSzeSR+CL
zi7mXpGAFidRNZ+rXQba085Okc1ZgoE0TICPHj80F3qrhVbBj8lAkzm3nYnLlpM3AO7BA3in6VXj
9AB/iRGC+XBrOmVc7ys2uDwvr3r+c0h3ZCQ8V+2XFZRMqzruL3yNjBPBqHvUihqip6z0af3KGI9x
eIWCH7jKfGLXndGFN8H9VpgDvUsh6UKcRNr93Thp3QoCMUTKYv98yMIHKpd1S1cJqKoMMdh8tXDr
sAjb8nQeGZoajnBM9qel1jkc0+T9KdscTdPfxshrd9AYLYQX1yldDCGOk29oEZgYds+3MBUrkR2Q
D16ndU3pMJ1Y1+f4PAVPY8IXzvJbWSShIp9EpnA/lbLQeAH2m9VI50p+PLz3A/ul14s2/v5RLkVc
3KAEq2qwXmWmy7Is3z2QhdKiVwZ1wO8NOwkOU8WGux5aHu3v/XpWIMoMUvjdLikV+OK5DspPG/se
i7sa2uMN/V4q71ScYmYU7FBMfvdUs70+dQ5DEPrY3fybOCs82sjhIB6EaoS6+QtFh2dxq+j+dv4R
8gHHbai7V3Ym6LEkTXha/4GBe4m0NH5OEAbH16M+3CmiX56c3eMwKV7G/BSEZj2gSGqxkLma8J+s
kGl0AoyWp1QJx7sTqr+Tc1XqaeZ47tz4Rv6nNShgePK7mY/4MP+Eon37LfEH/m5E4EOZ/68+SGsK
4IMT+nSuCb4+ohWTUDHCkZUthjJGY/1MWPT+wFT6G444cfMiK3uXHw7nunWPwpQDdxIIvx55NKJm
zk3TvTJSpEGsYA4mdnR0HuZy5h1pluGybpsX9zic6rinMiieA+Amag54lZ9h7Ecwm/IKIETzg8kL
HgAq2j/e0RtIo0t4s2ypDCE+wSPGEaURF3NcbaV1CZebuLiWufHnzqGzd7PspTZkex4ZViaELj73
IuY9FfR7WR420eEqcKva+ki+d0UF5PqVMwEs4JrUuDkL/fo8TQlF69ojGbDTQTLsZ3UVObsmbOXf
RKkbzk65fWPM7JiAQHD/utV6vCugaHaz3dTM6oK7Xedvo6Qw4EaWF40da8HEwxYP6o8+aijiaODn
KL84rjEbdh6vd/YwuE+JypWQWbg7HgwnwGwkiTizDlgJViTPN9FsxlaKG+9wt+wgso704oBlhcJt
mQ5hJKAB/JcnJSOwAlO6UxaaI96DgRkg3ZipWf9SbqotqzHGYXJreZgUgMMhXKnfUAWT9x11APWL
odovU/7GPwOWxrlSn1EBpYAYjn7wRWYqixQJ6IFfoHuW9kOPBdrTckxG4N+IFrwniKEVGZve3zd2
/Pk8epsTbyVK5fk0qDY5vKP0yxXJEvTZRp5akHKo0fblM0YiISkWcjViRMoo4fAmp1alALl97dwy
ZJ6/edNC6ej3vFbKRVber3DbldsjrvXcNqNe06wxBVYlbZMWPDynkYihCfbzlYuArF64Cp6NnO01
sYdLjj8vBOhfNoU7/olB8PxJwHQabcoZ3L8MkmqjkaEDkrECObA6PRDUTn9yeJoXfW6Px1w/gJbn
loJ6oWL644L6R2puZBaeZckytfzFy3S6p20ZsVHkkQX7Kz4J6C8OkgextMg0GkwrMYNoIDJpoOcF
dTMZWwVHjW8b0zLuOs9f7odWMonR7SXi85qBtApi0x7OZ9NzPwqOCDtiXr2FqD2fjr5XaYrrhMRV
t5tv5spEcq/KGoIc7It3eqV3QKtpZAn7a2mgLgPDi7S3iT1kxt80o3p9bmBV5qB1kebIl/qEJusC
9ZVjxgl1bfPt2rfK07SswvciRidINNkclhZyf5T7sTnEiHPG4uqHBbRFavzwU5EbxYO4nJdrBXOM
/ZGK5NHYxIaAS2l/hfLKi6fcbYnD02UD+GE5zk8E9MHNKZHK7T/OoxDxi4suho9fXjLHXPZBMii/
ULnYy4GxorcHDofup5NlkKWXzyl4Z9dkgRtXNDH1n0q5+uftbZMhokwthDs8WhjMIMFYc65xK0A3
A4dqiUAljzqrdSJCIh+qwz127vJ7LcWgp3iWqpCDfAxIaR7vLmN/SmvAGUEExFUKrvoiv/vR/3bl
8oP9GdvDpnG1sS8RzPYuZJxxxw7ym+DpY8d9oadCpJ/g40TTLrK5+FIjALYa8vIbZCGCYDqNMyJo
GcxjW7GDS0ziz2UEOmd27lI8eUtDzV8p1M22Vfxs1QGBN3L0bIpBfs4Ogcoq+gAYK9n42I1/rPPv
1qzpUCdymGw3VVXbz0SahmCE3pyabO3pYttSHPNzYsY0yQPtdzKqaI6eMiYmdwHaqs2pP4YnvCr/
7nYLca6MroDVV6rUSGI2JLvs9IRBn7laOdjMLYERxifD27jb9DbuNE7AhPaheyccT3aSxxs5xcul
NJ/w0nUVWvOIDZ6O8XiQbOrUmexCEmgsn2kf0rXUdzoFvDfFcIKp74PSEnvuVAlFfoOB5pdkTr94
YJdjgBP2DYYREGYzLov3QULEPK0aL7ej31VLARdM07Zk0WclmZEMX7EQ7iKGsZ99/tIrsDIPpztG
zALfyQBlzGKaazW+5VlRyYqSZiSYZbydrMhqzftDqc429VhvnF2Pd4knSMP/1iY7PHNrekbN7HK5
JPk7isW455gOo+Tt6yfpK19vOnGGUA7nI1o6Rp96fv77qD/pAG7va6FDZM8W6ZFS8G5A3msbZWNx
XSumXjeMousYIGSk1xYDUrxVZuE0RCVPjj8HdZd7g5YSIrhoV4akA4mHbpEWC+4PVAZkAItrC83L
uwZJTdYtB8Yj4Aftzr7XblMuvxj1n1n6+EJnzHxlaQf3NX2N7KPjwHnUeQlQlxAVkkIl7hIu6pT9
Sxx2M8X+msTlATsIep+8r1Mb5/IdH9IenzuvieMp/Ta33yhBKHMPuaDVuSeL1DMspqAlGrTVU6QK
+Dfbm6OjuLWHW46v3Pwb47qd8nhE8Pn5QreULJuxRDnsmT5D3xQjYBt1QW+bfCWyGnFnfUXdwM4k
5ZsqbJ3a4ure0fWrzCMUDhQYu82OZKWvGqhlUCH6WdWBSzodYcqwzAotEvbM3ozPpnhePaSTj9tR
wZvttOSb8YBfVpL7+yoJ7chXE7ZPgExtpLA0bZuO7jJqbzw1eUKMMWAlPDJGcrjFlPE6EWrUmiCf
xgpsS7Ntr1RcsAt8VtWQhzH06d93emDocApiUV1lUjiznEAJZw6i02pB9S7rPu6qjHC/RYtXdpnE
be2Upq/CM3fysGD5xjDN84S1/jg1IZ82FWhjlKUVdLZ3rI10Kt63lkqRM8ScqfKhUZkoXsUrZ+wb
7teYlxj0QKG1TknjCg5BziQAhiJGIQOTDFdX18MTKtbE8CGvkQ0BJgRjpQXzMI/CehgEow5r63fW
4Lk+Elc+/7/zfsjgBl6egcpWNfqcuIOcNHE9NXH3i9xFZ9TwWfRt9LQVv5uw7YyJ1HQvd3EjP68p
lQBsboOBhmMo8tGq2mH8hF7HZ2dvMJRokX/6BDgeni5HTZFEqPgCN4eHKVlH5JxYsgmlCjjmpcpV
tl6OCis3IGx732QCB43me804Fpim2KzrUaD/MHv0MIQDqjUQd991eykBJnmPIDO+jGCYbUOemFnY
WbQwubsXStnFJxHTIsqqWmBkJm/pZBS81NJnLWHJ/JyUdcEWoQFc3KckmPGMnCKPQf9Z24R+WKpS
vM6Ok6f5qdiL2WJ3++worVex06gUHCZmS4VgqzY0E4ihspHC5m4pWIXSKoZzj+KmsJvRhBGnnW7W
ONhEG95rAgbG2aJ5G0DGMDkZc7MoaP46T0R+oo1M5XDTjc4W58d9Uw5WklQbhi4qV6zCGvw968oy
1+kb4SgrhJiCLeH3riSlVsvBH+ZQ6FCckgv4rXjVacOcBKfL28iIzbvBM+i+Si9U1FgsM3O5Xdlu
mozQ3CjaoYFXgxUrcL7BbsEx/rVJaySCmxf59TRjNBQhrRBW7etOFJU8TBmCEUUSaPxvD9q6TNtr
3cubvvRYC+fNkhcv9SJhh+eKlkDosOkZEC20QRs4LG8q4bSSlMde1OsC97P3DyMjKaxSt4GxJb2T
Cx6mRVO3DwyUuzrhc1R9nqenro7++aZmlHMzqPcPBeQbPrBippfxBU337b3A/CGpnBmBl7aBCKsX
b/Jw1NcPsqpSJge7mtCLN7ARxwIkMz2MvjsZgBj2xSV386zX4FIbDA83Qi62GGBrOsuvbQykaOy9
X9yZaFaenbW3KN33JHqMPwYib46vmdrSlyVnKEk/5pGXjjogp0oSiqTI8bULtExOKZ4OXVPJPPwj
n8b3D9drf97x6fNxbhkrzrgcAvfZQrtmCb/kgwI++llJQoKtGbYgkVd3GUhdDRo6pq6QlNlBAyog
jzB+LiS4vNuDGhxGRsjTXZEvPghgBf0MkbEZkrddLjEI3gEH/uiIeK2gbLqWwCEdgfOJlMJdibdB
GiabWxr2WOnO88DoVsVF6EoyVknnyOdqUlfwZPvWH7MdIAac4ZDGv5VtpPC3kVICODoawtBqwj3j
pfJoC/siZkfIDB0PocFFUP0X3jaZ/x4l2k3y69ovFb4EnzeG8Y2IWT3guMXaYjoke4M6zzZktAGp
mNY9YWmrEKM++0nGTsoZ8iZeUr1kjjupGVp+SXATvXu446Xy+maCV1q/5lvfebT/A3efgeqrwJWE
/h7CG2bdEIkFigtyTTkbnAhfiMi5pPgVR8KkDIGkw+NSQ9cXAq6aOfMn1syFYtYfLx61O8crnPSL
3NG4z/Y2i/NV7RmbOBhvODCW+oW8bJEk/8PbAX8gRJhyLfmpMZpzTElnfEfgXekTDHuobXb5ArsM
0S+2+PAWtkNX11rh51+yLx7KlXarss2EkLsOTeQiTuaB1k1zpZtpQBL6EZWFiKOSYba/6vqlSnT3
Yu6LjJDgDAf9D836Z+iDZ1NU+o3pffuhWBASnZlFhX14iqXkzpUDgZVmV+gmHAZ4JjnbLfavIyq9
KjxsHuxCo33zCT9lTzJIyi8whRLKx7b0AmJfH8C5N9KdvNslioGreyZ2H5OkmOMpEWmZHp2T1CN2
GrH7ormXIMogamSyDSO5cjHqDVMlm9e3LhBYftDFzd6CeAmx86FW4HxkFm+OIzzt+f3XM+4zhMp4
kjS/znJOGcmmbN1gj1sNqIEoPVivTIQkbViGkda0jfuFVPRxVVi5c9JP2S65luAfJaDL+prUj5FN
RDnmXC4K5Zb6JBS6bELAyYNjXy0H12rXGvwaAlF8/Y/3p/yRxYHC9i5rwLHbdWHKYlSxndK1INdo
WXYZ/zfw5yDUgZpKxQYrJPH6H27m+mLoCDZeCTDHati7giWP/1UNVVanH05LfAvk+TqOCXuQDciG
INZU8LZNyHlR7Aign0PbX4ms6Ame+XqEzd37gb2jUJHI5qVStYU+HRvOiB+1fXw+dcMEFd4LBn8C
ZgEUvd0YxWCLAdF3Zc/7MKzjbp+vSRpWCY+icyfmIZpQ9yhSV/UabVc+lWYUqaLht0aISOA8/jRX
akmfyxYgffVFrT3nlczOp6YEpVDfswY/Wdp1jQX6LWAnsauOdIv2SBC4JFMLy46zAgYlDb4RW8ND
MCcxI0FXkBrrZ1Bxa1mkVqtQU5Suh2iRe+xcHE4CYnv0xn5bGQSHcp5GjykZnIP0XkyyrR9ckJnq
xBW7hSvy/89KGlWolWQ4/Rm7ljWw/MyiT+Tq7a/C0VdqUfOn8ErhPnTzVE7E+khGyGaSyBDuITUb
m1yT3AlUPHp9uU8Jr/5fYqrKHG6Ug5qm/HdNcpszve6iSpP2hRHFtI3D9H51IESXyNp8MBQ9g67j
V5+Pc+PTVH1Kci8AWqCZGJWJd0761VYa87D4lTE9rhTgjvF4zlrAhUxaGONbtZ/E5U7/FCR3xlX9
Aah+BLSIZQRADHXpCKd+TNLUb7PNezIt1xiFU+mre4B+e5CNEBgcM6K9wLQlvrd9NPGHFUAmBcyu
3w1nbH39lTumHoU8z3HbTrVsLx3Ip4kc2XTdfejNq5KwQ4MKgqBPByfeParW2pqUh8GJ/JxUiMXb
tcytlk2vb8b2IXG/I41ueVuh4fY1P8jg2zcly35/fNmki4RLDy2PA+qYJfWmRXAmKmiQRvzh6VTv
xctU6z3rVn2Vf2WF9bjwWhBnVECah9ATGU2tyZFY51uNbiAqgbCXz1KU4C5TxBG70Z56O7H1kY6Q
TISIo1ptJP93H0I7zfRvH2OTLz71/3C04f62P8B6be9QCVkcz3V7EbQSzAngKu4UUgutkQqah8jb
qwwyQxE/lkRnIlqIaldSwjAndtmJSxk77dRJg7G26q+UXv9zr4w/5QaA8GQ9XghFenaujvd4We3Y
gktWKbXo1QShH9hBEk3ICI3XIAqGFa3GpC5hCSF45q4Ov8cMJCx9iUQCtCPSpcJOMWaw6Xqo8e5t
nR7FDC57XTu35UTkp/fRF+OGNq5rrfeiAk2ojEZHDyBX6NWL07ZL/VYaMOkLeOZ+XHtAGke5+qCN
OPP73Dch+QsN2kWOkk8D7PmVUljMcfSgQsFu7HCZ41pP2/IkpSviVQ1qxGfbLA/CUGo21KfJdqg6
cO1bdJxhRvdh08tIXW0RFFcSawohHUrwR2GCJ8TngiyJp5ui9L5bsysHlAYipjLcdCMYTS7ID5xw
TmRM3BF2cpCq7jpqj9+GLBJQug+yvJniyVvK54PfjO1UrZbydsS+ub6QQRMapc0EvD7/niL9ZmZ/
rkhmf4IDpujWuLCB5ToN3udCZQvanyEf0+b0SkHEv+m58jvjQr8Z+VJRSFuOZSvbPE0CUt1/t3yQ
r0KeNY5RnHDomNLZIJkhXTV3OqD+5AjKLg8bykYrPI2JGBnNHc1Kcj3P5wmzBGlDhhXTis72Xb9X
77PxdUbGCE3wJrM9DkVJLMIvZzvNIA1qKNv/qxxLqgbnjnTc+ZGjq8L51I2rA+XOKG9Vo9pOK/RU
9E8NFKMgkwnfmiaE5TSRtdRWTNop4ea+fK1am+ENP/8byYjoJowMl6LJrN4gs50ngrKalDKeuJw7
90br0nJFZ9UzKUqs6y0P0HmOtTfdEWek7TmeBwqBz/2+nr6G88Ux/pjAZXJfqkCEZCaIxdLnTPS+
6fMtBw+CUdSlKhpydgE9wyUqqRy05Cq63LHzsUBFKI9nFh/t0Lnlc5IW9gktKURI9iSGtJOAi2+t
sy+iYRN/AR1StVsrxVcoinV6yv9T6Z/hM0IE9L3DeSjoFi+2eP2EvW5ggfHKs2P6ukXPiytziN1f
AlGtVoxcV8g2WWcvjccYtfOWKbac/B5FyNWDCq8qpGLdioWruR83pOxd4m+Z7KcVnMSjMOJVTNBC
DifN9ruG+4nMjBIklfOZuAThs/bvE5uohD2QWxn8RJ1sjW4RUom1dN9+ETFHbK8Y3yJw5HGwtGq9
qvrSciwti7vCHOvdhZsDD+/ltw5uYEuMnbz6Z/G5n6SSj6qXT//xtuJxYtlcJx3T9RX+h0ZXT5HU
rnIl1eG72erwCf4eCEUwPlUlnEdWdvOMoMC5FxB0czsKj3aaq827qyTiRVn2i05BT71bHNDsqj/y
EDADZv2wUMhLIiCg3FCI0EN5qeZ8ipvcOk/G7TNXDsN170/zraAwaPxMJUMjTl2z7lMYdr98aENm
B4ndUw4qNSxPAw3IkT2Fj7tdysa+rmAunMqa7QisE/rgzdo5Gg4NjYPIbbcMBpNv5MH9BY0nuoja
fsDJ0AJv/6ZPmnJ+Ky+G/YBsJyIFrmtWNm6egFX8Ta7riP6WUpVuV1WjXh4cANqU6h24xi+D1Eyl
iGU3BL6/dhDFiKBZaMqJPeyLXkShjP5aiaBPiKtlpJzWpgWaD1Hbu2Ij+/6a62NvKGcjTsbwfFsU
33FrjEf83rUJFRQRwCXuoLkfDgt5mWOEWiD8mVOfffINReV3Pz11BVMyyBQjYF8yS+8Jg57yiOBj
Hk78FHBXYnqxAuF1T8mrRMnoRP46OVLa896342rDel08HH7nHcWJ24cq1W0bTC3tCwjZhWQU4pPg
hbWbP2xV2xSEXJGcWFdfLzgu6TbLK9l0dWpsN/H3ULeS3vlN/ojwJLQb0X6rc5uiYRtBV0byAsp2
+c5RCF4Rkg8lEN7Npz31P0Kx95SJ4VXBSZX0meWu1c81HfeAIJjxhFrMHXK6vyZL1P69S3dpeuYm
QGLFohqjIBroKolBRqAChTuZtFEr6OgRaie+SfIiwyTn7K+Jcb0txxSolefJvXEQ7rL0peZCTByR
jWWV9HAN6HEQq+uc9kC6D/CfY8Qt/hOyCIzCPpSzCKZ5xwOzyzDAiE9WWar5GpMkcCCA0uFEFqKD
Oj3AAFrhx6qGiSKA8FXcAyU9FPOaNpGmylFMmNEAEp9RXC7Dk+BXXUOkSHjaa0yMh0N43HNkNCb5
XUpnO6Cr1dOjqnic1ijVdv7ohOErrwLk098FIOcxM5KwZImSlh7xd4GRfHuwcApIkVoJ7EQkjSim
96YTEm0ZWbqQkxXHxy4BDAM0XIvTJl4eHaa2MEKg40RejJ1clhU5lW2Wd16eWGixu7Bi4pqXVwBg
ZVRUVkbJah3WMDxPGJnaYGT2now8wuyUprIzXuWngFH6T9jETPS4K/WrnYKQORi1rZ2TyqbDgQcU
LYpUQ42a10oN1FoQINKn66Uu9WSq7N6D8PkbwVyJKhQQ/LDz+OZOKUQa4MUw0297/m0MZ10XW2XT
X+mr+ZDo0nEVy4q4QuJrAhbG3xMWP8rizzV+MXfvpFmisVCZVYQDBmeQclWQuGrD5DtcVBaS6pYb
aBveWjPmg7Y2jegfnwCkbVE0IcYxScbNzOR2jA/DEVm2w6k3sCkDc8j+SRwZbkLt7lZXZbQiLSk9
R7WBZ49RZNNVOHXKa9nb2uzkWClb85QPkiVHQYoh+fYaUfdLbvIVShUDaD4DG0W4VY0jixs5B3CE
185kVFn+a+8NWasGAlwoHR2hBvI1QFPncgImAl2DPMZvbxBjZfgMhXzhLHNfncRe5KLR/eMzlVGv
JWGVeAHRJN01E1jSacXer9JshbGW9vrlhvLvmRTfBEbA13WYt+wRznmSaY3SRxrQ/Hbf5Xp5qIFe
wFWxoQWDVuKywZfiU7vuWm7UtI2zEhXgYtcyF031NgaFMeKgKOddNjB+SWKShRK70oP11f8hDSvE
SYtWsH7L53CCn8UtWhvEvlxviLGE2HZeuMbOTOefRMkF1ZwQyn6WyAldyWOMK9KD3bOiIQifUDiW
BrGh3ot++DQx5PuXQAw0y0S3hw/62hXGbBX17CkVBnEflXRZ0Of9LBZEXYsxeUAQbYsb51FXDOO6
CzoZyXABXY8tjyTVT4uChX1WLrlfdIwcZgBrGtK0824JYpujy/r1ywigTrOKMxqCP5+qENP2h65J
9PmC2bejVTT2ZgfX1bgGJgiBQiJ+rdXpPkTKaUeXbuwKUxGPQ5PQQKVfhK9JdOv88Ogibr9sw3qg
MQmTXok5sCW/OYuerE8NnXh1sBD9a8OR4WVtVspy8N5UQY3jhQGs7BztdTUwwxWYO3mA8IFH9wys
3ynXHgvuj9k+byRpjan2BIaFPKCd3Guy2qSeIAuuteAsH8wg4SOm+YjL287JbjYqIxb7iHakPtTQ
3MMVGLd+FNSEccC7PgcTKnYHSOByXiPXkOhFgVWEtYDPV5FN08nVOZ9oauUypUj743qf7gXYudxe
8ObeTlHNIiFcHXx05PAYs+PFvFzenAFssKdCg3zFgyeCa/QunlCiWMEofotxHfa4jOskM9ciZFbq
m+kwGz4b5rsFk6e3wMrchLZJDXrNfRgZ7WtVfHlPRdPNyVKwQiAPYPsVxyglWBKyhOP3qIsCc6hP
mJgW9oX0kI7AIfipogRl5bPk4h0VwDAGFh3VPaQjv4jCC1SS7K2OGkYJWTMEwdFLrH+LboO7Jpt/
PShA/6e1aDKjM8tgu5KlFLBR/U4DPJvLRk7sCuEMrh1IeqvXREdeFf1oQ4qrcmOrJhnRtbzPBlta
F1IcCT05XtFWo3WL5zg/J8qENKqNiN9Ia1uYQSR5x0zRKVTSGLJMMSDDIJlssx/D2zUOsm6b/J/G
CJWlmpXBUBDJn+tfxtiOasHsfrbgww0HtmP7RHJ2GOcpqDClKqx4hb+Zw7cChtDz5IecJCGAAktD
aBIOYpWPmRSlwXyXt3AI43ZlaPapPiLGwQmVlRkOKjsSpzrO8MzE7Gxl6ao7McUZXehisRYSkZqq
8Yrdx6xgo/g0JF17lqwJOON2ySJ7PVxkAeVCVpWXF8LeRfEEga6bq2xUAurNKY6yCfdZMkHWgc5N
DJ0QLeywX6J4zfl/qtkw4IOwSFP5fEjAzTSl+VJEvxoyaGQUG1KlO+gEF5mryMZthCLtA5L0kR5v
yxElPX7l9C/Gl70ocjU0ItnDdmN42s6PTiKGEUl1xuC0cApBpW5XzyVIm40GULPjVK0vAqfU/KjY
kODxD1vR7QpKMvnhbPdyiMLnXetTOrzTUnlRi/1B74mTPqiTNceZFkgyysrfxIibJCUx/s/z43UO
TBrnwDkw+q8mPjgpOlfX8wHSUwtR1mEWdN4uLPp4QfaoyggTwvh6LJlCbExOaao5pomh8BFE2K8c
CRhc7C1kUneUkUzLX84f1y7ij9wPTXGl6zSOYp/gH04oFaAMIp4KCvpmIQWlsNASDCZWljiUvxfO
WK9AucTDw1AGr1HcXHAB6CPLcGWj/g+kerwsMjvshbJzcitov/r/fNDKgG85C8hVCzPlGdVEgf89
UjmfGMNs2HpYzMUWWnXfsYvXaGHua1QivQUKabe+RHYqBqC/n42bzuUC1/a/zL4N5FH2+x2usJGn
t3Z2fSkiaE6YOnZzizW46fsIjxhFdXl4IE2TCwAM8OdXGuA7XnuLvKS9OY0PnBsklhdmaj5TBIaG
kzAlG+dubd96gWtItC3mIRfW5HW0xUgUTB4rcFg9l0oW3DWaUMuONMXkUFE4VusRPS/Uixq45/9c
XpqP50jGkR5ueCC/wnqhTQolPjx+b20VmnEBIirRtZDwWHxaYqXpOT4EF9zwI0ReSbuuOirjq2VR
b0BevCvgobu2sOfkbuNZpKES7HLH5TSE5zsRWb3WGeWU85+U2Stprsldo3X2zN+QOQXIgqnS4y+I
aNz7U40/tlnlDUA696RZewZTX/8eYOQI64FLrauTq6/pmjeMfbFeURJkJQgkzBLKEYkiVrXYcOtD
haBx3pEBH1vMVi3jXlomBKOwPcmSE6P8EHH/r8ManhV7loGDukCi4OM6FHeI3bQofpLgwgap+0ol
yF4t79sF3UcUtTcdIa8EuIyG4NX1qaCdi/wC49BpsqBW9hBLiucqt5tH/b3WTTEqWmrS7lIPdDyt
gaDr1wI975uT2D/nUIYizokWIB/PPHQTLwQv3gIkW99ohfvzpYdPWSpnnd51KGtXKk4/3x6cMFz2
peCS5+8PsHuQQnaEgIPdDAZ+q6ygA1WSCkizGZ1djRNEGq1DBOwnPK6JHg41nLqrbarFM9/WYHLJ
qb/F7IF9ZKU49J3t5jntkNywJo+a2O+uUBwxJdX5D7VjpPIOSK8HgR4Y8szuvaeQeFFx3FX3YD8Y
Vk8eDFn1z+piODh8UU7eBMlmyVj+/mEYk/HkKeXI9supEBhqFD1NGmTjtGDJbPAqhdqV/zlSTmRU
lVTvvQ+0vbnrEWG3VNcXOnXAK93FTTh7yLDCCcgJFGnkLOaBRsYldEM+EJ6hT9bWd+RWEvEMwKrb
Nia7hwoscO8QznkvgIlbdpPMlUCWAlLMruj0nB1FeKBA3nKHHRFEMZq0NkHidv/as+i2aP7iBA3l
D7UzCYo1TLf7x91Id7t+59beOn8hBMkARc1Pj6v+4ctlhyzy5MYPsPbE7so68dbWXrhNGaF7sjAm
nqUZ3W3GoPX5FLiSQdpCHdbBrRY2p3cIOWC8rTYH9iifbcob263IgfFJ8J7Hi/Yc/xI6QR/qN0Yl
6zsWe0J7dh9dEv989HeO8oBtRunf6WqeVLEJ/P0UTVMoqMsosgahD9Zs2/FtFVEg+6W6NKY5bDj5
te+Dmu7SqtbK+QDhIS4oC9WVn2hjW1jjaLssW3ZSYCV/CWoay/yFr0dj7M5jDcevpXzQ61VXnqsZ
/1RjeeOHs5W65uwtt8yOwu3mHXT8I/LnJfrGTLtWSHx+IPWLS1Xjd8Huu019DVzSYVhhfFGoAb02
oUmZIsRj12sWQkbwjLivoIWouuUzdjSerYVU49YT2P2m6ohH6Tc1rrbySbJ7mCkuYiYB5v74hGrB
w5dLmhlXHz9VjLc0MTnnj0K8ipWOiIJRY6bcI/tr6GyEtBZaYuIPY+JQG2zvB1nX9PAG+g5YY0wI
xIxmaPnq5hmTsn+8ZZrS228FENfTZhhunfecaEDWYEHAcTSrs5xUxdpvPS49vQaL0AufR4/30Hbq
4aRvvLjRBsWnOpI72Uo4Is8eqWHDJEIJ+SE0MMYt6aqMcIIl4BwaMYNr14o6cRh0259ZAJ1pl1LW
vgLsKeqWF/Wvq5gpVaEvCg0pGIh7Pi+vi8aVWx4R2GvWQowUqZJmwuxxchQB+6ne/4K098FHOGL8
/Xn2d4NLtUkEo/spvxU8l4epK7p+pYRIt7WDZGs+rvfvLF5EGpa/EHm/HmbxZZzNpJATx+NH5xFP
uhKCt5n9QgOBOD4LSjEPOSoHCAcfxyPbIe3lY0tyK9C+PDTLNjMgNjCmv17yBEGOpKC9cLn8uqrg
p5T1PHLPM+40b1it7JW3iD1AjHIiY5pqZC5NUwz6eX4SaUkcOEAglWD5xFok2jFYlJ7Uhw5JaVnr
IGkaUyN7lOk85s9eynbzkONcXHyvmztpv+oNk5tn78EMhSDwW11371gd4Q194aSMvHLLPDeM5cgc
KcPjRUHfjxhH5aI4zj9gzt8S10ULGFdHqLVcjSocWHdkBv9riydWokoO1qKmaPnXTAirgFdGgBlA
86xg53nQFQnSldnPKypgncbRTsFdcpz7JZhGcCLVC5uck68W50sdP2vCKh9QjDH+Ijh/MFFqT9y2
5FFHV3WTtJnEGHh9sKe9m+b7KbPbLZDhQYW9bKJ6pHHtkrlqr9TBrX9Us0VzD5lOc2izJnbdyeot
KqSH5UzNH5IzKEvQc0LRzuTNCoc+FDeraIo/vhxyaOzIA79AT8x3ibD5sqfvhtpDVbbIZ2o2YaGF
dMiA5L7jejfynVhlUl9kG41Nl2PrnXebwi2MM1HFFEAbJ8RzB/6hz7MMLvDkJO7FzZ5FzO1hTMK1
0nsYWqfDr6O3/9+Sc7A2vtfjQjG2KQS0C5KbKq+Un9zZGToIx+Vp0vsp1TbJRDmzI6DSJGwPLsJ1
t0Ou+jsCmlcYlNNIL8C33+B3QIBhru+lW7TphRT0NNt/RktpSLJy6cyLm2HlhAwtGoxhnwK2FeCj
Zi6629cYBOJQCHKWt8Hegx4/mjRarICmhDJaj4LcN+Vm4kiMRlT3moPh0DvJOCRNGznqEoS2LXN1
icN/L0qJkEOjEEDbC9J/6FCZurGLtE7dO6PptkLxQO3qp1+CXWAk0UBwHE/Kqz5qGqS18GjuHvC2
g7evz0B0YgMBX20tAizSS2g/EPXrYwtPPuPoWFWOSQG49K0BqM+skgU8LJnOUzsQdOE3w3VaSJa6
Ip/JpZiPDmNne8X6tbZG22XAm7H1DHp0j9xEfFTGe8i0HAeZrRxB9Cv8R45V+U8PO741Uty4GIJ0
Z2dTtKeZwMUHU2g2JvAvifsJ1GoSfDri00ZmXjMIS70QjbXBLLN+DvT1D0g4co+n7RWRznKe0QgD
BUTYh5Dnu79Jcb5ODVR7IlLOEoGQVHu7WbNxvXk132vGJoWd235GmPh+LPv4miSm31xkZAy171/2
uO/GDbBmSrgWIXBRzFWHD+eBG2FLSXty33EHvzRhKg4EH9kLeBWiKRMzutyt0VHDihAVsyBVua1R
zqdm86yJMbQpz1t38KwdyhGD8Xtw/zeidZSfls+OlFkEdGFZxRDVKMTilD4AY36u646O7yvt1arE
Sw5Jg7K/TaGh2D1Z83nquGc4yoiwCuGg2swQ/U9+S/Rn16kBrbODlEZI6f6Yink+jHkzDNYVqUwo
JU7+20iv08kx5wsr4Ya3YKelHOQnf9H+cTvFTt2ysEh63CHK6iJ/gFJnNXCJZjLuoQtrV0qYwxR0
CUJ9Rdd9FSzY2wChpRFgx8+MtNLincHOvj/Wp1pXxPMbqofVhEHFk+0wthuiuWcdzJsdMQuy0OGt
LjgS5nfA6n6BBfnNB3DcNTs/urQ1xI3lmebMXZUkhYnseSs18In6ytLTvKZ91aDH7t/ENTEVYTnA
TUJNEtd+Tw/psRIz4J61j2KcIKoO1BNXAZ8l/Ml9EyE5nMs19VLRjVL0Mf8cdJ+JCwxXgh4FRh3a
q2pherdhxJx6HcVsJlYKZPvrOl5U5BXKqfNq4rAzsGHTbAT0ImFTorI62IoQLrLG7vIb6tjwhm4Y
HFc2pkYTb4Kv7rdBCBAkDY5x6VNra3b7MLDsxh5SgX5LdXlgbAKriUmlWMvGJhkEYqXTNlPqTrfq
3+iBJkiUAu2KcRXmJI6MCLm04651g4xWufZj4v9riO7toByATViv2rAySis6OOtwZU9vewtMZ239
MVm9yjNxT2ho0L8idLHIqQye6x365r3BluAxhujUBml31LNKUwDpn8Ibkpoy1kdIon2WQzQzuxUn
T8bPiyeI27eZwh1ZrTUG92fgpiEMSwu+DmWm9KbVrVOJVut8tw4Xsw5mSfdHEirDzUhet0T4B2X/
vCE748mIIzIjRiCQQRe+lMPIBB5oty/EETke/oJ/bmHXS9jfjhbon3MXIawps0Fq5S800pRGkxRc
sQpHAYRYT20VCF/hwidZBDvx6YXG6DUxcPPEc3q09Lb78OZa+zw3Lvcmez1QJczzRSBoKjgKyqi7
tJBe3wrlZyJ952fFiG+gBKR7hP5cuVBNIIm4Are1b/f0lg7jboPgTa0YrK25oq2xNkSNJB1rA3ml
pwckyB+FMGeZbJt/57826hNKLLqY55IDPAUGl2+76gYc6nqkmmux2UVmsOdN0oKfueoVr7DHQoBG
7KoVDsrWFF6dfPGo9gOF3BgZ6b9Udi/B2JaaX1Qbv4Ue7nxrjb3TokcPaL/iQPKtZKtNJnndfppT
BLr9duxBPZXyIfxpFKfZA4yfSgo5UzuGh8lJqLa4zk+s5VAjIRBUXlVvIn7d24f4IcpeflxY6jcG
K9aNMJydnnoC1ipUmDWD0TBE+ZM+Yj3PIEAKyhgPhrGoJvW/5FYCDuMBT8j4P041aKPATOUXSoI5
mbWv5zVBRA5tAJEleld82a7SY8j6/sKnp/EXnoE1Pn6b8iAJRSpo+aKbqQREwiG3LnxsVLXDtb+x
/uqpD4VpStDwZaFGE71Du6SFas4WDRn9hPxtvYTJnQvmVq/Lv9Q1rePeFmlRY3SC6tRqqC74uhLf
hf8/mpgpogtfoVlHcroUyo03AyUK1nPmrmEHdbnf8HjD1ODLNKPhPYWDlrIIORNiyqB7oCkCt6Ih
6syv9DDZ2KScHFV1u95LKXuBDC9r5CzxiyDvxZBRUkMsec/vUPuSYLtviZEBqfUwDCFdK75+5e/c
KxIF0RREtDTpYzM4COfpj228I2mInc8tLrhaD+ISKPh1EYmlHk6SVIWqzJoL3C4xQmztDNfMJuNl
0VY2m3MeS4VPwyR5ZRYr6brKX2U05FN4HQZ6L5jjXQmwApyrb+N/3FixEssCFp8kbBszZcv6j2DV
dnwCS9MLv2V/i3qE9yWSR7CIUywj+qzHIZ9BBH2L4hpOPd+Pu9O/nrDBHVg4dlsax0gLrMP7S+Lr
iV/ktm4gUyHCDSx3xQRTyzRMLOe4mlyzKX/0pjkdOtTQuMnWtk8l/eTGVFRbJWDAzfi4UzJOAqdj
VR4aIIO+EqBx5G+eYm6txCjiwxc/2J/BQU0Reut5uuKI5HZDJdN037IdMw7EMMuqRhyMsajFoa8E
AWbIp2xG0D9s/8xtxT/jd9Mvp6kLF8GAC5mi8YOAj4aMgXCGsnuhpsqOPUwBKLZe+wC/41SrilEX
sXw6PCR+zZ8PqLaYpgWsZXXdfIREAgh7VJ+0Yxzxh91bxtStpLA8QcL4QTWbp6Pcr++RyU0dihEd
xRj8Vu9ps++oXkCgf4lHWWGX26vlIqNYwl72xRUTTS/sbhLqfnlX8KekcC5zXLOAxf/LgSV2AaWV
HKGv+Rnu6RKqUE5sJ+bA0hN9cFS56qQ+RbnVS34W19w3qzF2DsW3nIDGjkBdKkOCkOXhBoTsdUr2
8+nLvWnGbvow2P6nZEPOcsZJ01cwXUoM+2V/FU9CGaQXeEhUNpK7P57497U9toK5HzvmfOOmC0E+
/bh+Z3akSq+gF2J7GopUIZ1QRM6fpXNaYpqnNytLiIRkItoMWVi+Imt+rNGWjXWosP69lj2tgGiX
IWY6TfvGEXTJda7111rhHi6SL4BdM6U0ZW5J4RQ8G1Kb7d4TVOcZ++Q390MHlcpo1e0y+jNw7m3D
5Sdo4JBWpn+ueGoeADgwDblRQnVG+854xIpOgic3OVQdWvDuFa2BRu0pDfPGTlm4eDpmrJo5qk44
ax/Jr3V9q78ANnErDF5efuhqnCdrwq260pF9TwcI+l/hRbrNKb5nSVzi8KoDxUzgBZ9VnEYcN1x0
UGFVBqgf1DlYdrT3F9OFha6vUunafY1/i3aQBs2Cmw5XBPF9lrt4kPwGQngpmAAnpH+B7geojNf5
qZJB8FREbfcf1SOBLin5idtlhc9gF7UL9fiZIp4PQ1D4wchlnECmRReEPREj+xc4AeD4CQ2mTZJV
4VG3xM9opRZI+v7e/LMj11nIvDo0z/eKTBMhb0XMMmBsLLAyOmOa5hbKrQx+dAmYLDCnWV3Gq414
SzXDgTmN7Rap0OLqRExa291Oqih86EFXX4+M2O07o7yO7fo7VXW9E7k7qSKoHlFf/UTpUfMJqL0l
7UpTLdPqS3ObigFydqparRMAZilyg9rsO2iIYuNvqbl5FmrFC3z8AI9wRhfziYYth5qDTC7CW/+n
EzQ2deK9E6TDfu8dSPnpf5CVUzfdSdP36iydjEt03qaY018eyNLWkU3gpYw9BHVr5sLCGCsv+jG9
knj386H4h8Wk2nkuSWjlXWvmeLgBBccxi5EgzOYXucEfw28p/7S1gfXKt9rqNaHDkr32JjNfESvt
v8cinbOSve8u/kdO0/llzv8gG8XuJ4eV6RrdsLyKtUX31s1tYrIwVO9qdpa6QiSY7YtueW6uviwk
kH1tM7ApwaWlbRGnnEe8w3vETZN4GkW4X/yJzWYm9Em9yKP+Y03EZbiwNyQ2gRfKgJ0pNntqbfh5
Bb2wJJv8TCZXcEUmgjlhw5FU2lhYWCy6qceEuhXbqSvy5M/bDxey+iVRAyhDDNbCq3QanB5Fd/N9
OO4iwEHcasi9sW7PMq4SeIT01uB+Ui3aEneOOhtt9j9gwKl2k3Lsfi5j2gPSe63x+4w0E0ucGcUG
hHSMMhruvkYkeGUyw+WBEZcuosawsdL1YxKqvDAi1CXpwjHL2x6uVmAVA5VGdxnSjgUuwAuMJHNC
QquotUgSI4NH8SdVBBLNQlmrzdqFLCL1nwHIr250PSN4qRQDmADBTKHWd1za7Vi140v7qRXUZezc
A6pWnFIyA09CWbRISVCxjRYcP76Mfgs1GLjOK0P/QLIh8eujiI16GKnRPScxhE6mIylt5apPW5oz
3R53PUOubrqwJAAylmzWB0mJiDyJeLdvFtFmr8lOk/g2GMMpRBOH9E67WHSAhx2IApgGML5oRRh8
evPnvc3LkK4XoQkhxSj+IkJYN+/m3LLE2Ne4LQxZStL6NoTMty2Tx1I3bTcpvmHV3blYKc8i8Db5
0+8vDtzQQWtStvtZowv85QKndBNHvDs0yd5W0PeUYwWc20hbWGTE/9t7GQRKiOqMGiUcZHns2kah
R22fTGYXB9TQ4YPp/Oi/A3ynNzCqlpBNwSZil7+fqWah43nzqyR81g2snbvFuX9UrV4lP65G8MPH
aDj2HN9FFR8JjoPXj81s8l2eVyHink4HnAeLM0UHMhM87Sppwz7FDSuzrzOZQRs3XMpqnQ1WeUDe
Slian8rbICGAJstjoi3Cb6NWfIZX8m1QwzjiDa+sGqDPmWTLvn5dwlVe1KvdSvYvSfkcX6ynZ++2
T9xUFpbl0jkjmFuZEF0OhYd6rs3A0MdyAwlB4P+dJxJBk7DiBrEhincltv0bMeKxoY5+c9kFwim9
mUmd6FnX013mRMHJCMwetdgdbSZUaA0U7n8X+w8mbjYwa/VGWu1lUf5eTP1jJJKSmddXPrTblHzh
iV6VDPDau7uy4nMVZ3pgjXNEqXllmYvZyFyjwllpJxEjGxNlmqDX4WrGHtRXYARMTR/kao8rJa6D
nidwmRRUskK2HUmyu8IDthFy8s7GcOK2o0HEbtg4VpWgNemurGpTSiyu8YGtHFdHTH07f7Bq/rr7
0UQr7FjZK/FD+w9QElwd7vgvPUGU+qk2iHQA25OtbZ/CasJiU4/1KCUbZtOQVH5ZlhQnusB30DHM
YqdV0wFexvfHXdExh9uacNtT9XYGqTfRB/N+qIoa9g77gYIfYuudKL2kjgR1IZ2ZaKXpYkRyj+TC
eirbRYQZbZpGjNwB6GMHNnxtT4BkUUq1yd/HcfgmBSlhpnr1+GxUz5eOx+z42wTzjzsZBTr3n6ud
7y7kVrGPEIXq+8vvgYfINCi1b2WK66LNI3euBZ5dqiBj7cHdJWOxsfe7OPzzGPX4JOnW+F9eztv3
pW3ZN6gBZ/tXb83j8GZMHvyoy3a0The2Ua2E/Y2wsIvp5apFaWLgmPqLb4+3aY8+Y8loi1BQUrpS
TrAhUVExu4nLLL+3z6M8XF0rmhxm0eUiNOpc7HlwNcaZypqlqk27PnG6lTEcB2ShZVX6StEvZOPt
6A8SzG/vz/52CdebuOdU0j+yRpPe9ELqCbl1Z++Hqvxgw9x7BG3MuY8kb7BBglJboTuYIg7ti0DA
/q5Y0D/J9tvoxp7HFzz0e4k+C1H8uwS7DwtH3C9TO3PvC6DjnztIvLIxfOWGTbmrQh3c5pBj9SJl
mzA3MAhZP+7u8m2dv9/GKEP278EVExb61MXRa16naTS8mQLmepknt7DHtDlWh7NR230htMmiu/Y8
/HId8s2Fw/iGXlImkBCwWLcz5bHrKqfPYPWYj77izvXJz2v+uwumQR83WEbpj1cydX6ERUIM8sWo
YLlLO1zbnp8YE6Egcv88uEo6GL6Jl+OK6HH22Wzxz4h6e+XQ7pXVQ7N/6kSgFMVdgVip6nCT9AVp
2tejHu99YlCzPUuuMVNXBlR1aZqS/5z6f42yfzzufveeqIDNpuMFI0d3fgklKDRuLicBNBZV6nZC
Sq0r9Bvi4fMnX8JR+xn7mvyTcuFHgyHwBKsyiok9AzfWmsGbPhNy1ctnIsFhh6ON0HA2tK4Y9hBY
i5BCWo0g5RXXDDVc7NugDLYQ72EJw4y3zAdB7A4QPuMOi3/UMuFL4vDlmHaDcfGSV8uLVMp6sFmG
B0F955fqaZo5Ykn7Yg09S8QZvQOR481L24z99QAGhoQmJbL7AZttsfVC0tBS+XAovYaZ7/4TTL0c
0Ok5jwfZiR2tmnYPJdYBHUeJ/P1/eyF8CU32o+MkMRxfxVa26N+FqrqqSrhr3RfQxKE9BkFAZDcy
hwupQEtScdAKwdky5SJ31HCOFkDmNpx52xpTvHSgvjBV1F0lqppYgmVzrjc7LjJrhxMVVDLa6/pR
90uyh80L+dF0a0aFPqNu5bRtNXGEZOXKjOgUJsYPr/ot9hE9O0TRr24a8ynuRkNmM4S7SB90qlJd
5yCoN8qKk6s8t6t+dJgH4WHV7NNeYVpwM0GbY9j8QF0bidSkawmWnpIHAgv2qt5jyPw9UTcopgbI
SrG2Shybaoxc4fsqjJfmpXYdhvv3duNZ11y0M9yWkHaqLRohT62qc8PWzDNG7pjbkVoMV1FmLhsZ
oWugqNuyzWsvikvIoMHyziizOucqRxM+FquMHX2U7aPcaueXyuslG2Wd0GEr95IUiDcN82ujku7N
tWyOf5RZkwJyX6UtYxgmop3PAER47DdMdUc6LCzdtNZuZ+Qe4IXMvrjdUuUsgig8uycOvbBVC4p5
9x/fcUxDoxRNs8QdNDdWktcFuT0fBEHrLMoO311c41eIzFZLLBaU8pf23XC5gThpBZF1nlbZeviW
jn917sddFVto8FbqGYEcBYs8x4gh499+ccFFmdN67b+Yl/yQcJ0eMO4dg4u6XyoU8OgL6wx8ZqfD
//QlQEyedlMQBB4YaD92A8rY9YKtamlKSO01G6o7J/DR1gFElcivVXrwUIZ4rsbQnCY5SXvJ4ebP
iVDn9MrTGuZnTc722ckf5fBaeDf3lStD8ZL3hGZ9QXKog7iO5S30cL7f/LSzRklF0aFm9jFWYDj4
5Fov7ckwHosDR8XJb7kq3TvO9pTZjqomZDshtvhJ4chlZr7zlLwPjuuWyQU6EjpXi5uy4KPJ8OXm
4A1Wk/uDZSq7T6U4MdP/2Tzg8zFBMhblvHm705RnxbS9VYf6tADtFBn34rYMJgl4TOd5Axl0+t6u
vELkOltzosnYdIgsSRm4ocgKQ2DXknkS8rQN/xyqIAxVGu5OTbud1yUq7i1xh8geRcVTOGAxirHh
jqn30xc/lrF3iIlRHwBJJGu4NSuNxUCOP++CLRTW5AHFb4U8z0sq+kqdfTmATYfsN1P1a7SapX2f
VuK4p6ELFOyMm84Zd3O2kX4p6HYtvOLA8pB21RDnWAR+Wy8+xMB7xPN7L2bIO1SmrtF/OtFH+A9f
Gu6VfhxxcOUd9DJH5KTwlpXzG4+/kb+uQNzHtgrEGzMbZYD2tra70V8rwMJOef/xgdKjOioaPRQF
UcEuRskNVr6X1SeU7b47JuJxwD6ZsJ87D1Jj0hdFXnso6HRiUcMPGJ83YDc8Qbv2k3ZNDvxLNC2k
qEihi0xnuHAY+Qk3ztY9ba4xu5UHAyD+AV5sb9XYGpu4W0pIguuPFHJc6zy+KHP+4qmpHs+M0TIp
IikMBb/sK6d4wasYT0rXSoIMxxTZ+hr2+0QgMiuXOJZFQwhC4z7bnfS1Kt8icHTvO8HUwFhxqKZr
s/RZdW74ku8tGZw+MY6SW26wEqUJFTRBhoYJrjvAp3Ohu/XFSdWwMo/pqGWNSMF6bQwRMyhIGnD5
pIO8NzroF9qC/aMWRIZCOTAgKTKVBDng4ESlVLo2WrXGlGVtkVkADBvr3lbiHXOxWM7o626sHx8Z
cw0mEIbzUINST1tDMkWxtcNCPJNk4/hQdois/uh0xZKdwiymZyBYExZz4TT/sCTtowQpLP6PUjGs
JBQDziruZmi+ePXcf/PdKtiVrDFf+sS28NP7ofpJYl0ondcLVnhB62Etesi9sk1K9f8OJDKkrUsy
NgzXfTuBv8em4Sub/5yDeXj2VQgnVHJjhCJRuGzi6NlAL5A3QBzpnTwOHJSq/fPk7ZEJkTtJ90YG
h+j+HEXVQH77LziBEX7PXU2atI/iehnK35tCqOH1qHDGXqV1E47JOtM6MDemXfoVxceuf1eG872O
Ed9SM902lQlzndVj4LUKzb2Nn19QYz7fyoX0TFbhVkQcOUMYh58XQNqZOfPP0cRSjk5MGc6A/WMt
MMd/eezRY92KSm0UfntzKanhua8OqhRuNcYQ22j79zVMn+sh0oxvbVpUgLH9PMWRVo6Fu6E15TH1
WbrmQQhzEafTanXOOqOfkOidW1zKKW68Gy71POUHiKyZQxGZ3Mdz3mli25eC+rqKyImLyMkxmGwy
Ra3llWyOdolM80ypoJ5VJG24QzE/tR1+XjMENxdfyS45WRrqO/MgAtwr91aUD2WPMUSjQ8f7/Tww
jGzB6pvIMVhfnZsgtg4/DwF0Fl+NxdrOC0z/3Jku2buQ1vW8ij5UWAByGDPe+FCZFcQKTlu57A7J
5PpHSCiA0rjbLIeEmOFUyIpoBwN8yqJ1qAKgIDr4dLXlGfgelcV9PQqjkbF1r6Rp+B2x+vqYTvkp
mbg/lbVSKIZj107BQEI9JHGYQU17CdWKDIry0RlzKX2a9dwlrXyDLWqmPDG/9/y4/0rdoGXL1P5r
Ih8ythMc4PKVaMb0J1JIXf7nrrIR+cF+XbgbboAMke6r49HjsBLd9a2fJKrxB0e0RevUBvKcR+4q
pDLgZIj8Urg6OsuK4QIdrCorc89CcJrDq37B/bARHaNFIe+XBZr+Tz8KIa9pPHQQnY9pxqQy0Qqx
8NIlPdeEXlDQHWbwWiU4C8ez9aPXsSa1/84/3gaag4GmkwiRQeCLoTmLpXxPU0DCFrNAbEjbpkvF
zESO/lxrSfJTwfnAWMOaqZhrbOls/88SJZLHtQxlacQnodY07/OqZ28hxt8DZtd6snEFKX4FcyOi
BhZtbkobwTMFDgJtqCrd9w7HQPDFzAmTxJaUvsfThV80xg3ffztQtc0IUjP9XtRt+bx3icwGMMfd
VFGJZ/GqKN/BDXfLLdYNoCoAd2V08ZEepmjxjYr53VzAfs/Gg9OGQyrYuO7HK88LOw5dYbVSLIRR
GT29WKqfh17E2AVjVbRLaJ/gKONH2aHKuJfJG/3jDpL/FjhTRHIiaOc6YRvMWbyBVzH4wzgoHkAN
ZL4K7vg5Z20LDPiAb+oCOM2zz1qHqX9knLlMs+CbUc5vE1wdQD1o6ad63q60w/eZmQvttyCh9JJn
sqBbQAXIGQ8/C6hQQmWI7X6sOOVz67QSCrW8JoPU2XOAzaC4sfk1ToDr19ig9cIrgyH/fBeUgm52
hXeSynaNx98VlpIRFYRdIe7LDbiI7XsxtXi2su//ly1XaCyxuZe7zUr5DLRo9HZIODcGeRT58J9V
bh3njkSV92wcxtU0f9trvmMqxPR73siHzYVlBYmTNG3vSB0H4bvonPOQ1IuvDgVfgY7+X0HXBtsV
hiH5evVLLScZ7LxuCwkxVARjgT8ehHPuor9C6jNMSC1Szxdz+tQlfUUMeYzs13tRXqRxQEprevUA
CHcLd64hs2uQT/f3nyl7iU3lXn7jc/8gr6CS8ci555hR4ItMF9ClNaRszfTBIiCWHWzvLbAD14iM
F7DzSkHuRw4Pkp2Z7OyjHrWFAEL+Cmcwb57QTsGWV817xckCcXUTttHFxc1zY9wwnKG7rhnGR0vt
m+1AF3IO4bEVJX2mlbtHN51pjidi4Asq0ZfoPLF/F4M65EYhUTn6qldNMrMn6B2oCJxSpvnU2fKy
1Fmzm7x6WjsS0xlDSJYkKx7QSwUSAPHcxiKbv21Ik5lVKBM8oVfSzKYC90TTNjEpommBzxjxrfby
3zlEs9Na0MHKK1khgtw3N5/jgyRpV3LWIrT3CRyiOAt1NgEND52iGk9MNBS+/jyNOjP8/l/LYg4Y
PoXlBIa8EAYKFjRt6tuorBXuJ8vXO4PXlkAezf8ojzbrFwsfehbnZwNyEFElAShtVUtjASwRYDq0
MKKMYXbLbPqlk5p8I924e2eik9f0BvmdxHZldxOxBW8o0Bnhu1Ds+AMW2juFx+L/9Cz9uzXJv0R/
DuE69FjTYeG6cNjXzZSGj+b8vsTaKjaFlKjSH54am5ovB9c7k0jmSsrYeXY9rpHG3otbFXnXmtAD
iiBCuhT6l8dEvk3j7d26JfulmZ+si4GSV3BhoNGkt9WzBXwrwuKM9FmIhOO0CO6USI2XnGEE/rpF
XmHzI5AmpOmVitgkJ4G1s+juU6Sd7FxOjNL3d7vHn6CBsNrGMDA4NYnHIp6d5YSyUqHqwx37RlMa
3/wf8sCiHjWvauvB/xniNM10zo2SvLdeFVOKo+gRHHHiudoFjVGeSPhrOBOpt1ElY4NQRvHkuNYl
XJG9m/j+C+tLw6t7gUG6ouJ220i+EAzbX0lM6+noPVCKe2arLOYrPZg+WueMsSXusQteuSxP1G1l
5zqw2G4Hl0cGzAe7eF0Axw0XkGAGfM6EbgKSP0dbM7sQ0wsJ1wrIX62zKlvJYEHcl4kywlwQNm6D
91VduKjQnJhEL5+/z1aqw3L9lte2YgMzl0EO06uP3xL9bQPmFlIC2gp5PxjqudZl2k5IkKZevi95
jrePJc6Eh4AMJUw3BfjI/s/BKMt8gmh4YDQlFplafLOZyUxK6lbcK1Sz6nHTTIDdlPY0kh6LYfje
2nUbbdYGkF1LyyQEQbIb4N/KS3GuTdwgh8p5Kiu3V/qu+8QwEM1MPhPA5JScEFG7Tz5w1f/uH6sJ
ozOX8VXG49EyycW3IefPDBseC/nXGlKBJPF5f2lZXJD9oNXoops6vUUywUnQ9N6W5yNcTl31fuWw
URUgFZ4uJo1dz03fAI2X9cUT87iPNN+6zIiQ4fZDbnXevqGwkO0PlLfhHF96lUwfmVkmU3e19T0M
Z16DZn69xmqnOkshl9KD6U94xsSMYzOlrYGNv7QJzM2acDusRBRcXZ01MhLXH8s8FqMFg4fFLQ3a
ytTlXISZ0r2r29jo6WOgw7TvjnAy88hcVKvAjW0s4oJwPM3uiQJi5JssI5YuZFpIuiy3bhFSmG9D
CQ6CnIhHcYMYzXPi8gGwSWEYJhi0rfihTViHUa5y5znqbOSK4e3RLG0vXp7quOTNP6nc3zSHkaeM
2G9kbyZLRJwud6j14I5mkj5PLEDXFF60smmIoIvLXOwaYBX4YGz+yV+G11fdsIXBg6USkDvitQWr
dA4rHvJrNUAzW81JacBGIaXQVtcLD5QuqjnkcGF3WYvt83cHphO5KcqhRn1WKmd5tNA+DlwpoRSK
g7uaMcjg+TNGlOGyWNIUGZyzddVzM7Uls6U/3ug9xv08mgJd0UcgJEteDVpa0BMjlmRdkMYwA5iR
0qOTeFJX66ZOlQF766QGLFiUvh2ytR+h2JGhIRkTA5i32yD0h+eyARD/VH5gae8FADxxudwSV7dc
X/uRTTU9lQRwtb4E8pHkm79ktTAXOaeHqVX/PCB5KfOZ/cBI5EJ2IQ0EJfUueJJ0VpJY4MLiTOku
XCX8Nz/xJ/AAXDfy3XJaztV8QGhKCIlL0UCv+ugy9Ndt19Q9SvAJnElN4DBmTyx5i9SPkD3M6C9M
SOlPPGcBahE0kMJ2pGApXQE769yaKxtoWJBGFLCWV2xd5WcjLc8M0+CZioFSv/Hk2kSgKNBpdILD
qbyqwOOq6eOyIygsly9av6CZrz4cQUUFNSP1HDFCajOuP8jjCVhRoAJeiyZZFwobQLTB89Xik/+t
+YOz8O9iESDMgET6y/6x9Skpz9ION8M2xBizdUmVanoETbLeL7OYL12ZNNFDBI2v9jWM4PGpMWCB
HrREXlyAF/sYo8AF9rjRIdiROmDapXJkXZzpkoFfVH6UkD0awRgJR4n4ZmWgaNaPoZyOuZUWWH/E
ownMaZ9kc3vV1KXj5QX1k8Yv2I0y/6oO5YVm9fhj/ySU87W/AUuWbayWvZWSLWd/veQN9pF/LGlM
8oiaqxYmTH+E06NMJjTTGvSukhkx0a2YI+/taDoq5VmfslEsxvH31tNo4iFkp2xS+Xvf0BCvKhz+
KQvqlyvlAHJJScCAy7AJkr2tiMjXjCGev9g9fOdFQJu9/ETRkAPxbbqWN690Bru4UyzV3Bm8LJzS
Trn2uom7c1PJdVS0uVDDSv3RTIlx5Dh30X/yLUa24SqFkSLg99sVn0fS+kN4wx8xmRXI1TDa5HzM
RH4icRGDPkoIao4enjWB5DiaAgUQbvSecBFqmtk05JNeFSZQFNlitq/vPzRptSxeq2eaXs2lNK6V
k9MFC2t7D99jrJD73luH13LhyL9sp6SQVPIKq9YUDReRLWq+fMFHFDhtt04PulQXVFO47ZMaXrfc
3maJbU5L2pCGUQ0KhB/fe6biHubG8ECOlLRng9adFKf6+AAIWpQ8pwBCWivusbGkqJFRDqWFlxGq
UlaQBfK4IkBmH592zUIeMiKD1UWzamK9yanfW/gPb7llZxS0WNC/hshpBNnxJChPe1Qo/kQRlMAM
Y/EGaFF8j9/t6ZOMG10q7D8xYQI6Lem8lYPNs+zwwi+I2JbHJ67S/5HrtYciVejivNHUzdSXUk9q
u7HPiVYcGxTRwJkyQECmVkJRWK3qx4If5YqMij5V0e7NDgzOhh98ys3oWlsTlD+Td7lgNdI5skcs
TCqTqWe6ZjNXbu5wjbHvfPbwRhWuSVCee73oxbQM3E//69lH5rvI2JRNbbtSQIEsppPk5uhAQSqP
2XCRW5f/ZhRLJIWmhemZ+pUnt5ofxgteoYFEgudt+/7haw0Bh7SlNmsngjpEDtLVvC6wefeCpN8G
imJHWm4AiXtb7qHZE4tjIkA72NYMnMOMJrscRMlJJfuM5awGRSCs8UZzLsHuvkThYOS2O7m/Fexs
Mk7a5eh5lqXpsTHnthBeJ/y+PX0ojQpXqNejLBIYi6Bj4J4HmUKy+qAOKK5b4Wa6mtgllJVzddL7
5eV0lOgKnoVVYbLZV1e0nOaQ+sB9Ue95kaau7OhnRe7ooPHqAjs4NdxMP+5d8Ewn1y6CKrtjFr6F
o4FQnGuvE+M7T+UcYQsiQpG4zs16yNKuTTofE1xpqHIb2oizd3Pq9RYOTpvQVS8/ek3kMC1VMhn1
6qdZRZrdJ7ZWf0GySTk9p7H2zYtJ5ILAgsqZ6t1Jeru65qLoAm3SizMIolO24HLKxyXz+jL7wifT
QVFOl7wisXNqmpSSLGTFxRfJ+RNxym1CQMIq53ad6ZeagRox/DDw4YN/pIE263DXPg/XqOiOpA5v
2k0lNMdlXJKmXen/f4nT9z2/0DcsxGoiOq+tk0EdvSXt851fMhe49QnRA5THY/mrYdd7nuiu6arn
RONBrZV6ytw5XefB8oWqc0AmNgYxCGX7uWHMixgMH7DTfIG9bdfrdj+A0HfjFMxGfUQYz9Kv5YpJ
RUeE2c81OK3WCVCz5ikXF4Vnzm/9QIiJR9WpscCBOyoQincQh9vrKWQDR7yUZzwFUgoFeYvbG9UA
U01bKPUWKzghHmJWgK8uwD5iF0lw7aOjNkDLl7xSC9C6SQK9UD040w37o4CbhoMzw+LHw9lb+WWc
Y6kMw0UtVAgsYgW5MYWEJZ1LgrruIWS+EBQbxeAxT4fkk5K+HXldXFtK3ybf887Vuo/0okCjpmNg
4BHm74pzC9oElAsDM7oicm1owNAqS1aPanwFD1PiaPOcHtBdcrInoOvNWkE/NcgTx3VnhCHSgNDC
60H1w8mWItvMv5gA3dkDdVxmOaSKcPQ8bfLlo76f5t0A2IIMzw5KLQqlR3SFARK4qCWb5IOXhV5a
G7tpvpXxAc9pVchsc7SMFfsAbBY5Yb7nJy5mk0ZzKrTdbqjgZigl/tmGh28y9BlPcZr2rUT1OvoM
j0rMSsDNvbd0tnx2cudb+IptvrOSMG2I0M9X8kDqNK2sjxsXmwNEbdWDv1zqfDlHxq/73JoEsXC5
vs8R0r4w/hI5xL3/YJC+YIRiaOEcaSvntquRTgtUWB2C6JzuDZ0Dd/yOeo3N/0CL6PWo7dS1VuL+
AhRxnJH03v+VPbb3u8CCB/OwxUWpMEXxiFhVFOkIj7Py5hrciqH6GEqOgPGC4B9ITLkGDSFrdsDu
u8HRE8B4/l1YQWYb044BSpyxyRC5dTrJHnNqvRcU70khScxlKS5yV8iVMbH36c6Ltyk6pxQXr+0g
qrjIb0Id7nrtWJ2pj1U0VKmSTe7xeo1VDDbg1tno1P1SxI1SDod0sJyVuJfG/AisHcLJt2qJWNWI
9baQHC6xqga45tAF9a5yYxGQGARHjIMEry/PqiK6Y0X+Q8M63P+/THLAieLuwr+iADS9goKISfSW
BD01Ta+1nlfZFZc2pKrCcpcmmFjgD8rVAX2rALBoujuQ+Hdgzp2ztkTDOPg8pOdcC1Kw6h/kt+fZ
/NiD+kQem1VNJ3S85xOYG6Ca8OKmBmHZoqaUorQZGTgzWbkK0Gq3pmQvMI33HxBaK1KgmstZb0UO
NPePJC3GMdgVvjxXgfWf5RHX0Pb5INn4GIYRS5beNzXkcFOnJvDbQ0aMWUB3LnGl/Y2j5nixZh85
34t79eyRHplpGwHhA9QxDf/Sj9z8UWtRZIul4pgG35h7YqTk8tvU6fGb+YKnByhph1/3N6eJYFuH
YYTiASComNhBpNTdSTmsMyTOUbb7tlGGzH0JyaxLv4xrn8YgvGU05V30sytw/AUxCzPVeIfJzfiF
/i978yLZsmK4Ag4iwvYnb0OJNG7X6GorhDajIGY4EBxpdQAw1/D9CfuDA/Z7xvm6pzBNmcbROfN8
TPmcwaN9GHXQMwNXRsWHz+MmPTzKb+0AiVnzN2H0ZS8OsPi2cOjxEgMcYKDqiKgKdGbCi6L4X4WK
Df5FBgFotXTiEMCQgda2DM5uYsNWhxbG23MJY/WjfnEJyouWUrsMbeCibe+H5bpIYtMzHGA+bpyN
GgNJdPu6YR7eXJpm8V1JoL2Mbs87qgQ7sIkRlt3sfoOP8a3hw3Pe4f9BQapiXvJGlVn4a/yALA3P
oVpLiWc6QjFfeKxixAMlJ0RCr3qRagjkFwO1R9pgdM0bMMFevaWc7m5hGM63k6YLSNmEM2aOQtff
Q4CcVn6vZhn6dptxW1nglhlT5mk35Dwoi6mLPxYshKRusi6oToEBoirM0rhtjUdezGVkAPzghGNX
vSxM232Jlxq+BCM+qs3YBJ6AN6WyI6OM3md6dvLymTybAH4WqxoKA/eiT+4vbunRy/Rk+abdB51i
+zwwI1OENf2pL91v0hVSws2/yOxcChCEBA1oU4PSmrOSrb4BZ0s6Oabo7h4Y7HQlVeMD/14BWdFC
wagnLVqT/81gCc0myk5PwhPV0OeRLVjRGCRFhRgtISdntHN42Lkd+hwYyPH3AZSm2yZtGoJr1P9h
luhO9kcWPy/a3q59M3HztYFD7eNrSpZ74aUXiXRmovcsH4GTBJ3V1JlylnZNMn0hdAoKPI+//yrN
aYJJlsDAdYBzQ9/j3n/GImoQS1X7pMkdFTykdWblIgmVyo8KFklOQpP42hM1mLwrxIF8ZbQTJIhB
rUokP0aC1PHPk4niCQwbWlocxjLSBEm59lLwMLk7pTW/4LHQ9bUaMsGeTuKc75BF/BNfCEgm4/z1
QmrGKVD2pK4DErs9EsavRkDrtSou5irukv6sLEk2XlH3knXQA2+5YjZgi4pNplN0EVmlcv2bKkGq
9NBMgn87VmJz7O5RixjpLeDHg8KUth5PmYMCFuqeVEyQipcLf6paxZUpRf/DZFUdYBN8BWkpRy4f
YHJfjiiSMHP+AqEDZp4T4hsQFJX8D5lln0ro/xQeZu6Mrp4AwwEtoIw4cl8d25c8+frsLcLR9tbe
TQF+9q+zXcjxx6ROTkLvDTIjFWpR5YWMVU16lEm8mBSrfMOYeuFViw3Ug6zoDkrEayICHrVK0yWm
wlllcWA6FTAJpoZnbBKWfXrmkdxNHxZhdIuZKZ0ZRTAnX9q655mGFiFn/PJfQqZhywsHjhW3vdhf
+0MSJtFMU5Dhuk2vArRkGZle0sNNjyeFkvWVUqSH7wGJlrqlELXTzGqXzFOneUWd0E6SVwN2aEM6
FvJCEfRKsoprya6HFrrqZcCbpwlUbKv9T/K1bfAx9KJwzBawBwk+VYN3cgIbkl1H1xIWLkvdupR1
jXgyIFyZpViSPQfYkiQRT8QfEVLCvnBcyqrsE5hUSt+YOyWzPvUPvPwhNxKnagoyXckOTwnQNxEx
dEZM3WcW+PGNvoEXYPQPVEazfZLFEFNhJKtiCPan3OwpKkmDvod8R8WHtjbudWWZZe94RAUf7qqT
yDkfREys22zt+gc7mKeoLkSGyhiWlBBXtJHOb5+bKd9Fr5V+jMWwGjnYI7kRUmoIEjnw40HAXjnE
TkJUiMBSC6tfYN8KvyqY/do4JNi0nJnqBvAS6ZIA6CTBxRKMCes6DtKaTI/0fiGzevBTgxNsIAVx
1EGho1zkm/tNtLnPNbZdumRYnUI8YFiCvGhczaid5Etm1feUzDK4TFu1dEG/gcsBudoz90sRjizV
niKfT2AwHH/ZZ0BpeMnz6j2/Ojk1Ks1tHJeSYDUYPFaYHV0IQWb/nQcOfn4fjOIJnzzAH3QRhCiD
dgYnH/VEZjp411OKAmaft2iDETvx/nrSni7eAzz8nFsRHaWUEWh2SVNxRlc83p8Q0KVZQUpfMY8W
+wlyHD3++BoxmYzmpDuU5SdYmchQIt21Uyaw3hJlzw26QRP/xPD0iVOCPMgBQoIUJHGgqC2F1Jy3
p2iE9AgMZA+uQV3YcApQXpiBHQzeHXnz/U7S2FiqB0dW16Cf0VN5ukVHn8eOMH2enGAdVQwDWIlD
RZ4a27m4NxK9M6ATC4OMTlGJaJk+EgyHuhTMNNmQpCaAVLpWzyL470yyaZIc1nWFWp+YlZCkMFyD
LLS+5BzpgazzQ+Z4H/BcUWjudsRqqiT+OlHb77/1M7+ryjR0YWwQ5MgEhqCeqPxhrC6QC9c/PmhS
9catcWDAOQcbQHY98q/gq8gLLMYNl0B0y2DGCfINXR3tWwT66XL+nMWeqSaMfHzw0q6dGaI1g4KP
JXt2S9FkOSCYVSYObVMGoYwqN04Sft5pVuizOPds70iqJy7kQS3f1ZiNfni+y/BCfUUyjDafjb4h
ulppB7ffuPNZb01EhzQkRTB8K2sUbpXA3EjLGc0L3gAVls3uNuaR5G2c/3vaV5XHEn3aUzqroeAd
6Yr+Be8XEeqM1QPXKyWPvQ2pVCDwOBHSBgfZTxbA2G784ymLo3yFqbBzZqifnl1yc90HtWEW7Rd+
37bnC8DsRtZ5ckYC28JCtG4ttSZzY7ftNwoiE1ZqqAvxJ9ebviYNwI6C6H0Y2bX2XAc4EPEyevkQ
A2KUYiSnrxL54ivHWM8bxsS/Adt91FDyieCoW7Jr8VsGnQcsHCb56dbEf9YDT5sa7ViLwt9sAqeJ
6zDhOHg94gO32WPSwmmbqPZpkTxDmwbUGv+yjRRHvwA9sJ7+AoM1yfvrTKdQTU7xwwsL6qO4sJn0
vgs2N4+pHVvF4zCnz7AC9xc/eYcpHeBmrzvbug7zsRrFFz7tG46CmMmQCu8z/GTsu7D5kGiTUwdk
aUuHn41xzWA/1yRehToFgPbdEV+SSX2YGvTBs2cm7ihrVLRxZ4v9rKPEMDj++aS5UBET5xXHPLDf
BpIw8DvtMO7ZvGH+XSzgkL0XzgmY4WLVGhGzYPbjIKARZoO/UEbQs5tXd6uLviKiSFzcVZowx9nY
vfRA4GVxSmLvKmZ1BmKaEGgprVdJADEX6qwAw024lRV8Ic/47dtF24Fmuo2Mj3wA/gK/u8TAqHKB
PuchUixddzF7m9XIb6sRrZHidP033ya4jssLgDUDvfB2p9eIf1hQyvdP976APH70EisCVAGyOokQ
Gq6bYWASNmkR9FPKzBeL7VXswsOI/pn3ZAV5Dpi9oYbDTXBnKWrnA/jjiQ8kAY6brVOqlE127hlY
Rwm/CbYPXpYFMW6u5YuINPsfK5Ldt8kG5WdTEUeFm75XMMh96uqFlx3iimDnYiq0nkmnWhro9bhy
V0Jryl96HZV8NKCxGD91oolZUv7a1aX0XNBaCsL+3koCDXXOGA3Hy3qWfoBNkHOTrjS2cpTph3a7
f6Pz/tWKJDfJsJXT0nSuCmFVWfItmtOHLROAJKVG2tw8XpskvU5sssdbB+Zsni0I9Vy0u6dLldj0
tIGTlQzjbnahZ8owUmnyn+xBulWLf3LnqOb5HbjUlVqS/BqoMS34C2wHK8ySXOu7tGWiiJwLWhuV
LYVuWxoQMqprmiFRkmbissk5o+y+1X4gzYn2blXOWMG7PaWYVMMmCYDrTPeGG2T+JR1DxxNG3+DA
wMRtO3T5rs4LtVhd9AZGH7N7ToJoOI6GOf8alhmsOwnJUYMHYkd1opT08lPWi+8Mqd3Vh43Sa7AN
H/+zivMUMm7US8iGduU7aIN1sJ//ztudht5pFVye14DEUJUNdmYr53+O49IyEFKFi8zEvAYNbiPf
ECSA86Xxre9L4037+0CO0GdIKpBGcvF44/PbH/UfeREc+kOzJFAyLpd/K06oZizhJSRrKhVhJzwE
2lh7XTVwUXLblnmGqCHcyR4EfB2DNXb96hOTQ3XiLb29ZI46r4odZm4enrqxsIvSbvonWGrSb2RR
ApzFrfC1Q+w7170kWkFRUQG2/VnLIp036hpeZOlSFiA7xPMTgw9R5JCJgs0N0XQSCU1vEeM5+ttk
yqojCF0eFzHuyH0EPWFh/ipxlBGUj1DdZR0MXh57Cr0bOiItkwnI28kE7mgVmaYEzfhFheMHvJxD
56K6Jully3sbJ3NVr9b4NNeoiEUOxKymoloF50+mtU72jMRGEg6DGVtbD3aAsbx7iaioC+PsWyty
a4krepBThhriQ+ecsd187zoyLHiDWfGu3sHZYIM3T365oQD1LOm9NH2jGUYkSGLib1RUK8Xh+IY6
wdSqwFgBQ55uQaRbRmzeO1ovkRFP5i4n9Q60CDGYYU3jh74u008wj20Bs3EQef9DUrBWZeHQAPVK
w1X4yYcr3+7CEsJG7YbHekC2TUWxS5F/y1CT5OE8/RHC7LOvFVUeVvITBRi9Zl3vG6YsQetsuKQF
MlmgXoF3bQvpRm3x+B9561bxn2QqcuP/ikOVMqaUuSGsQ/G4E5FBqFMBk4EuJ+P7Wlr1rDt3G/Bu
ZhT5bYDY9kodtmWiU2pD8+TkX6zzDFDnLa1aY8y/aPhUic7HXXrkVpXSOsYUtZuKiJ5yBV/RHuC9
HqAVYFS02i7l/qiqGM2BufZk6a69lUzFFS7R/x2YvA3LEMWKZnDo9d6dg+xba1ODqXgJn/mDblAS
DY8FNT+C5pVHSEmehpsfAWr1dx3px7r1Emg2mSC/xmlyxrR8HDFzM/O5beJTjR28GRjRRRk2oQ8u
5sYRx7UdVPTcS2yNCpzP7Cw6in/Lrwbrv5wnzq+w9sqnT9qUc/APvyI86G54ZjKDXMHscJ2Mb1ht
6P0nVSj2ImfK6JkAt8bIXYBbbueCBVjPNc8QnSB83/cXUTQp9KfOEC2eSXKj3EYiejdaIWXp+h9P
NjvDFhBeY1W5ks/9pIweVFe0mSoaeOHrMhwKazRobTk2DhvXt0gyRPHrcAy7zMXLVNd3/HKfYyIw
D5bt6ROX//8U92Wyfbq5ygba844psaV0Xnu/KA/LvXm5s+ip/BsS+em0LCtVJyXDkgCJBEKjevXx
OQp96iM+9HdEaYfO5t6uAd61B/bGn3sLrTe02getoSjIQX0UuQ3qzzRwKAexLuUBt+Txx7uKZbOj
54BxnrFBIWxTG8+3sZDoCwNh2BoABcAzoAd8smZPR2P+H8ZLXVDyzQLuWllBVCstHBMmcYt0a2wW
EaJuFXkG2oCDzIwO3fSeR/Eky6Xzko66d9wYyTcTaMyovo+HN60t9XKj1QOr3W2on3jk+oLabgJH
PsP4niphgrKPU1J6gQ81w3afYUaMmJgGEhjCtxVx6rrWsNNhQ22/83keUh2ZHmoXqFTwv1Qyc4Fv
/khTHylDm1SW/qZ38KATlegegWJQGSrPd2wwNskKJrH2fJKWh7M2MqMvUW81f5sI7Si3RGQzja5f
buEZ2y+yitoyEZjQipV0hJh7d9qxSnfH7UkLbjrY3tqdX4QC8GUlqrOUxAnE6G4ADrjhFPL840Qv
Bux7Hqje01Vj3UYwIrHajg+wBby8jRG3mM+cWS7NuhVlhDBG2oVVG+5JOsjLq5e2f8+u71OjclpR
sQ9CHl4lapBCw0jcvNIn6LwH+ldbOoJeqrNlFGlVXTnzAs9iepwrOAMWHk+/ceddAG2/2B+pAFRR
F8P+kHL9GpOm5U995X1c8Ygu8sjsyHh4IQdl7JqrmvFDxdaVdDpG5ksXs7IZcwt4dSxPbB4niM4i
jvOdLUpKuOdZCy/Duy2KIyHOLDD6MOsPMAedWXJxGrX/qEaif5hR3KCvHHebBRgQ86AeIufUdMf8
k4Y6xQklvWw+VwffYqWi2f+x8LwiXkWXHPV7daH2yq+m6P1RhMsw7UVF9/QM1U7dIh3W0WfhMvrr
E8E9BpvJknmqFZlRHf0U137An4juOA/pERMVnFBkf7612s4v+nBz7ejbBsdyqFKmj+J+cOu2hM13
LoCNd+eHMindeETBBgCPzYmymEtLuY2v07mI+IVd/y5OedNgJLzyhWliJ3JPBfVTp7FL5ia36Vqe
XqzJvx0VD8aBoD9fhdhJIeUwBKTPWtvoB0s1TEre686+9y/0AjR7nhXD+kd8Ds3k6F6qli4eoY03
TI07Mez/a82RPaROOCfdhSOiBHw17sXh3tgOHIqxGKG3/mu1ycSN19eKjQjcJPEQ6YxL4PIenAda
5LhpjlMEuedRIKwIiXfxkKdQWt+Z0Y0abgbyd1jqKdLtIEiAW7os5tJJbxVVsO8OlanX/acDCYs4
TvCCAc6t/VpJPf7tYFpeigA9hD2pw15L14QnSUtkLm1bW2xBfwHjuDH3LZ88pdJeDv3C1FYm/cj1
cN8Q3kdm5CDr/ze8zudgux+vWxINuiiq6ni7b/oI8jd7A7e8a/HfH/6wMRmuR/Fh1tPlTJXpb3jc
83vqFrXyYVktnwmdete+wS4a8NboFTCfse69/nWWAvBYFVPBoMBk5d3TKRYJB4oeluM0SV+tlaNj
KdaV2YJxDMcobC9c8eBWsZXrHfzQIasbK49XrlQEJdp712qtcO/oX0ghk9N88M64uiKiLaYT7qhG
UwDpUAlCFeyDq7QKLUKyMsJG+XWEld7ugztMmdhZR9KbTGeYdPkUWpLIG47xP7cboHLJiEKkR4qz
f433+J7YD28k+TtmfhZf/3NfCL3+7uDLGCeLOzGA+m/5nnm7zNI7rXCS6NGW2l6n8DNvp9uL5CvQ
vX5QpfljcyDH9HzxaesSaTCAUnC70S65iLmRMK9XoePPPAiVl9rTzmL7/+bBf+hOm1W5+5zWg0pw
atFkAAVhrVgKB5HTPw/uARilL6vN4Gjvvm8ydV91WlB4ut4r58X+b5qA1Nz5dBGNJI8n7de35VTC
Z4pnxriNVu683dtwOqQwlSuSJ9xgV+yu5fd4Lhe4MwJwamSIhuog+sejAITy2OY+Df7geI4w9Sqx
T69ozzx460A1l0FytP5MToQXO4EbZHmH/i7l5ubw8jHgkGQUCLaxZlK84XjUd+hPikpjwLbC+DJw
Ypy1JjEedZs9voGQFYck7UZUf7aX3GSlsYGwgoWCVzIajUVDDHiR8RUX9XQH7um21L469YDojKlV
JPak6/yOtkD0ELIOrqH99T/ERHcqXrK9t4XigvZqS4Tml1e3hYzefIFEgk55YLXOYbEA7PzRu6lf
961qiGXwvOoldL5PLL+3hVl9Uegqwcq6ge9r2pn04JodSxXtSl89qfYfBd6FRsiLVT8JcDB+S9xV
p93S9N+0H04r30wHD5vi5u7aNTM3YY0u08iiRFtnjfTPi/+xiuEwI9Ux4T/Yj34K1MoSwH2RigqQ
GDIWdWsJvtJZHBba9dnmFENxywkcqSKvJ6TouWA7WzY7yZ89XSw+rCBONUk9r6hD6yzAi3GlhmZM
57PVrv1g4ozwky1Zd4vyYPs5xeiSHpmJ5pI4ePFcYdKXvg1D2wvF79QyEkV56u5fxktTbXvLLFer
ae72Xs7AIbGx6a49ggUY9rCBHu0Fqid962ERV9r2akhxKuRbLfqVCfl7GbnbS3sV1cFAaKuPviva
O+mOP3np1DA6odHdLyGOv0uLd+MiHp6OFs0rjNBHh9v9ANSP6+uUxeyO+/g2W6LVVA0ZyS4qGCkp
vVVPleELLSW0MwbUsAbkC2OBxUvGG12viuTfTuhTbxFU5AyGMRqZBUIXuuKS0PBF5jKq+lrpH2D4
RiZce7Y9tB4n6xe63h8JCRHPn2ec/oTQjPyXFIpVuETmVuxQz5QHSKjChWjG92YX87e3rT6VHN31
498wMtIUT2Y1X0tqSkuAyEt5SopNvzZIjD1nXTxZrdSfFHPcSoxB6TCg0e75AnxJ1Vr0RinhDA5j
IssCcJY2rfDN+az2W0Nl1Ttv1M/zB2toHz65YMM/ScDG/OrDuzXCg3l/efB4njdr6XTWGu2h0pFM
L21JK5KdsGErbyh8pEBCHda2N53SDZHu8FNLtjlcSFcaPNuyD2mLzAd7gNDYSM/lm/1M/USHvSNN
7tBZTFi86XYlMNqdyfqjbOfHo8yKsD8f6Sgd0HotLeNPT8CtHdEPvQRN/t5QDEoJjW0GBvy7johB
4hftp0e4iyjQ3bVx0nc0HkNoLGgokqVBrlfcxeTfBiOoLsFF96d38nUFP3/GXrykNEMIpwY2n5TZ
PVbHL+xOiWadVbCjpGzvYLzvsbaZWHv5sM0sYVYCAv1dB7nZmtDr6Y8HpI/zBalR1ORmfiHH5is+
zVTxTe5JTBX87vg48pzUrYXvOhWnoN1YoQWi9qLGt7aFI2u6JH817lgM0fH+jQtWqJZMzFMCThXC
KTk/64lAQd8gO7lFwVxnJnin5tyUgtsoeIcwut0Nxb2d+wHGC2rn/G7J6nE0cOxCc1W4wFyIy0or
Uft6UT1RyqekB7mRM7EDZpUMdWPMkTdIU/XT1ll9KPzA+8gqXQ5M4keLQARlPAz2RrIBOzByZ/Wj
dBVQb3maBGRgDNsfNL544i/YMcRHbul2QgY5GXPEtVNqdt3zz8t5nCPT25dyYYWrjMsvH6hUYsLW
MX9FQE2ojU2/3hkYgi6/yT/9cL/S1IlEGhz/UGUcYFw4gQRZtSLYiSsfxNnZPDc48AL11+rABIGp
1yFuuLT1BTPb23OKqlIAyGklnts9aOuTuxmnUGNVr2HxH/cxFsdEeUaKAtXubmxE6jc+6JtP+x44
zmJl6Z4mbkAd6kolNEawQOTeLHqMlJw9wK0cmRiVmDqHN44DtlvDRX8DM/bCtBMooEM27FnDDwik
jTxOkatZvc3BNTTIyQ8TGABeUsSUo4+MAMZ2fa86Yd78jmh+X4xoCEX/QZhcTfyBShx+zD2TYyS9
45Vv5wQvGyNVB/YdbNFUw3yWno6e9fzCC4v9lTZoo0Tz7VR7WY8XoksPcjwo+BwiApy//k35mW7v
C8rcUnAvQXLMgq+qF5sABTygdvdOyWgLbbYSl+hqS8s4kFEDly2Wlxt8NYZaHsloTQcBwDccjEfG
akDyCN+Q1UJqk3/ewn0Y/D2sg+y6hYmDGkPhBXmLcaBatkV5r0CkeWCJyxFKvcbFuPS/IlnJ2UJJ
HJvKcObOXKNsD4UraTZa4jJsGYVn6TwcMLPYaQhdGtHRb+HOa11ix0+Uy42X1IAHe+qrnORpx2nA
2/M5qf7UdD4UJhMTzFuFhjeZgmCpLd/C2jsbMSFeCpLJrtv6xyXmOQGjbZhlMU0TUN65Y9uqC0BO
AOvKWLZp/dw00ngih0ug2MWo83NM1v5Vl1LuJFUqxYc0CW1xaCsugVfaHE/+AhZ0BY6PIV0S0oaL
MraNVS/mmWIzhvHXMtRdehqwalWBPu93w3RWwksWm6I072gRCSlpD8j/GxFv0yZhCDCN13TXO8aL
KAB37XqTLPOx9gLh7SihOJVV5vc0DGQmO4ZLZe4tTcTYFcAbYIR85tqxND4oAHmEEkLTKj66kHQe
nRvjHh/fJs1Lb6AqvKWgY3RK45or3eThDwnG9CljgW3dL0mebiUaSXTEA6hkngcA/w3Raofl0SdV
vqUTwUkpdeFDp1G5aeuD0O8N4YJD6AByYnkf4hnxJu1WNDdkj4+Snpn9dEzQ4g0PfwjJ2gw55ioN
RLUswtOUt5ZKX21m9f7K8U1Ii8owdeOah4k7ksCyfhVzTSS2I0i47ko9caAhclRd6nJ7VUuvfEM5
3vRxiwfkq9ChfUpo+e+LMa4orcGbjBifzEpsKBy7dqAE5vvzd0gXyot9873++fdImZ2DZWAlKe+T
A84jCTUe8ZQH9k9RK+lcp6OHjcufw5ss+hpEz+aCHEKJ36SAf+6VIoYStDbIphotIhvLNBiJPWzY
VIe6zQZNoQDrztp2kESG/9g+NF3wZf1K5aBdroGKLVXI1cZOWxL7eYCRcZ/1aIgFTCWdVexqybRo
6E/PAdd7+ltRgMwbgsFz3sVW6MoJ5bFzwhWMnfimzTR+N+M3wyTQQg09XPS92jHjqGwYef9B+Ugy
y79LKMH74RaG7CGSIIdiChPu4QWfgRncQgTtfshFCKfpeOFVRUXRU/99AFFsL5fzF4ostUsMKX/j
DttGeYFmSIXvxjvUNFiFNesRFXpcuM6AaFlXZeUdq743kxgrd1J2kINHnhQyEE39GXjhZKDQBdIH
PEzyUL8aA8cAH8RX2a372gmSXWHFo/MVdNC5ryjhI/aClxOCBs6ErB+z/X0afGFO8IAS+jePaGpv
7SyU6aP4jjCR0crGHsSzquvboZpkFmPfBlz0u1VbuowKV+D6xuKQIywhrUDfYdVzJ0+4VIiVXjBf
TUlud6LlYmn7qsG1Ij9EK4/7LDHc6k3l2WiggQvoNxKcjBjno9aQG/0RfAzHTHCviuHGVkq9qN3h
z14+UCOPPB5eFhm8aectLCUC1D/tjaUneRF3JTix485qLueKUfvc7Vn3qqFGEVVnEFZPjRnoTVXL
u9ruswMic13Mi882Pcc3aeRyzdd7bWgtl3RliOJ8qOE05u1Tk85MSdo+GnGbYJVpSYUVf6g1nrR8
45xNRZjPIYbbsxdNjrrgZzhLrujJIc7nTiDNxA8Sc74o0hXoF3TwCi8xGx/BlMmk4oPyBvOOrZ07
om5chU8bKOgVh0DGX9m/0PAbhrgLvDmxziFtji/IZi9wdQrymkIOsIy7pm4+kfoowxuvDdgAN6TM
Gd/SkmKXkfKZIuhu5iGfqvcpUrFLfXtdQNkv4617ztzUS/E4u5kg8pc8WVUCt1o0Ab7Em2kbp+oo
c1XGp+ySCwB6RupJ/WiLikLBwWRnUSOpRhQLCUs44yNJLQCNKyFhPnE3gxcz69rtgLEU+ghaTS5A
c55czSBB6573tl9AqrRCPjx3pmWLEz4+rB6ItkH8ahyIPNWZL/4Tk9/jILwSwbMCa1A3nPIUNrQA
D1lcdYhvfMiazEOXCYs8kpAvNbq7TV7W6sH40eTu0IpUMWpXdLXEn8s+rjdfyMrpEKescp6Cnu+U
IhMG7GkLEU6+5mAc3b+Hhkdd/pcKp7ILTszUcTsiJjNkSb5EzJuu5hboGSGOJT3PaENQDlf8DYqn
RNeRBNasHPcagl0PwC1xIWv+GQ55JiA5LEjqru121CP/edgJPoXBjof23OIq1692GE2++xtACiRz
n06d6H45BZdDn1mrImmXl74xuZsNv45RIiScLJ6EqBsTE8MmnvRIjpqPx7w+4kcx1vwfuQYaTnL5
c+HA6DRiqs4O1vZZgZFNn+gdP3nuEr3zFXL5714mvSHbbhNTpROjOM4abvOldD337dfPtM4h7EeE
mYXjlPHnLViiLHMS7ii8LAOCGml00eBqSAX720u+wf1Sz7GkAmy0mwu3f8vRX2M2mPbiFRuhnc+c
oYXU0vtb30j7nKENfc51aHK7Ze3JE4jpxPiYC2ufuXEx4jKaZG9k+VUy2H+ZlEtzONNEEcUGl13e
FRSJGSryhSpm7W158VEeIWoeVVtvt9nXBWziOWgVZo/7PVFibCH36mLJy2qWn+r+qGeF6cYgBGi0
uzB7hCxWyB5ZJdooBbuO5EdSVtNQVIh6ozFPIu6Cquz2l2n0eGLh+yhOOC7ccBEaGj39WPCmXhGq
pi8zRQ33W6lN16YHPi+hMSNIYkJWQksNYcmsxj1AkMkSro1BEStYcNR+ALJZHJqvsRPMX6pUxfRf
8II12zLz+fPkc3djqBUGuo83an/ttogVbZ77RWC4+z8moxL1xPJDPVgwDtwRpxRvHdC2dy5R6MiK
ANlKxM50ijzAzd//2ilT0p6NvguEcAiIdF3lH9g4x4T+IYyGghjwJqdyO99r8xqN4aObzxX8Dc5v
wxded15ZNJFmqBw0+tlrUnEDWs2HuI271gs1ku5u9XflDSJ7I/oYI9+YeeQAJ6YPwxv/Sdy1hY/8
8bkYGKkQagrt/syBHioPbH7Dow3FQSGo6YMvPhwTuNOALV9uPzpv/+KEXuo4ZqjZD4u2KeEUnOJY
EC6/sBItZEFP2/I+f+ydNfYcur9ICGg8I+iUHBOfTjZ6f0e7SeNLz7HTDpQgrglTjQtmMzeZkDOu
bmw5WJcB4uymI5vId8KwCHOythdHoJbuiLBoL61yLm1t55EF8RaJMG4UUf/UMXGuhHlHbuwRy+Yz
rCkR4ol0vgxaaY3eVAyXDhiiIKzAbbayqqzioHip8u0BXCpGt54ZPt6UY6rRznxidulXZZglhOoB
nSZ0l+EFln507LcHV/SfhLG7eeBhDvYFgUiS5AGK9R3rYUESpZnJjjNdco9elHbG7R3j+EPHnNdJ
k63fZKXU73CDkSL9rCWP3/rv0q4okgrma5rRrR/+/ENJqqJAP3au5rDI2blQpZSGgsvHnxVGMr1x
y3UN/OH8t1t5E5xnANVWQ0iIm5c5oCv7cDb//1345PfWQShvM7FBwQk8TWPhLWK9kBw077xiu/YR
2BJEpPDTiUSnnrzvz0n0eyyZT4YeUbfxdixpcqMY4Txwa8XqfKucI93FLrWKo7X25QgZga8/FKjs
EKJ3arL/hj116ahh5EU81UmBhOvn8fa4ucNP+N55oQU90IHVNuKhuct3R5Xc70LScJ17X7oeXr5O
M0ZFrXJZDe5zyx/ujfWjY0nK2SQvgDT7QmMFppbEFIoEGhGGST3S+8gCqPf3FKNDdR4q7IwAiwOd
B/tXOQNNmHwa9muhlbQBw1w+n9Bjg2lhf0mUOZVj9GQ4djaSqqTy49ZsNLoxHg1gSWWfr6YXVq/w
ba+CXPiZOMgXANh0pY3PsN0PS2KCP1J6sN/RWWEObHrM3d8KNJuL/V3VmNu9exZTNo+cMlDIMtan
cQO1jsxT6ETTpum/S3Ft7dGxGup0FMji5yNlRA0gD32Tl16IjjsAbghGusyiHEAHaD+IpkH81geH
FEObjgq618Zu4WdYyt3I0s8wcWUe6KhltfG4TWWoByuOzWWmOHgox9KsAQMgm7ii0r02xfv9OiWP
ehGS8K5wCLYfHCCik6+H7zrdDyYTjcwD/hBZcHkA33Gr2cmTYCQuMFxq4FAkyvprTLZsVsbnLFXP
UHInzLnxeIpyX5mglWJv3pKW9uUS87NSYOFYvXsOpOgLbwxO2nYRDY9YnnSKsLviU7SgDMGYd9eI
qgEOQ3/7aj7PNW9D/zM8UJEsMV3AuU4Nbp8HZbfCGEo+KmyFpBkyfL4RUkESEVUp/3bw2uuCr2TH
KuZK3Y8kMOssIp3X/RJ7g+V0aQL7J8LEOwcC+9I43AA9ZpuXhsD422AEpplXi5eb6T8x9qnGn2J1
3FSaIPtddmu00HU9xFwy/do5uYhaRH1t4z+0eImkTdwh9y9i/M55qHZy5fqDItiRHJu1N7XprUyX
ON1iE42DM/97T9Q8k/PUaQ/Ef7dbO1DwGxa7yfGk7Q1Z0TBsi2PbfxovgewwJsFsykD6yKLd+b1l
H0HF7IHeFvabPv8lFAAgBCXrT0ULP9vgVifk526+zNdzNCjzXBsUVO2otPOUcRiOSgX/WYjXMSPk
LOUVUxD5R3gPF0KcEAFK4emon2c/p+VfIquCfXTJFJs44eHWVIpwBgCFNHbhk3Al//wtDnifwya/
LMKMZl7xLTqigYucyS3hJxfhtszIOYQctw/ZkoTLIPruuGZdRLo5HU4A6nk4m3+dGRat7n4Q0HdF
WnBWA8Bn6tMigOmCKDOxyzIHLpnAk4GqkGOOP5JPwEybMDZ9dZaS+ahzau1YcElRM8sqbiCNYwk9
9a9V9WCldzjnWrg3x7ME5KJwmg6uEcmhcvuvenHCRv6Y/MHntuqHeEZIVLxuNu/iiS7dWov9qmRX
Fbk8ifCiTxwKLFOtTtVFaQQbJb4BtvLSJieB2KFucU/IPcCwJ4HhcLiQbvnroOPeb2FCJ/I7e/0C
BmPcopSSC9UdK3tQO4cMiyTmM4TMKzOEV/pgkWenR+/9BK4lqp9Dkjllu+PZ18fU9jS8sUicCkNa
77mzP8FQ3P3/lttSbvR8gN9h0L77OPC3FzMZPuIDIc3+scrfUKeQ37xdi3e6JNQuhgGpEKgcrKDc
rFKBGI0S2hPNWjZuzZ8skYLeHoivjiJOHP227ndv0UF7/E/5Z6hLmDir6X0SprJCAFK79ZJISckT
ndUlK2pt+59VVhjoMStcMVM1WbwKQwS7DgP170bWYm31RYN3hhSSZQjW2/J8Bk0uxVu+7gew3NwS
zI4vALEttNgRjnIY83RFRrOZSjrN1/5MNyy6FaXHMV7P0wGrN54SeZ3DRhrag9RIuuyaghr5Rygh
Xi20oTuFLoZI1FwS0Sy0obVAnsq2TGljtS1+YaYhLhRC3M8vKxGaS+aILIjx92o2ZGARzE8Lmhq6
UhF8cW4pi3tlIRH6ezCU8v3YzdcOiy8R2GTVeREgAU3e0GuJ+LuLbbvX8v+85Wf1yrz1JeMCchQu
mo1IfiuvB/9CcyfVGMuN0ygdlKp0+JBEzr/nJ06p50zaxkuDT2fNPmnAe7ucCL6ttzHabkVXRR7y
S+/6aDcOeyAJWELUFclXXAWCNMjKHedpj6dZK18C7oqRRzitwCql43ZeAKvf+JCFvCUYOoACVjGX
mbpf3uSCg1IPYX9lzLITgLjlV8D401IQ2KBn/21coyzifJbNarzbVTfU06UPybRC0NJ1S0vbiaRW
+kVzypLwglmcogQdCGbKbN3imBcKRzxjdbAshZqrigPeCFISJzhgH7Sphpo5mHxRSLsJzaj+hQRc
KCjXCWVtsgFc1ZIp6V9C0jsIP/kC0jOTZzGOsuw67+shdTteeDbLchPSwZZLc8ENQPvSRKCcW0Hi
h86mkwfHnRCLdKVBIbIEv4Yx8d4FNEi4LXpekXNuYZ2GSpXwZTZXb9xVyW3qhDtGQdp+0mgLSr/g
OplVXcvWJPaZ1+YzYXmcgVIIuS2hRHCxJjYyBsnnTa3DIzBD0K6y0DceS+e9GpUAmcnQXkFbFLay
Fmd7vja7glCDaEJXJh8jZU67FrPYm0uuA8TiCD/140B0nacqyYbtXpPhFGto59DopvktEi3ufF2T
DoF3J0nQefreVxTBnMfuOQjzDXS47Pqd86k5oZw+JtC1Ij8A5IKezqwQI8JIf+e+0MQzWfrLBoEv
Yp8QFHSauSEOIxOGRG2I9bw8Ft8QqdCDUFUlKATVso2Cr6ILPQA4BrvBXz1m8Qi+zDlyGYYJ7Z7A
c8RRyWgqjXupC3bF1RmtK2FtOZMTsgdaYrI6WKAP+nQVzt8FoTycBYeB9SLUngKWxmrDF62GayPU
d5O/PRruSyg9vNXvG0WSCN96OvXQg+ZKYsjgHT2zOWmVJzvXkFjHAAe1jHwmhDCTHTS2PWeiX/AP
euGczYXSK/+a/GFLnXphqjwdsmQASDwwDHByiEaLG5eHJ8oKwUFMcC8SOYqzTc3ogRagJASg9iRg
3WiA26biZMELVRuia1M8aYX5Fl01a3874fEJff4pu1xDf7FeuF3GDh+AfoOZYcE7sjGuIo3KF1qi
YWeFqnv2n6+WXRmA4Hkf3g5FKY4JwpbciaElCGw8fcIcuYuUdbWq2o4wPdn+j0tJOQullN8JHXuz
Xd3GhZdX5JOH4rIIavaIJFD+r8vuNfwMQMvXGTq6K/GVT3Rc/EvgzDYKBNGCJv0HrGb8cxRLOBGx
9l+GlSzahXAiWNP0jn7mX1Rg8TmYgp3NKEtGnDQ5vT6ykaW5kgqKX1vE6BZ1gJtdOKDXS3kRVhsO
qCsRxH8H+IELFlpZ8zTOjLuJwarkgdjUkHmiQEbdjovOKmlH1JmEQf92Bba7yXdc0zy4Ogo0i2Md
b711xU4IEThkBbCgfvYdTc4MXk5AcKVYac8+0wdc5hIVJYmbnRWjHbVoghGIq2T/68kWbeKeMhHp
pST05XAWyuEI16slFkdu4HtFp0AQgOMgJkcxz61S0WwxCUq5hYJbdBBAbJSsgyv7ynb8isJHyU6S
BzPLPHhJNsKts7++8KGSN2tWn5C2PkJDef1yMdS6QJpuHgMaF8xa0qvTI8u6VW1UFE2AeNpymr50
cz+RZSW2R9a38p7nMYwunE4AJjMipJ2K51WFFaT+mrHpyqZ/HnGYCt7tyjzndbB3pCtsHlgpuyeK
l2ZYrmiXyKqNnOIjNw5oFADpWkDxr5CA471yg7aoVD1wT8LR71X++Q3WR51s+a84xa+qJ/60bnZH
J43AyYGhlxVVFwu0sIHvKKafin56gheyJUb0vDeLTGFAXRr3aiclCWd5txL2bszhKj5QN6/e1i6c
pzfvpAkljsFGYn/V2SJnytHp9FRPUT52B0TGco+5v1XJDllqKyic6IvUTiYvT8yHLXCu0WkXf60S
E5C9ZVWF7Rl2b9dcUev1e/b8tVNQtkHV20I3XJ84AWpFZozAVZGJ/sCM2mAFYq6cHGufxEOlefed
T2pgqGPe2ROgcmTAPtPB+r/HQ7Cb3qnF81GivzJSxvLUdF1eY88Su7QrShvwcILc2PeT5uRNAwPf
1chtURAFvlghkOKFhbUMkvxr2LaAcbYTpNt6AfWZwewvhdCFXq+hU0ZVThIisqnhSQYTifajPrkL
Zv+wpELHwx7tJfoIFyBWKsazFunEXGxphU0unMSIKU/74U0VcO8gld3nMjVRQsWolOA5uXHOUjr4
VTVCFn8cxQn5d8jD3Dyp6UMS0KTkt0qoW7DhnEZcWJ1lLQzrbVwzcVynv6/1QQLXUXWJsHaTKdPU
Qwq/LV2vqpQWnI+mFi8v2ZApYUlDh+3SSpmMuF/eXRV3vsx3ZbcY+p5wFSOyvVAhlblhGqwmZ7oT
Uk45bMEvMk9yqaqzGRWJ2Yrkr8QOEQGuaa0ATD20a2pKPQaLGUDFwe+k+9IRfGscFkpxUMBhIRtn
bhg0cadKuDMHnHQ7SsjztHETK3Y8GFCMUeXI3nDiZaPm5J1RERK9m+WWV4Fha75wy5WaBS6yeTUc
ksBn7FlUT0nEI9/2d7pqbNp5Vvw/hAbmOaqdZjxYRI3wrGPl+UDjxwFljTHsKlIeAadL9AZxMD9w
3iA35kR/02T4OuRAcXHNdukL/s2IMewOF9gEV+jqnjZWYITLLSRV267/gxtVP6T7q8zRs/i8SXzD
PSQPKu8imNxbZRH/9y346O4iTH685P8SysC1dVgBsz2R88YVipPpAs+UkT1PbYmkAV2sPddpJehg
uKXL7Gm6bawEKn7gzF9FnU22oyly8oKviUlhijCo3Fg01EMbBc8mKcG8MPCvOx0iLOLYYK9kac2l
0Fy1WX7v8VV+BrR7dAi4RGk2k0E/NTQpxlMa6quYiVz+vio1dvya8sQCnxvXxJaKW+JwBzyYbK6J
0L8gAfBOhwCRa86opihkjcqd8382l3xB9dER1EEXQ/I8oWLiGx7nImipMUY2ZrfrXcc6yGUgqdPR
BkWsEJnH79O5OIRzOx8HdBv/w98OLz0jPds8+sy4v2rRkZ6ZrA6fzjOzOJmVXnd4PTNM+YlXE16k
pMcqzgI/NfI4qTMR/eq06XJOoev5+mkswqX4kuWH/lbznAymlxL+kBerVneKKmMEYDIVXU/2xfPD
Q/kAQrq9qbECsn7QKsqL0GPOuCvHe/Y1uW0U5n/pPysLfAJ7jK+0WSQL4KVOQj4sEnI9mIYrb2Qd
tcQ7i0mY/Aj0gt2cKqq1+Jh/+yrGVxx3r/eJXuaiw1EbLwISzveFd9R8W2ETAOJr9dZTLUXfvAzL
/yjyQ3MPcHSMrg9kp2KtRM9hqhfo2gxHsXJIOnAl845Zb2p4qMnYOAKLIAMPQfdYggz7l3ijFk8t
kMR7qufaK8JC2URo4IrAURmicnMno6knyRKxRW9FGSVDtx0EocVIqRNNNgTdMl+CeJr+jfXg4iCR
d435Fn659CoH89tFlOubMnN26L6iwNZJASyOTvJ8vCqWBtb+0sttOy/6hn+gNnSoLFHhBA+p6MOq
0tt909yb4wpc2fPdphmoq5txwXAF9qv8j204fuL1WaiF7bW+uKot4yVp7D/fKxDm2eSSBiMfNDH5
DdyjLMRvAretlJW5DIExJfmEn2X+u1Qk1l1jSKUSs1XW1DiUNRo/6A6IbXjGz1F5k7CbeUISN5v3
QWRUYSFsulMBNJeE7O30sY5LcKUAWAp+9wKRoPaoODHxrJ0YyD8eO5pkQjV4KPqAAeFkTa/1SPgB
Kj3fZfyolgwS7n7O0QXHwBnPMiJANs17G2fq6GcRCCzRZsclq01b/Ome6atDj/KWgxregKPwdAY9
HGD79ZFZPRqUXRBG5W88AvwEkOJdCSa0zrXJ4qJtWzomLjp/B1zJFk4B88nP+AeYeAfW9xpV7F5M
dDu9f/z0pfB+zb/7uzDn9TAlyWcqKvxk2WWJIabpFyb1gHK1FAj0OskMIeOsZNuuDeNotO1Oy7Be
9eJTyuPL/VKMwkv1EvPOi+TaWCQhjF+ftLxvSdU6QoqZqK7Z/ecrOuosXWiG8zUZueKI6aQb7VSG
a906BIjX2Ophw8RBIPi1ZeypTNBU49iPkEFzPjRZTNZqOjllQ8/+N5cIP0gCybG1IGjIMMFzdNkk
Kqc//yHt1rUr28f2Rty0PVGf2TCd9/wXK4h3dvbJjeJ/rjrNA+bL7E9WSbZu78mvfS+4foiQRWBD
PhoY/b/PxtEu4XY8+cvoGUTLKtVYazNE5VElw4gChpazkGvf0WAbdDX5GUfpAX38Po7SGIohMLIU
umIEsJH+lQkotUGkeFvcx/lD19cbHVeI9v4T/jimK+1xoBBJg4h7XCf5+6y38B2UbILoaPh/N4RE
1IBggEIYjAxRsXuuSzCdNGpt7gRJF+5AdH/dFQKzWqNZRZM1730ng4aTK6FZOzTIKBOYPoMMGrpD
4xrmyM+rWwOYq4hDPGAuxSkztWoMqIY8dLZdv9L9o6EZNNMRlSKEBEFoHiJreikHCZuNOEFGfzfN
2cCFK0YqI7d77ajIwdRt8rEyKsfg6zy+soB4ws66Uxd6NMOfc++lp7s64eo/ayHfj9QjNbcU3PLB
W7TUDUQyp32BPPW/h5N2ScSqK2hKPSKvY3c4g2lseIrS8CWjOKEZM/9mA5I4AaYV74w4LawpdH9P
Z+lZqE1K43sPZqci/RrmhfSVBOE43VI7/jnam2YsJthp0VvAMVM2AyTCh9x3JLo6MNG4OFR+GkYa
qTt2Jk8M+cd9KyUnjeCQAEeP1OIMbc3IOLg+MBFMJ7tpwg+IK614Rr6Jy2kFQ4Sw59+5FYL55wTx
WSoTSXfYAflBl7HdGqMAyGeCGdjwHPqj8PYtGHC4J3PKSyOVE8jrbH13MtrM+h2M4GdZp5oIQ0vW
YCax95tOefSmEbr3mtm/YTrXgwfA5kfh9ldmMtDzslLLoOK0aAh9oni/8Se+sDysQTUp4vGhttTh
cdyL0dj4U20IQ7bFfaHdfD4MLEXjbnus2xPKeOT1mpb7zteWSTPejJkZd4mgumWXNzbdrY1kxl4B
X0b/YdwBkJSb4/cbnStkPW2FsB+g2XwDkN+R9VDmL9T9gOkwPi5em1bVKfUAfNu03IdO55tCO+bW
BV8aX6hXxlsg4NDB6QofjlM2cyItAf96lihIlgjsv9C9AMMY1qydzOy+e16zJrYihT20dIegK+0d
jJ5FjK9cE+IgqnBsC678sgTPm40ydhkWLZs1KcPiw8MlbgDtZqg99dBumkfCqV66rky07yNOmYQx
eQcUtm9TbbdzL72VzPKeJT4YM2wLmDfzc4DEcLP3uxxx5qIv7hfiKIFV6Ftqd8c83ky9+Xv14lf+
xSJmUHKx1RDOMR6YIY9lMy8BjmtBQj+ob4cd/N4kIL59oK08A90Xf6By5jE6O4XvroOFXn2aEdQW
kriNggTIhWPFeNreZygeJ47N8kSRV8XHZLf74yXEoWPcy6a9zl6PJC0+V3B+5zohZs+2KN3jn5oA
Mzpfpoy/1cvXo03uH+91lNqC/Z/aRwisfWM9pltZZ7Gj3ChMWileCIfSW6X7LjreUO3UhoGdHUyE
WH5BvUQeeKxxppQo0OhWxz1wqMa+Qs7kHttjl6HFghVjrNWIIf3V1MQM6OFRgBpCb4SfOd4sO0Yb
4RcBaqGxJeAil9panvdZDqf9z8iib+mwFoFd+XfuvVKKtd6fTsuZAWU4zk24xGsqqEt7Y8JrXLwY
39gUlUyrIpXoX5RrIfY/M+KBkb0YdKL6nqhyhjOTvxlMgePtBI3Zt1clq7ldsi2UxWz9IKLdLJ7/
zQUbqeyMVVJacu4gutU4T5rEQiZBRqgpFFGI2gqobBbMtMtG49rK5lytUZyvzk3seDLxUeMnkADC
tQagDqxL6NwZD4foFHWsRH5SrOIMs22diJk3YAH2TWlZZlbvsxqf2zk2WO0/Tl25hVeFqEzJaxIN
Q6HTO97CUmaGU/90taJhA7KOMcaMfbbnVWXsWsoU2RVY5tu/v46/F2M20Gdr4tQ4idPi4KFCNuT8
a2mEi9o8TLX0TQNVENJ4DzxFZq5q7JUCgsxBwfNRvPFpbTjTEZ/4lvBSlTBTTJzacv2wx5LsB7si
Uck64/zyvjgsLAfGFtSaJHaBd/E7EDKgf/aob1uTY1KgaDNEBVoArNuSsAjcsJghQ46i/3clEBK5
PZx/XFue7J0peamPch6I6I00SuyIAKFj5LW8tKdxRfAQ2rEalrrkaqPuA2BLpSEADFnYc6LNToty
80ma/Y0mts4Xd2gpl10qW2K08vr0DDEUbYPZi/SRslThl2ZT5qnRr4BLKFEdQ0ExSTas5mjA+pTb
Fu42q05C8vd4kJDKzZfMLA3zfNcvXruyCHJNfXVcqdaze6AH+C87RG3cO2lnETiCfdlAo9P45Efc
RUyziHd+0d6Qa4ew25crYeH581O2UJk5iGLvhqgFCErE1YYPd5QLmdDA/G/Ma0CaWYJbwTMLV/30
AHHn/BpmbTON/gPN+MzHqv6mdbGQJdvZnrU/O5MEXljLpD3G+wfyHLRgdWuW4UHxS8cg+k+wYmGW
dFaZyHPzNJTd6epDI11QTUuI2MoZCQgI2Z9V7MokucTg9jrZmfveFK3BttFlaQFkM5r9w99AtvPK
ttY4dZOhkmyx1MHVbeiJSZ4w3aIeqMCZ9CNu65N1vmXLaKffx2GwEOduKHhc2aBB6xPJ+4hthCPa
vE7G50VKhiHcs48kTdagj33v9C01/2LCwcKWe1o51RR38zOYjA+r8qO9wpAtzk5sllfNbugHAmha
L/JuC6/IXwaRrHEIIcEv/cLGaKBLJ05JnNBRubEXbITDHku+WWJHqPA7TbrEdda8lcTRfV3blWGM
/7pbSQWKYk3EN6oeA/wt8pgg6KQRjPnySIEzD2lmVrbgQpdO29Zh4DBbUkoPpGQcD+FcwcVgvC0U
AYzbwfzCdl4veBjdI45w0w73qlR0X66LtHZxRV3KjBUBycutJvQuvMAwT25CeBKf2DGFsm21+Tq8
2id4bMy6/rYqGr8h1mM2M0Wq5CZUURbCBmOo2wguD2kXUPrxplJwxVYNw/PeiWccfATUevnbayY8
HmcuxXVEGveudWWdK54zRngh9fNMNN6aZpjKC8AJPWpT7KJbINTB3XF3I4dxdNH3mgqD7nGve4mh
qe7HnDZ6SmHEFyaik9Rr/q2Ykp+zjTZxcVGIYqOqGXiO2tfEIcMCPqKZPB1UuJ4fmpzZxdnEGRab
N7OGWrntNIJbNauRYGl+aj5Ivoz16v9Kxc394nLHmgXapiJWtUl308FNUXH/GmIvveu1DSjJlzQu
XrqzjIifLAM5lP5ZPEEhhTDbe6vIEpB3srGY7jpn35gk5ub92nDdUNy9nGVG3Z2bNECgj7e2b8Cu
Hjf+GHRMrCw8xz0tUdDjS8OsIYR/6bzhImCNweH0BZv1Mlkz2sB8Iz5RBbCb3b6NhkUueDwz5dJs
yVQPjmNVsjwUluZeWP547KmDr8JoRGiBethMyB5vNkpTdZ1zecy4HmgjYgjuDhuXiSL/C0Eez/PA
MtflWiLy8I7un7OF0hXUgB52/pToT0O2x8llMyczAv4cMWzsJMU/sgt7LLuXRL1SUnVzpxfV07X5
BJI3ZpG+CDw75iFJ5fQHaLL+xaYOWhXitMbgvdtkBbBZ/0QiXMBVkqsdy+OcvzI9Mg2FNbt6d+fA
RsdlMtJLZ5GHWYrT+WjmGsj+PgQanxfJ9/efn4mBa6dTqzqOPHmnevs2sy3Dek/EOl/ew2f6U5Kq
rZ8UJoSjuUR5vHRZT8aWMPTpmX3y4RL6Zp5S1ttSV7xXpGbsBopr0wpQYUBIHwTgcUfrdBZg5O2d
KaMxsrjuGPjVTzbcmxUVOzJhOLqVXdiIXsPBc1MkCxsr2HiF7e6v33qcXXYXWdyMkMhS05+Kz4QY
CmmZIZV/SygZXdXskpp40Ewi88JpnEPGvPk6b3+QhHM4PNJTc1m3P0Nel9GjVdE0TPlU40GhY4RE
TCSaLLse3kC7lu7KTAgTop8xsqQjhCFH6xUPfuGEWE6n5cbWRxCaYsORG6Tojps3fNTEdH7YKJfO
I85Rmyi/UzuvNqY4rAI6FVu7DEfQhkzEIELscWlZs5vRsSiYvbKvcDozBdQmbWWH5z4GgNn6zyKc
5DyotSVzt8eCsjmI69MSG2vMiwBWJnbArbjUBho9y1Qp54YfoqYrW2/LXPiMVbLZFwV8ZMC6hVAS
9gOCwjVfIdvqTTnEGXw/tT04ibTnixwGaR0PjsSXMzQYedQy/L2u3RR2U1Xni21K8FfiVa4cIpUN
hNDMDJdxZm2IK6VNkvXNnDkRNWxMNb2Rh4cI6Gr1F5kNC/hAp5mB+2dVhsIKzfGjEucfrSLF5X5x
G+BcT5GMo8+5Ev/SwAyLRYeHmnJHHwFMWI3MwEpP2/vZZxnIAK8ctFYDQdPjW6jdPDMQKYg/83Kw
p5JJAuxLAiUEyPNo3rtxMaX8wNONYlRycANVvRiAHvXRnfoZaxYAMFIox+IHoTfFg8J9oHlMa7D4
juJ8YOzBkoi7sfQsIRNkwziB0gfrvYuUFVjBT3iC/Drl8s4YxauaZ7d4KsmEPcuzvRmSUGCO7+Z9
HzPwpd6cZlbASmSXD/2UhWAITe6v7nJrso8cLLtuLHPMN1hxWv2vCMMkI7eY4EsyHGOWW/lbkPHq
M19r5yUhSFN/3YS9pf88fFZtNRuArgFeUblaKiwpD3yWhiI0LCAxI8Gauq4Ij1PGsJLcXx5QaLgj
Ejf+izQ1cjMOuRVz92zvmVAZgH1OxgMj9KLPqjByi10/wempNaMHbjxVAVWbXfHq4kmfeUd4hW6/
NIfR64uUfPl+d4K+1zO/FhyMRbCFa036CbDB2e9szphNYf8J1ZwaIiTMBdxquyo7IzLzLM4iKmYk
8H4ko7sbwPQWqeTequ2831smaLBC4piY5pKgzQj2tI2htglChkJqoeL63Qdq3vDxk9XjhmIne5ei
wGyGexfh5KZJdNJkdfpUqPEo6F35oGX5F7Wv6DMjE/LQQgDhC7mLa93n5vLTCOvlSn6nTaJNJZGG
CcQmdiRTfffoQrDVODlCJzqK49vS+MoRlE+Z0RTMb4LMMbi24ngsnnkh0GsRaRIWCJRHwTC2YIfh
kSQqqGChhHJpbffYbaQ3IEKLmVd9+Atov39Tmq0quHMF7sIQ2LteSqN7Q59+lGeXwnSUZ9ia2+gR
pc+/ppuGh99GX86Wz0DrbUPsAZ8bHsuGEsYzaczas3EQViSTm+FLaKPEvDhGqfuaUKyXOejuBne3
O2CATf4iMmAUlBosMXuztAS5h1GYSB8izvjTtnG4GUraj3zSgYbFrAqJTjMkngNndzdN3VnzBDvD
ySpaKZniMtXQ5ZauvepqIKJq9M/qL3oQBqSNSbOfEpjPHG3L5YXqYSEdwgf0XoVQZtxexImxz1SV
Re75C7Mb9ITXvArmEWMRh6ughxOlhF+bhxFPV+cjQkwpg2Kjq9dktHsi43EOhLvld3aQ+il0fzEI
aw7DxmlOfqSjUDZHp/4czWDW9xIdTV4MKkkedYqWCA/rKfmW8QoQQl9z/OegJnhksrwJN4wAdsnI
D64lTNzF473ywFrtVGOvd1rD8XOuM0VbZDOur7UfJzQFsncUK9vtRHazlm8Ociv96xpS+0wap8vp
6qsWuYiME9oc8rWWLNUE58x/ZNpm0LW3qpKXBpnpauOQXpzP/CBbIWmkhYXQV13K53PwSxgukC8U
1yx0vRiyjYjIchxK/4S1TNVxJVrL8G3wroHYx8+ks+bvqWHCfn/OeBSSRtKR3EJEggteClhbMuz2
Ss9gejUZvdwWAvNR8hd9p29U9ox6aTnQMoGNWWfgBayNgLM6dBvqBhJSFXrq8go2BJMLcH7jbMxG
PRA96TnPrvaG4iP3ZMXwDZpnSSYA2ZKIR5V8WXwAYL9CEm5QA5qMl7f+uYdNNBxHtJGYQVBwL0gq
4oKv/8eB+4pJ1dchvayRFZvI/hJyaTkhdw3xLmCl8rkEpun2aqEzJnWyCO3RAuBX0IAPLemn1Vui
IF5HsezAHBSt02hNJPEnItfkGM+bVH8KMwc607mUk4h0RXIBl2KV0f2QGswr3RM0wed5dTLPc8sh
P8QFsqGCUl8AKMUw6plqSHFUW7ihC2r1X81xnOZWWITglSLavlLfryYs1Iwz12xVusBu/I3b7lwi
rBhHx/l2IXwB3jyDzhLphR8v9jkUs0oxyblp9d3OLo+Pxem3x7MrbEde7TywiXPfiAWdNpnYlfA1
wudFeeBPiKAoMC3sOq6bzRnqpNJjH+n4luQuLuH/TelyKqhGejPyawWbAKoh7oVQGV9xPXh1uGrb
07QgIKWjEi8KLlNw7knR7OqGnt5/ZuAnMIn7EtmfMMb+xYtYLc4QAYrZwaAm/QHUZnjpdZ3N2iG9
9clLCYrLi2lq5GOT8rErp1sIiYXq2AeAWwzLB7ead0zouyqkfleVuOq8NZVmmFRUllZajj0GDE5Z
p+/F59CmOfS07MCooxq4b8bgs4H4SebFFVsTE0wttfx4NPuhDWdaW3jH/pdksx/M2XsliNS0kX6i
xsT9bMBABh+uiRKIyXmRTwKD4uioFC702AOI9u9KMzbpPIPNp9EmJJ0v4xzMvA2gB8QAyUCTXJKu
la3EXkNKsy0TY6fwIB5qWjWKc6drpIafjNEi+PFsTQ7MZGBXDtm583mH7wVRqmLaF/NaPneo8ToD
J5wWI3GPm3EGyrz62CDg6HlBx2JTUr4eh1DqObvWBMM3jipEnbs3ugftuDs6cCsD5epq+M710AMY
aXfw7vmjOAJwzhli39HPEkRLVOp0//wZ1ayQp1IsO6Go7lNNxPlnBN9MMlystyiTc0hxHA6I4v7O
ckL23oZopTRBwSJESUpY25WVkM+Hj7EyPuEAeRwMKqlMdKXRSL8GFMB8uQzdZOFCsIdtabE8HaGx
/XFPclzhy3DxNLdWM+G4AcHi5h7XSlWDIHAXDtd7eQbm6Ck6ySkFT3TYsQoiVpXK+oqnc2ZZ8sI2
waU9Qq6nbwRXQXwtNmLDXG/IQcWpEffD/UV9fDEI837sUPynABrSSyankwpYQzkts+0wyKzk4T2/
lfAsWJLwh6GMqia/w3ClUYYtq3ooTpvEgR+lkHrVRrl66G//JSm6vI7BxSnMj7LAcO2u5pDmlewV
K2pfINauP3GBWMe0S8Ft4P3+rGPamzm8eYMvmNZiF7SUS+czJyefjfekd1K04vThpWGtDwxtV+gt
1w95h+AEENv8eT+vXg0NFzeb4+BofTTIC6AgNBgXBJag5Z7ra2g+H2pkzPuYSXbvIAvBeAKEPIpr
8tzC+6Qxec+LpjqGogccw5aay9B/2jpDU0HlUvbMMxs8jUGT8b/lS5kceJ/G6oQk28XuBGw0zkEU
sn6HKJGWcu6Ka+EjtxYDsr9Yd9Dq6yzTRNm5yjE/adB+dliw7JftbXJVOGaKXPjPiFnmsQ1OXlly
eCwqdV+3/ZDWWDwp+oAM6DSaKVUIdn9Jo1MStSxRx4jLBXsOs+Lx6sqKQEiFIfwg5xDDtn/rdu/C
0TLrQePyFOCRVVrL+WjLab0LN1JZkoRnSf8Wq53jBw0WTh5Q0w0qSiaAlHU4NQnN/Y5/eMF+DB5R
WohAy5z/wclXe2yCs/Quhwm7lmBas6VtSkVuIu8iHNNnoA+H/SJ3jZor+ZdZMgzoM0HBnUwEMwGf
q+cJ+B9KKT4PJIHBg7oX6oFgQFZrY2zxjaL6h3Sr1lkZsR8wSG0VsAUlAqeDMSfAQ7e6kuSTT3QT
YMRWZZC/NlmKWb0pE2smRyV8jRVcvVhsnOdrKIJdpbgu2bkeUuFclePcVKcyLTuoh7ePrNMcLvDq
dOIgCzoWnYinapQYNWkPJbOE0gGmsE0rhp6eHyhmIFrNzQDdMsfHyTXl9sMIEuQ6RrLLJNQ/JMD6
LKu3sXNdXR5MP/V8sYUvk3w8p/Lpkml29owk/0e5PrTm5LhLp8d3EtoaiojxOsWMwqMgr/S+ar8L
psgeEgZjkDxTQKEeV1Hf1ThKiXHD54Gjrp59tnhH52xNxddkb+4BjwYIRW7/wBNn2LEn3GpoYfsw
Q5bnINMyC9AkBMFL3k6FEVbkpNcFSbSYPleRwfCo6trzHGJ+LOs6wzp3ts4I7hGnbxG74L2nMoc2
lI2ZC8x+CpjvhKPKu9YI5UHbNlAy6d1ACQXtx6uEqJMmFzH1DO+ctRJJb7PNrJeQO3vnTB9LJehZ
/YD5DzxgUMGv1xtj52cxQLQCmGYO0aUYjqH2lTwU1VggMmQyOk76otTUVv6cAiUN4hzY6d/v/7nb
OezL3LFPb604cf0TL2MU58svCwEQUxGCa6Ubd7q7JW7tkR1S4cIFzQSsDNTiLVOoYYsuwUuE1jhh
/FJNPAgpWCEqRfyFkBnHlNNAdWPg3VqZEyrze5xxMG1SDlXSfusSwm2eKKSCVOoE9bwiNgo3Leh4
dt/JXnHk0YZqUtYC5K8Ee6dmLxSOSfz4DA+y9VabVBDzg6HqONaomMPTP1GgxS2nZZbV+TdN4v9w
Omo0kQgfoNImTeRYxhzxBUabupYGG+v30jmLj4QStp7/0QfqwKTBzH8dvgtN+X/ur1iqVsikq5K4
1/zGP/0LvOBMSLjZZpZQgyOOt2urVnWtAb0t5pkHNHUY+ZPSsdv+U2zbfYC5B/8FMAHcV4FG3JJC
ZDhGSw6uUbkYhYG/JMbYeuSP1ztfVRpvxZ9TcpD6QdQoovtif9pIj2Ay0T5m7AxPCdLDPxfKShcR
K+ay3XYZSkWv0pUZIcUGuI7pZUvZrWwITgzGYr/oQanFd0yUUvleg3pF3CytpW7QPtfkvg6DVyhM
6i7UbLIlTfEly5UZkKup90yZhdRm1ayJ+m14LO1fWD9I6KZW0w7VH2YKwr7/PwWlpUs9E/gwgMpJ
wq55N66JeWP2BzGKEZhD1GL+nVTOlqr0Bj2Er4nDOFrNrdKMGHCFK1uqO41gPeeomKH8k0VRGQ9o
znbYftEs6oEt6fzyS/RaXiYs4ez17JIqsyWZhSRltyTqSMPCLGvtdFR9K4kdnhpCzHVjHreyr1Wk
BS4uLE43IPFmkNj+xjpjy1cIFF7ZB4WrlpdBOnfIgRP5w4DrV40YbcMJuWoKX4V06Ft2C2lx15ZU
lEbfR2yCPGeDQAZWb6FSMuNxRrjl3v5wfI3yaktGG1vjXiSaPhfni/sEk2YEvCvEVCQwrzY/PShS
eTfQeCb1gEN41u5pJT5yPerDrMpfsODov571j6nswQT9Db8V1c6RL17Ask+xyWaw1kVtCKpc0hee
k33AgFNRjoscqICWrJ+drObSNChka5X2LDSUFRkzGnmeQs6q9nw20rciJh17vnfS60o+zGQAm8c4
bahmJaPP0Rk+PZ54UT9njASDEHOsJiUVLF8MBU5+LW6SEl1Ijb0FB/spyI4eWZVv8vSRiMFyqheQ
NiNzjtP7hFeitbJzIgbmvHLxojBLWi+c9Oho+51ITdtreSCbxEITn+UbLbRMf76GvIJ+39/h/Dyx
TSv6seS8vmrkkDCbHhJFitadjmL0Q1WRt13cuYm42pQdXaFqLSnFGKn5fj6nOFqac9La/uAZalEb
NlyhoG4xU6g+zSwt+T89N6SUHI27W14EX1R8gXQU2YnHlIN4b8ErkvZcHkNXEqUuqLG7qgmqCk57
uTb5ANrETnpBGoKWmjQBGXG6ytk2i6pvraL+SgQRRXoPSyNv9m7CMzRAmWtG+9G34HjVTaP9qVoo
GKODPS6vQ6njeZPR8l43YSyXy4NuXbCDzY4ibY5UQbdJQ1+DKfIQxRcSIHDOVr7CgL8FnF726p45
YQQjjTjQmUoByfq4IF8yemk58fP6h8wmF0olX4IRqYrn/hadhTySunSJPBxZcMbXjZrqMOQEdEw6
/WgjLh5q3dF+4X7+GpEJXcd++zyT5S6oLQFts+JzrZ3NLYSsOnzkf1a9o8DeRB2wfML+A/WtXKBo
H+Z1Q9OVpA2IRf6gmSiYpcYccv3M1Xg5lE/zkyYlbwFrSgJp1NGmfowaiyKEHGqx3pgcmGgPPybu
3d8Wy/Kl/JORUCr9H/YCmdhsnYP92+bOUySJmlA2nzbAGe59LdNcZ/FHMQNzYetC46IA15sHO/Uk
7FA/MdIfbZO2a+LOhfvX9fAnmMMECddqfpmvZUMbi94wySbnQVqqwhag4VuC8esS3+50at+w/nuK
niBNM9WVVMeXVIdeeBCJrO8NYFxcREopXqoi2H+JBGcdnPTzcluTqdEEeLGqnm3RcWpHuNpAqMU4
X3MTL+bhrsJL9OSQu2V5df2KStOmKgUbjkIvwdu6sgGGhBU1z2xcVrKeKSMKwKr9WMH/QyNc7+6z
RwHJR/puAIsntlNfl6H4BQDt+aVHkKkeSpawXDoJNKZIbxZfuLbPdV33EWsyLUGtzk3X1pYMOeYE
LtHvTOTmPWhvssMu6BloBaWuGtgOnYinMXTBD0OsHKt5IjrHgFaNBM3C2nxGES10kh0VS0SvT/XU
dHw2Elvxd+JbiUh18yuMnv+OpbXbs/+3M70Gir7tezD/iFKgrzGWOLPIJd9s9RQAPrCVYDrsMcqU
ZF7UshGceVFXKyXPEf/RnAe2HwnkWQOciRKyKl8BtRxbV8aFzRCbUKayeh2iR3lGwIRZTs4LxbzZ
wBCyCYWp1CYuEjXk4WAapWsMkJ7YcbXkANFdxykn17nQXm5z7TKxMn4NUfTpB/H4PXYUnOtJsiTY
w0JKl/POyz1C1ti7SGcPrizVzbx531az982igH/cTmi9jXWgSeoJ+TohM6qHADgH2buz8KPZcOSN
gWXvyeE4MuF19mmy7stdYUrt/axvnP6XYkDTyeT52ZM8D+rZ/dQkOYW8eMYsZQdsfTDMOuBQVVHR
9/257Lj84ekLCTzNa9Gv0ClKIoUVvhI9N0uEr2MdoPdTI6JLiI2rSTwu+onDHWDXOe49D8I91YzY
E0uVawCpeZeSR8WFarM09kKrCcjF6cmPcGNq0DUB2whn8JGx1KcTdf+9ZEQgdFReLNOK/gBhCKHc
p+zhdikjxIoL5t+TXNjZ/5h0DDz1f+SULNQPVUYZtxQxVAo2IdIvr/39VM4bL55JuAwEGBCp3nCp
klGpuWXxZMbwV8KIE9zhenNdxvSLA7SGUD6qDU/pFxJKCW3Ni+2Ua9NuChhbPjVjdRxvBKt8rpEO
KqwR7AwOocwAaT6oER8zOANSn0/qV+IMV8+2Bej1MkhfjhjTRjD0aQLZRs4lczAox5AtiErZX6lf
1c3Shv4csHePOiSm5keh7FK77VMIa5NogyXarLH/BLaRxpD1Yu2i3taaFOdYwpVHzj8U9KR7rstW
GG0p0cfzu/SXfbCgtDQhwoaFNOndN5G4qSXZCVFUF5d8PbhcS+9BcoJIdxU2Zr1FyDrgWOok9q4q
wW1aHtopU4YUGkxqGQiDhCztgOLph4Rw9v/u3xHPCyyFSNj0cOc8KoRVI+Dik1Tv2cZqOiNBzk4Y
30h+eYbT64FTSpQW/dIYMw5JMVY4niEXTUI/fGzMQYNbi1k7IrcgSR60hDDur+R2NY5seuSv9c5S
0WIM8WKJRKA39intprXRsdmeOHKdusAq00ndffhzRTZuH1w6ctpclZTZd2xebwnE6kwG8KAvPe6L
m48p5LvJ5VE4tAdCoRiQ0M3HmkmhYy5b4hHN8I5PnokghViXQmfjMj7D/gTxXloXpaWr2x33jNdp
yAJPyNn2ytoPDR9H0thcPyerb9lRDmlDcRsuzdSnSgHV5ofJUnmw1APtH0O5YF5N76Fcv+uG155Z
MvBmfJSbnHuWduGfCyG7p+gGzpLXv4OHSpyBt8Sn3AS30PZOdkuD4ST3qwhvMOTqgd214bDnTcPE
PRCTd2wMbrF3yncLe5HZULy3qoUWbBVX1QsAndNxR6BaJD/tfhIixDrrEEyfGTgOh8KgknNtg9S3
o99aSeknvxiJ4T/feTNEiGqT34BQDRH+AXdbgDlbfLIwNJc9Udt+ea4sLvJjK6cLZqgnz9/1an6/
yQDxnZpP28iWMMzIU43hTqI2Y0iGGKgWtc7xUeiSemB7xVNBYcG68mUWE48M9NdxuRG+6rf/b0cb
yFBW/fMKMNfXsiAheIziBSpRoXfzxKxzxlurZSSuSNcRbVWXLTVu6wyph2DW1ENt8rktyBlUz50M
C1Irtmp6SD2HTfVDuT8Bh/nchdvjG1NO+ynIA6KX1MP1zhvPeYEuo8gjN1/N/L9kJch58lvC3IlS
lS1lboD7R9iUXHN2GMKIkSS0SsE9R52+Vs18KhJ2QKhGho+IYjPJG3zTJL6eOL1zYUKUhakyYywM
sFwVJpa+cqxmmdMD/EbFMj7+4da5BNSHyaBYdKnwV1hRqU7wqHd7L9oBrwDQ52pXXgQdooZnh6f5
/5QzTP2BeyVvqA95TAwrFpoR8qgvSID5msXDCK3Q6kAr4pcyYf+8I3b0dIzJ2yxD98/rke1Ur1f0
JMPqe6yLZKlvbVKLv7qSkT7L2e3yJ8uiIj01ABpud0kCsTjc78MIovXvSpRQCANDk0s4pqacmYLC
6515XO17Qxq8+OXQ9Mrq1InhFSkkFKkPt/JRmEPxeN4mOhmU5MD32zX4vpVVFXcHE8ATHfmv6azd
SzsoFnZCgsTbn+qgBoeOK4pFU/tK05fhAK2sX7xLeuMgu7mTHz0//fBPoKkiINK7JE5dfdaTjgEL
UhLognJJ+lAM6E8HEV0sL+2r4bgGMiQRekUopYHp+lHyh8/KqjsDQh8boMfVhyxRi5Mc3VwXEjpB
bIlzRU1WlOWe8x3CozkOlgBi3nCuuy2Kd46CPpSIt12pWWlRorHCdSTuM0yPdHA/MaRAzsUKz9Oe
7VMnLEZslw9RCiHyd5ICLFL78IrMdE6fPOh37TpWKXA9Hn+cVLeNsZLp5q93XzUnBP8onnBBwPyb
bi280y4iA8ukb2oC+lQfj0a/ABW6Uve1fysdiYU0FK7Bb4MSrm3UjleUfK7pRbMUFJWFadC+6Ju9
hAbenmDiFHUCrDS6z0TxqcfPY3hS6elW4jmOTMx+ht0Vk6mxC2N8kQ0hGXGonddx9+/g9TgJxwTn
15TsAmE/GpHtEjEbrwkb53vXBllQSE/BBMkwLjL/4W52+Cz13zf0LQ3NSCKK0qPkgzWs8ZpO7rrK
dKGRBMXGhaMq/T5p4Y1EE05mHGSrQZSlYk959u3wPNi0IOCFkKNfYoFi/pXISVlVHvFF8axGYlbU
sUXMQwBLfWnycaPlvCy1CkpeqSj1NuMhHx5VDZSYvK8GGXmGjlNOU0lvN1gfDGqfDZXRIE/NqUeh
sQv2iTjdvU3XSG7HxqF28PXo1AjdwE8GxGXtcZxJ2bOfO10VB0k7A0S3ZrKa1YWGcRkC9nkJamRu
lGmUXd15VuWH2/8ezSQBc+dqGAkuQsP7G9opxyI+CnNgHk2LwTFuq10oO99brci2/VWIbV08sgqi
7AJZwZwiab9ij47QnuWqarMi34/HD2X16YKTMfhROinCp54OpsyGVmdlP8KpnFGSrmXwN1PMj5rL
Cbui1t1+reHV//MwkhhKxlQmCjKymr2AwCtYqdPh73d5ZslLh2/njmUeWSUMc51e2RtOGqnsmarq
E9nRf6DdcRthG+nWvodaX9Iu7wR0pnPR72ji46vk8BrgEQMTennGi2Le0+mOG79UgQfiH6zVk8UH
T2jgvZ7AdzBdpYPekYRfcJXJ8Ku1sse0bCTxSmnxvPi8C9XUFImdDlGRuuPpjSeSJ+D7N5KhhVUD
89rBeIAJ1U2377eE1RgL8X+/vm0S0d0PLOOH7zke0SbGXeU8d6Atmg1wOfeyx5IsG4zJNzwvqY1S
PTgEsPOJr/bUeeXhdS5vIFLNaAftb6E6y4+MM7DxsDpYcehF04+yE5lncIUOLtSfFAp3NpZrb40D
i6eN3TWehexwcnb7tbivpnEc4wEk+kVU9A6pf642AdvCA/Js+63B2faIyYWMKzteXTyW3Qtm9hok
AJqsgWBcMWbVFJSDXZsJHCbpnZr65RlGshgkFuGKAia02bQqtExUFN2I/g9yHLnALtdlBqqidT11
51TC4+fy5Ac2S8GhoWYfvs2FtSPp+6ongB8cDyV2e+gwndbD2vmGTl36xsCIYwdHvhUmrJ6Qal/+
zbYA1+7s7mi0C2eB+kwYC+arar7p36MpVQkUbIkSoINF9wrX1CEmAOTVvMXMPec3ZjqWsFvDP6gq
8XoeY538aBTwNgep4TdDjdj1adaDtsqjAJ7GAdcBSRZBbWUrWwe0HE9qpqBT6/SOkXzEO/MsIAvW
Xuy0HSTO9vQEw2CKWQpAJmNwCgFQg3hDTRLS+tldEV4Z/EuJ1jdO6o960D+EwT/7UWmQN8FALXuu
CHqYklWOGDlWImd/Qm/ai/5Yioi+Zsb+OF8sLykUO8mNiVsBPsUWwNZkHvn9+wZLNFH4hphk8HGQ
+SuAQlSFg6CEb0oHqnjW2HRqbhRt8cVf+tgHg9YLr4BdSVix3Yc+jAIWr802eNrFJOq1R4sO9OZo
HrObYb/g+FsXRwkQj8NXPrpxyjO3nj6fsAcpi0bmTCBdlEySwSVCfP/PXFbv75jWBEPpUsdgl9+b
t10MmMFYx6QMyMfNb68Taok5/FZJKV98NMpdWXBrfUnNCOW0RU72YGT7CHmuZGHOmNJPx9E20kXC
wv1sh3QaNoWvjKKDQHqudEUZVQEFh55tBMI4E2H7JuhAFsNnRUBa/ezU/60hGSyfhKIpdUNYek+P
ovR/l8EB5N6cLSqNb8ozr0qZQe6B39LPHWOnSdUVDpnn8wBlbrtH4T3wQXMBc6rNckL0Wo8YUxDB
60EJrU9KCdJ0bcH/HAr+lpqmKISkoMADqnf/kixh8k4jhwz2w5x29TLreYdSUYZRQbAEcnsUpmrR
dLVDw7UoMVZfuEL3HkNYxgXf1dHb1mTAc1fBR/RkcNYbkm/H0dRLeWtFROyVIlCNYCKFfEaNGxdt
mUqWGmeV9uL62CqoKgbze5dl01NPVr7RIHrWJ/nYR2nwCH1Og5LYTCfWmj8HcPJ4J7jW1FSJOEkG
s43etxaI0AAzwEriKI5n78qKCSVGGj56L0VHgr3VZyaDocjeaEhW6vBtoRcR9Yf4+oLLGX4eyBdP
ve7VJ+DDJhA1R60NJ5nOivE4bwCrlPadwCM8T1AtoVIKhBDYf/oC7JQUKVkFYHzJnT5eZ98bK/B8
2SUDFuKSNV04AefUZu7/XMRUr5JPjCLxJdZPZX9tupiTYUvWQZSdlyT4h71oBl40ffOJ3JcoAGew
n9XgsHsAvpquyTFfrG+S6zcUOqxm9lLTxcYlS5ZXgswsYB0e6kXQf8iclR4iYputfXII8IwGJC4z
lgUHpleA+XOWTklMAQkslqZpqEb0lq0fe0LNjashc1DELsv7qvgbWyrewIVtUpvMNUoghM77I/3h
4tTHJDmxk0QwKP5ja+hhx1GjnrWnLS0/zrEONsBP//nH1MwRJ+lzqF/Lyom+V2hx+wQH5/HitTcL
6m0fUpGyBdBbGDAy7k2nKy6v7gRWuVBqozZIy4+PtBwEzDVbMy2B6kSGuEzoJTE/s/J7ReWWZWn2
VlbaPagMd0DIbGGS1kw8GEzmm1QkhzcvJJZhlzrs/4QhPsrrA86loEwnBdjVOcf+zuRegxmsdj4Q
TzJKJUliYj4AbQvVDMSbLY6TvyD26B3YZ064HeWO3xRr0Tbk2iEnIW8awexxfADaQEmNrP5hOyrr
hRNdkjaOD31/G5Z7fYQP3+JtzqxWxP2THq2pfeB1aXqIJIA6ekEiyoutzF/QD4wNYLZ7DPJth6AC
TTS7S+tWGI0+lXSu/+eiubCla1gCIFWwCryhKYwuWu+/1clDcmGY90ySXeDZ6g5chRmFtfGkVbjP
cHKutCjsi4x1AFCZBVyZMGY/nYajoXrxji7uhvzrLJfPPSuAvGwncNinotb8tK4ojAH9UXZta2kw
MIMDkqAVRUEkH7+ZnHUUVeaXGcBb/MI0LQqyKYhVwUGY3zl29VRzD1k1B9qxtP7iNt0fxSVgLn4a
gt03FU8FGT0OTFR4BLNT1a0kdC91JKxvaT9LjIzUpyrQyQOsYkmgf8/BCCgyAQm1NgzFThArKoKk
cPdafrYFdDGRcYHwK0MnihiNa4pmPJBlISEQUY0G/1jgYU0jSUPQb6wYsfamS0ngI+6T1YxR7MNc
cZ8+oSNxAg89gs/DI3B8Q8+Ne0zqg3JAUNSvSz1oK42XuC9U9UVa0s28W62CPPfwOlcl3en354Et
UQIN0NwaB3c+0uY1++zmkrKYwcMa03ahn7nU8l0iUYcNRM7+ytnYOYR46IEx+cdOpM/kvfePA4qK
KAmb43bk69Y3kc30vAfJC2tK38hNSFfiG9w79Ohpy6PWcOH1mTCwWTDeSiSeIOq7WCU90V2Ev8LQ
86+fKYe1GG/diG0WWPFCCR541EvTnZTebOrFW1twk/Wp6RQ6byZcVD8MVIlpfNKVoef01zF67e21
4aMMpdU1VurgBwHHo/Iwl75vVH92HJSxCu0r3KTd+Vd1EntiFp4UdRywpGk7xJmYaAe2Y7IKfOVs
c+pWTmWDwRhthkRCV0mdTqtCG5zADMNl8jNfXKAqk26MUmTmDsyeCCIZSGwPI6E2fZJtrGvsm5OO
CiW6I7ELv4ga0YcmLdSy3x5ocR7FNFKUy7KeZCdJXAeiLC4azCeArxfHxIVAkrAsOrStkX5cnHTX
iaCyq6lUwETqfWUz9aGdUcOuahg9bSetnI8iGougcTjgGuFoaHWglPjfKhtEPkQLT15miryN8Gzy
faJzYuCojWlV1nTEt+Fu+JF2Tcbahsoyy9y1jzfx/N0geHKqkUmnYzrPKL7rmHn9vOlPjp9tn0Hg
4lnp1wO5umwhmsjydFapTrYdBwJL6LmpqWLphuNBk9d8D04Ne6O76l8DeRiCO8VQGgIiBNtFhiR7
fkT1MXp4ajsCaLmSfQYk17ObXJcdSR3zGs0NSNd4GPBztSghjW3hpu7XwECPSpXa8ljMLDciK6+u
Kn3/RCtfvzAWNJqdpt7x8aRNYVv4aOOdTNq7X4srCiq9dX6TA8TGehGZmtTY4ju5EBFq/aX0mnNz
6+fLLbBndByOFvvjTTWeU/HI2JPc0dyYNIFO42+bVNoQT+i4kTGOl8A+cYuJZWl6UrBXRqV7twxK
QTG+5MNT75hPHWWpDgn38/FRYFwoNN6a089NN2pH9xIA0HfX+9hfpXpQp9qCpmBXLmAmVMF27N2d
iIALsRVqeDJdsSTlF2yLjQDycCef0LAuDsfefCNoIsrW+KH5741Qp6D+ZlEHUaVPSiwh/1ittPbB
6CcwkGe5ugSW5cEFhbZxeYLWSm3JHBfJtc2pEAA8blT2UYX3LYpsRWc3+iB1wIcTPFbUx7zSa4R8
aTjaGS4OXhmmWps5o6Syy9d/cVHN/CdLrEeQPYzgoVkfCqUZsffl+SlGIiLNs0q5dfnTrBwhb+dc
JWuJ8dVsaBK+iLxC1WbQiQiwzLusjrkdUCcMLULBPLMGIYzlyGNCe1Eo9ZS55qwKqBadUWD1dbu6
mkBK0vWxHzkuDuPGza6hLyKFUF60MbOVJ1ZGgn4bAaTVFudKoUjbNNDt7rgbRtHI/xPY9P/YIt4j
r8pviU517PheJSEdTXfpYMWs3WQpmMhXJO/bcanG5tMxkaW8YMhOkr8VZL+gMUNUGAWhhT4fhNj0
H8VNq5p8Hu4RDCxEigHgP1Lwdb5AhO35s2XRwIlzihMtMuSWqJirJ9YobEHVppQmvyVSvwFVvSu6
z+RVz4JqsPZQmtY7x9wr5vPf3LXjVSyQcbCf1f4XLGAM3ZWWufxbJCllCjzPsk/ZtJbiCoEMoLz9
r9CHBwItTspOLo48jFLnSxUgyV+JlWPEceown0u3dJiqmUIUvRM3N2iXOKigcnrxvPHZ4F1P/rmC
QIfUCmQeB8j3G+hQBkpsB63oIyJIuOts1RM1SEQgxQDzY90UTnfEsTHobew/h1G7UjKFRyWwCssx
6+f500M/Jm6f8af5FtuZq/Q1stJxAuZJQ9R1sWJ0G4YIJIu8L+59qFvVsemVDJbLrxnIRObRBjED
mghE24DILr65R9KcUwWzZxWNmBzQ0+CEhjII6WG4m/Edtv48MQrzV2WeEh6It2uXdyNfN3VwYPD9
gYEN1xcvtvJrXf5YnAGXHjV3mQJu7y/3OVDFpnukeZzBUCLWBj9CcEg/vXvC48D59fFGfAINkHOL
ddoe26WUMoWSkckm/ZQFyi7hQnt6jDfADy4r/t/Dofz0uRrXkZvd0MWUfVr4EpG2qjUqMztRR2aG
bTIOQIk+nW6qw4EdQckMg4x/isp8yUpEaNrfrUCd+4Au8ZTQaPDsudXrfZfzE2LuFKOfOdI488z7
nOwxtsdTm10XXYkAeiCQbRD1CrJcjpo6QmOrOUvyvCF97TUONFdFshU900wPCeBsS58MuM7eJALx
QwGx/rZf+lL1Tdmlgtv8VeGqPQCSmtnxAdl/9FBw3CIjuX/Lq8YP67qWguF58u6QPXXE7y6V/SAS
fFrQqYDjXoyv17/Hz70oaRi4fibPYDZv4z0p2uTE9yDQpbiE4JiMuacS0U5yCT07fIud+m+y2jtq
kxpTWavt226dQJ7+qv8gIexK1RdQtbfFIPQAU9tPqo8n1uctY+6G15lrsnkFFRCoctaWu2MlyX7t
5qIubKCSl9J0agW9zOaoMnEWRQCaV+HlMvutaWxBfcj0dkK0w4cfExyQUQk7xXEk0R692LQxrPds
7Lh5a96l0khPkg+knxvnPTCnFD8e3c5nQU2iad9ID7bfCPbXBHmoN5ZjBJLg/e0ZDO9ybSARSAhO
LyUC/yJ+uO3FQa8MbmCEx/bAbcoMzmXvC751mMBuCPcbHjI887CKhhG9GzhHfPOQehSB6NDMIYdr
0HFUr98Xaq5pQOu1rJckH1lPehw+wWcZuWqAJDnqClzSa6j3xEs0V+BYxAorCJuvU44/lNkoupHY
hsTY3dfsPHT4yaivuIJTTgXUZlViWZ8l/pYaoUOl1vkcHHLRcwH4qUT935t2i9pN8rVJTTqPK7oO
Dk6GohewN/qqpqPvuU3F1UhJOfXt850J9zCEyEizmBebLEeQHrlxvu3AEND9g617N7MB7+jHUZ19
d3xSdH7AdzWn3CT8kATi6WpmtkxgESw2VhEjCy3ebMQ7jG8/xScvwTff0Gy6kWZhMN6eQ3O+L/Ud
Qb+xVkQgZErfEUtB5FdTVVhqpwuOtHYLrZbBgEDAwJJ33njXlZi+NZlWvXI0n2JrCw4xBdolR56h
FEsT5RrCOJLkzRIU+QEFxBRe8mtWjnBNABmPEtMlR9CfUfyusoRBcvarvGP7CSRJPNf1166ndtzR
tqq4pKmXXpqh46cCcveof88bMr77fDGq6GSwyRXZ9stV5CuX+zs2yXRex2YcpXWQhBbjvnot6KSV
2dZWgscQM31zP4JFUvbM9RxsunBN/QAArPZVU/9Bzk3TxQH0cX/biJncd27nK7E/ZgStmzUPD3XX
rYcj1YKxcPYzmx4aZ0m4jK0tKaiPCZmEeD3AI6kgLjFNzRZpzcGM/9UvM9BBmo8Bu3whwRh7Dfqf
sGzGH57hqYJmo7qIA4c1rMBEqJ5ysZorH+dGzaupiZt5bztZHrW0AmkbXC4ovnEtnnv+usKJ7OFA
E8GTt7vs5NO5h9rb8vnHgV8T43BxKQghe3WgMMLuBjq3sLal5nPRHbraT1QYEGqcAN1EMuVxH+wk
BLYJTDU/k464m+ZuZArmJC+CVGDaNyfprGnRZh5ErDi8I3uvr8Hkwie0zHxBP+e8c930CGzhuT+G
OhXeRv7dVE1Peql2CZjZS4LO3MFvyO350XYeBg6XQJiIRND7dXbrfaiJWFmYQyz5fnLkA7lJLD1j
57dU113/iyHELJxBMRDQp0UWqeZwAFMAkg8iJMt5tI8QfAhIQBMNVZCWhKHJj/j/dKx8uvrWqsKe
m/88bd1S1Tqlab3NixPPvAZB0OSvauT2bnZ9xsrJS467bDzXveD1bovyungSmQ1lkvGaELVtcWrh
Hmq36mGuJVLJ6zc7aTZLgED43HtcVLia2rD9N3HbNoVcQjHajw5t5MM9cRgpIlNWrHfBGNwUW9rC
fTzBmUhMd9CVlpPpKLCbF9gc1zfeCrhM0rQO+ApBcFkFiQJANmBl6BenVWmyCtkNmhBIljv1MoOK
mBrcCdAbcQXvNgHyeCaI4a3hyqwPBhTLbEbx7RIFL0S40/YhwaIGfIxC+gDPKWRVpPE/xCPgPMhY
D40SO1c5hw3EnUQBRCZ2j7Y/ZCvl1fix03MGzQVpPU/mwo9w3kRO10BTEs24mtvHoJ0yarOQgkc5
i8VZQCcEF6jbJUFDUJ942ufXjMYBgNgbY2V7kriuBF1jW7WF9CZS3mGbKxndzwDp0QeVu4fojNAY
3FJ8/etbOvUCRM07/lBUsflqihZHW2Qa5Ne8nY4k42zfMuvMmw7YCRteUShwKvt3ydEED/N3juiG
jhWqx/iU8wK1ILo5OW1/KtjtYW/aoE/Er7B/NN1yi4CmtI8MeiPDXq11Oq/uq3+p1dDgGBkkBnvd
9OtMJV6ikuCozMyCarDhvhsaNpTlMoP5uAfDdMsoOnEvS7x0RJ71R5mPJtSzO2j8E4oempTzYWml
kKk1edOG8DauaByVbZNvhWOTue35SbWcoBbs37lR4kIF4tKeM//b/W4Lj6mcDMyt87bXRS5XOOSU
HZdYDsuI71rwLbxKteL8NjweQYjRNtBarrUL5X2rQLRfIyb4/hNdH1boBUaEs/DKDB0FkGKUuzWV
Fhgw6ojDg3QH4vnUlSrP/Lz/AKxFm83pGbHziQEMhTNESrRqA5aORgnVbqUy8ZZTRK1TQS5sVQpg
NzkaZrxm57QLUHOvIcNyT451HbC13Y5IrEwBkIy7J3uIhEQ79mAgDtU7mCC8awFIj2LO9efFO6mL
RtfeUhSlpz7B6Q9HxmLdj1xFrkLeoR1D6hkQlOp4YfoCitaS9NCdJqxEpbXMP2rQ8NewUwjLtQrq
ShelX5raiDAhjdPtotY4zwctqofgeYCGbmhzj5U0YjsKB8jmyXvH6C0N9ZXHTpnfQ8XD9m6cLRDt
bCpMLz0QVDlUgmEN9ChrmTjUtOnaEsotvk8jsmnVfVlyehiGel+a6/9JIhWhc8nTTXy+pJjiEjqy
yCjeqCAFZ+ugOXNJTmez6LWGfzKHEC2E24aCHdS1OVw7K+O1PU12ubrwsD3oEqDnVqFrghlBqerE
nU5SyHWohCUsoT9I6Pl/XbFjp4q5Onz3skFPNiBNjBGd1msQB85LkhDCSlMFFkXUs6goGvhevoCW
XCBRerFMDVU7IhwBc20qboTeQFaxJCtE2H88qZQfUnpishuVKxHRk8NDY6Ohjdy451uEzcYg7D7b
3Vbt7fCdC/mhmVCOGfNagHJK/znqzlaM7F/Iw3PIlOw/w+WOoZwuGODKeJDYz003XZqLoNOeAvJk
9qlVqaosKai5PUsiY7sRqAbfhs0/eBHmp1gLnwI7aAaJRnD91niFrD7xvkOmm66JtS964lKFtRO4
x/5L+wbwAHzoovpg/BSocyRGbNRGalhjo2Yn0iTv/5I/6A8GyFGvMrUMN9byNbrQr1A1W+9f8m6f
P/lcXdMDx+7R6XcwsYFvMvzX1Xj+eOiuKJsWs/TZKCt04oopMursqdu0s1SzKf5mNpqrkMGkP+Hr
EYKlIVKysjaivcu2FlsQKg93P57hi8330HMhCqUR4czLVnTFbGzbjF7MxQz5A+iP1NLu1YCX8OvN
qXSTaXvh+2MqKKHDNsztJLkMFZUBasCR+GYyjUI2E0l3dh8K0ci1vkVEsYpIKzIFCNywv5rdELO3
lfpfPm16lE1P/GQLWZXdq/hTxOvx/1BJaTUL2Nrp62Tmzl9S8JYCItT8rXBHzzbcLekiIcR/LJmZ
Wlo8T7ABs6r4xjnQPLgOuTexr2BpxVrbD5VYg28aeITqYeMVnrrAthTd5913t61mOHqhtHzyoR99
f08FgBZqTFPtFz3/L8cd0zY2nxAY915HASIBS64JXVY6rOCEFQBSCIV07ZL0jQDDci+MDp+xEBeO
YZq77tGft1fz4/VyJosQujHSNZFXWzlh6qBm74G7H6gCF5E9/BaJ/PrVraFmB8Jq0uVzHL9Cc4pP
Ax0ASQzdre515k70naaCzH8Qd4tIdgfMc6zmDDqdhe9iXMwJtfMBfp7P4Ui93vZL2cQ/R4DnUwG7
MleIDDAq6TQiaegIlwPMdVYfA2KNa5YyiHH1ND0QZJa0TRu+thw5nDxoV2MCUwK1LbLJvjI7qy4r
Adrce9BqY+H09p0jOIxnuC5Aaf5eY2lTrQn2RhG0/MPI6iHcoyJKS9rrNnLiSZ3rlzb9QnFlQ0ea
R5UWvdS29XAsg8rIBU+eidoNcTEhFAATVrunUMzgWRFE+pj66A3oSjuUa6smjRlOzmMh1yy826kD
9AlDminVYP1hOxKCOv1qSnr/TGtBqHo7PP/Qydz29x4w0LfJIgC5hK/WxvW1sBWdtQMw7FL8Y5yS
PaSEBdV2GvAUUMGl0UHEVG3/4DDAnt6jIxnjt5eblofKBTAbboTezpPXFheFp66SGuB93DPIukNx
NnyADNByzD6MbKnoE7taDcTBzxkDEPaNmCNHmAau31fmrMmP23/2DB2FW1yH0p286cYwMik849/W
sOzpKnIiMPS52/HgJX3FxF+YwBZOOox/ji8HIgwf9fKICUdK8EC+q2N2F+xFf98v+vdHeya44W3e
U2awrjd80cz48TOm9eFbBq39iIMuL3iUWG8Mm0dfC6U3eHnLkZH+74BJVzHYdzhGT6XFhJyLTQpD
WTjJ6+5K+X6bGUdpNSW6CcXBvxVpAc16Pp08eQk/nKmLPdh6offBqyejEf2idisp7dt2zynG4h6O
YiDkPUyk5Yti25C+vPRzbVHXE3ZxfKsV8O867QgQEsMLfNhlCMgdz7L/eIs9rRz4ym3jCTfeOvHo
NznEMuq1i+cIjptpHWCM68PeyC9Al7QWsBSo8GZCrKe4ezV19bE7G1ozRowLwSsyVGyMh9VyQv3q
obqyymXnW7/J5Ikbn+XZsnFdK+D6xlpOWf10nLXhkZci7rbk2pzjHjuSXuZCFR9oBIRGdHdn5CER
lkyz0vPdsYZ/ExQf0Q+xK5FNFNtxPjM98qLPVslmcSHocIy0epfNmZa6RcGjG27IKBnQMFdNN6PH
8/J4lT0AqKckwRGPRlMM7coT4OOOteHikv2+4J1NwZsdtwmO0eB00eaWCD4vde4+zoG3j6ZwF78Y
Uo8av+9fCBXx/LOVSU2bBvZSm9biA6L7ffhJMl+KHilkYpKE5mHhhaO7Z83GiwppnkUg+oghnMoL
xhl3vm2TiGg6NVs8D4ES0VpmGWcIo3obC9s80TS7Rs1BoFrMpdeRO/FAYKvtkBvFRofwQbOgJSII
51s+L0ZJyPcuLFJoxN7FtDjDLF0/JkZVjfMXR0eJMqy57kjH2YDyt6AWn0lWvXKbmg9is+cif6/V
fyAiHDkz98NXj+2+Br5bpnKUAZS4PQtx7rev3kYbxkvcdXE0U1XkBJCzEXnquCwxjwQe0s7OYDgN
EaI43c/HA1uIsUzzoZEf1IIpoKzN+o9M4NLimC1Lm/1MQWkI+h59q3jID0NSBx6RYPdL9S1Xq7Wp
BEwNFwQI2NEn6/3g0j/scZtVVCaiO6myXNsbHIOCpUF6ldWbqYNtysdtw/BMfZujpaT+63uJ8hL8
Ny5D/0i3XoM/4m4G2NKQ2k0UxaoPGFpQivNDYlIMyZkqBd1ghNGfJgkLG6/+e31bcP/bA/1zUFVJ
yW4DYTA3uwbosfw9SY06wvii1ibE4qiwt+D5+kmu210aB+g6R9CSVNaRG4Uu5GuybdU2ZF13NNEk
D+ET/hcJBfmP9xgNgF9rzfbBErVyR9mus3DlAhM+0B2X1mW2y86f0+CA2UpWvJxgI5ium1nqAWLP
Lwkc3mIkNs1p0vWQOld+hnQ/htPTWXw5KZ8U/RV9TWaboIo9fkfT0RlaADIBQIjvy8Zb4nBVFJtE
7u+pGrNlEst0JiWSb+zFhCXvXn1HYJt9RfX9UPm+z6J4r3Fw6N9mfE/LqKJ52nI6vwWU6iIfRoOx
1KBpdry5nsR0iPUCXN0zyyVadMTsxx6j9Y3Z494FCMTPJkD1n0ISTtHsMnQmvI0Ou5/eUdYodwyb
9LGL1/iJ3WGCjAW7OWFvD074jol4DSlQL44+XBe9zoe9VSeZLqQ8XOjWINlAmh75EmrEIlK2LcJT
zrSvmSeh14x7Ig6uM3tBM40rTmjQzmEsFi3Xy/s9DLzCdJhrPx2uJIDHbSTp27vfoGB1fgYWI+UO
HRtELg9f5KP9XTrtFTG1RDbOUImykGQ6yLoIXp8EldZiQ950SNJW3foEcQ6qYC0qXp+FDEvmasRJ
HW9taoTSDqls5IlWvB/3xVfh5D27TtZQDCv9KV4rCfGs0iAFCs+pCOl4hfJ/coomjsmzoL6BUQJr
92WE2AVtA7PX6J3Kz2i6NsSth0XHL9kiDr+wSlFI+PEU6nQTUXj/vyh86vaNBdoEQPFKwku4ffma
zB8NpWOtMHts4qFdZsHdB6jsWAZdsLSzdIclVJChxbqpQ/YloxRSimaBQgVHa/BiUvqaA8qxj8vr
Doz0eILxo1wa2wpSRL24qjvtIZJb+ZsG9wy2BVapL2PGumLEc1q+nkzjbl3B/k6bvMIaQU9lyGQE
PnJjNk62IwXSx9wQVY+aeQRO3ix0hYb0rb75LuYoAoQbWipin+H9awd6R44eqPUISNd02LPP7RTI
jpFjtTN9gBg769hAo+7stj7O/9cVWLqEjSuzPapCAcanBnIXSkgbL3nlaiEXE5Me2b6LBZL1K9yd
HvknO+ORxofcZK8Yq5KZFuYU0pB8MegnVh8FDZjy2uBVEb+a/z/LzngNht5sYJiJv4AP34QX5DNp
mP8JdesEdGbAy35KtFZFuFJ/aatbkaztTq7BsNPJAEDRk0B+z3GeOs05daTdyT2TP1r8i4C30p9C
3poGcV5kvjO1/4cQOj25Lf4YjjOzEhaC969FysPjECLK5Y+NT6af7CM8DyeYfOH0WHSqhNXxgr5R
8MtXjhjNX68AltNr49lxK4ZzjsoLogwDpdpod3m+/BTgGqUlliFsPZh51AIDBEOpHPHeGU7cgD1O
7u5MXqhACxBtSqcrAROiBORG8uygMkqJ66Pd4O6l1hY4rGAMUYnhjAP/dxzEmq6nW00o0roRLXTB
RiNBDzVsLBfxKVRcl/T0/5fe1wa8+lWM6c/G1isPsiG8nPUsBnIWMCBn2TqUKQ7W1xWxqK5lsbRi
zi1OZm5u5a6ULllqDc+5SfMjROfXy56TYADKKV01/8JsyHly/w23gog/14dJgBvCjju/zmOqrmVp
/q52gTePlYy6/5sm4E5CRGVAsBOYqurGayiR6aJJm8CDb5PY++agtn+Zh7cirL1bYzflzWiTzuA+
p72wBPamEE0a3IYtxkPBnHPVbLa7wJAwUgaQC4GBDFVSFiStAqX9c5SkyXdTlS6cQZ4dBbVaOxVX
U040MvpdVD3eE/36vJ3ucVDnGrhIpBz8OloD0bFVXng+oOKCmV70O3IgUapPzqgbreDVClldZmMn
UHSt2cynEELfVUnrdk46GrCPHY4MAXK3forgAcMEhVg5p71gvgNxje59anQHWs2lZ5zMQJtt31or
nDjwZxJJrR8JsY5y+ItT2mGrBA7RVqWbDMcmQkpj2QRw4wpEiQxMOAbpavkbY0cHPnS6nMbOGlS3
HOfzLZU0o5maEUGAIxZ9NZWAiKr71mj2iIyAv6GBQZaBGg8u4HJdidZs2MnvPyEH5vZCDAcAxUuP
aWcRKFhbFlf4Mx7jrRGV7wdxBkDRjieWfSiVrN9qlb92bI4j4cbwi57OSrneDgrXVkM/7Yr+R41r
1LcZTfvHaqqu+qlk0Am8c4uuNk56wq1z0Ct1uYQx+/gdOLpJOJay2aPLNxb/DtZxIPW9xX2vSz3F
JNTgX6TCEheTHuJPOCZ4bodmoXKtx4oAgGzkhp0eKflOHWtyArUduUKRkg8yZ8HCT1RZAmYaVt4w
pPoCI+fwL8XB9a9N/6K9PQwI5ADJN1T3oSO5JnzdkP3oIei+NbKNefvQaFIrXtEYMLYKZ0SCc19R
l0XGPEb5W0XksIgAGHDKjVUjYpSJitu3BgLkLUvHOpI2kwgtD+/B5BWe/F+fkJ/MB4UV2z52rDVD
1wQbL7Sm9H8NMHvT9Mie4WISPj7yTRWQLgQrTFIdgQcnm8Pdad0d1wGYAtcUYNru1zTTZeoG6TMa
ZmWO6STT8AyeVxKl/XR3tiVq5kXhW/ksW25tJLhz9anmwCxevVjgvl0HxpcNaABYFibMD/eFkthT
3pgx8ndhmcW1C7sEv+SIQJ4Jq46S6C84QFGVuC2RDxLtxx/aJsu/lnFSduMzc2LDqTLhDsmqwqKh
4X3hgrEhjcB855GBuz78mCnkeFEBH4lkxJObDJ074UgYr8+HpgaNQHuvNrKp+Cb70L4aKBFefmzc
KNKDH5U5eq3cHsUigC3aVHIYXS1FowghhXxcsB0EMhx+gEDPhfic89R3213ZJ2cr32wrIMwDTEPP
pWR+4VbU0v0+ptMoKAyXxIQIWVVpQ8smG0dI71YP9XA/nHNyhowcIbTMZY1MtNl+H2M39weHd/L6
yJM1cPg95KqdWJdDvhMdN06iGYjlBS46ynJLejLegUCzo8EM71vWqie0N6SzfdW1bugjW8YkfoRu
8Sh5gx33C3OEm/c8+QwN2OWT2T5i7PWLUiFLaxTrZBy7TOc/qoTaLor+434cOpYj1HvCllfYKaUE
jSoewbu2xBRDkMmN5xVTqW8Hqe4zALTwQr8HhTfgSe3otO5VddyRANWM1rnGq5rBx6SASt2OG1pl
pDTkX9Fd95L3nQGFWZp38BL6HCfOWkRt4y1sgRkuCV+/XKdQBDlMpKYB+if2WBJ2zizX8X5BjROQ
lwEwOKDFO3nfMb0p2Pe+8DbsOhn+lzi5k5mXhWLUeDElF7vYY4IoLj7xyQJxdqBWgErv1UhtGK/C
N41zxNQ3T/QVnXpoujiF62IFMwJBZ/2k8ucwcb+Ulax7II42zumuvxew3/8fYkLA9WAkbPQ/Ihve
13vo8wKK/Q2WEOD+YKObqqO85BsDtHXSVFMF8KuMrYg9iRiHsnuYAjFzqGz9aKrN+DE45AFcNmrn
HVSGZRI0mUHwCE8Yn+RPVTQlNJBZRT8Hp9UJfRz18Wb++trAYbg/pk03EIMFRiTzZ9WfNFk8r8Wk
D9yz3NCqtsFKZ6mTgz/QMFQhIE4lljdWrqUiS96a5LRe6OhuMzRIlJBuq1Nx6YhBkDnZBxERfAAB
BceRZvCJPpqbN/K71ZGSfA+qq2t4xAkIyAmpYIKZbBAQ2oi5wyzXPXyEICxq921nQNFHu61FeJ6y
fSKMKL8Qi3lINC22aPbHv/zclxb8peKS0Vj5P7DDeBL7yNjY2bvC6bw3HA7tIjacrrBMwncyT3rL
Ynhx9q8/PBsqve+su5G+RcpGVzglUTwPHdV/o3AiCAiXfQSckBZ3LiB8DElJyKeR+a66WNWgCoc9
BuKTNGiZORyGLrQ4PVsqpdpZnjfEfNuPfhV6rdQgFtvy41shFDBXoVmQCdcUcxEFAErQATSvBKKV
qve7YR+6C8xLr+sKfr+caL1H4pBdTKzZeEw8kjLoKJpJxqcVAxWZLSIdjbBfJibmGv+kLKIYunJi
+g0BSgHImn5KnjBM0nCQGPHnDIkbzeAVYmF3gdxmApDHe79J2J2wSryA7ZQ7Yb7KfovVNRJbuM8f
99quol0Gm+1NW35hKwwf3MyQhQtccu0vf4p71txpNG+EKf0IyjzwW+voJOILTTHPNGDWSJwB0NNY
3tLtDETxgO3dLgdm1eshMHzVEQeuLEQ5/nvwwFo8CuCuq3D7574Q7IXRfKI2CBBCa1YGzXZFJrTq
bwiF0Rd6YxaPI6Pl+7R51Amh8bO0BlwAzDnE4LmOM4WgaUR2K0S22vIaaRKPVY8qb0+6t89aVhOI
qGJdcnDVu/vN1e3jxANyiho5CUZLMJBTKqhuJa+fd2fZ74d1qOj3egTYppmQbanNV8TE1E1h6YxE
6C5Hv5Oy5MwuzGjFx0pQqJ5xZmNnaCMxr3aLBmpXmf5s9ajhyC5DeP+F5x9CZbqfYG7WP/JL7+cL
QAvB/uPV5qN70Mpj2oHZe9q+qcmTUC/0MD22EW31bR8iHonTrcZzGyueiDSL2ARgyCSwBkKM3ydP
N4eKr3doJe785QLj0U6ZJDlFIt2ztABUuf3pbwti+J4EPW2nCT/AtKUsXpqVBUYObLk/zqw4jVQe
H6ouNUG4PhmF2cZ1NYAeNQhp5a+3N5/eXjiK++3iXxDqkxwXEFLAxHpTIkE0AdC1j9DPvZxHt1WG
XAdYVHIrM3VAV6H0TZHlw2t2T+kcbkrYKx34ydyNx2+5Ne0POsWT1gIhGyG0aN8U+NF+/xH8vq5D
k4wrhlAUQdvppJnDEgNXOB5OETS383ZyawDewjmcLkuB3bG2VY0H9U3QI5WPL0O6IcaFr1jJ+WYa
E/6otncr10n0Vqs3kY3vu7/sXlGGLYsXLGXYLSXqj1OVE11ykhwze3Os/HT/BTZT/U+OZsD1bY0X
EvkWpR7Ng8Nkojr33ugLDdh4kCQrm3K4hpJaIuWSllrJzBdGQs4FtSeydEMUALljtSmWQ3iKduja
Y9soExgvT0iKnhaL0NOy9fhqdGjaQ0lMmsQ5CgHDex1nj6LA/Ic1nr5sRGg085yZrDzRcAzL7nkE
HsQCxuh0fdiG909R+oxnY1Krre8tVm+5jVfJarFFNL7pPb19MCbs05AMWIzWY+Iqj11amIlaVaAQ
CKzG5obXhOT/pVYyZSGVreIrwEYO08B4nj58UVCZf0q2cYink/qkNyNjqpv3ij5fcUuXTvh+CUx8
7b9ohkdxUl6SwrBDvYs5wvFct8EuUJe4P9RlBe1N2egjMg7VekxTQxeslCxhkWaelOKk3diijCvV
DijqalIjDkejZuVa8eXhpmu2LInePH/acM2F1HjLecfnCnOtA/eOwDFgGObf7LAYTS4LKpJHX++h
0TnCu3zXmabfJz7z9IfSAfEM5MIL2tyDZQUWSiDHJiVARTzSYynaUuGV+pUioSCilZ6jONfmZ6ev
qWDwMbH4U4rusQO/Dwrf+pQAXjsihCuF86QXcAy4v97o6QcoRH/t442vtqb5In8oxiC9+UV4Jb0h
9q4JqoAV9i7conTGREd6D+bA4GRuNNuoL+MVqhcD5iepcI9j4E23SywaEqpiP+cKR4ETFMiB3afe
jMoGe/78WludK4HF2wOsKYx4xmkpE3PFKLe6Ui0/xvxFldKFebnDGN5ERrjAj9cM/Coh51YdnRnu
X9SoDNNbu53BhCLWZgH0t7T96qL2B5W5JVrOWIaVhNAdOX6hFSTMxenHlxlhfV0CwPRhec+Bv/ef
EByNTyntk013P4nTdax9EZbw7eBoaHf4sJLx1m+FZ1ZATInOui/comlz24tBPWUyzvG5qfmUDlx/
toO/6QDpZFjL9ODn1sS3uWXediLLHNXOvlqfUzSTJUzWi3m78WAQY37Blap8KO2Pm5ntUElPoo/0
HtrCRf5ZY8vpZmFjY6ZtewKxXT2hQT3eh9DEH5oFZA2Xqj/AOqHm3pm+/GF3FvjvbceioTjpEkQ2
3fFjDIGQbhAQG/VpKm0RwxLASCoz6ODorV0sTmsO8tcJquykl7/rqkZ/ANA/GQLqfMAplQo3sUmd
7xYBpxSWXtkwlTlYWbhxvN7WnxPnt7pRi3MbI4WZbeO+7l/t5EDnDyw5yBsl150pLc3nxGcs9hCc
/S3zEDhR+4zyV1Gt5IcHXkJ/O7F0BR5bvZTKQggXIpfvijQ50arLx0XZH7hLO/uHte8WvpZFQycE
br1USRwhOeYt9XoESOsnRX5BYOKYCIgwBd4lyU2DpKJJs4pT2Hmi6ytoEsV+OEciHylpskfdnH3w
WNdY2uYdoNmvJx02uf05JVzLxfS7Zud22FHE5BrDV9SiHjxvYf4NqgRLsV9C79l+NCjY3F/kaYsz
1UF/NcVqLTB5GsnArFoRyBNQ1puQCtuOcKHNsbC6RkKZ/XXeYY4m8rpHp7ZIQYqx2KUQKdd5csOX
CIMJT9crm08ZZ3tBHgD0WG83fH2vbFkDlUtZ9dGiz1waMDLcVpzzIyHU4pl1HbzcPzrIDj5FSSI2
7mK46xadTLCLq+8YiJyx+FqfnmPvI25m9ZXZhC0P4oUoqYcD3YBPJJt9yqGMil9lX6L/vbq+m0Ae
NHiUyIoJZbHgAu+Kq5WQLKplXXKSEd+ed8tporBoaEiQ0cyg3rKxXQ844jpql7RnrNuq+BNHCjDK
sTZrktGOtejIhoib/r6QN1hJSVuhJD0qg2FVyE1WBMETqz3wCHtwtBgSDMyE8D0II2jrUUReP0KE
K1KnrhLjtubLUy+hPDFwBTnefVJv7Y7dYUtEl+c8EjN4tbcps4T+mYmWd89WxB2d8Ql8CLBm4rXG
E7LuWWeHb7OPKZMZp91MzS/h3rrvk/oOoXWN9vbJYURcTA9KM/FaUyqWo18nHnDT4R7mYwuG0Ms8
r3h9QbMt/QVFsZIt+dIEkmLkXQAYjDKT9MMC9j86Gew4cZ9tI/aTvLdUWCLl3raDwrUXgxieeEO9
+hlz7+FhiDR5KgYK9zfa4dU8YTREBqu4fyf7KxJ4Tgu/YRDlZf1xKpe8wJF1bzxQnvbRBaN8PLPW
CS5aoEY4pJ+A4SivH65fADmoPSMFciHsGzP3MMZdDqvlUR/JGsBpauQ7l3nsC2+ToyqYPvWdcikm
a10zyHnxQQ9Yfx4iCSr8MFwetKZN22oRuD3okRnqI/lI05Mi+R/JAuCLp6iu3qiK/shqk33+NBLI
9VwNSVhMVaVasYnWSypjKkwrckGt1aGQXhEG22IAMoBE8KTxfQ/pF+Tt729OvSGqhEYjO5Nnpmsl
sdt8HVaxusXWeflj9PcIZ8hM9NBd9+itXdMSAYE1kDlcu8jL3M+dGqpjfDmEUWK4o6Ul/xOnhwjR
V0jeq6qJW9Oc4InbBNC9nOGwMW5HB67TDaDzIOYMh0exFr2QQZSryjCIqDmmjQM13W+D1HX2nFIx
UaCJyzzAsCfAOxosDYP8i5Q0+hB9D2nFloWKxYjwZYd6lcgi05EyXaV1H91BqSuo2UZG1tIjjJAT
zkSB3iD5SyfHfRnZZgZtFJE+v1UkoApgYh1ETG6yz6ry56GAp28WUtkjU/VjQ+6amYGLntIepL81
2TacKKV5w9XmqC50bIrvCWZkhayOmkDeOgGpJA3Xa3JeL2D22gwNy/dk1L0xer510P1FhtULaR5K
tNXzndDKYD0agvEQV+CwV2FreuR9j9fHbtsOBt+ivQPMtznEkK1eLQk5iLjLymuTILcxshLBxYIf
z7eHrNwxGo834e9jb25MDks1GzGtPP4aPH5XnZyhMfamZtoHf8ccCX9EaB3Q6LiU5Z+m3CsbaEvQ
XNMZ9bSMdJQRas5P6E1l7b4PhcRf2CdkSge8FDXn7Ux67t+nJZh1pkrIh92+ctPJRnHEE0OVfJDy
xRGVtHBZstbahXMPkgpHw8+k6+RtTBAzUqa9T65WbjIPQjgayLobby/EqxNXEzZdIoxGhX5FJ3K6
rO/poItEVcshyO9N11XIFFpZeIQz/gCYmtoz4wGxr2yJwNCqj1cmCH4mENG+O6QRbbfUGtTDcyCn
25QDHdp6HCpG7Y7gw0FEUvcCvdt9Dna8pRxzmmJJCUC57s4MbUjWUxrM9DmG+iX9hunGXF/3Ymyj
xZ+GhdNCc5a40DN59og/2sN/yR/+UTlWjEUQh9pT9uaN2TSYLwwCz/v3/9G8D5qFdjAeGgdyoqcU
HKkDMZXIcEocWv2cYNlsJWKWl0pTXbJ5LXV3FMveU9ksrNlxfBGsmZvNyjE+Nuibb8YCG6wyKKoY
ooHAesrKBJ6az5McIi2gYY3Fc6wUtj4ETGVuA9pNfvuVMafLEy58LEh8gMSyH4DsSz8pQq1fyM3+
9w7x8vMdsVeG/WH19KOlvljdEXJyKvQQ+E6PCofa9nZPBfOcKa2oKAyq6Qxz1z8/Ff4jGsUp00tR
fTJVIdXJ64oqwR0yOfdgdQw2/DcmI6kUU9K09/rj3dhqnXcozHKve13cPFtW6hq7znfHdAwabHeT
hE9BzY+drBLgL2XSoPPMptbdIrYRmSIfMHm7bYC8xbCQPbKyuEwMZDMw0hJbnhB7uL0Zh0e+0Tp0
+ok8Uh4hvZ6rPk4A30bm5kDxYztDUXKhGYtRjwCapX0UQvwWFtuM+e90WcGfQXaZ0cCZ6IqPGHP8
5cAJLRsdN0lv6mM96Eip4rP6Xa6YIQK7QXOmR6DolsPZkn0vz90pOi/GJWRaVNcCfNdu9wYeFtCH
o7HeOWsa/3hHl8gYvnVDC4/pUYhQHzKGMibUxTE45WUAMzGgzU2CrzWr16faWy9rdGUMN4myol+g
qmUDehf6T+YtE/HzyAss/7jEAd2qwU+iCA7TARo1CXPGHt/ND0sQhm16UrOZHF2HDJOFfZUEFMJm
WXBjVkQk9aAAoRnhZMKUwKVVtSgbyxruTG8t9p1hHeh/vF+GgYUOFsy5K51qHEdCIfTZnAn5xfq2
Y057A1YUy3/aksJUFo9HY/p5ortbmfwzxq05l32GsZk8ETnWGK4SN/8we+qwmAQ1TwoxEf8n2Pk9
phMtFNqLHH978ZUSC3/0ziD6SK7EZskhrUBxc6RBLiHe9j2X3q70ZEN5JrQT5vhIOgldsTo92yNb
f0ZtDDpKPvS3G+Yxfn+ixHR1gcoeizW9qjAJDmCAq7LCoyHiPDv9k5quUhxsBsJyETAMW8Qrc9r+
CsZWyf1H8G+Wn06YFJmHefl3e+TO3/NMl2dWk5P3VIRIV+81fn9I8Jm6A41fjPP+9aq+Y+HsbshE
MXmTLctQiwpyZt1GVDATxtG9Bie/rn8DHrlHSyXvNnZZzUNSB1ENJf+L/ITwcTNWfHJW9GssxJ1I
umPrqVZwcRbnuDEL6uQhX+/H4qgndfCSAG5mc6Tuox4zRR9//F255C6BHisbF7RFTNLaOqBZ9MzC
ZoKIHcoBFskovqZH5BVfauciF6f/eAPK0PQEWIimTPns4+nfUq/QOcycWGAaqdp0dVr63p6j4N12
Z3O/Gqu3tSUVUaQG8tCqOXRrv8mz+EDR9wAT0HGOPNW0+VTjYfYzYlw9kZ0lWYiGOlgT/oR8D6c+
GnIjrFEt202HlULcIbVOt+UXHUdoerAzxFX7TLGuNhiQVVhi0TMyDdz1HolsoDajDvUI8ghvFU7G
SoJ5oisQzvv9sHUl3a1m2j+KEi6Ombz9FNp01A9GORd/15fL70kgmplptOP02E6OnJfRx9p5PXBW
yzByiDcTgYqB+iv5roRwDI/N+r7uGgSjCEAuj0J7rETQd4hjYxGwpkVUVKWSAGIcRwtEqRfebLIu
HkYrc7ipR9Dq/YIbzqQ+Mb+rPrAqymbAjzbyS8URC5ijEVAqcQ3ydhTngTixm/syNHPzEIwJujhW
DcpWAF5hVyvmkO5qH/387iB6i0Nu3eCtEUHbz+hkXoQuPZ61QOOb50LnLBmYWTXQikjEj2qpBHc3
la4te8Og4LKfzWT68Z6NXqQ684XQQjf7kAvQM/q544rzteUXHayqg0mpONwd04qpd29irc1ZClud
RIhxHeM3FacCMvJB/IVMjavKRtmc8weq4366z2ZOguWBq79XJuAYY77Bg66+EL2a2D/cbvZPGhBw
GxWRp3S4YTyo/GxvmQWa6oz3omwQ6oQVZhrmslib11+opcQRrYC5DUBcSDnWKSRDuSvCGgbhR1Ns
0DxEElJ/kkfl7v7UJEKSR6HKOZdOgfXQIxLvUwpm7cTRsPOaDZtBW8JY0v5hbaPaW3S2dhz9LEao
CsKeFFqYzz7V1ySCj+Xes6XemeBCqKyiO2AHXIugAtwuR0AYxaMJIjkOW8zadpjcqsKd7Ao09AUv
ZUY7ENHT/wlfu3jBuhyjVRuBcu95eq1Nm5/Ub63KntlCWYzKE97gqxTKjlFHd6jXXQBNxrhdCu7L
F3cstboUVvIuaRt+FhLSa68+nvRR2Gqz4n6wLQ/37DWiq0YeMN7GHHfl/hr5DvUSzfwagwAiFWdu
VrddqHpb2te3iangzAO8Un3QTKIIJpQAMpFIGwgXgOTT5ouuMWf0KisRIH1fYKCqwIKXdC85N0uQ
c4opDbQhYYTZMkrEC3EcZ2+SVvTdXgiTjfYqDtJTxyDt0omHplbhNf0y6FE0JTDOcS6hy9vk+xur
7fc6EsBHgg16lks57WlJfxNAztpGdK67xZWGFGePPFm3hcTx/1KP2PcJg6MLZjQtvn3H2CNABqDx
ZBFMMZb+hTKtjLfU3G4r20G3Bt6r7Bb3fxvUEWJwuFZ6/Fo2f0W4vVWppMb5vblCnMjTJrxmtdkH
c5Ead30CdXb83204nUVtFiZtOEJczjU8Zf4XIVoAPc9P+yCJhmgpMk7qhyL6q5eVyj8lVYyhB4Yp
ApxgVX1rcZiRshLtZBofEM7yyccnIAY+rXjEGavTuxoUjpw9EXvolPfJZcbn1e7oOQVZ8KfqDTAd
pj6LVljRULj03rGEVJTqerJ0nzU/bnklixk1bJlVSMQ1gX6rSVbGq5qL2Xa6bbGj+JELCwPQB56z
f8B6niDROmrYWf7f1c38uW1YWv29drtu1Gph0EsydYwHTLpslp4GJFUWUvui3ZKSAapKlmM7Ztfk
53z2k374rxbbaMFIH57l4hvvC/vlYPh0+qFQgxY++9VB8CzciMAK4+VD0bZre3doq8fiULQczxYc
wkGzGw6ZBhxX79A6/G/Iv9iB8BQ+GPRBphiqLw+6SE6CqWlCMe4cXVh7EsrbZo4BGB7gcuB/aaM/
jV9nhIQdAHsi+FVNcaq59D9j45LaDl80LOSwiBklHgH99+WAP0Yo0To/idqAbqCRUAfcyP8vWzD+
3gkDlxQCdsNYTrlVsIIzvkeUxAxS1f/HlkpMuBwCRssj9wIP+4PyUZ97Zr/00E1P61TJXBaGTL0u
W0yYoLCqKx+jGhFbV5oveHiMCUXl8W7JUFbTz/dTZh5nunTJ0kfuPNG7DZmaf15CSOTRkmPJ+jhh
lLh8An3MJcqLDSY7PhIxjx3bYKpFNLQBvOl95BzJ5O31FPiPFohl92b0yjYjaoAKdqEZofZRKA/H
8Q8Qi7r5hfz13+QGY/TDJIl6FeAJwqovMvgg4YIlIW4Yc9JFuSDoqExQfFAysqbJo4YdX51gIQZD
I6PHiziPQxUu/aZXt1d7Dul9HeYwtcF2wSiduigiXlxi+8LfRmANVnv42gSkNvPVsDOZBnN67qw3
vD6ArsR0bW6Dp9DbMBafddUdzm+QXO0DgjoGgqUL5R4frCdF5Tf/C/qcFeyvcgqU8X2dgo0s49jL
k566qf7hRGeQs+WZ1QFZWD2fR+Qe0ztgJaMb0FV5zZVbhPhCws4S+AD0TNNcmxzIfaPaa6X9TDdO
tiS3ohtKtFInxWpphkwDRQzAfmg9eaxyV5i5z5zLF0OSgbHichELJ6rjDHovcBdr9xWDSHESF/n3
uuk8NLFCYW07OA2SPnAFgFmikzEP03xBCwq5MCW3qoatMi7/6Nt2FCLxZmpUIy60tEu71j6E9XWf
cu2dOSP5nj7B6AjQaOyMlRR2P2qyNBrHfXOYlrEk59OZqWlvvAL59DBPDDbNAA2LYzfIOYVzlgyR
RlP9ji9P+3PoC5UYws37AN4PwdIIq/vfwEDqSKl7qKxb1w8Smxxq2A8tNskwAVrOgK5TcuPy0s+E
yspVebToMmGre4oLifrrtSbyEKIE3gGycLaf/0THS6aRewKeHVFuYtbAm0rYGeosl0NAJoy/QmP7
V70bVGR3d1BFvBTd0CuB5H5JJ8d3rta66YYIGIL+bTf0FlBRWAOM8WXCiIpufBf/ZA9X1h41xNeL
squ9m5Cwj/yVdmdTvN4IOhgKKYFQ74syGX43KK4f8OzgyRopYg5ZQigzN0+64LTq4RgFQwB2TiPm
kxTRaUICq2DO62bxFrg9eaiPlhUs7wwvgMWfbiCSU+xdCCA9axhedtNlvWKRRnyb5pcuFnAdNDS1
jz+kZm1+gXrkA+7e4LX3vcOrnU5pEYPUkW6fSSJ+V20K4p3KmjqKWfzFwgSDq/xeqf2HS0t4Ac7l
QB7mcsq3Q873XBNjubFu1n69mMiAYkv1uTFSKoaFJMd/mTgaEjMVQGTTaFA+z9UoQMinSi04qoxT
0xsw/KShs5wwEJpK0f36/yCIPl/g7mwOZu0BsGrW4ttBi16z3KFEQ0/NJUXJoNXvv0QSLwyDKERX
U5wRs3hN+W0h88Yzv9vLg3hy6HZUyn7IPDyS2/MBtzrd3x+1QvpUIMaR59X2bBCowF7FJGdVrMdo
i8TjKU+b8jyY1ci/b62MMTdwmH9cKtgBx/wCoGHB7G1A6v681iRh6IHS+MapuJrwLrUqMqXm+UUA
pNEMjKCyaKpQdBpDwnxMvyousrP2JwA401cC+rZSjryLIsVChuuqDUllKloYyW0zsDAuUgtRh9RB
ZQuxEWQkwcTol1KXtTYgm/u1UeIzt5JxHNlAo09H4i/ckZr9RuYH7se/6D5MPGf6xbVZdNNoi0xw
tS5fku3ZI2ATg2hByI5PZgbjlkPPp/Orp79eqis75FNfxYnk6u2GUxdliVvHexq4oxET84fA8weH
9EA4Wg5tu6U9wKQ8d/kvmYLTraCd+mWyzGqYHd3q+JWGrLWQ+MP4t67N3SaYb5KfblR+3niXEIhu
HigLt6JyQeH4jrSXlzGR8n2UDPz4XikkbjtiPdM4f1E3+IUqbKnYRiudPbJgYcQlVpDJ6yYax2Kw
aBVlOJa9O0bie/U84gZuUujjneTNqESFQUjFLqKluXF+DFSxdDhYhJ+LpapManJYG6b3oLBZCrH5
lyBlDkZVtN3GwpbCem+1eNj6FK6/2Eoy2GO1ruDCdiPtdhgY645atwu8MOExptwGsJNM1hMmkJDF
P28AIdiGOyXY134qT7Gs8syW191geGDl60iPWqkcvWdAcJ8xHe1jKGxDl5zMc/dM23NG3DoB8405
cnOj+vhZKrtVY2CooojiuQS2rWNZIVgJ2c28BZNsXCnx/r8Gj6u9K1GuIorcKUTF58DAimKcXTm9
wQJY0bxtzLCMU6cuOBxF6VSxvrfkj6oDukw51aISdKxxyqs+yXQFpvTq5I60ysj5saK5rjZJscIU
2LybuOOz0/pRPnw2Ac4VltSwK10QU3o6vMenZPIRd11QhijP6XjIPLIjTBoC0g33hF5CY8tUVVd5
u3xVd69LihGaATmlgcbfy59k76m8HW+OrQvrOWIXbA3+9in3MXXJJ7VjwQx4pZtTuxkvFYGCKwm1
63xAPVy2E27Y/u9QzDB8iMGIrLimlpdhesgXhc2pNxhHX5BYaVs4qrk5g+hu0D/WD8GypSsWkTs8
25AA4hUIruukdbv/KFJpkIcFWCRGTmk9o0ITXRWrmBR0LdqhET3/upRw5yMYnQxvAHKBuV+F5il6
WPpqOv0Xr91t3I77KSuRdFzyOmigArGqXyCrNWpIv5NC8BYTFnpQbTZWVZ4XbBhYOCD+ul0O+/+P
I0+5Hw1wd4NZanx3JDe+P51PHXjFJGTccQ77OznS6umSjuHtbAWtsROa3+QZZlV25m0CCv82zekA
GbDsisUE5KxSScwQfIHPaK/dKNYUGNO3aa6otOo3TltBs1cgSBy7AAnw73Ma0Kz5Juxj0tvxWJmw
/rQUc5CQM9b5ElqnhgQ/NKaU7tTqB5earpwSqBMWaE2IYMdXVqUAskyDRGZigjcHY9O/c53aGeDB
ujn3pUFW8BVGqelf+ncYfW9ndZmVPZH6zjE5RhUuaH4yqOF3BW7bi7bZ07GWbQEECLT2Opfwcz7W
l2MlNDexir5CVqoWYcCZ3cT2ZpbW/XLnCMVtZxdaByqC//xVn+uxH9K/aTFtLruqTzfd8zrzT36C
4/9E4Ztiz5SLIDl1dUumvwRD/G3d2aUrvjmirFaDl1Jf+lX5ZnttiXPsHl4JeD0CtiWxcM2NE0eu
KDerCXFKxYnxd5C2TeWKkhr9Q2xHTTSRjP88uaUz5EbRtCcCQb5SHQjv0yI5R1PHeZsYxZMW5qtP
UheGUkTr4z1xkgkM5w8vE1APgD/g7SQpeI7+WBTZFpl2kDFnw4AOhPPev4pW1pHSq6envjHofPp+
0SUoM04xJ8MwImZ0NIdotOJd3jCCk76KWfgS5/XteXgoFEQKeo+GBxOPuEvSypKdqJ0sCYxzbWTE
YXjbCpG0jv4wX4u9BLpKUR0JY42S0UtATn9AqUKv/wZ2FYPSF5fC9StcpOlQba9RzQQEgakiBSVR
W5I/eTE2Y4+1nmx4hKY8+yZNc2YkoyaDHLIDNCONYkB0EHot+HboHfFYl1Nb/dbHEGsGRyUNzH8V
vHmXPY8v8k28PNAIhtib3LcRSKyLjLgf9mh1r57/0kZhzKu6T1Jz2Wc1ouNyBTa4tGqiJXTR01OF
zuUaV2GPGXvrXciccZa/bVlLq1C9UMfyX42r3TivLKC5J2BnJIwaEx7o/Nxfut4op/JCjp8OOB5J
AQQb1FGN9E5kM2+DE8QRTSmvmWNFgS3pX1DMNWW+dVakS3v3AHTqW8PWZhATpjdS95lUltQMM3Oy
05medQgPOiTdqsvCtEYJiBhUoRG+NJC+pL69UiME2fq8/O8O/+ty/7ynJiyZG7J2o7WbCVCmV87N
NOeDVamHzJFl4T289aBBpuo0Pzky7VTeLs4Z2/XQrp4gCgB/OSKSOuwwVzXVz81olulngDv2m4MB
RTRM2lR8hLq/e00tJGdvbGlYJ0ymJekDKgJDQ8EFCjTM0sJIACPa7waee/ZVvA1OFjas3HNEofpZ
1RPjiyZcJbWvyHcy1qN7O5RPSWzRlgATtHC8PSGRWshez5GMeJryGZ0R5k4qPNllI4Xf7YmtpI9J
qUOXJGhfbigv4S0jSQV9zOr4EyuD0F3wREbn1/Yc3dzDh4VwVmsjeYCPgZQpV/rdJST1GoCcycwi
INjh972kBDdKEQ8jb3FuVz3js9RX2Xh7uWHhrrgzG7wg9KdvrIbP/58SJyHaeNE3vup7p0aZFMng
opz8M90PPo0ejb+bDkv7GqqhbJH2BqTZSxsrBhuV+OWCl17V9DMgwgSnyhtOeVC5IgLFm6NavGh0
xAKRJKiD7du1oBsK9WUWSy5B00DT732nuggGWboCvkbbyNEAiUdci5mePogpfWMaBFYoJeMIK7B+
4Us0lmGvcDWuIdbgUhCrGceaIVv189/2nN/xr1uJssIgqBvXSA2oMn+m7gacXDHO96ZlooVeYu4V
R4xf/ZBSBJNAzKohDQ25LM1SzqLVIzU6fW03W58UR5nhV/CeQH2GfkMqWIkLnO7ASjWzTdTUz9wE
EwhXUWrngrqFTbVz2/p+exG6O1cyt46Q6CeSyVVKLZA5hO1AiyH9log4QIac/HyU/TLtFT/n15ju
IiG0abcbHHQG9TsLWyWCGugL+zD0DAhbVydtdcpapIK1t3GcRJ5MSZ6GKyipoG5FQvZhjlWgCziX
RtNeEAr2l8PBr2XL4H4m14acap+LZZJNTxr8gIhgrGS0EujOMQwTm/wK+EIhYaaKWKKUemn6J7oo
v46uGutMoYzpYtWik9RTag/AC/MrF1j1Ie99r9gSiWyk6vamvLYPGyyilCpCE0CN8cVlfnnFklSK
4SdrSPuTmrlUImZ96AE7P+7s4fXRGatGfOqbcoBVOwlQResR/KYocoOJ0BJnuHTsC0dQFLWxPp8F
3WGYCskAHt8AW/lEOHIoDz+LJZ6qhmNiLZaSInV2X6fbI59o2EMOVJeEV/GfOFBaEg4i+2jVN8KM
8oKS5vpQkXz2u84pmBSTiseABXp/FDLUVou1HsMNA5q51+nIkgj4luNPWciWtI5kUOBlNoSV0wPJ
OjQ8qA838uKmRtJKF/SgBLbVCL+fug1QKwoutGmlIfNshMkUiUyawEnjnODMuf4YG0LJTalcQeMf
/lGReSHukmVscKKdhsZDS5EdTBx6X9lKbDPC34SHp7W6T1vJsS9AeoA5I0RWWVdN8kaL2nk6P6tr
ioak6pomUmMgU10ceKJhQZiZOwsGrx7duKgoX80qOyiPOuKeJ2ZjOdJbngSk4dJlIutc3Y+A7sy3
iwI/1Lfi34oI1DgrhQp1J0PmIG2r855F09NcfO7dZ7ZkOvdKw4JJO+XRHPwusPWfx2xpHBGYyiQE
kZOVeQGUVK+EYfUbqLQVQFH7DOZTSjVLWjgiEYqxHyVaGYgLrmKyXiyQUj1J9dQn9DpLsWKLT+4g
j9lYRXWPIHHheHBfTkAjlUdNVYs8eFW/EYzuXhWMjrjL9k+ixOquAFnHxtsmY9SzaaUkgn2iNa6o
GpTbtnw8cht0csN22iwyiVLl1tsAQUw/8aAQGk7OLa4UuFqNHLi6nfgtu7gAHuMYdoCg/VMFADlv
mX7t8/7H5mNPAbhY46y347I0ztVRtcTWtbzFMifFTRF6M8iVDl8/Vq6zdPAEO4Jp+d2rvKW2Lypi
S8vCa8yhHVFiYcqvt+1A8EWA//PdnE/Ygosz0DDS99T/5OktAqsNwJCCWAV+hK/jTrnEWTmlsG82
EWR3sgBBzi+kpTBze7l1v+sCJTimKaF1hcouwuov+Y7lVM+EpmSNM0uKkgHv0jMMZwkgPyXhfu9e
MX3lC0M28lJBHikz8huSTpK4Rh7eVXLs/bQnfKCkRGgDm6bdtp6KEuVtoYN+tBTyjPowj5ZkJstp
h0dQdpS+DlY4/nDMOWP9cWhSJMMCedEHJRYV3nWGoDqIUKTdew5m2ud3jKA3ayV/vo7xRBdsb8xB
iLpEDOpSDW9OZap4sfm98GaGOZmY49EL5S3nnCERWienDEngwCSxSj+YdBcHsPzrZMDiRwUDw2m+
E5J42CqWkTfqLRoasPnsb8dyX1vELREVrmTtfTakLcjmj4rQg6GC6NesJD10q07uW4mN0LzK/FLJ
SyOgRBevLMipTSD7lXLsXOVPN3nRd+EHy1j/ie7Hs1KjTX9J32yU0tNkut/FYgfz/90Kdiy/Ycey
GusIRFl9FlCKIMN9tq2vz+WWjBTAiS7SjKLxWQW2BBLT/my7+xTfbOtuKge9v6xUBmBrjNtfJdKN
N5F4nDV6+tmbsepAGaOggY2nS2sEZ8Rc1xa7QDMWArdWh4D8Nik3zXjhzsZNpiurWM4eDLc3SvBQ
EdBR96HY8zwp73Cs8N9gyuBikbjPjh+ogXt55NDuCTj69tAPZ4WEDlQJyryckprTiKU1RzNw8cUO
P1AJZ1KYznMAu/nOQE55B54zfTA4bp2GfHY4Kcxh/qIzI5zpT9xB/E2nNrQoT5x3KhNMeMywl7ET
jKT+2XNvfdBieFgqkQ0ecZoyEa1nQhjWaX3sWDIl4O1ZC8yeWpNvEP+82K8mFNXKNLRiUmnfIbF7
/ZA+5+dDSLVPrWOqWhsm0U0bHFMtdOGS/vo2p0ZnWWmPLWXLwO2PqEL7xvPk2tga7uDec3PBE+78
LQPq19ge9lyfRRo19mPGL/4NjZ0yVZeBPDCzRWSZF0DPyfKPn0yqXwgq3tKHrW4XRd6Ut5DZKVfD
Kf4/EZtXIXrI7C+DZLzRxPY/hSbhPtH50j+32cEzXl8uu3ZIYeyLWnUAvjatqHjzgyIHpFuYlGLu
ImlW8wTVRZcEskaO0e57YTgnaToZcJNPio7xU/IDDd94+3Jq0lxO0QG1qEsNMOo4ZIMazOh9jWFz
ctlpd/s5FvYjUgeu3y4/yFf3YkHxQXI+7ckkUtxPYCxABdR/y6LHmVgbBfYpJTCp4AQfRzv3oI+p
8/ifIh71X4k4LPSwmMef3negHKQIqYnoJv+tgU1txWLCOAV6goFAnrwJFVia8e3fpKTmb35MFUfb
uYrDq7OC5GjT13HbZsS1wSD1p44M7vsS04Dct1XswhTpVKMn5CLz6xh89rEvz9wVxNsYZ3FxSq0A
ijjBSZVeEZevXG+f8B1ArpdUNj3uWE9eOcocaghZK0FaaFrOF1vXoAiawJZPL0eSVeLpibEF/jC1
Pj0aXLKlLio+p9Lt/vwGwZVEEpF8NSksXgJGGfu4V6yu6/mNl7LdCtVdW8HDnVpZb5MgI3kwtBDT
UBOckmI4TC1BWiKsPjrGdO9cGIbEF9UF47GGlzf5hjtyi9eyZ7l6TnAzyHDgpFExYNoGYbvZ5/iZ
gdKl6zAkDDClO/qAIVkhtlNHDAzdhO3wo+Uea58/pN9kf5gtq5vOsjy9suGXWxQs7jEQmagilNtf
fX2lJiZbtE9JKrot6Y0tcgnPPFmlu4P2t7vASQcSrlKvYtFXpWw5KQqQazmd+IZnSpD8QpBTQdXD
wLzEd+0t7nMtAkWmq03jWEWF8J926dSx4GBFocDK4KGPfDEWjjS0LxTZSQ2BywEtXAI71UXIB32K
EoWiP5sHItaqcHdq+WSwPE/LgTlE5Y+noagMo16nauMKVuxTWjvme/6wzIvL3StdsOKzdMyfRY45
st6RRleaOT1lHujjbKSBMCZw+vyqNDNIfFmm5I2R579SjUYBXlUtiYHocyTGaUbde+g9k4KP2/PY
cAYvIBeLe/AwlkuS/uzxvnv2fXHijFZVIxbwdH4FpAaWIMYf/2BJKKn3yYxl7SNzd/Wtgy/Zv4sN
v7e8cMusVlmScM5x94R+MekdGaTjXitUkocZSy/aESDZ1lHm/5GAk916jphEwEaBLHiRrTITmHmr
GA/flQZAJMAg3Ja4rRsa1dH3O6QekuQsdpdcw2/I+dNcr4JDwKwY15MNZ9sGCtha9lqrPkM8Q19e
blF0BafKnq5d3FF3X0adDI5C4gXXGwIbtloy4i4pT1V6m1WCWmHU+D+5/Q9ol9XzR/fvL/APexKg
Y1uHvOEWF4Zc2VE74cXJpQBHENVMMzWsu+zqG1U+b32MvxBMaSEfax3bSu+uW9PWYAWrlyrVP2xh
6m7B5vYlRpoikad5v8wyEpRKnGds0Boz5s9+qCfMKGqRKsvt3aRuavdZYimF/IorO79zsBASsKKh
NG5RrAPXUlIc9O7+0rj5lcw67w2FX1CV1u+kkHM/kUr0emJQm4PYd/0uxdgzG5QXdJcC2vCyTIaN
Kpw8JMO1ggY68BlXKlGjOnibgN90CeFw70CRjXO7HMjgodu7DsME9YsIFO4b4MglGjh0A4diiACx
heHTaX+gr5uxzDykFIMMacEhZoh3HOS/TsDBttR+TMhnNDSEkyrmxK1+2bVTEzIcmBFGJC2YT+sB
6JrCbibILpXh6JZ7O6zQmk5at+aQGcWZpQMt7VqJ8+P6l7QGSRHcP0/ntF8xIhDIq48enOpR5hX/
le0fAkE+4s/6ajhDt5KGMhcViFraC9LreAPl0gYxtbcYEmWrrQyC/HxfKX6R5WveZmwfB2GK/JRl
qv+T/EJMX/3WWCHVr51s0iB7Idyxuf2iPgrY8SAgs41BfX6j1EDlxpiVzSlpKk7RMnb/PtX9F7IR
FX33hrcv9zfa4hHQ/5PXQeOzhp5kHzk5gjByXxavoMmT9PcBRm3zea+iKPsXeQTV7bzeWbvfItoH
VfNO996ine3OH4uEnJLgbOP7f4K56o3CUJqUocQNjW003zPV2+2Z6Ss71zXklha7fILIs8JyD9un
kvNTHIkZesJj+QYl9ttkHLWYKV+xVzJ5J7og0S0F+WYt50JsIY1OkxwY+g5CsLmKreESTdhREKjW
UUMQ2+Q221m3dq2jB4MiMOQQHojjLRN+8RkdSGFZXjsrnW+dbPdgFAbff+uPgxwH+icp1qttYlKS
TTmlJljTHYgyIpFz5rI+xf9H9Xg7Lk4R3c6ZsjbbcjAVvfo2kye5EddMLjA9Sq7eqKmVEAahIlqN
W4b2GYFQ15NBj8FnU8yr7BrGkYX3VLBDzWRMBBx9RyFWCmfD1RU6/F+QJqOcnm3Xk9PKPb64LtlB
UGK1DFMTHe8EWavgmBPkVuwcCjaPYXCiBhLdHkRJd7JmEN3xRMoz3sQIbRAtvmU7q3YfDCZMLe90
zIBT0np4V08DEeHKMYAwjE6Rjcnj4lX0RM05giycur2P1eKOd1R/akayFcCS67HeRe0KBdJEiqEK
jNLFItpq9MIzwkRZXLUdm5ZkeVaqdUpV0nOe0w3YEXtYZ0jORqadGv8U1lUdnqdLv+z543Uwc+qv
k3GeTgid4mSvV3BxdLxyu6Zo7t60I23+3PCrpPGVFLF4eI48y8YFEHhKMUc+cTsHSd6JSsEVOaPC
aHYtPbGpJmEqyxJ6jAow5bjwDdDwhfunJW2on3W+xmFdcoe0KWIEvT/2WtZaH+l1x66ufl0bincB
dwzGowNYKQxfj1GXv2c93ezn6RGXn13+LyeBX2cRzlhdL5WsUGKlrGJKEZslDCOoqLtBvssqlLmz
ODO1GEEDvLPYhQ00QUB64mQClGmJfiNNx5zlRKY5JDf1kwutM4rfvdP0kwslNP901QBY8jNVuKAP
aHwPNMYlCvdIENiPNOgR3Tr4JSY0f2PqDhS4Dz2vLJDkS72DsEeHCp2HRR8oBFmrLZjWqHGt0EN0
hj3eI8hLoifPvGpM5mmWX/iaN71v7zRrYnDZSfKSR1Kp2VZRgAG9LKVOAvCud4nq9sCodUjLZv23
E+ErvMF48z4LZYdVecIrPOMQ9bJ7Ty9tWpmokI/JYD21a5tGjCYKP7lT4aLeo5MPrjHUnAz/Wuhw
mcl+4FkhP12AKNLtPsdAdpnG2/bua67CszYiRrVSXr0xGzoFUv46OllxCjl9I/+FVsbxY16xaufg
l+UxpN7oEtiO01tb5JVmiOPv09liPvB77IiuG3kW7WBiP9vq8amVOJ5vJg3i7hlQkWkr6VYKX+Tk
GWSkQYDizMPK3JFpHnz6vi4asu5M5g3wIYNZhe+bNUdvOYg2ePuC0ReRJp95+otcBjNQIRyNxm1D
9gN/H3ES3XEfN3ALuyRuDHkyD0YELFoduTmLM2kbYJ5VELcSxKvZdpJCcwQaUlAQ5Vqd54zuy3W7
E3f258Ns3U1XAwqF51Enp0C1dQInzTEoMa6e4V7SNYJThjN0Soc0aDLD7BfBzxVdmRK87b5Q005k
ejYLpiwTAHYhPPIAwqTZ5Id1qQLnvEyl4yJgHszNNRsByOydRlU2eykyPLW7MoudxkgiIGZl83wI
HQFjgkNEegyNOYCRGXWMwjb495IfS7VBuxBG6KitCpEzo+QaJGal/sQdOBCN+jP5BHw1AOzEodid
2XRoOe0OoSbuM+s5qJe5Z6lRE0tDrIjKnz+2W3yAgFRzPMfrx8Sk8i56HLpSanJiow1JutmClk2A
Cd+iQDYn3NexTthsGReVWolubEO25rkW13hjMPWXIZBqd1vOTr66RM0V7AEEC3EIIQTBQiTcMa8z
d09r8kj/uzwLqX70c3pCZJ62sR/QwpBVP4sLEcrrrhRz/Q0ZZywFzpS0BQgZAsK0WMasgfR2tPI0
NTdgjVLo/HGB7E6UWF0YYUdpUb5fuZrBN8v8pdwEBRZpscQL1uCAXbEKKmqARIKcYeH1UuTX2iSS
SA+3NI0x8+6raWOxdT1kRveaDV3b402TfBS6gyJQC0joNj0OAnZ3F0kzXg3noPa+OZCFMuhMa9Y8
tqEDrF6SM3g9y/u5iwGDIRKzDqL1T+mT4xwct/8bvpmVc/GjMYvlm5qdVYR0H82BGZBF3TWS5nLL
6pEhc1NqQZBBG75qGNvX+O9AcQuuu5EQ5kAC86fTRLRbA8rN8CCi8ax8JpadslisxfVO76sGH42G
92l8V0jrK/5Htiwr4bW4qHCkIjxi5KgJ/UnADZXIlaeV0j6HRc11ha8etTycpLukzUsF4wx04IS+
Xe8gE6kq1zEE07Uzi0COhP354KjzzikdZKN7PbfLIKcUBeo6OejilU1VGQ0JqnfnIYTOEZPRn4Eu
LlrLBmKx9XhUKqrFquJCrEu/BPb5uS+RQspGkX6lx1Yli+RTmeDViO4PFn/6o/FWUxPxX3m4ZC2I
K9QaPteH1bZGkZPTy1SE+d50HXKiQm7rj/e0+4QI7t2aFJfjbdA6VpmaVfnv0HKQnKZ+AT2ndReX
MjS6HpESy355pIQQ+yLVZlgr0ccbhM866EAvaTVIMqTb8vzkwjZuTWlgHVuENu1RHmOWVxPBVX5Y
Y6C6YvNDCxiaMfMdWmLHZt61x2+YLtt3j3fgq32vyhGifl/HI8sKRl2JLDNEXlCjoZ+kuVOye1Eu
xOqZtY2W3uJXd3J0xLbvLPnZUn5ZfHojTj11ZyGpXX/dJZHNM+4Y1fPhRMPJjvy/1cm9b8YUpNKh
1J7NcAmOFBxClPEiu2Bi4GpIjgTDTktr7P9mk1/mIfaI/ovoseuZU76/srSfZUhFOsJ7pXKEACQZ
VF1iIi9ql0Tu6HihQh/Pe4QQfCt+Blt+7XTIlt3YUFod4GupL3LODdHBeA88IJE5VzJzBujkUdCw
C6ADuF87TzbFEBvplWArrkLga4PriIfgT+bOu0TpYaKISwROpHUx1tpjkS76dL8GgDnpoKOFXVAl
/lRGnnq36E0FVONfDwlc2Di4HQWgJA/8VrBbwwwxSWjoQJiVzl9EhDFSTmQDVvYYGSEzMTPDX+nk
rfOaRlJYHdHXfiqfuZuILkINFQ4d6uvL+ZVD8nrJWE1mE0OAHrg39Lo8In33mddhQv6uhj6Qviyf
YgMpmhlPE8oln0+urP3LRanX26jkpKejcquYwJTU9Rr06S1aamkoAERimaNHqoqnm3Fq2Jej4919
XBaeE/bQ0iaGpsNC7rpRN6erOrxiW1iiBq8veqcESjwiwdZKT38uFpuDEOtuW51C2AvcnfOf9W9T
Kq1rleaiPeXES4UaxfjsqC+OBX1l610/4ZdLtJqhmjSYP2ZXgCl8DvwbGMjMqzZLf6s7J096IIsF
NYCGWetu8rr2lRWDV4pc/AtqqwTcg4cr3p3Gu20ybZeeJ1iway+6SFqIg2n0U9JjTxwUx5ZwAHWm
+opsGarcnRUW9i47NbXlAMl7dIleO280UiRW+khB2j50ZUa8MOhb1q08Q0YOi8VL0J984TCLbjAK
h69LptBw8JHjQEuGuxDHNrl+UkRF4ihD4c8o1VmUE6rtR/5D+k0G5az/Y7uwoqgXLx/7FbXFZjNX
xjOXUElSQDcKIB7pdt7lD4k4GCPh1ZmaJzEU5pzpkxlBHKEdLj3/pAwfEIYWJ2EIP0PMQifK+mq+
RV8wBTE2QIHs/LZtb6iZ6TgZ1TU0TiSYc3fiFzc8ackt3yjFSIeLsAw7/GOYr4vxVPRQ0JOn72De
B24lDwuk+SnHWzLtSdIC/mheQue0ONeHQOIq4qn/SrwIY4ZsIuOTffD6v9RK3rvJK3yyB59xwwBd
XYQWBZyG3YxSRkTQkLyZ60FPNZ/OYDFy9ZI4Foj5o9Fy8IoEKUmMsvUIfkOD+0SD0rLo6hDTmIpi
Vj6ERmoX9UsQ6icmDONY6AyoCAM5IHfbWgR4dluXe9XuvGC6RKRyym2pA/6TFqWWlVViT8rRgbA7
5GALblMrShV79MVjL0pbFtRxG6QbPb5KSvWlPnMU+S9iVskfX0YNAYttBWCcW5GXYn34fIVKt/J9
kvFE8KKpnfjegEmTFACADeqO22rR8NAeWaNfsqTJd3iL54m9H37cxHB1nW0RcHU1nVEHBPICeZ8z
H8eZ3ClXp/zcZenJZLU4K3z4Fny4lDj7iwqtqP2CVwtcZs6j+2Hkc23KSm0EvgdCrsamWyC85ISJ
PbG/yNgwucRiZSUvESA282B7gQWbdBUGCHc29q6qyq3cd6DQEaFNoo2kf4Ou2fGKqwHaIta2+ZP7
nCdsH3WmU37kBGnvwNtbnMBBKi1Fwb1nPNAfbPZJjjGnAyiggWtOWFEBnCbJF9lIb1WUv1B9heax
zF3JH9hwGHW6ZMPqmP5TASrW671xhrulRYKqVxbqqTrnUDw1w+TcVHYyKN3NiTKTmIiDJhXmEsf1
NgLsHiGys+faXdoSsj6lboxGKTEd9YYiOTEe/As67sEm6VtlNUoI1JsUNBfgxas3GcoFxoEtw3Ec
1UcQS4MlD4yFkkLZt//KeO0FflwMGvXX0cmaphG06TLHdvViIg9vXa02X538FKQRJ1Cw2zV0FXzP
D10kYrLqikyEDpC6VPWrcTTYrkfR7sgZDYBClOhVzBfdNzYFuHOLXBaRMwmK8yQn0wtJgHJLbOFl
+vn6yc2S/z1cWzPi/wFt2L0xoOBoEFSChJRbM1wrdMS39kuC+GhEfdpPHAmyeFjfjp4z7eXqGaE+
+Ys2IN5oreE1GCJKXqCypDmXsu3Qd2XZVP+R7/eCEzOxF4l4/0z4KwwNywjzVtHUA0np7avdJlMu
xpJyQwuIU0v29rn58MQKNq7jK4LdyoyjmRsDumes5h3SMWFiD6oAp3uPcm+kxo4714KGc8388rsI
RxZdvmTK9w/BscyS56VzBx0EinfRXFmYlZzN3MFKtLCCm8Sxpq8lj3MjY7Ntd655K4SiYGMGCAwe
UKa77b59qTZdPZFQLuD+o7P5sVKLNH4hW+3ZY3yESxS/SVXiGv2gviMRLYqqDipMur6rVHMVotWR
Xxg4k8sdSzBrwlkZYhuKfjVUmXoMWjX01mV6B9O4xK3dzuS+EDqDvhO9iB31SC8vhF2PMcjnUflx
mQxVYUaQlJCUVR5ZybpaRRRP/sRKguwCOK1IFbb6AFQ3/silAHrMjmd8i9OBCJvQ4vZqe4j9JXII
jEtSoqGtTPDvTe8dzPgSxShvvIF/I0OutD0F4BahyPAx+vVjUIU9LaZ2ykZBYvWv0cI9Ai6rDZIQ
Dwv4yiuqSfk9KQBXfbKN55XFSeTvzxo7qyjg37bh9100n/uT68jgOU49kE4P1K5hJRtGHTH3z4Ee
czu/2uP3WYGMLdLc6/lRVimjNB+b+krgZwYov2InamXCskuomHZx8sEbD9TIIoM0u+F91HEE4Q9c
83B4YkGjWMC57MfuD4TpMd3Ncl9WYbsdb50lrWhzyWTORaAFcGKD9J9Xlrkvqp7bX5FmlsAlIvwM
sQUgnuI92dQqMmtxgX7G+0zn2uXBPzJf/OzcUBPjWB3CcplzWQ8qh8swj6vMXBsE78t6mltKfKGL
vDdZdZQO7n6HovKtYz2RdjRqJypgBaEsab0NUJaMVfuMW5j8kuONMLTMo52GtiFWHzFX9DxE59mB
Q9eBVNLtT/1thX8QeSb5BOQvZYGcKqVHZr8hR1DYPS/2BbhQ7rArFs3+l3lPEMKH4CCAiWdUAqEd
hDo5+QFw+UtNmVvprc7JjmLm9k2uYAJSmbvwV5rAuX/UjiWHydUYbjGZwMwo0ENtsTqCGeJpqAPQ
8XucxQFx1Xg1DpcUlbSO2oHeoiQbJNFxx+IcFN+iAnDyFdt2C30XWBFXSbJP/BYqLdV3pmdRZz/Z
ozTrOKd9jV6V0jy8XLqBMScYh6BSRgSRi8Y/gVGJX7Qi5ybAGdRPLF+9yuVheCyM67N/eaft5ZS7
XUueEI0bizweLGtGOZi6vgqjGZd27ftLbnhH2dfbfXhxFc4+1bD42BPK5krXsVqIzXOkGHxVjTT5
Ddozh7FiqmceZPUTBIq2udhcRKvXHijUowzcSm1IXDDPf6agvTXDRL6OpzjjPAAqjC/lrYayroGE
cD+yLpRAZ1mNV6/MFn4PPxlrA+U+dKtyA6y5ydf6Eo8oqnCBw/a/LFdNZvDJb2pWgk7krsqnx2qi
NdPOzNdU5yR0Haq/BpMo7cmkEEX946nVCPe1exwB03qmrLnJO/Tq3yRejrUxU8jd9CPJGaXQWyTI
1rMIVmmnkXXEw+pfWvX0SPYLZL74J6IbP6R050f9mfdELgO4pNAcCR4GWRd821zmcPnwdr/smEzd
wmQiwetMhlqjnvGnH4aY103sSzS23ltdtklES6Apk+pUhB0/2+nqdyK3seydsh58z9SsUygHEX5h
w/A5ugPhN1fBXV79phTBWLEbIyE0yvABLbuQlBcl2A98oGHtqK0CoR2C8k/Se2XnVEePl98hNd6y
+IqTHYKtX/q2aiShWcQUDecT6xygUORbO81/mjfwmx3wrIbfA5P0wjGqtAvMb5SdLZ2U0QC/Du3i
ALKqO02Q+NfnWuGKJq4ZXvUB5FrlUwHi9gumYdFVU6QgoPjUSxk1pnMwvFqhqa2B98jzhdQaCXEN
8Hd8zDulZCds/gs/m9I/CVmzC3kgu2EHsQBSI34MOplEf4WOLUuq1oC4fyFXdy+thxZaeXgpObNF
9rrz9g8b8dR1QkJlfV1ckZCxZei2un3jPFHC59k1mN41LU1aV54QtxQ/Iad/t2XkucICMwQRZcY4
cQYGyqXN0FrViY+s0fNQrsP+VmfwQFDUuH4wws8aqzRdjPOf4PHBedXprzm77qEPhq+LBTIh/zeH
qCMeYr4btHxXK2iptc8lCkkzV2/mkl39c9IiSNFdB6nwNSWkp7E9fbIIqPF7J52QLaty4ACDFmv8
C21JZ/LDoxbZQz6aGxnA4avQV4cv2n72VvpjPwKJEyApuxhDX6o5bS/1QGBLmTZ7iqYhw65Y3SWO
iw4/eowM7YTxUFDoi/rSMlKBPwFunNrO9rns1T2NYtlsg4bPVG9U6MPGeJgkQCxhhXqfmxOwbCDh
d/Wfbqd7EB9NNQabpXV2p4MUUCPAiRntqmyvT8MT4Gb+gj2RXvNydqAuRTw33Urh0ZlTtlYCjHIZ
T/oyMdHMfFwZL558qFFmRa3C4Xgz8IWVaTZCcP4FzsfeU+rB74eLiRwajmsLAkB7opAhQM9JNreQ
ZgjWGflTwafisI8HMbzEeov0jpRg1CsqTjS8TfOlYRTvo+GN3SHgs2ehnyriJqx8t9EM1X4rpuxb
3bFWmfOjM3IQUwl4Ndbl+KwatP7KIGxLtBYJyc+VSspyTN89wn0nYbjOtD1FkwPys/QLIdrqhhc1
VEwqSE/cpi1811eahT6qIwpV+CR/6puUGt150yvpjKS0r8Grr7kPfSqMV2qOZ0WNwNheaXFfKnUn
irGR25gE6F6F+3gN+UfGCPqYHBgkZTiw/42Sz0WhDBqetskS/b4OvJ0YCHhXeqS5DaqF0HxQueeX
7xP22gdPBGm7SgXqIut27UikJOo+yy8bF8IGlZcuRK+jX1KDBWX/SvGx7Xvs0bEdap8iPAWUNrj7
8v2oV4x/3fKUBoWanN4nERUuL7wfWWKjrbtq7DZL5p9VLF5Bmiv52Tx+evvBqSp1tXNsRPyNE/my
dm1kFcQQQTqUuIGD1fwC3YjFkyyH+5CY+tYqnEXMt9j/kDoWWWdf2kpObWwXjh7rtrHE0t4+L2nI
gGqODyWM/DMnN8Qj/TIGQUmzKDmYN+jgDZ802TzGC0r0M4oOM2s34hqw12hRJMI9ns8jLVT51wLw
1xMALBhqBZHarN+9ChFd7U9xEcdaojPAketxt2QQ2J8tbNSH4AmfjmvngNQuknBxBkQIZKYU4dQC
x0LYlEYFlP0NYKwI8hGDcHgQ7Szjwl+m+9h+G9wL+pkO1hLdzAmgZAgy71hvb6L3rVqs4TfiWOmR
L3coviP3z7BxFlA+zqJyl3rtHOkOwMI33vdd6rL3VKro038rVgMg1YRXpIn3g2r7L6D5pawtOpI4
q09wCLi3ayGx4kzSLry7YPnbx7KhOwp8fYEKckMV/8uLNxdmUnpVHG8soApZma1W6+aym3Ukaocy
PaFXsN99chM25eHZd2pydcnlgD+v1cful73oOkDT0S4LvMm6c8FmNkz1zj4GNOOVur9R5GVXLuDV
HjXSWzcYHW9z1sk5FJauFbqWSuuYueSTNNThu48oYez9m68lQCDGnNjlQFBbF+jRIO3+jds/b+Na
TqdvFJqnhm0ojslJIqqfxcrw4FHkHdb37FeXVRDbe0t2IpzLEdeEfNVcpgWbkJjrHEOgJeIRoGZw
ve8UF5zd0Kpkedg4U3D0jDG6Fo/W+nI0UPszoa/OG9kWIBrAIYW9X2koW1enAuf/4j6WlNYFiiax
7Djsk8dBJpWfPvAUWBHnmJUbaROyLhQDdGGG81loZ9NeQIGGK1x4VGXrxTtg+CGD+u2DLxVBViHL
ph8xid9/LTMV1kbkxbhmKJv9TmY95+xjTpbGmD0QnLIR/Y+XiCl8AJZnaFJoNN+lbgA6+9w26G5T
nPFel0k7ALGfnlJ6iveWuK190kOIsA44VyZygCmbhyEtD3jiKl67BojZeGSoHZP9KXHsfsSpJgXJ
iWlCnqSlhzPFpu2n+vfu7ID3hOI0wE6menlwlQc4jGiXfNDzGwsUbVof0JvqSyL07VmDaHdP0Qnz
qS9NQMdVOFmjg4HIMRPAYMdV/XNn1Gl38Lknd/Jo0by34ew0vv9/g8O4He1mxkxyZM2CkJJJesVB
jhh5YkDY8e0YljAjauRBTDdfmM0YaG+tfoa0SI0wjsExe9ZS5k5jFAowBKxYPvbIpyroUCkg08gu
7zwS5HeJX8Zmr3KhvFe8JcsknHCvud/SEtiHg70Mo6+CbrqUHa/AvR9V0jXNTba34xM+r3IG+pv3
3pMpXuxMvpS2iIWFBuM4wksz/ma2lOC2LUeOMiO1bfEu7naWmFK1eGnm2XPJt+INNU/KWhxuiTlX
f13/DAqmBcDb2N4oE6UEcKS7NlW2j1mSwetuDss/Huky9cQBJ67AMBQDqKHnMydW5IKs48NU8/x0
VuOIIyyZwNgrineaXlAbAG478IMHyA2Aj/Bj9ROq7JkCKkKfAHFXFnHks6ErM4dLIyfwPo9ledvu
EV8pzf22iCakpmjNUgkXrd4JHSJyfcyCVAM7bYXrVAgZPyOyoeQT7xYQnWi1LGT8vnNPAPUdQ/WG
lQyGO+ozAUE9I4SJ3XYWh7q/uHOEVkWQAr5U98CGf/kTQtTinhbusKQSsPjsbEWtEZB95LnLxp15
/IFM0WamWMRC8kIEjSUPUD9yyet5+BBRp7M21apcfBYv73G9QJgbfnRHW+nWpXsmDP1DUiswZA8J
3hGg2kuN8cCa8MAIwUvlqE9fjbaRFtxKGod0sM/6cmwKfDz5LJltlCmsxy0M06uQzlxlMstZMzPY
lNhKIfZtQuX06ycT9Wb43b84DtZUj3tDNc40nkxJrBjMoCT2F8AzSYOBb3KpM+NYelE+s/R+919a
rzDlarQe9XLXGIGyVeTbuH3bd/DJN7v5fuR93pJkTg9JvFmh29nQTQGyu53St2au0ayDKFaNaFYr
zJSG3mlvuExdUKOnTrx/FQOYoZieE7a/Tp4qdDeJEzK7+RxmjkFODs2bBLKtH63xoxK7aEUlgK9k
W1u6Orlg5ZEs25RZQunt3cibxPAGvsRVmOdq9aIAr6A4cW664Zf0op9MJAKnCHjdqCWf5Uwnov3a
fFNp7gCkJRIa/8SodCAwb5+wD/JbAGjQuzZlL+N6a5gs0XzGQ8q4L6qQOPqDZKa22RfYNDlbJuqF
opFigP+Yu3L48pu+NEGz5bTAbu2XUDHS+675QzgCuRoIO0E/G35oIZgxCnMGEhhP3uR6unnCH+eE
W2BnrHLkR8kCHES0rf+cfNBdnuATuW5JsUH/cgiPwMda0wft51L/vazaT4vR6fqa0Uyb8JpypoAB
QW9JPu3iZgi5+I4n2QIN6VQqoqqq+IGHLBPoH/R3ifeT1j/PKbT3gJ+2hSkT+37C/37BikMzXB92
9O4O839NBx3s0yDc0jD9+V7Cs22qP4WrxlbjoSB0yy5nAogINqcUABViWRf14TMMKXHetdveSLfw
TSbqWxqDjQxsMXQIv10J8JzBBk4431fXi4vODqGDd/Rd/T4DvefgrO3WSRavWvoGdx1KGVMRgOLI
jcyl5PBt3AYRUTeWcsEDy/Wk5HS7DOl8jLQKfohWK5tYpAH9LfSXOuoaBBgJ405Ri3iQU7Tt5wd4
yemiad50UmlSc4vIO90HzoAyUVTIn4+p8OrYqScQl+VTKUyXKf8IDld4Gwp5/km+7XJUwtmo8+1k
lzIJrpZEsK9PjJmGVfsG+uz5xMnlH8Mrq//ACpHIcK+v2jcpB91B6T8Z+uKVo6jMDPtG5Jc3DdW7
hULyfIIbUXFeYXn29C90JKEJlBnFAqi+ckFwpdYv3FNUKLqfXPmRSmliB0mjDf5YWrO5kSjmlCm6
oOnwy6SBIzdGzkloCnCGOENbHryzwXkobOU55VAfsuG9i9hkDFX4Ka9aMHjpEGQQaiZvpeh1R2xo
Pj58P2tDSMu+31qrO+UclOrWZuoA67l3yvmnEAN0VWff/V1tuUbmgpxQj2RGNfsau4sU3/On0slH
EoPHuz9QRzEA/qfAtQAabZmxq8gEK/HMazC2FKdc5W7Z6qpKQijtRJUArNmUXhGU5Ba/iJFaNlNK
3YiScxDPB4l8vY6qtHdOaxYdVbcagvogU7Pl7JrUVpwM/Mc9lrapyNWAOgYKjWwJwN9u7qrW30dY
91yYpbyA9rs8gDJHNBUv9tLfL61dhF0j7VISc8ic6/aNhNyl4z/53IpSm/loycWT/zUJh2wZT39l
53oUmaLZEHOR1OLq6fKvN6F8AIjoCtMKTd77xATxH8vyL96t89W68U7zxpW0znCpCUbN/wAi7YeZ
gV+nYyQHIp+dsiUuhD8MUq0VUrAGj+45jV4slXi3ovcdKiCHKNH2RTgIReLvYetSWfDxZmQ9Aa2Y
jL8DSPEIb/Itp76Rhf5v/Jt0D1N51hXwFP6E0uTl60AJxn8xGgI3gAegWdifLRBNps99psopQ0C5
egaAfEzBPZ1dViRIwvd9Xv/uV2UHa2f+bzFbCOXwY39j/43dJ5ZSZzhpVWIMVZ7DXy/3P0fagdwt
EVP0FXnkjWJZi2wji86opX2OAu826TZT41KnXS8eJIlb4+cYsWF0hVB4qwmISeIh6CNUeHaoACwF
TQcNHvQcQpJ+YbIcn82SA34U0J2ZSLcVM+tS4o7ExBbYVHGuGmn4HqgVhNJuiRPCqD+BcnKPdISz
aKIgwut+qxE605135QpOGGBwm4F2drdz3QhX7ROgYUstyv9jp24XPFypy/Fn+d3v7tJbUqby8uyB
3a1quLt8/l+uT9uWPDSbu4Y1AjPPrerzu0jkHBle2c536HCw5JVIPxQdktml+jY8P4W3fC6p/TT6
oZjTJL+cn3cuLVnrGvs/MmS6HxzPdK2h7rMFVas60RPPR5+tLD6NfarcuvHhlEXivKZNtH1HJnBH
8KansKllFljixaRgunOzZWRRXfbd/6ZVoFQHPi6/jHsT16zcyEGH1AhOBse4XN+fGbqY1igTr39h
Y9GQ2q6l98WYZhwB0dByTuAuEnpaCraMccmKontO7UXqNIJnk4cSsre0OmVToPA0C5SLYXzq4Vi9
BSpiJx3JN53epi9/P1uQvAupCyN2OxV/MGOtzKzwuPv3O6bXT8kaiP+ExGOkkF1LsglB7KyJp2kf
XqfTCixnDrPJJMGzjDmCH8zJZUzmU9jgjNtzYkmmtoOPc2Iw5VvzFzXpVuvJMF6ZwgwPSnnD7FBp
bMqLbBqOpo5A3MlWGR9q7wWott4WO1E+/Bxj2AqSsK2hLe/2gcPJFHAPTEjg6xUCabvz6AByTmIO
Y4kzVuST2TSBbWGKKqUR0CW5D0uj+4wqNKLmet1oFnQ+eSREf6x8hjW8LBb9nTFEGNh0YF5YdewL
boE6qR+ZuSbaohp5jIXAzuTIq6daxVn8SYyVptHk0O1cSZYbZsGRjK++5ojTNzZ+pcESs5abmq9D
2S7KlThK3WgvCO9Jvx5tFy08QFMYZS40xm6E6VrruqGaHegyi6ZJrI0g9l+TQyoC4VZsbHdAhjw1
B0y72acg6xpKaQ7sdOUAWW7nQuFtckqXX0t4AQIqSApuRTQGRv1/qL17oJtscSg5JmOMSk8QMNtl
1T1E3Jey6hMl23g6oWouzXvpyUiJb/Yvob53dzWS3Q2Bc2fd4ER1Pta8WNc11qx7ojqT+IiBnLxE
c8D4ZAZ0U5X1Qjr6RiLw0AAIA4wIpIR+Ug9laEffDfXOlfJCc/tZej7NWtPzjnem6PT8zInFV2uR
qys6XemmdH8PlA3NWNgoby+XTa1oH/p2b+d7/7OAtoEIdogXzMxFVxv06+Wa3yKGrqpLeKJlymkC
Rf4ktXmvWpYtsUsd3v13Rp/4Dcy5w+O8Mq9b9tOlMsh2vw4nT4DkfihkNRJkRHwyfjP7E9rz+Iwi
2AANdpbIzaa7uIach7wN9HC4Gq/2QEdZKJHdjcO8IBAiYkLHLGdZ4ftpkxMuMuqTWHQnBLb0XRv2
gojDXFCvsHkkjg5yPnL1Np/zCPOlAc9AG/9IE3i5Ukn0Z6edEkNmPwr9zDT4/foKuzUuZ/UNjauh
g9ctHif5dD73Io3wPdppDdRYyOjpe0CVr7vREvBxwh87KXzpr4/pBSMB0FIPv2b4XWqBg+TNk/ic
DonWj5M8a9H6UdeoEa1FkEYS3PUDY18EhGC1hbC2s7xVTP5MI9mMGnSwnmQds/EMVjFl0f229I/P
pPaENfPvLguB1b+83MC5rvhxbWIUA8NdxH7Ewe6D/5ddC4tiLIxlI73aVSnCMg4/Uw0xEmtke6lx
p21NYftzrv7T3mpEezewbnXTD0ifZhoQntU4CMuJDiTOJg7yDi2ID5rAgOn9/Q4HheYShDtLaj6x
IeUs/rqYutfIA+9ljtU9bKgdSvOdn2+hHMiKOs5vtOc8zExE9CruvzietDDJbNpqMdi8GGfDxBzV
uLQK1tICXUcM2e0DZPtMytPQV7LAMOZdKKO/9FXFeIneEXrsviz7L7/CD/emxnTjsLmgQ4drQBrL
Bh8VxKLvzN14e40TmncOzKljUMTV9MBD3D7ANdMk19QUPSnFWpdAUaHP0zRu1QFs1bImAXRp9yt/
bszzUaco3sSuP7Tvhq+qDqt+eX/G79BtMGSQpY8DehELwF22hKYD8Lsopo6PqdV9itOz6SVlVr+O
bNaGk2JzbhOcCO0hB4v9JPxjTo/jMPtlXRxhv6oGUyqv/X04i2zeL4kZL+Sq/FFlMZeOxTYao6yb
Nsoe9PvegjrQKtWKqY3WE5fEFVPYF8oEO12zsTXFGPk7cSLcqX6h49mMkfwLYMhJyCLS4AwYfDbO
HS7LK0JWVzh8yaQT33ofpwef3IZWn2axxlm9FEKuQlV9RGLAWPCUyu2TlvCkIqIsASG5iBDdsgRZ
Xz+r405BUJRF1VwM1rbbZX99kEx949kyyRTEPdrR2HeHAOWvmrNiBt54m/pxPHbjEkoIMHT7NXLW
yOk+HXo8avUf6Lh37jHtQvMhGKMNvuLaZq9gh2PtnGqPErQ3pYARZwrHyCjPeeJrN1cH7LMl+/oE
TiUMgNci6qSLBS7cVnws5PHEN/JFy+JRF9+hkFBS2e/diXi9wL/dNIVLfCQJ/iS+hA3qhieOTtu5
nccrsFFSte0Jj6xSiekPwAkePcS3HneUsE4r6BkDY7rr5GsCdfyYcieZ2jinY7/LpqS81mfTkgeC
BF81UlnVKFLWLEM56QQE7udY3cyoDzxjAuXUbR2sEqXuz5EP0IjtxmuEG6yykKT2VNhXfIeutUj8
l4h6V33NX+YcqViCtZfUWjGY5KLDLDJB52s6JAMs20rit0TjWyVEe0534bC+XzILW2zmmWzD5ty6
/Ln+M44Q8eYN8kVF1CrbzAacGPtrGkRpkldKa64w0mPiEG1QclZqPrRHxa4f92M43wKX7RrLlcQ3
9hvTiWiQnD2FDOW3ZsM8cUIxAYdEBaB3b0nUrIG0bzZG4jFMeDcTw/UQwtsKPH7ii+Ko7QGXudnb
DZT1kiQlN8KUmO5KRHNBYU3HvZQ3KRejR5BWfjM+/+iqV0PqbEbmHeO7HrKYtwEm1N9+Fb85hZTM
XdvPi1JkOCDwxGY2WNyIkNbaRy4e2UR0DU8GFh3VllBZXHb0hLMMBe1WemgzvkcbOedEN+8T+QfV
vIWeOkn3t1HCD5SKrWkzJws04vBAk92ymmQKh7xqsSx3nURfZoaAPpd/9L/isMWIY1eN8bNoExRX
tAKGJkQAlwYJxZOOipnYKGivvxHbrLf8f5y6pbyE4lF1h/pwnon4cRUZ94lcbMHFo5cEPRV0Jxvk
EeXS+19uD1tBg4Ym67D6q3EaIEjE2tEaPwpQGqNwf5B4wBQ3CHwWaLMFxfjHvlDOjjuXlkInRDMg
aviBCPt2Irnf1QXV9AL9kdQuZK2lObi0H2ukJfE+TJs81ONjb7ORz85e28hudEnhC8gSssqySJu4
Is6Lv15L1Q8tEvWvNcS0RUGytao2urShfjhRTG25d01CSjg+/jDJvE6KXMmmypyRtEIV9qwPDCbc
900BjR6gRT03DqM6Is2Y2E2HqZd2jGo8emgioHoKr2/8Dm2ql3QJmYJ/tT8M9HFhgI0HLtLmMaty
aG1rZnpW1GnkE0nFu07jjvwctEBOvZJHokiVPM6IpMgWK2ZSlmREVUUJiVEzOeq4RrRUL+mnC/S1
/byFMdDzSquqY4bd9qAbeOGTFrv3wOxi386HIeiHy7RqA2VwsyXWBlqvmauqNfUPREsBY3cO5OaO
1e0g9YGVueMP5v+qt9+5Gv2pSwifmiajJ2nImPmev166ztETlVg/tonMEpiEmjySUs4U8GFeSEYg
HxjDDB2Q6kLuS0kl7zawjaONxIQ0+qDnvEK/of/k19GxL6JJP4Zcb85bYOBc5wLsbZO2rnRHXvuE
7+D06cmNREw3NSaee2UIbVU/KiSxnlPaR1iAfHMQx5VE1i2CvugJ3KYRL9/l/J+07jAV0kJFGh3B
QjuSsBbiIrkmk7t/zEnHdtU7cGa+FL+DgjzQqEC5qZCDtsydrthi7vHW5Q0IYpYEWsY5vKc4q9v7
051609b4dTPTvdxmLBMx7aDBU9xO4pFxdjdTDVBIe9zk64XnMK2HzjtlXcQPQek3ZD++6f2to7Rx
2RqbMjwXvMtH5gyP/a8/KdbEdf/brLlKqds34SgUT5CsERuPqNOy6DR+1+nneEehsfYD+cLh0Nuz
nYwriHknPyBjqlKeGy+9Rvnk6EaZAoz5eVOcDzwT+Wv3RSdvFhwvYauxSicX+xSLfaL7wO4KhIuM
zMstvEF1p0+n3Hfc8h1OCfVVnhX53vy+LrQ+KmaCmI2mRTBVyeLqzQbpyuy1xwYW/22f8JScfm8B
MOplLX1to8l4ahAJGCAfgRgFZsaQHStJHPDUF13bDvoIcS+o0uVEuvxAvrYpJ0/IBv5YkBLFpU3m
7C9rb8S2JXWkesq72o6vj3NT7QHDVGClp5JDU2smG+BJ1+Ptes3pWDgv1ZQXP7DHTi6U7scpwXTn
WYzQFFf1sM8K25HKxTTzABkVI5Q4s8Z9KUW4WxOuRGJ9ivD2mqdInERIXJnXhylQ2V0JL4otnK+Z
A6I7VVwbhF3dVj7pgtoAXUcV2D7b2Uhc5F3OrjoKtPUDxz8An9hWYVy2tp4I7NwMopik9bKaZgOb
QcyNjBT5bhx41ccRAJsgKvOQXkLAhO++mNGa61rv0l4YghA2c37Ml6vs0o7CyuD1Umo4B8k9zJZU
eNW4iQK1irEg9q7XOCLbCcdlZlFAmLjrBlNFJChtVnAidGntgwjJBgZYcbGcPKVxlFoA5bctkDYY
C26GuL0/+/YsVWIL6z9xT1CqcA84jTEvc3VIoq5OARX2UNamWKosrVqyHWkvFUBkm6FsUdhyZbWt
ZalY3VQik1ToElkSSijzDLl8ruQpxmex5kY2oQOPKbv2gmWcu78vH1pNfc8t4eDFYoTg/QSRjEs+
kSnCG01fQRJWngkEoRd+Wzxf1UM1SjQv7XRDA8XfraO9bIQUqbhth0NljF2np8GjF7EhxbUHdCO4
/Pc0hVnlq4XHpqrPTikUQQCLLhzWYzvXL3uR8OOBpS7HE+gkOxfZzKTNHn82iZpNLqpmyFTso34Y
suV7CTMvt1aKtRZaKMT51Y4oTWG9DFr5aEmWOThtg0Ff9ZKVcGRK3p2S/vW1PuYlg2+0xoM3goSa
9cuAStmycRsix96inTPNuE5UQsNtHRl6GKAHm95kR10cDtSaAZVCfRLMbhqP3we56nEiC2/cGpQ3
+GvwIRXLVrHMMdWjCabwnRmXdkK0edGZSDP0Q0HugSEvJIJNU4okfGsDfEbCwmE1CdWz7wyVigrZ
qsx7kisjMPVJbgP/ZEM9sexbWFNEAziEH7BIHWpzee2tyhuXbQng996HBEdTU1WUlfFHAzqRmVXq
EYWKBlIssLdop/BTHZIVPzDVDRgRoD+jRPzgDVdf9WmAaQmNJrwSlhPaiuqaHHGJpNnWJRcq0J8k
ex16KcEXZQzeza5Lb6fUTd+l8BpTkx//41G7T/n1A9kSQFFuYaw1tt0fr0duGsyRO2iDtjSQ5Ned
uWp7GEd19aAIYtOPpNtd3vFb7zLQSdPDnGzWVlpzHTJr42sqiA0mqy2KhHwbIviWLxWOZlQosNKg
1EZ5KRQMQxorC1re0b6N+FjsLGAbbz1W/6xPxTCttye36udecRJvYZ2VZ3I0kFB6ra6zdzZDm6Jz
vuqIPcmDR+xQs4l6/kvP6G3M4GMa2kdhLUUfLrZyo+lO2nmpceNi6nZezVezyNRaa7zhzr1Q9+FJ
ttcfRw+6PdgK92yWDXNwcMM9K4iizaT8C47v4qXqn/rcaiSctdWsvpXqD/3PEeDtSOOWLzpyFVkl
Xo6mAZ8az3ohn7hTh8QDr+mMUEXSTSRB4pr/rmKtId8ukch3MtJ5Xae6Q8Sysn/NL0fu7v696Kih
BXjgl5UQcuxsLGidnNFXM6ta6fWf8nIB5uFpExKC+SBk0HmmQN+V7B7bAiZz5L9yatOhYDFlPTjo
BPkW3Cqdj80ziGj7lmDaoC0DUXiMWVgJt6JNljzG400KfDzQAThYkliiUyPhFpVK63FNcYRSCLsV
/QNIECZCv47osK0jsi7RTl20LziZ7qqChfoAuB2mxDqXzXied2jme5ihW6i03rgaqcs09ZlfmTwG
gOondH5ijRQxVHO+t0fcaW7oYc4LdwY7nQ+mbtCN5KpNI+l5yHLMOpQMu3YgT4cl1Bi2xfQZ4yo+
vs7a57IoROs92TX7043gFvG742mEPipR+ipw0qtROs+v7QBEmAE8AfnmvlSyu7ZoJweEF9fql0J0
KUWwEhENHisfLFq1Vkh3p/e/Xb8zr7Fj/OCO+oDy0Ph1weCGleD1AGAxIVMdejPGzfxGaI4RYgwZ
KXKeKwNfU4guqnWLhkT24J3n+sEggGTTRdqMx9vgufuXYNp2oykblYO5p7d+1l0rQ8uP/XhMojdu
Mvh33Cuo1bPyporCDIB7NKUX/M/BaV918dHCBM7okD3E/rZ2trSdlaIN9u5Y81/wAP5VrPCgs0h/
4m6/KCPprFsS28FLrx6JJEBxEwIOL1wWxTczNv1lp57pOom/pmVMkdNm+pjzFwciZ4KNjRHz3PsB
5Q9bi2NIj5C44OMTaxayQiWi/ggv5PU7kIwOpfxxrD8JJ9gSpjM2ENVi3uC2e9lgMxhu03634mTd
sjVqHtQE3Tqeql/JDdm/+qPbd7AqcZoteCpTc8uY4JY6dglZoy46pjwKvduwPlZ7ak/vONirPbbG
Xw70vSl7KgPcUlnAgsZVo2PWGERacyjZ71Hn7vtA7qM+UG83QulBJZAK7/G03xFsl05nt4405tlG
ZzajS/rUtWZ+iIqsFSi6ZTkb+COMoQTEr/fm9GYRbTqFJofhYJi3EjjbtBuXgt+jRKsAVVkNj+2K
mYpP9719KE2v3Gh/pWTsr+0DC5lQK+RoKYVLU7u+7xtXd6J9dbxvOuKn5GrjMfEDHi0/id9DryiQ
veqfkRhxXumiXtvdIPlQy51ubIv84fu/6HPUsBiPrJPKxPF9XTiMmZNLJGn2dykm1MQpFNA7Pt9L
3tVXPvqMS5f8hIBpyOzbJydHcJdRdLcrNzQXWhVLLZglIFJFEnDmiS3oPla44Nf9Ouyp93HX7uY2
mnqXXh/Np0TbpblZ4L1jLGYOWydXpKRUKj/ZIivacRI52lmuOIkUL0nNovdl3dhpZOXHQnQkat8K
9uqBthnesOr+PsMVtSaP5JmwsU+s8MHxSbuA03VIMq3L3ziaTJB7hoJhrD0fTWfbTN3RCIRkHvEL
DNCaGQ9BY7rhiKaQS91cz9OPyrxRSYbPtBsKdEQ/ymkwkWbgSJ9iqYFHULbkXlyXvqwrc4Yka7Hb
wBzQtOJHILBDOaNfqL7ZqFTrqhGmIV9Jofuyq6ghMh2oEAAiNHkrevFkY7+HG/jcH7O2I1IeNcYg
v1tpPc1AQFp2Fm7+jC0VeQIDv4MNcd9b5VVMpehAQChc5u0EhYKFIpk3T01XLgTjeDhdPfiVWWLU
9QOM1uT9k3SoNuLHLiCynBm3u7y2afDMUBCOnfJcx6yb9AGWSbkmNg+320zG2B1MUmhsZ/laHTMj
E3GuMCG5so+nzhJeVmUC+wBZweJiG72qFsJyfjRUuR+yaYvRv/1KPKOAqXiRSGAKwqqid8YDhwN7
Gqfmm2Tj3MPdzhhZT1D7rvv41Taput0RyP+OtcVQ3ZQQy0KtUmSSfevVH2VyGDl7V+DvNYBOlIue
OOYC4z+V1q4s036doKesPSOAL9wbROUtO1Km2Tp/wx6JzAQAyjxnrZBk1hTgCUJhVPLrFXs2fzh3
R+H1MBnc7+ce5knkMAQSutqocAgSmEqsorzAPxzNiGdIaBtYIuaJBKKhV8vNR7O7FDiMJ3KzR8r7
5MMePZLUQ6+XYcXJ8KymstDuSB9+/PG999CkCcMovZTS8w0nmfGr8ki55TUlxK3jXGqbz2oxLgIR
PrQdE4s0L6k4AL1USZfKS7sQ3Dv0X6fSrV6kF2Aw5nXDxK18+hShFWhUnXetzuxq3s4MSGp3279Q
LHnTgpLLx/HA7gqb2PWF8ZwwpWy/U6dMLLDxLKEzHFFchW6ZeRb6wvaRVXXi7L7SenhwFv+8vql5
BqvAuvsM7dYBT4ozTnJboK9iw75OgQojIVc7UN7KN8LXskVdxpI9YMb3/OAreVmudsx1fbOR97/T
Dk1ZuhQzft1koGex3cUZGQ6ikYMLsS/N5TVK3XCCQKOtO9tsH7KihAp5KSqUS1ezV4TEOp4oLNuW
pfdorD50XugNW9sa6TeBn4yFjcnQ1DHUVUb/pv5qcxjO8WuqCf5i1satomfGZBGXAL1EVo/3NiZP
v90HM1KaYmNxh54qOnDsbQ4gVuZIv4PARwoSk9OaIBM2sDJRxVm7nqmlX1iZ2mGmzYzyj2DEyygK
SdGWEnAS43Srr/a/+FJYMedyC626SwNKH2xHqnVwEWg2eFIxwrXYZ10zDACznUAzZYXB3+9mMD5I
EXRa9kdBQR2TwGDKHidvkeO9MCNbRmmbZGpshXwF2YrSSAH9mq2vbMI7Z3UPGAdQPVOJCairIXch
sA3llHH4gUsfd2n5mtkT35ULrl1667mchI5UR5wHgGLcVgPZDBJDVq4t1F8kVDkukixCAwFjJw0K
cRwYdKoLvg9jO6/Q+O0oH+4GBY93ANfIDSvvzkJeLmdfqtxnRf4AWkkaZOXGPoYVvJuSREE6gRbq
rsA/VApdhA1GKfMLu9razahjtMmxgCIYbZzkWZLdZTcxWdUHfYVzIWlHHiZpbsZzwHNHJ93xNScj
5+pikXt+0l5o2KXNLRYbbAMI1FHCjApwBx6pMkLCJCFmg9A+eQwDbQzmcEjWZEm3Suh/jk58jPY0
GsYOBozxEMP6jSsEIB7mwDLFHcUdkJ/S9+PiqFvydR9Qxp9av4KwhRAOT/p0+Xo9X4gQ4IBySmyp
+nEEJzLQLwU7KkRz6vKhl/vK6s8XCGP3M+PYY52Vc0/IL4jQst8YvQrHsAClqEP8hgII0phehkLR
ewecrlVdF4cx2IMJlEH41MnFJzEkDvdsv4CjXyuFM+bvUCSKQxsbE6CyE4NVp46qJj94YATfIKt6
4S1DS72Is5tpWubLMOsQkRMA8Rb0ROgUKGGDpqbBRVp8dAal3r4h+1dMTt1b1+dAIZ7DwK3zirTk
0FHp5jJ0sntxnPKWP8ZAyjqV1Pk8S65xkY9+hn7K6Uz0DOBsNsMiQD5+dJRm5oIHoHxEYkKYIRGw
C6vYI5hEFQkCUfWEtM39Zzy3iLzju4jvZbWaIPx+vsrB+P14YFfEtbps+PJp7zlNGGiH1xHgrlj7
36ff0JK+hVmueE1LQOW9ja0NLhi+3JK0VgdKgAKLk0K+vFKHVwQAQ9SH3zYMHxh/K95qxi5a1Ro+
AIw0n5ZvqWVdMoRxjpDTd1P29A0Rtj+MzramvVpe3f9l56AOMRosnR0qLXld3PzxzXQxeQK2djA9
gkf0H3VuAyrGLCYcosGCmABbxJjIbo2lS/AzIg46xzR2i6Gb9Lrcu6xt9LobTseGt1KteBL3B7Ve
oGujt4HSzdv6uF65Izm6kFStGpGe/NvZUVToG0eWV16b4tOYamJLYGpVRXKKyD2JaaBlclzibXEj
AK13bu+e8KawLLc41Y+MfsZArLMmh2000BP4TONlCSgTyL8fNITSggbzimd4DQVhSwdUywe4savw
nxWcoiGMjedyguQOV2DkoOmAXVRItzjxpJXvd5VxAJ4EaZFpQ9SkDVgd7EyIkSSU7bRxwSAVk2Uk
UlyD1655T9DmFnXvnpgMprV7k/E5g5v9IcZt3mW7cWWk/kcZx9nJiZTmP5uleY1Pc6YgltP3oFst
WmY+5oEXPP8uQ+2LMRC/nBC0MZVoREa0NgyQVJJEnXvPu+oEvVRBKMdhXSgAUEiqPoDWPSvi8oTz
LAGrZ39KSddF6EgHT+c2mpEevxpHXZqf+sj3sADzUXm4VheJ0jLDcjtBQPeNqyF/irvNHmQ13F/N
ogv1BzT4F0wUt84lyRvWELnZWujFLkFlYXnZZ/PRhy4c2yz1c/Jq0JDS/DjiX860KQEeBUO5WauX
y+dUXqzbMCSWdb4e1YRizN6An6NvKKrHwHUVh0cbn70SbilQ5JWRNnEcPtcZG/iWsN1EpfEUvGwe
rAQ19XmLopI0km/eVARnfk2eEOd+p3ZTfdi+GVWUaNyYeyV4FcMezipsErQ+2m4KyVU4ehG36w9T
kG7xGipzy8sjP1Bz7MG7cb/YaWsWq6vmbond2GzsPitWysiAWkzZJM7NVbGa2vYCHfgYRa2GQ2rx
otgokFnGQvT3iwsuLbEqLseWHc28UrzciFWGAPHWdA9GlAcNH+kc/yLuJCIjzUg5TS3EuAaiTX3q
kWSVWexNaFQwQhkqGZF60TWNLl6ppD9dYp1eyePBQZUTW8gQJqz3zlttH7mUfPWjreVaApY61eYT
e5HxsGKzy2aEu9/qwNd5F3d14fA7E+zOyxMu57OS12noWkgEbvr7DMGCyRMKYMPvtjQrMTCKOyry
XqYl4kmWAHL1sS7gljfPNyq2hNMOdWF8nXNuR4xvvUYOVR46Sx1AYgn6slza04SUJ5GCofGGo6vr
HFLf1br2imYNCpjasPMdKPxkvU68x7GssqrVAMxFiEjp6FPOHP5inLk0h2jPmx6f0iaiZoJ4ASpB
8Nx1bNGcEUguKQ5a4vzDy5ssHeZWMdqwhyPvpr62kO0rwISO7Q9fEW6QyFnfoei2n1857kdT1F1o
1S1bGjRlrZRwhlyM7oj5b5iyWtpvhGtPGPrP2jCm9AKrtkNYeiAE3Nvh9RXDV+ci+ylZPcgFIyJz
1NNrVMhd28Vqhp6NItSKRLkS9ZJgA6MHTex3i5Kxxl9Hjh4a8YcCwi7LZ3jy0gWfR8XSfRvFXuO4
AZG9+Dv1qeedkYXvGOIIUbTgijgt6Ab68uS3bHNTeGvsWsfA3D+QyYOLGN3gNM45Y6Rbt2ZWTuAC
PtPsmbmJ6UTAZR6PJsp6Q74pwE1/Wo9obhMD3ZcMB3GQ85n5vBNbhMc3D5qB2dCWq1Sv/yVeNSbO
IZH9lBlDukW8hoQVDet1bwbV+IVIGTU+u7CimHQ4xE9oZD9+SOT8FhAP5JRy5343t+qYi2aJAwFJ
v7CtAWqdrS+wtiTrWB46mONa0M0QMAw7nu/XnORDkYShKyWwS0BgUJa1/L9aBjvCo9vmo86pd1+t
3l93hTag5uYUZ8OJfruZYAwmE0PdlKsIuIoi1s3TEzjirTEuLTFYu1+45taIjs0suHE/xp9pLoHG
H1rjy9EwjRo1sRvPmkSj9F38zpPe7NNo2GRPBBadhvQ8SxX5M22sZNfdJkJ/ka040GAfej5yxr8w
wIO+uLOrxazoODvnRFNf43cDmgPJD08T98FsRaWIv07BI8kwrKgcw9YVoE4FpH50ZVyfezBsox5x
Lieguf0SNfEhtc5ybu9Yi24jRpgdcPWsa73RO20EXNHLUCvVXIU34KnyryV1UjLx1aF0SmMD2bRu
TUbFAYd0yi75BrKOTQBQSFelyWW3Pny+bbCrRTYqlAHkbG2M1wNGvIPbqV60ncL8VbJm8xdDo01x
5VNgFr3bwrO8MKtOpw7hdy6yQAFvdtkWEGtH4T5MGePSdjQi578hIu9a8uh0bHGqjCFibVWYoyoU
1hnJvvTxF0QSg+BLMnfMjvZH874qpeKf6Og2uTk3dIxn8EqMZS5Y12F6YVVvbRUXkLye8AsfeSN9
kPB/4B7cosa1bmAU/WGF1vGRi07bl98aGO3/ce+5YpFA+NnbthMODgb55uHTNhldHe3KMKDLkNBQ
vGlm8LlkjkStTzCJ0XrqOdSYN7hLHFid8K6wxUFN6fvmiA2fP52W6kyhB4uABpHINEkn5H+8aJHF
QLFuAIMo3ZGAd0D4/F9Qe1+YZO+zxDKxg6hO6+VAtc8ZHjA9b6F/tSTk8gnBrkIhMcz0LgOnEKOO
il3FBiME1aO/K1+BGWBb++ibGxz8Fsk2Qi3q6DDkRInxcK2NeKvGrbkXPhcQmdHDgZpDVak4h2Tz
yXr+p8M0LCJ3p2OvIu0sL6q4DMUhMLVVUpoe+5uWjj4+KJGST2NJwO06wITd6nuV0EzY7MIeogR1
O5F6CIzQsWS70I+8tl7QcfGTyr+LvST9CuGJtB3A3ZJhzjMmdzRyeM9evhMhWnrjP8xpOiVaJhdk
FJuXyPwrKb39TBn5RgE+7XHfuO+6vs2Vp9YBQaRVHSgYg1zWQgpYPTgCWjkwy4d0+1NQ7beKqTat
tfrUcc5mE5AAS/E78sEwQJJgyFaGD5eAl92+FBM64PC+t5GjqVCfm0BMhinhJBndnlVrP4hZ9+5Y
5izkEZe2Hr4Ob6qT5ZO4VgMC8Yr+uDDnPMDO7uqzT1lqKxJrHNmm2g/vXxMP8NuULXSnn5riRTXE
RRnrYkydKaoMgidKP95b/fhXWkT0HAzC0eGsXn6EQ7VxzJ7IINzqoMdyjQX2Xb+HKlt0C/oCPLiv
eWweP4gYzyV5Eax/r4XMjO31VPwVExdMI/XpnngOxyFqek49XF1PAiC7KKJ2nHdHvPj9mlZUND0R
GliuAs7962onv7jP5RvyXv8T+MI2hmZVMIId4J7fNoMRCejbt01f08GS7g/qhUKOH8UKDZyXfcwS
KJWaqcGoE3YMudWfvqIW6/0MoCDB/Oxhp6wAEhxpxPM8bPDTj5lrR+MmJWDKfUBKfw4NL7nYF16f
HY/RA1OPihQW6SpqTWBdCZBKq3+4lUq/Xj+LY18pdaD5FzgKaTj9bAYYAuvfrIguFKU6YMUFJ8pf
8UuRm2Mqg75/htoUBeisKuMWwX5JDnDbKoz2Kh1pZLMOx2BSYIung+KptEO3bq3fL0+tmQT3UXcn
m8zW1bQIgrtYc7hdJt3wrfNK5EdpmqpjGGzX5Q0LLUrlbMIW8c96wBSw5yHDJY/8PQjQIzdQSGE5
7CF/awgbuXgVHZMb67xI/4C5jdckgvnLbZi/O8fXl7LSYUiiPwzObRun1e8UycF9Z/pWpbdnCYJ7
2tyDrXoVbJ0aFtXqrJFWr+m06Saqr1Yc4PsB86BwgNaHrn+9KPFBjT8BA6PRTIMFsHEOUrkmrqOM
T6WQzPcY/jHAtj3/odEjG3Cl9+iKumX+Cp9Pu2K6xdq7oF8u7jCzlfYaewGFY/0Vkw8lbWfHy4qv
ZIl1oHFetEMWkORmLdO0t6iMg7DZmklTUJD+RgSE4QCYJrB5CiyEqDxUKbsFqTIrZNhMI86reXZE
cqQOZDCKL3ZObLmnHJ48n98BbUrpUy5WkZbs/1qN5/s61FG4pmshsmxRFRBAxuYDvJQANhBtNVHs
HZk0Pt7aJmMma8CEAOnXumoXiJ2dPf0p/63yO1wRLIhYWqFnFEts0nDp2/xFHUy5CfdAOUSyr8JF
+Paq+a8Vw5IrAN2jLYzMDUQB6Yb5MNNkU7jzSFhyL9DfPw1KSje0rLq33jSx/si6QEBUFBLgtsHD
PogUdBracA1AHvcABcozidPze6ljtKngfthK70Xj7iH3SceRU7jfRtRQSm4ug4uUDgpK87Qls+jJ
b89EOnlstmxnIS3hIkig5O2OiKzlWA2pnxe7Ojk+VegG6IgIWqDOeFOuqOf3H55pto9M2rcVEg3Z
K5f4X1//wuviXnf0fDsv/nH9ic2qDO0gzWFE9I7vWnzaIUQXHlULd2aTqnqOpWTQ1wk2ciLgrzWI
dt1GSoY/ZzsOf1pix5EmeuaBt5sVgfDkTIG9uM/ADLPwWdVK30MuTn5omKnyPdln2wRx3mNwfuk2
55f3SfqoOH0g08XItM8LB2Jz8WLWVULbtiKTjZvw2oeZP29Dv+7TSf9y7v/dVaMZACZZSXCSNBQi
bDMoAuZ/TJgLXyJO9AjE4xjbnYgtZvFFrKWFrBeHf+/Cv0OiJOqUbmOURXfAiMRSRMy2AwqDGVJn
jeKEcudRIB65BGuOjNhtCTt4iwp2+PMW8Wlvn+EUbJo1QXqkbJiTBOKUFgfaJAxgAW3LYTBKUXsE
RFuvoRQ1Z43KLGByC2n3k6CdUXV3Glq6IG8Yz+1UWsFm6UtaNmufjZdQjoJ53pP0Y/DguHSRZwNj
tLgznrTDBzw6oUI+cbnZ593g4Zo1cQwUB5I4jAaAfFDO75pp/EKluKvjKvGHV/koUXY9ExA1iWFR
Doist9d5l0mdPnZ42Yu5gWxEt1fi8b/fscPcs0785UDrXGfV4LsIv8bU1MjgDb0ghov8Bi7t1/J0
t5a/COSQOQ6WQ3ybsqPnR+z4Roey5ysVebkBwkvcWXzDXzHGEhGkzfV6RNUFEx9+wTufE5MX6O/a
Qwg0PhoXnFNZU0f53e8pW7Oz946nMnVK64aqbLZGHRWp+TdnGtSvkZQ+lwuxaKrNFoVAYDxjHLwY
UoaftvmW2weob3EvurU6DoM34xbRTOSt8h4vCiFJU5zssuLtAv09zX7N6ZTSNW5YnA+kjUnTfxz9
05J2xeXvcxDjxuY2u1M65gCTrz8ujtl/NUXgg6jbwp+QFhh/8EgP2CUdsOuJoOx2Xrpm+968FyU+
IZ8DvkutfqYZzt7Xgd5O2ej2iZrjaKTubLMPbwzaaEgQMd+OCb1ATUD2a9I3t+vT4uPysaOvxCIJ
y9Vh1K/dYiLnUgqRFhn3HhwhRepWTf1N+ocA0jX+ZcZcoPi2dmMmq64AMcbuunNRB487dBQCx30P
hE/mNisuf8JRawPXdTxBInMV01ji2r3YFNDTg5XWIBH3tR7IGsYYVz+hO5U4vjz5gEEbMmnaOjGq
MREgfrAzxbOgUYiF4KhMW71Gsxh9nWgAUHIgcwYyZTtlixQUWKPlqliuvBvyis20YY+PlRuZ75pw
tUNMX9/tfEAh8wZYp778ss9726i5D1knXLHIVIbMb7BZP168sF5x0MO2HF7jKgDXu3vWeso1qwTS
1ld7jj6ZDaWK0DJkwNMKwEt+8eu9TriIiL6xDlA7I+MoQs6jxfGtqn1xJCqugWQ6ROLUFVb0gxAT
Oys6vxpqJkW1lpNKPFMFyHIqM0pTy2m5iThtyX5nMP4oFFMsr9Guju7fGjBBQK0djk1jkF47A6bJ
QRrqTOwAyoKU7xmEjTvHWfeREM40x3O90l1+KJCpHRsCbzsQHX+Wrh58dxgHAust/2gE1qxiGGBF
z8el2ehLikZ3OHTokrUlIBSGgoIbMiGXZ1IW3PkiS2xJw7w4ArEBI+MBzyW6omDLHUxUFyvQd3XZ
uaQ0u6iZcavaUdsJ3/Zlq49EMk/6GjCi49yvLD1VmkaOQNFh28pDfK9S+ih0J8r+b04r5zkNx413
vTbsrMXL7lpUpC3VJBmmqP/kKZH9ixLJyURxwPfYRXeGkRfsBiU1Pvc5TZrVckM32TVgUW3JxqJD
DgUHRnYYFM2AMHTIE2FkARU0nlpAGc8bEfYYFYECKq4CvyPjqiahy0Rbu/8WSx1G6tyQZ6kC1CXN
wP6USJZr22WqUzFx1xKZgSX+cM8oDbab3yJcljz7+VBanSxESF5QbyeuMIt0ySYTI9I0TCwOAb0r
HlX/4ceHo4ZEvFEDbDcrdT/vnoIKQY+5Ha6CK40d1r+VdGbC/MGrl/COqCbsHCH7mzwpLz8l8C4w
Agac9grKnAWo+9UWSDKmfYNP8eC25bRSP8G0IWM8lAatcLogBSQ90thXqjqIqjqY9H1LbtcJ/a8i
20unBPv6fY6PlozQ1bmNxJQszWMvOVoak9ljCsGhJdG71jdDm1ns0X9gSfcs4pMWoFwCf0CWCc5Q
R6dX6xmekLcX84eO+WClrYwh1O11DbeK5qZCrl8KgPYvVbWGi63Vdvf7DCkSKM9G9Rq75pKe3OAp
WdJ4aW9ewC0b03F4bazTaEVRBWbAAkpQDtdlaT5Nmab5EKtcpor2fRlyJVE83HNSC9keYKB27RDu
N56vr1sCXNcaVpFVLs2vLDHlNm9qn36CkzFbL6h/Z9LNS3R6kDy523U7/eIhl9OlLyaGPRXcuWHc
Kc7XkRgDNB5JgVx1sEq6NxNcHK7RGT8x3V7Mfy+sjk4wpZiBSxBX1JMYPOoONAE78C09g/Ca+oTt
PEH+8IqcfrcKqWnhg/jIqs0OSEZGchQre9jPQmgosmal9gUOFosTQ8P6vbSyo2kdGoI5l2R+jmqT
bDWHVpeW2FKFpLTcCdjg1zFLB6Z1Ix7IdANg2cbrXjVanx+T+wI1E5TiXMpCIK/Y/IDCTfO68VEv
bZW/WaXOhD3yQyEY9QMStMN3asCkffmF6/4LQmEs7ZxIqQX/mp5Rt0jX7mp2eL5Q335ZlAMb9Btd
rSPc3c3Br5EeQoIa14R9M9wjFt9tcmeQC3epIO/L5ne1+MvQokrNyIbpoWQip9/FFvEPT74zeMyO
UWZ2cQZUNegsiWLpm6vHDIuDBiSlN5pubSLDXVSdYp5m7YZwTbQQLW7PUwUkPvqtCOVEkR/MPHdY
quJqCW9fbo556DZjA+RMscGO7IqZEx8Xo0e/at66IX4xLKTHVRn2MEcNdKCltjk82PEmIM9NA2by
vD0NCyEwLSuv0y3F4NW5o/t0LmF3vxvMaxQSqhfw9JRTPrV5WZUgWi0hERWx98ZVKqPIjdCGJmux
retXTef4GnxuT8Ted15jO3J4MkxcLE1GeOOeWHIlFxHjwbhbzM/2abm3h2apN0hQ1m6SVfzU5/pZ
rV1zNnr6LTYqCWvIyZPH+I0SaQ1tRziEhb2/cwbgCr7L9lh/SnMRudUV+ImF52LmfQ1qnvIeitio
GlnB9g8H1VCmpE68bKQknRAi7ju0HLsqXirSmiOQl7zxhoFGv1qYJfZ/m067tybo1uaYkQdWSHNy
hsBSABJPNSbPJZoSXqL9hQdVyaV/ClrVJTdJvwTmvlKxoFiqcYQD99f0SgYRAG+MyaMKgkChT6Z9
y9CDtTOvzYoQ8UnX3a5ILGfQOaHQi8M8im+fVlJ8vPyvf8jTrJH06+b4YvjyjwCiD8h0wZhiQ4B4
CQMNHAMfRCPFChIDQHvaswf44BakJp/4b78wsGX9q/PhSVj2aJHgpvjewcQ3p5ggnDDfLeUbkh5B
xMAhABccqRTWnXNa4vkUxcaxgJIe8xsY/+sKpI2tnDsKHkcqd7d7l7oUqwp462kFxaLzX2oKXKBK
ZPbLiDFUxrEj1oacUuOnyF3w3V7+dbucIU4VEYtWsHoiVnGbmp8qrxf3fpEeb40u18czHgXFxqhq
4CGTaGheqbLSNbIBeuXl9nRQ0A+6EgFNNzamihS+J9YtSyHqzVJBO24Y1qxIDDw7p6zH8DM8ux4M
2ATirozzRk3aaENesKzQfvkK4XzF0o697jwT3Vfv21t6MISMaJjOAfBx1qN8VjYhUlkmd4prwffE
tje8BbFF3X/k7fQJJDjMkdO/sDk0r6w9rUavLYj/4CFlBGGU+9T4dN3EmN1HW80eoTl2Xk5D579U
fviAc5dBDKTVOdB6DxoH84R0K9WFOUA+lDzrIEuU4quxeGVhwq+VCt857jU5+0iMVOYPCCR8+Zi4
nTKAEe9SxAPboL3brSUgONFcXkyBQZWPm3go8vXc/ZMZAUrxj+cvk6n9rylZEMYaalUhk2oHw2wb
U6hPPdMkhnewaVsYR05chPVS+3Dfl4FF9Alnmpm6gsRLN1F2bU4+QjNajh8bYweTgGmsxQmBnxqF
+CJ94zXSqJieuaxRTo8/M5Vg6ubfmBvDvaCf6ctC7OrcBEcTFfh71hvGr0hWL9jUzEI/mUDGH+S7
2f4Lr6cLGqWCm+/GWubcaqCF+sHp30eNsA4FxE2FlB42lpB8F/FD+WmARfQQ6tThv4HVhj8OB2ba
99Lb2Q1vmQHU7aqYunWGErHYtwNvQobdBBXUGa4mPfzTqgBny1aoRl/Rj5S/0N9LmEWrFJ8IHqRa
9rppkaGR2YwzxQ7M3+RqXRLg0Goh5T45nNTq8/G6OiwNDGt5+cdK00fL3WnmUcgltcfvp7/ToG2c
wKKKFR3ZyxGFzqd0GgiWvkM7IXJ9e4NcCwJyNbDpZnb4ssyDjeAUIMcXxBAbLMGpmTnW6eU6b17c
1Cqcsj1Ekzn1xkPVOrbxj+hAAWe0iCiKkwKZC5d/hQoBOU9WY8GneCBqNKyxNO4WD4NN6O3C8Lgx
LkJv3msXRUaWmFWzgMAm4Kkyc9B7fq3EeRK19XtjzAWEWekD6zWjBYd7UQbIxhnqIrtjbAlGx0NH
FOpKhuI/V7CJY2mzRLakX0nothOxGf6iGc4N7hQnHKVTdpkWVGGZO5tNFbHyhvxikwdc/+N58mjX
Bt+CJcbcxit23pHAR0PdydVq0mSUsCBlj6JWHN8qBxlGVjgJzZbnK95C2P5WfDXmtu6zkn4bZ90h
/5kL2yFGLJR0PDfSF99cTno36rg/17R4hXVcTRnXU0k9MJWKasVSVqevjxu6jFVceG4udwTEWtGM
Dz1E3FnRi/PiGKK5370xqL8BC5Qo6lyxZ+ZuP2XrdmFcHISpjrK328VGSYF9y1sssUpeDZ0rWg5n
/G3G8X8jqs62OAZwlV+5oPuBSLryffeX8qv+LmNLz7hZKx8yeaLdit9l7tg2F4XtO5i3bZURgSlP
KOBIiAdQfCfwBQ2TS3yg/xH7b8pBe4wnUNxtqGRgmTMdVcZUGfS57sj7J7cld7O7XvKFCUox4GXD
byjt9G6HB5aI2XC/di14BECuA25l1uHQo5/HgrnMmn6ewYbnEedrrRGuLaTXtiAUYl3KL5Ms/P4P
8ZrN49j+UE4y8ZN0epjtr2JwMql70nQP6KNRCHYMuR6QMy+X1vZRSatiVCNLlG86jsAeLDPze3Lw
pLmIEnD6UYKMRAqQxpAKU7EzDFa7V5ta8hAPSaArJtxKE3pJqbgn3+PXb0P8dLd5p8USXSSQ8WIa
o4VRWRwPklF5dBSflAgNZHoZxA7NMK3ECRDl4L230DXEfRimHqirTRcxL0Hlh/BcB1jOm9fl32hU
jk2qCmvjrujSYET0WeXJ0Q2YFtm/5ynJjaotd9C/8cli+jBO8udsgZ7Qp7GJJwzAoP/AWLrhAlZE
Ni+oLuIgzYo7ek8q/PwdzoCdvhuIWv79bG+yhSBJLKWzbzxe0BOmP2ngV+hchHrAUMulofYUvNWH
ueZ1WavZRxePq0ombPpwDEkGIs7DylRKfb2mLsWo7q5WuSmvtoij9usHfbd8Do+iqXfVctGQGGEl
Sgg89XVh3blhQAke1Y1lUvkt8tSVl51MVTCQufbgZkVfT9+FAwh2TKq6sfH6q1qwOHkU+JXTvgWu
W+57tq1/+wM2F2HdZ6u+3LTwKDL0uxvOOnUppuK+BA7VtzDnyNnsn9K+fJLpjY5ULgIxLVrSBjUB
VxBGWr8IfUffMMVbIYIDHJMbHAbqYWgn83cY3GAHnps35/dCHXEMgDnWfl4hfMN/r0L7mdvvKKzJ
6RawbpqvIzAlyHF7McRmAGc8z/oGP9IgKEhaetrVrF1c3BWyvX/EUvcYQZCGItTd5FTD675N12aq
HeIZ2i0jk5eIPLRZDVLM/QwbUeW0csqV26ZaltkCghkWGWQUWTHqKjnCrQjHhgRLzo7srjnQhVhM
RNYdTudBJaASdX2M/NpI/HDlJVAvcAmcAR6MoAjqOX/IJGbMv5G5/VFiRi8Ye0L2JCke6wbmdcOp
Szw3XGmkqsfIend0oXSRSIl+xz6XlNm0EVh5ayitM77QTUIdLa7z1DGxTRSPq7eCBP4GMQUe5Sen
oATz4ft6/zzSPmXi/p5ZS12F8DVx7s00M/k6Grs50/aLJGXuXir1DCD9e/RXmlDxfXR1LyNuye16
wP1SH95lRXMqQObuumcOnvn8uSoWuditqv2bRjbc/tp+OPLIPn9yyNOxIrvq52kvdeSin+Uk2NwM
kvU11kQtLV6TAz6sS6xKwntnGeSRsROEKVk7R0cY+lLeE+guetRTr4G8tVSV65KCkzE6vF7qK6qM
O+zgCGR0VNDPjv+DoLYfySXMtNOsG1YizI3CEM2t3Z2srn8idpSlPHypRxMAK6ZDeGxnMEWe4R/J
aqupk+oq8nwWdJuBLIsprQKfJUks3e0DI5mjhy+aSC5c7D80IJWai5Snp6Omu9ZrVrJBtHPfiQS8
EUhYM7d0bqEoou44rWsXvP9JknNzLtuTnLB45qbi01eFlZ9MGrzgKPkIpxd/aBYbmydSTOeaATUb
BDFxVOziUZLf7kwBf/gZlSnZQmD/j1/DSJ/XAxv/VVPItfIL0AhfP/O4Yng3+suKIpDUqrWljRja
06QE6CTRWb4qNo7KimPDVsYwHSoSsBtm82n0HUH6jc1doOBQDYXeEuK3IovUr6GEEQKE4ZhFLtzx
Aspxo4VNXMlL6AcwJooX0PNbbyagbCO849Fy6LDmlclzOPN3v8tfZnz2NGPNgzIinD20Xa+I9KJm
e9lemvswF/q8dT4ZmSTCHsJfwlTVgS4ro6JFK+B9VqZT6DXpxgQmTR1DJk1TkDdIQT0eJH0URjvM
cece8b24cy0ygT/SA5oUhVhSQhoaywE9y399Jomb0I+Urt3acBboLHF8hdfVe7ra+/1ZbJpgK5Tm
GC3ySBzoqQ2TMt1QuNq6FVISBAYRs6eiYfIrVgI6ud5TNVjQJwDLDWHuUiHL5z4ExaSXitIlpC7K
CuwqZ5S2cKlM1SZOFsItGS7HbjiqmzsX1WaKF2b1ysPcApBd/W7Fb84scYtQz6sjhq/6rylOnlu9
jgRz5o64AXGVwhD2RL12jX7HA1SBJXITzVWtzHHvfPC7IZUoM4jpxL4Ikh4W7GX5lmkWbw4gIh+C
H+gzC5wo9IZeQRXFLrtZIfjrvpry0mQ+gSnLGUB9PX2EOi524f448rtpKoeB0GkcztA/CSL716SE
ejyWqPv+f2caSu2FsAaHWWNwIifqDB3ElyugUvsiccnW7bmh+W3ROQIOvt6YT1natx3N+7X9vVUv
jao4CGEHQvFyn2aSu8FecJfCebK6wO555KhmfYByEeplckRl+1tHgktFpoosElhjk7O0i0e5SZjk
TW6lR4O/TfAbN6NdRonO8g702lRK+riBvznuwQRNuIvwhHGOXqtA71qS1tZbp06yEXWDXLYWP1vK
TIsZuHBQ8l8x825orztPjjR1hwteE8iB8YGeDI8rf6ih0jYcO4QikPvjrFpPm4ABZHzxBRpnuuQp
3pmJuQZnqFTW+hl4xLW/WNrKIfgkFwXimQD8j9yRbG9ADQlO8LEtyj3N7kwP8gApl1pzWWqmNK2L
rTyovxfxfho8bHV8sbAMDo4+nYj1f007A/js1anKcBUolVnyoWylj7zdRAxFwLksis1FXnycatmD
51lwMdDCzJ0z3GGpkNrRx7x+8KG4bBVlWsohQaVuUixxpTiRzAl0qIiDLCDMLYCm39v2HI9wX0va
DpedwNKtuh9PKr+/SVEWrpWn7QE92VN6x7FUFAabbZ0f/WymjY7q2ZGZcZJfYjpU5CisnEInrIgF
+yeZ30cmK6/zFA7L3f6/8Zwcdol2YK+qJN6qEZUWgISzwWyvfeydOZS5o3xozuc5qre9A5Y1IWlm
aKoCfWpXCO4neQwEunBs0u2LmqUpJ4wS9nmUgAvY5qvlqifeUm0Z6WrYpxijxYc/491B4Q2CNZZ+
IVEcP4/yaAGEPeOo6nOU7XIg5zy9GLgk24p0trF1tNvT2EkFb7JPzg9tmU5S2yMp0QSLyLkW8x2d
tksweGAqPBnF3PTLuRIqkSwaSYCpsCi7u5mrWxSweE+3mUCVNOAGOUsi3uC8oD7iJcg1F1lRsPkf
5orqHzt07MKQyDq+BaZsxr0mFtIfsw/+0Sntftmv8C1khKlt3yWVuX23uwS0QaVcUJq01XM0Y1pD
GRq5WWaCZxJ6jFrKl2B0XJPhNikc/mxkbxhwLduHkAfzLT7rU4/YUdVf0bIB0lEpEWq+BBZYrhk8
DPxfIWVW149MUyrZSnZqdWSdwd+e7sKUWfDjSq1mjovI/5JFwOLFHPvuIwWfQ5N3FN8PwAGwn1M4
TYAGFSOx1p0ekUg9l7Skhk2MuEojIp9cR3Hcbg6G34MMZ4FwGV04PhVdUQ5Wumpvdoo9dtNWcSCw
F9nvLIBp7r1tzcwASyN8kv/JRx2/QzLjePv9MJwOCF0MvN67SEka/w8wUBujczd8uscu34mBYCif
6CwnalVqeJFmJO0O4YpT0T/G/MNJYF1GAckZyh7NW2HIr4NqoG5zjw+75OEXYWtZx7Wkj5HEgiHj
m2yvv/+cW7VnxfZ3+a3wHGBnxvcUT99/YmqdcIQAEgufS1+WZtLvpjanuSgVLRCe3CGJnxT4Z+k7
A/K16ZPGFJssYKr5x6mdiGJh1zwnfCmDrHxdE5c9DGfG/07eh2njGes36VPKPUie0q8qH70BeZxt
0g4MTAOxDBumpTRs2jeScjgsMXEsQ3eWfgKWl5YOBmoL28EPsk8EEjFbTyQmFGLT33zwRa/1MQ1j
DdL0rn7DCmUgTwvYw4wWK+Xk3HvCBxfpDQAjcRLozxiYFfX6JYUSxdYe7jDGOZVLfpV61qZ/AknD
4lA4PVlAyq7TJ0ZsdGp0av3ZhWLW2dbw6dUAjKZhxu3rZUi7J7cm96XrUOKHd1qiR4auhNp3XRw3
FQCreUUQmx6k8S1BlKAexJnmbSDNn+plvjgn5MCI+c4kaMiCKVEYvZV4IVxT9skJ6AwGJeiwlN2z
9wTgeciOr4ZhZFvED/yjXs6BRVcC9jwcKmS6b2dfAx+iadaR0QODzKxqKhloKP9/poxqooHv3St+
wguXn+YcY/ee34rgpGxrVX33ieEFWK0IfKKVzymSF8v/KF2zVL01pd1WvEYoaY6Mdr3A/pF3kLUK
smwV7J7FpbcwDZ3t5TgXHTMnrCx0ZJCohdDKYCX8/smwiTDtuHf02G71PeYjDK4zb+AeiVyZ5EyM
0Ec+JdEtwsIuhT5eZSmRZy9XHmwAkCIrbC70VMxtCnCGf3KH+DX8vY/lfr86jCcaCCiumXpjjoeG
qyUn9OO5k90QBthUY2tK9X/D8ng3HvffNAlPJV9hTnoynWw+aUczV0NvM4uBhFlKpErafLo38DFa
9IEgrOqw5nFWhXsPUhHMEBZ2lopn/hTP2TBsn0/sNjJMhw1j1k128aDywvbcPSF4YZehduwlOKod
eI/quqTB5kUOZ20BkmXmBQzd4CZCrYNcxeHonbCX1Rq2IEfUOzozZmQC8QyAiiaEqFnSKivoG/8B
rk6N23We+XLmc+0Wm9pNKkxdiZsGmZ4h08ecQUDqfGhL+S/ZbQ5PUC6rdQujeXtf0nkfA+UEUpz9
BPVSy0atjQQS6CJXIKYrMrZ5ZDntWY/zQvJspzqPAubVD/M2QSmFZra4MGjhMGRjMDfSBKyYDLOj
43e16fkly4GEUYQEXiLzisZxImrMiB7O7k+ScdMILQJV1sYmvecIiB+ymGKZQxRrRIy2FTQS9Jt6
jyfnD6IoLg0UJZ3JlopZzJRV+LY6ytqc7YIjQbLbB+sTYq8IHAZfbiafDLo0uPP644d9wq+9R5iR
F86N5eHgJMRCm3BsjLEW39BKEAKUtvbOZENKqn4vXcJgxf0D0EEKS7MhHe3sT1qLEBM9rkAf+1SW
4XEhX6ife42F8+FgXeHjDULpP2rGbAcizorvkhswoAf4cwx8jStG/J+EIzT+nAF5ooXTINbQf2PJ
piAtt2gRR24bTzO3eF37ESZWiZXanPQz5Q9g/SgQSyJqsMaPzHwGxaRxMb0gLDhlaf7YO55q6rPK
jeyTHTsm6RK89fVnDp72b2pTYa6gicIHc1hLXkdDumVx8Uoi/RMMuWgO034Kw8s26veJG7JiR8N9
9uaL5rkj6QjFw96TDzsCsJmI26uAWUZ5Mpk3L3wsf/OEhuNdXuitLFSfwW+oIdQ87K9T8EL4a55j
AulxlPep7Q4BR5oNaLSc4Gkj1Xk8xUD7stVwwOhDDaeQxpmqXnFuyglmpxEF/8fOXdJJQnGxZi1a
BKDZG6tucPt11gc8874ONumuxqozSrI5gxV+V8sDAVOZ+Xrk0iXr0UbVncqOZkcMk/Ng3kQIXsFE
aNtNpNfmhD1CXcszFHzRw5kz1uJRgwemdgFRkewIq/IRyrzjbCB7knBgC2S3/ls4O+i29QXcF90e
XPLLDaP2YCSmEpT7Mc4hAVXWQEhJySzP/9jHQ57UZ++pQkJGMB+o0ric28+lEFLciJdeHFEYV0if
9mFMgDcwFI7fkyDw4M5/u0HHohVq1d9izjkt91zfl1/D3OSBEacfgJN18XFrTZ8xS8BkVavRJDPO
FZT5dJAwl3kaas+OD+xjxI9PVgv4Dce56zoylpEJy9HnzsFRlXV6Juyxn91ZELHIP5dHwKyzP0v+
xroQvsTuBUw6YRsYAewcO0Xkj3WPBxw7wZVjrTpc3Rqfkg9obw3GcIewWpvYs9VHJ5ecFspeuHL4
x1oA3xsw7uOIvNHN/3XTUYIURG+NtEsiupykzCeX3RbL/UIq+7xFxVb8Ak1DrCKnAz79+V/1u40Q
f/C8GAVNTcscpDUiykphU9ULxVq3loYxhAtEcobUOaUUWDV2u5LUnXAzIuGv6Eyv3fZld26zM7tg
gTHqNvsV1VNt5VS+0VnnzfbgOKxC6jb4tpnnjP9PVwHtir0A+a5M76zurKF5oKvJk6JePExa+vmd
bDfNr9mMkHDJp90ykRWnV89o37p7BJWT0e9DHdtmmuS3LW9I9wW5zXPNovsyHXtrIjXkcaw814qZ
mTUB+6vGua2XGOSlUq+fWo7iA2I0BnFtuw0wOh1jqSEKVQTkgIcqss128SlevompzfQkp4MfgAXs
JDb4YwZVgAEMBUSUWZm0vYzpSfgyB2GhFvNTKBFCnreeHKskxMYC/Mos9CUfYwqw0YIZkTMsjPMW
I1ET2iwD+p8fZyKHbi3vV6rFCQqzn7VbBb7/1GUj7MCbBdCTX5ahnwJ+pv04ExMc1f7dWnnqh/pX
38CRArUTwFp3tyFlGJ25t5ir/67FkYGeZePOXL2lu0MqbsB13p3nT8evLTOnhQE4bVRHeA7hiB08
yyA9BEaVJzeiTGMXbd1KsPSSRlovhulE9+aGlJ/C/zUd0CA/mFiLIA6drk5iUOByPAGwqGPsptCg
Op/AV3bTJ71Of1auL2at5KrwYOw2cMLdKN8a3Lr+JNOHYq94C8Q1SMw/LJmQRre7dwzmErdTZGTS
F3e/eJTUnpy85TapAgNUXoM73AGllTkhyV7OEkO8yDL3iNGb8LMbtnVpQQpPyvyyhMxQD02YowI2
mE6ZyGc+73x58z6PSgLmSHAWmvH/nfsDafpCjENrus04XICMuMb0AHR1rZRC2AuehoAM/LsiG6mF
VUiv+TU/Pup4mSMoMRM6iWHIXgSC/85R8UEw/9mDoTRfbQ6JFezbMSVN2rzRZy08+hqWUlOsjfaw
AIsh8kuV8a5Nb4/m8rSomTIftCrvwf2FNGpiLtqfBpk8UDMpWL000wNL9CYyOgy2mISo0iVxbOxE
hsEK5iH1V9lrgbL25VccbIRFZ0Yspnj80P7iX1djD12DQ+VyihEtBZk6PvbMpUmhKp4yV2tXWUtC
E2tKEw9aZDasS14WhBriG3buvB/2JJN6gy2k007AVc1xpoQDr9h4FCiTaR7lt2adxwP7ct7DAaYH
fvK3ms/0+PveukuiPY8Lspq+h7Y/i0YF43dwZ4SlIfo2CndZS3SkaMcWbIQ3zMnnbbq724KCCKK8
5Xx6nzmQ6JQdq7r+UzJeHtCThS+wUbF6dQRmTVvtv01kFUTTq6ex0KeuQbUrW4xZDuW4y4X5EoTN
thRS8DOrev1mWnt2Zfd5eqA+RiItDiQp6v31m7LzxfQd1cvS2D3gOESyN8Iu4BtbHjB1aXrSuEro
8U1JvJ+jM382J/KqxOgQgcord+X2udC/Wv3938DOzmXU1vl1bsHvu23FQdumzwjb/BInolYclPSh
8HTB/U6icaa1czniXgmUzcnnzEs+hYZZb55aBwWvKcT1wBYO8dSbDJGlY8ie5T12Y4rWxw2B6+Dz
Z4Ahm1uns8Wt1g2eH3KiR5u1t33Rxo748wCK+nSU5DJ6fETwDgkRaW7f6PajA5y/0a3QfRlNEvpT
4kUf9+tUEI9QSbxlgzhn9vumtlfkpvKABo2gzCg7XCxlUaAOuVKb2jjgoF1Awg1kAPUyQhU3tCnS
PwwNCzheylJF00FNp7bRgtq+N2Uzcwgki+NOFmZsLNDckMWChvFRiHvmSJxk1QphZmkLtAwGYlFz
WJGaHY78g1YrVvqU7S4DNphR+RXzAee9TVEphJvKzCzkcu1JwKEQGk/5SQGOXCQ2ivKiihqMpzwl
rHei/mAezrfAUieYx3LNWcvzAuX9ldW1dKFvnsEQZcf+g2ohfdnFJ5TwnP8FLfmbnnSjjEVP4vOR
6F9c7P74kuIBFkReg71hWrXwEv6/xbj5/X3fVkxq5HW3pC0wXIU+106nH+WWTVBtB4gwhVwEqKnu
aP7HnsEQXOD045TYIULTnWxVX0+Rs212Wj252mPBk+L83OCpLi35e1A93GluW0Yq71rCQcyBtYES
cZkV3OL6r7jVDnq4jgOh/uSSuH8m5dX97w6Ptxj889amYigu/a7R32Ibzg6L6cVxRWRvX27yRsbx
c8mNlp9E8AsgWKXB8eMUHV/ywf240efyuOK27+/bVnHmIsgS3ycKd6VVBVdC5WlsrlM7MWFPKoFU
0t3TPklt6sOjnDvPssxS/eLwVZC1cZZhJ9EMOQ/z22ACT6ta/4tqb0Cfn4qSmOD8V0c3nFDPSHT5
1mZNw/yf1XVyLGJovEgNtlbPdf6ju/7NShOfuOhF2M0Ov6AzoRfctUv1hRBN8cwumZRn9uAdp3Nq
o1nq6xPzyY2K5wueRiAxpu+xTv93nalreqIaYKIWd3nK5nNDyb/FLW16dGZ7Fb15WqrlMx4/bJWz
pCqYyTU1hUgYqC3eGFnWG1NBWxvCavBAUjW+lBFIHHjmKsmBhusB/PrMDJrAFvmbaXhhh0eXjfop
VrfMr/Ke26w6E81cZMmoV7m4nPYPUUT/U36x9GbZatnaTFktIt/8mWBUaj8NmP2DFM20zM3MrMVP
P5e4BmC4Ef876idoiyVNdJ9tmwnuVi5sMSJKZopnNotMRqu4F4CVPIWNdIEC22aSYZltnm3qKtPv
cbo2uRsCKPJnx6k+pNB65GauEM4iQH/kFbQka/op/4wgsg3T1BIbVo1qfnXjgdSByUlKC+jrM7rS
dUrzJQzpvOOZ4hCZz1GC5BVzYY+NcNEc3VXqiNSD8cJNfxsFkEA+UREQ8PdDwJ1E5mO/nAJcqNjV
RshYAAIc7KGxG65BVUgHEubjb7/yTjr1h6u8rsIl4hpBQKzBcQmjyHkgOr5lxR8RB2ZQwDjVSI2G
/yq45MgFvw7cuH06Z+JX/KH5JzI71C6BgYGHUXoNWpCATSlTh2IeulJ3Z9TuLS2cqmBsO5xTiw/e
eta7iva0qh7+TwcubdJmrFNiblgzoTr7kqa3CZe38KhJU4tYPXGKlHgo4bIJwcBllgfGjfwzldys
WPRDTFAkcYvCx04PTXn9c7TZ8UW/qVdZ587jJN5/vrJy7G3oWJwiVHfI9DR7AXRRDEwJsbi2XK+S
WiZrww1f43hhpze9Vj29QfzKfF4KPopwmu1jPKjcjeoqNHQbFA62+B/6w4J5jzyV5/0CFkxWc8ur
7LJ87SPVFZBHYpgqE8FwBo3kC0Lb7kSWqUd0f+FVwGWy/M0zUK3NBrjFWa8bLL29e2KGc312L2vH
K2PZPG3tfagF1kx4iQW5QozzJbR3e+hWbpbSFGymlqtQpoz2cKqFfaiAtA9Irb8ICaa29rz4D0G2
0wHyGV+za1QVkK8q6dh5v0Bl12th2IJQqW1taCFlJfEXUhpK9ID3GzYfw29VEjVSxFMCLvab/+U3
/EWR4RnCYmpBQQxN06AH1yEXvtk8UNloUslGzoao6vledPC/kNanv/M9Kjof8J8KxaVRTMb9aCMA
diemjzMAzW8/RqZG3t/Ldn8QraJMeEKAGQOLAU8U6to0mXZ0uQuKIu+bhY4VYLurMRRGDZqqGRuw
YdALJ5xIcnHDRpPnvTKulfKUtc0dyK+WsjjEbTLBhYVpwsE6bRwNYSO3i2fCN6pwxNE54ASfZoNL
Kf5PlskZ1ORY9cTWOVuqaHWzxP5h5UwrPon1MDofWvAp9Kk2DH8iMSfoqXHpFPCqDcB2J9/M62t2
16oHJuydqAjbJ6kHcAgqleLzv+VoC/chKd0YngrVlvOUTf0PkOQZiFJ/TPJNeyaoD62U7NfaQ54U
KyXlTDaqHwpDkQsmpOCg4wW5/FjaBHLlVLU/H7h3yVncEyoI96UVFbTLC1Vkf3Ise7cG+uTc+h8M
GtS7Cz96E30drvqbv/w4N/lEkVEejn6mkN1JAX5uGaGoriltya7EVtpjQ40xdj7vvxVDIWOtyO1k
0dBxeuzY6/Ja7pwn+eZJVggNf6mhqdnmlnQ/jkLqKltwtmhg+itUv84uNQN2Z6M/VZ5xFQXkMcIm
IQoFXb0Hb2OKU70TkqJ3cyySj7E7dSbjoomcRT9/kp0XxpeFxLSv9v2f27FZCgUpvYWFVPvs5te0
9eCPOz2/jO6FjG4ranY+BURRfJB9uZTzMDWovxztw6/q5Xf7pzwkRFfNHpAuYdUHPQdW4DpmZoes
J2fRXbNDYUQO0twym7ieF0evgpk1Spd58APO4z3evro/3ZgKYXrYrJNBQSOwwwSRCo1+tFq9Ot49
geD12jBqtO7UUkr9xFHsHbTsJA0JAaYfypSsIIDnr0efehurFogBN4ksrL0Jl0pMp+RwzpQMlasI
vr6SawNqE/JeSFlHtYh8V9Gln5fC0PhQJxj6c/2q4kR7khPXDY7SnDH2MXXKX5aquRyRFrEWKkYt
FlI0S5I0oJxG31SdoJopGDFQYMUKGteXM5LMnqd735bK0pALt1JKuXRWZ42rr8zm4eOvMeT3JgKq
8w7omKEyOPbqh2ghZfHkgqdfkbQ4gitgfmiChukhaB3EiPL5ODyW0D1o0hdNI5rneaEaLXmGP2Fe
bxyvygNWSUeuckL5dlnBSm8XBx1lfkPnR+yTnNpVl6xdxQpXnZcN+JHUGNiJRXNpQdPEUYokExsr
wqlwEYKcLuZrdp1rtGOTINwG4SXf9pzjYOH4382XPeANexyR8DCsejakIO47igZ5ej36U3LDWhC1
PxJZtW9+cw0ZnB8pRN0My3iDlGUbUaneOvN8MNkRqv7ohW1fG0UzKydvAzv33g1bF/+5+T00YQC/
CKPqful7Dv/yXZBcx/N6Q1OmYBaPUKmGjsXxkk2EEB2mNYR/eNrGKuRFbWhebc25OzeM/u592JCl
oIUKMLbm2zdPiDElY3coxVM7ogVZqbnG4FeoInyB8UIuLgElnWfAkcLOUTXwuoCSpVxBf7LE6iBZ
FNTCdvO0facOc1QoYTDUkeSWTybK3evO2xvdSmm1jJA91CB7S1qDZZ1lWK1shuPXpW+qvX/P4Xbm
1WvEEtJO/o6L71uRPeYb5jeOxc16uxSGD2LuKwP0hNQlCywgHNDA7KqYIEx0zTTnysRjb8+vDDZn
CYGmDcvv1GIMzkQ4M/CJnlFUDe5csH+rpxPSIOrxIPzs7Fqn5ULmGfmlil05UdXTzhnYAGQCFy41
l7GrbwElpWPyukSP4kJeTOtUmZUX+0tsY5bttAsAJZAEZer11InhmaaB9LaZdGUnrd45zSs3BV51
qGt8rfsbx883oloFt9wo+0SU2ZaJmp02Q0bvf4UtOrll47uDxsbPHQrcwlgDowX4Udh5dLAFLcAD
tBodfh4sm/SVuUsMu2exQA2FmTSl8COg0z0bVquPNtG76phNFyCjilgG41Gc92BzKwO/s4vU1u7C
+4VNkQd3+iH1b8SnqbA0fpfQ6tUrITn6Ry7pNkXvi4UwuE9uqrAiBNANC0JazhQ7nqOfdqxFkao8
82um4JxPyduV7fM8KmsOGVzphMmd19/CPi99B6J/7+cCvt6/vRKYtflJ6Eoz7ZbyZ4zZ1NFsApSA
qUX8MvH9L/AXHmr4UEo46gAx2IL26XvZ44LI+UT46HoWaJC+kvCzcPZE0jUfcH5rVcnzIhtZlDz2
8Hgi8Li3Qa8uRdmsCtkEhQz5DNPimm9aKdJRmPyNtNMqmGR6nU6f7lE86PfO2yia3A2ApBK2/UlP
hBFAEfUy6ewjd8tpuJiWFzAiYmMeoBozzUHEi9W535wGvjqaEKDX8vIt5bjeOYCxWcKXXxVu3QL/
exANHZ3q3ReLPm5roVFrvt4j81muCLIK+vRhUsijv2BBzNyl1tk7w4AwLZkXootvTNwkMwO6b0e6
RywfOxafj0kLFHvfGf6ykrQLsdPX55TfaOyTxDJ8tCnakJJxv3Sau30BBThkJ/v8TQXDtSp10pGk
WZFOLBk1zAKjUTE7ySJj9K6zDU+jNaH3iOcMOVCW4I86/AYa9o4OBQkKsnmiO/SFw2JxRrU2EfrV
/C5r2up9MiiQ4uPBmWfvQvqTb4TBtHZds6YcqdZxgRFqt3qPg1ni+Gj0RxlEjahQBTH2GH9biJTI
+zOWKv1YpIQysUqbQD4/nw3ldXT+Hab8V8FreAWzhy8EDx90I81B9GWMq7jEKLe+qDmZ/mgPY6eQ
UWSwz6pf2Q1cp1NrzCWqV6yc6gccX0KQGMjsbL1IruLBueXJTZLViqxBJ6njUU1/HJ+IonFuWrjF
Z8ajHm4UNAX9hl8n84gUlN1X56b0irPUJCJQlyhW72PAquJxeOa9weTIFVpBLsxuQSAh0JaaeehQ
mDvOUnGNaAgCOBVcvM/fjLNnCxcrcrg0Xfoh3K8gxy4poE52Mtku2yW8VNPMrkZeodSewHInb7Xw
cd2++q6e+ue/iVN2BMTYodN72Q2DdmWcwfRMnVvaFPKfqebW6DM3tX33wtHK6Ze7vmGPZ4PCBuDv
FZy2YZor8t+JIIJSb8huJ6Uz1q0Bxq4cGsj+WRGwQPRYrZxCdlhTqEylx0J1O8RjDJiBLTcNevzu
OP9OypaFJoVR1RIcyFEPNJLNr72FHnzWUbzWHTgHRoAzxVzHlOPdtfOiGrfwmesHe4UWO8RnzGwT
aiD1OSFAtXoHuMaOdi6aueRnuQwt7jbAoYoVpgvbqjaPE4olSF4yFBMbG13aNOM6s1zckfGMoqKl
2/V16Sqi0paUzCyWb8C01TF84v9INIIGin0o7U8P2Zeswnb7vVIAjEv51JQfXq/paBhuHQPkCmZ5
Pn5FvVlrhkoTVhBDivvuZY9JAvScAmT+YKEN+YaLhlhNvNrBfebET6kqmVHqRntoZo9kvm41iWY5
UUVeJKXRS5hI6GH9bTHsL643WzoiV4p5oNvmMbRhC00WsVD8bwZrCm9cfSRZ5p1A59F+px4ZZHR1
XkbbV/HFj8Koeoj6pq76IlbK/u2H7IFPPDZAxbm3LH+q8O7o62BqqednnDTpou/M3PamnKLKzHsi
lGuv6KNa9eOKUiUn51KNRm9UxIoB1yKuAMy5jeTE+J7uYRBTPwLnTrMtdj/V78IF4nnH34aFaZUT
b72026fJtgHPs7uzfV/ORpM9Nw5GGFjHoZ3ql/Nxxf86X88f6lttRbdyaubeEDgFtUTc3wGv5Smf
k3GJD9GB7LGxYbCzAEr59LmZ682dBpQVKoBBy/pxZpKcH06SfGdSiFn92RujwLqYxwpLN4+OwzqE
nOvsjrnn6TGMY9zcmqA4AsZoEH1WJNeSGsbw/Rg6+Sj93ngBRoqoXc3+UrA0nzBKGbGnbMSpRjyP
sY6FTpN4a9mRQCthPfECu7ABEuSlLtHIEZHNXlj/MnkxWvN5wRWh4MaGS9ZSfD0jH7V4ZWuqxyAY
ieyJWQnD3ZJbtRJKNfRwuv0mzXgwB7YrmY5IGMnOCvcP2gZduDfhnHHbQxAIxoOV8Rd9t+F/1wLB
hmpKNcAaD46Gm1mBJqvqoVlORGSZ1n9+UZqUNRSRNc+m4E4Qe+XGWQ1PGWKk8i+9fIj5WX21gN7b
s94GhP+Xev1Pcm9ZFAIDtgcoxN2PrKkZ8JMm8HxpUZDXmAOR6UDhu1rtHSg5VfYIL2Kvp2ozgdoV
v4GTp8m+s70oZvRVCbgGbbSBBy7zfW7RawSZPv1KvYFVgqWdfaj20WunFH+wFucQdOOyJbOqp1S2
luUJNIitR7T0qqElXmVzSVYo3XFomuJP2+0+0rUI/h4dWMHpef/qGu4TFmrhQVh0dMcPrNMr67RR
uqQAU5XslvwNGhmmvxMovE9YXgoBbRbnePltu/ZaNfwt7+9aSgwhvnp/p9OOxwqxB3Bj71gN2Lek
9dJNmpidw7Zf7qj2sto2+m21NCXqshYzz2PmVYVomLedl3xC3N9HuVPykVXIAobEj/A5Xi0cmiMG
qOpUg/7aRSUTnoi4e2mhUuhbKJQfxvdYqW2Dq/92VNS2FnnC6z8CGjXn5MMy7gBpnFcRIJFxWtnf
mjiVInCQUvu0QITecu2KZzQNTWmc/JKpq0e/kM4wxfoVon6+I9JbRqFg2kI5UqsMvgjIkJqceSIx
W853C+bPfmpUJkAVuyMkgidrGyRv4ASLioMhC7jMA0oi0xpulBmUxLdjIHmSCclNmWySsJtKQmPs
PEkN/aEATAWHQbkJKtj9ufquwDn3HjYt4hfS9cCDcTw+KcPbpoRdMcL1PYCeVJ8eC7/hMqlEnjN/
hYnQrVyJtH3I/npgGaqEsxYtQg2Alcx1mrTTc1bUffj5kHSvMFWfNhNcaZCAca9I0dqKOJxMLk+N
3TgOx7HZnYJ9lIc7AbgPpQ/TYQOu3eMSNW0KPgdEJZNMHXlHmGVX46xAuI/0n+70seBYaiD9oM0I
VqxSbA7btLDymgbZSilgImXxlc4NtxUwEE779oT1NMaMD5d5hVLQI9JKEM1wuwczTI4Wv3+cbOhp
ESzjfUIG82WGcZux6jFxQqxx3oDo1wMtyNGIA3hWlnL/Q3dsBf2QI4okQ+J19LMu0xOHWgcOn6ZM
gykBgEKpwL3+u1QdWIlHGnTHShO6a6/OrIdC9rhbdrIkanwgTMrEPOqrd9SuuIwwKTcC9XvtWCMk
lgBAk32KO0z1KdJWQmOidcsK5UTleecF0m1SDlz4wgEZDAejp0rFpLsTbiS9foD8KSn9Ik5T243g
qPJjDFrXoUcDXfJGHnuO3fXFw5K5jyRctNGogrTOgGXYtmz2cvp5/mi3uDAsQ3rq/Orgx9b0113G
o+AXUH8/ObbGrFs6ITPFRQTz53vGZYuvexrhg5nzBWzBhtklti+jIjWFROUlE0RCn7cCJ62a7gNW
Xil89NgotmvD+1bbOX2zwy4ssTNfPElJ4LWp22mIksVIPr9WlUCwfymkdz3ku1gYZuSymAunpIcz
RfwHCwGOJQPTp4K7UsiyFtiVb3A93j75rW4u1/XG8enKyCgHTZRLa8Aa061Z823rMT3sdKhSkkSR
79LJtrvoAxgnakCDbCHKEByFQ3URZrsbcI/jhtjjP+kyxPTlb3udboHS1WbDxuGq8VNCIknALB+S
VUXrepCvAxHF1lk5Na17j5dgBoOH/wG3/X32gXQ2mF1E4Z3Ya29z4oL5zJLrYAQZQEx0fyYjYY3+
CF5DhCnVHb/umw9uSapEa44KPxhLjQYXHTGbj0xbZy4rry5P6Sha4b5V77hLfjZJhiQLW+TK+Thv
zoFEotPDeVvYDNAvANsf7aJQe6MZ48YpgsqjETLebWA2jUsdCu4HDmPyEpLeexr0SzgsKJGfMTjO
i2BjAoI6+bw0WlK4vJkyhTHXYVgnrLRxOlmVL0rKpB8ROWZuAUccblknKe3TapuedYGxwNJqLoBo
hK3hoUjqiXKay65PF3P5ehRo/Q6oXEBI8jgZsnD0aACbpi6KSNOSoQno6d3BZtdPCU6ifYBUU29m
FS3EcQKXjVhwUvgujDG1YE8GSonIyKOZL1vSK7HNogUapFFE5e+b6H6sraEFzHrgA8bKFL1xofzm
fmEYp8moQ/i343j2d3CYvlSECCzOZ/nZMV1TUOXlNFP2byBQ82e7lsLA9RV7IT2zPPGRFe3UD8vp
WTl4pMR9gw4nVA805i42rNPlGgbRbAQokhlEoPXYIh9BRP4lLBPLCATdc+puG7uRi+SDLw4evM7k
utc9+dH7iEQ5Ks5k0Sg8HbCMxxf3h1stv78jw4aHTAsWBN6QJp3bMFSnVPvW4oG+iZt9z481NYgj
48p9N22DDvDMd2STCV33s5dnS14/ha+n5QsHGRRb52TvdlVGGqXpgsOSqPRvNHbsLW8B7Z0u/PaE
VZ72lN0/3SdAMmVF69sxQxlA4jBFvZ62iHPHh5pCg78qnz9HjTIxE2OcPYqS85RdvrDowRXSsUJD
UbxpW0Agx3p4OTaaZdEKg3EaRAs6WspYEAwnMpd3hqzfNKUoRZnhPQJ4qAGC3yPG/qihwmLBsv5W
mRjSurOCmn9vBRoFyhRV0s/xOjSO9SD8Y2ZxSpf2ZbwLKKYyUTacRzDHi3BSOnofwFX8cvVLeXl7
SGmh8oLy96UAbzzW3gzHT9z/m4jZPR61IOBJAoOf3+N93uj9FJAcONxxKfg3jQ/tKB/RmAKnOSnG
c5h22bLem160us/Iq+7moj530NSwHQfJwQ1XXqLP5Kigk2tSa5fR/3KQUexIxeGQrZ5+4syJPc4Q
+8qf4ZGUm/GOnyZE6KGcbDARzKSts7t8ryJr5vZoABwbOZ4RQpNkSjP6FSCK5uQGHIMv9SZSoHi2
jxJKs5jzPDyNbmXCQXOfeRwkhattOF+jd/BTPHM3yE+WvJxp+RVLWtXQZvfJaeg3iym3YoaM9A17
l2y5jm9SGeGIWGJmpcIgpHTd2uhfF5OJEzfJUZqWKmmHtxN4GCmIDxsaD17t/wWIwLAGGluK/Wre
ePQx4omZ0wdQPDmEvBXRPyWXV69BxFpUQuWn0dJSxUoxTLP4bnvEmGgSc3KGx3yhp93nOA90Fjc4
UVO7NP9v6vhIgOhmxdpf1fIaMilXYYjlY4OGfZvP7fLZCuyOsbNrMFdKOaIV6R5DpfPOYfCW1FWa
F+oP7XYDNPe0zt7wd448lnGYuX46+9f+QRgpXrhfNtAxYL1t+mwJb5TEBTj0nxt9npiLRO/E1yuX
YiEeyLPFW//xStLbCiWHUye3uNpgngBXUrbo7p8dtgtX1sl+A6AgLqfIbBXNP2ZqKxhHudte4j8o
6U0913fnrDHqm45MDyON2CwaRCYIeOrsARzYBDzKnu4eR1LXE0wtWaYiQQHYiAPozziG0A943cfX
OiC6T6A11OaZIHEavEw3+NuQS/BN3oV3JGxEtWu0NqyVfXVHDHjCoCKoyD5KuRk5HZSsig6qhsn+
RXUB3Dz7a04UXSUL3HbIkOknv3x1gGGR701luYGfWJFVsV0Vc/9RsjQaJ+zilk/i7wUcxUqmLi86
t69eH5iVjD8Nv2OAF0WlBrd8X3hgUs8YW/bJX6lD9FkBdFuidAjVciRG9TcGTfxSnbfH/JzXzaXJ
aIqiB5ZW1bFXQQWjMnVUDCGkPu1mzYaS/Fa/AcwEAyNKMVIGtoVCMX+7ETBrlReqYnDqUoAwvqMu
VEnRHfk7lDoHkZjhpmttNz7BWeXqL04JJp/VRU138kG60VDkBop1kipvQFqgqNLoPxNQMcczoF0o
50YqDnsrVHqM3iocCkmwZYIKEz1bH/t+c0t2Tiv1Eriat65hJ4FHNudVXbsuE823ISeP4YE4YT+O
GY7nl4q6uTZgHOc09bbbL1oVuMxz6MGDN1WiY9mFE5YHbk5qVCtT8npga67FPwy0biiutN8yRl+G
tNlIT2Lrao2U2Bquow2LmdRhHBuyVBKlVVNB2LWUMG5Hu+ahp4E3roSeh4UuPh7z8zCwQN+xoSM7
dWQDvmVUIwvEdGyw0pYUgmBDuOYBaGWO8N1BcqzRo5l7Pd6LKGgolqcuM7BAnqB3xoZY5Xc145TK
w9GG97bN3Erb3VekpVS1VVwY9C2mA0Ip5XMjMksq7aj/SAKuyUL0JFaa+JR/EYri2ShZwIs2pk8R
fHPFMknBok2swL1NIu6KEHTlQWzkz3c9WbFTfVUky8L322kF/j4NZUJDJhakiwSgx+ha4WDZ6BXT
LmiQs34UxrzgDkdjXSYPODM//jto0HJBANduqwKB6WcDDbFvYc+zO2K9DxNYBSutQM2A2KsHCHrU
NrZofp9w+53p6U0m88la5i/SvOEPzTCp3Vs8e1s8v2p3gM8gDH49qmGcQP7JFwx4/uwu3tHmq/BA
jHV2KXJ3NA6nHdhNcIMLBHvq82XkNLAeoivATVGfvXAXoTJMZr4nLpJxRt+jho0R2W2YPAU7JkNk
6CIFtx1aZqOME3dih0O+LYuBJLcYv54cyzHirMxskpkwJc63xy+5KXmpj4sgvBr4vVbL3V3bdhZr
ujbMHFKgJRnvnqE+wUSCqCtEtE/dafscK7tHzmmTmkJQ9KDuDRXbSj58ANf0PWH4VusC+MZmTZfI
Y0GQpwQZdwzv6IntMX82k1KtORXkT4wU8tVr5FzgcXqw9U9yYIJrc+535xYnCde9fKNEaeA2fn8E
EDkAUcMMTJhXOVA37X3ZGIi9lnDbYgovg5yymbNJDeObm5oYXwK+X9k/cy9XiG0tn37QWUV3/qDO
uh3FY6bpA587Fn8efYYrxaTuTIP6pHuI02GoIGYDPMA8DMKIC29maf/Gg0S3zXTbgR1j5bLZ10Zf
QUvPjsGJ7hKnsJEkzmYjk6lhKVBnE9B35Seyf0RIwPmrU7IicThs/EICtANqCNlj9y54nE0+7+fg
iIuZsuAs+96cYrQvtGVFrO9/m4M4C7rtbhVCniR6Cy6ELrJesEq5fuXcIHA3CzjrU0ptVsNHs5tK
JsC6i1aj6L1NvKqfkcyYelH3QsLZkcrsSruSt7r9oRbCg2629MXC5TfPXtgkj9a3ZMZdly10av31
riRJCFm94Okks8s6suJKL0OkWFQ9y5HmhPahqXOW/syw5A8pj2JjVSkTbsfAg3NZvxQvmOXFXAD2
yez8kMUXgxgxgGEhnjltn+gMFMc7o9Qg9wHbq3v+iMvcjvgMOhuQB0UIz0LIycmIqzBreRTn4ryQ
lw6Ms1nGrFUNlKR9C4CInYIi75JGWsM/Q8RpS3wneY1+H3Z9FUHYGH7X25hoehU61FElE4xy/+BT
ByXr6iWQLKm4Ai8ZIUT6ncgsILUJlFa2C2iBK1txiC+ODt2vwXqA5z5XxbLkDJwcTyCmqBztsLgF
IMG11ZubR5hyP9JypShWITx9vSDWqvgSonX2Cn7rVR7VdUdgNpJBVLLwOknwUnF5QYQTXVUQObe3
r7y7fCrbV+1TKXNWDNKAL4Bq1LlL6sf+24DFb1nXuEeqqbwcwpr2MGHRypDtlajIkxlLUDpkei4N
rk3UH52llngtpUAz4Hh8b5E1uItgKYoMWyvJtI4sBl5KEr31HhP02DrbMIKA+uJVno9H7+hJ4RLT
upgpcZiIxcE8URkaereSE9RJTGLuTTa/VanrVtxHhbuekV8dpn/OTrOm0NnzR5HiV49uzjR63Zck
oyfiRvQY+wipo5iiZM6YVKuB8qf2g5pt2U1sshRlet7znnD6dSB6Eef3gDbK79cbwUBIN8xB99hn
dVydDdeSzKdtvR1L9fp3BycN8us/et3pQVkPU3bn/RDA1A0fD8lBIagTM7Hy2B9Mdlxfq6uwyr/P
XfbsDZQaD380eQoGS/PLLpCEf3E/Ma1CQ/SZYhd3I4Ze6x7udeu3ECFHT43EWHoSR6VtsZ8p5K80
fOquK2P9HzFgAyULN20uvoD6KtmgaP/9iKu8tZ9Qr4SrGdEu9621IBm0L5TIFgCBo/Lb/8pAUGk5
NPxtHvpK3ygqUVH7phON4JcU2LKDydqAVya47YzFjMfg2V0yVBvbm2gQA0eZ+bvnd4vd/uzjwBv/
tOeQ5mIX76mtvEHrtq6rWMycE6RKWO5Mi+HMGpC2U+4JGn5CiMBhXcOmaZ7Dai/V/NKtatfCuf50
sYRnBN//8aLlELBMFIuNJYoJEHpXSaB5eMAkvm78/2dttcfA1GILLLQ87DeGYrK0oNKo3n6/A0na
KcJ5m8yo0a70m+fdCH/rKpf4NQWra0b33RwOquJh9R6ns7d2dqRK9YQFPEAj6G7OI+ub9uCFwmfs
kSbHQ5IWnJ3Gx6OItlgdhHOJGQD/oToOBxnADJz5hrG7CWRjkdOtQgU4zkuR1QQ18knyK4gS5Ads
ILfDlnbhjNYsYYdQ84dCBT7TIFA4rPWY54JFqX5WVBulp6T88750fyCjZZq7ednc/oj/hatptEFW
LMeKmVFDLVfAjK5a/TwNh9T//akFZyzA9H9t+QewbJ6yzRY8S8JUaWJg4Fa9it/+bQ1nTzQ3VEIl
SUyg1hRTmLF2LA5BOkl6xAHpNYnkSm3kpnn9H9ffKENs9ohHoe5HOnPR7IXf3eEqYRN7enWpukuA
76YGn0pScxPB87BNZG7Z1oOAEkC+/nZn3RDAg9iEO8zzmq+tbW0H3KA8ioBrWATmJ15H4CG1gVea
uZ7+XFsCMJM3z+1PpowpdBextX0La4hJhYpd+XY1xzyXSjBRTbqE1xhk1hiRDXdGzi/QdZECOEbW
H+OQrzrZ3WYx3rU6Nq8x/qPiv0DWEz7kXZvfe0RnfPzG/MIJ8wgQu2ZD/egFa+NVNRZ88BiwCjKR
hEWGr31LLeUS61SnqP5kzO/2EdVSbq0Rt9QoGjoOc3/KTMQD2ANfr2YHmSgMVnyUWiYyHNnPneO+
xzhhQHhwgD/vzaP6WaqaohIMKN7Be8chkFYkyYpRMs4d0slV2TRJZVCSotN5+L2dhyullG4xew1Y
oqGf2qoNX41zQ+DvN7UrOB++6BdDvzy1TS++tBhn90Ymd8xZ7SmnW34SrnrS2eLbnzuBCrzMoIO3
Av5bF/ukEj7EDMw0y6I+CARBO2LP0cg8j7Z+tq9nyg2+814HEF3caZSxYqzMLqMAY0BsGsNxnDR3
q/QRxVnMC6JIHPraJJ7yI/fjvCxLppNciJTTkoQQChjWsMXzRo+FbIimL2jtgrWmp5p0hXawOqe1
fA42clNWgLfflryfMYvkcXvljUqLihSJ0jRkdDAu68PCKcRP7xgXCt1V/XzeMc4B+nd9wXro9Bmf
XeQS10ieb032NTLO2L3VolSXw7IDkQM30cOEX7C0Pnlx7gFpQBheLAKpGdkaNCOVt67oj7FQTWwe
jqVqKJaPRnJ3Xh9QXBryDG+zS6L6dr8q/3GJoV9Tv08korAdnxLuyedIsbJlSCs5IA8NwRiTyf8Q
PuzUr4/te5hvM2no/i1VlksN+wdX7q1P1lf2veV0HuF/nLvk1jRoyqWylbXgASHkj8k/aDamdf5t
sAh3Nn8ucyveViQk1TaAiWK+TW9zvO6z367yzSMcvtM8bwYOVUi19it0GAqAxnPIh+D1C6/I1SG/
olsDyVZNGwYeZ/UUCCE+jgAypI4qDpDtfHvW0TEIWRkOk1k5bEuenD3O2Lzi9ztgQVWtY6KNb1Zf
dqXvTZQtO7KoHXdGMR/FFKygkgcfVbnhv6BJdzKl9zqL3Gxr2OAxDPFIcBP5Z5nmhQH2oNbvOtc+
TRYmepFEUu20p2WnoWZcyvEbp/bsBixnNtJZG0wcvlq0RxI2ZCHHWjm8ahPpd29Nv16f9e1jlR7j
n5tVzGzUOU6e8Ue7a+JGlDB6hdp0AnClbJSRBhBONZk8W/yD6a3hngM6pnBCkK3RHAWVqpa8xMVF
Pe4UGcOBWqXeq58nVRTlbgsxlyLj7vIJDC8y8Bcos3S2C+8vtbEcWpH60s65ao8KZShxMNFpCm5X
5y81RhOcBAUZy/T4Q6ZKfq+MOddYcNrHyVvpR7YpqjuL9FEEDsRwTEXAmSmNUpmHB5nH9+1zwFCR
1GKdQpDN3X80sDsXSjwR0qbc5frDQ+zlwtBQlu3McgbJCxtPm5kLz5Ffyo72S9QOZLoAz9EhTIc+
7f0SQHz1IzMPqRAeInsONn1ibeMECdVV435FLyaOtqFpbYlDJ5WpRE65vHAj8QPSXN/gpNv62rYK
+hjv6xlvaiUYCBREVbpybEXI1Hy/VZKrsW16/5wByY9SLS4Dgel/Yqi6gi3mAMKq8Ey3jf73mZXK
7LJPF6HkstX3Ml0XBEcqqcaoF6kb70vTllbp0QLGJF7g2i+wJYDBm2kazBk/t1uwyZPSMv5aRiVG
Q1PSzWHQMgxbQxSRmLY0o5wVLmikNtdP/pkk/xxMgVOZbuDL6STEjOfjma9WVVb16CzKLF+VryV4
kc/yrGr8EfSpiuTggcE6ey39nXtjc4+oqJ+lQUOoPGyEbSkW8FijkL6DR7Qvs8BzAmk9dqhTtGiX
ZRboL+m8OdzHjLp2y/vy7rnnIKe0E8OH7IB95/XHrpbvvV59tFb8O125mQVnoxFUFO0HCu4Ji4Ay
JPOBXhLzIKgcPPHlMIgWzCuuSIvIuOEtbjlUsrWkhV+93XHgfJUD22KRR4O3MM4VqY11yRwvMllY
O6sl7wDoCItwQmdm0c+kaIKxn+cRl6fumRtYG3DJrRf6lpuNpShXAK3wGUhTFjJOdmcM3Q9fJRoh
HcjJJ7lwxrhmdYSjzDBcooRidnfsd4cYpVEE+2b3C6HLB9uBBmVd9hTKR9X3a6zf8/oiZrqt1LYe
Vin0/NgQ3c0uBc1DgltrIgHID5wqoHs5oQnp7zrzAI6+PF6O7e3/VLbihkFAPoQsC06cT+yaJO1k
w3pzYuiQjOd2nyXpcWANOemIILM/vP/0gu7qGbWg4VHHP7/5EPYqh0KE2ucBVUQpDwNRRe0aOdfv
Ke0QPIr4nTSkMNFpYst65Hb4R//WbgTvWv07I2f1P21bljVeOHhSAvLMtNiFx2nJ48jC3Rn4CxND
NaoBFbXYxjLopGizhaRtRk6Kg6TVviJQaUu0iceedwVW0b+yH/21wtvbFWLSR9Ah7EHOKHe16CuW
O8mlbdD+9QCzIbDhZR9BD26WvgMURtzd0uEjKNzdx9mN36C7kZKgDz1BZ3GUsMS613y0nj3Sn0RW
jDIHODelD0fit9LXlIplgZZFwhZEC8A/uLi4hhMGPrA9BdNg/Nc6FanLuf8TZ0iJOjaIE+lD+oSa
12pclB0NUWumJ6im9BFOOw6GjapAh4dwA4UQmdCp4hGO20f6EKBeZbwNXQXAm0dINCzSylLHHYRS
Bs4eCxYQgBqmicwgQ8EabVVBaT/jplNuSJLemk1c2LDyHFRETvO7Boa5BqVn2HvUuaNyoA2PN8iM
bykO1XYXM/93+TyWBYr2CUkYohWQZTNadciVq5yuNL7m6CPtv07yFM1icFTkkmUsLLEKBkQlMFln
MQcg9rhlHTptpHsBAUr+9D3lBCeVC4IECbVgJE7eRd/kBrmBUYuPnvRJvRU5HErjpAFNQfqyKiXT
29Mh3xyK9J9mVvWc51gSXyWBkEdDqjnOJT9cnb7P/ad59+DTyJEmVELAns1uWegPrnEoWuTaL3h4
hP6W+2ikjuE/xKtsHMJdOTterx14qWsi5ocC6QOa9Ie/p3KiKe2xAlMOJAQ7+5byN6VzO7gM6YMw
of3yy6v1wFKxvDJMyh81gCYWLe9snJQFHSA5KdOZibMRWFApoc+xDvtthGX4M0sUmrKazot88M/k
GH66g9XQ/xEM8f/bdLscSy/8uzSFo6BFCwF3vqyDcZq3dlbgTY007ye11HHVaUIK0RRULKrXGphT
s+E0IJX0A0U21/ZEXKkTFWzOL4OVy1+Ff616f2k0oYmrmWkyY/p1BP5HPeJlegRDv06pIaFlmeMo
P9hQEnKNCRBh2vh8YPzuIYgP5Qn+AlioCyV9iUZq/LCFtFBOXsOi89b58rRiqTnB7IHl0KwpeGME
TXQETLHedkmuhs4LpNzKK2TgnkPpCikjW3zCb/MFZIftRHGvr0iI8U229TD/xCLQThT9qtzYv8i3
Dp6Udo/M21XhE6ITxLjHT24FPqNMVVHXfcm7KaPjnOWG7aV00xpdFKmxPnDYxZzeHo8RralOiNdT
trs1wjf11jymphcH8XPxTkN2GoHQj+z5jH2H1Wxi9n1OZRdp6QWXxcGuzyrO8whuLWe6sRdlpWjO
k3fVJDnLgmrxhdwk6dyYK5+Qvw5f2vI59M1xnIya/J8gz5Ojll112B354sM4fZqn/lkerIVohTnc
k4jTRYeQ5cOVuTrCcsidoLeoIWNfvKXIVSXgRn9MqSoew+GNFscoHQNiGJsIl13CO4n9R3bjtb8N
DuL4N2M4ni8tBCVo0wMr31OI74yFs/WSIebdMERJ5FuOitdHetOikrigAa7X7vS8XImYpek0PDIy
Um65jqjJqJRL53cOFxHoRk8RRkYpWX5lb677PtSHL9WayuEO7Q7NeO2ivUKtUjneApYOjR9RrirN
T6/PzgTAKtUj1flPsdRcTuzfFLtqwC126bs1bb6i//vIzmorNcMu1RVYn8oL2ZfYFJV6GmW47UxD
Tg1uvEoRnl8VKRcRQyQAcklv4vq187uj86IdZQzNQVoxXI2WPnoyayhHsCEYLT3wlRM434m587XO
7mESlGKdVac3cAezx0kZUMLvcS8Zx+UFUsHENJFLb0tF9y/kSwzTQ1KGawy897XHR+iQCELyLC+u
g5REfSTB1lQ9AstudBPinWCBt3MF1UO4ZemsEGijfZ6JHpgbMHK+A/EURrnEImK4fnD47GD9hDrv
+zU8BfnQrVZNDrNPA07ao+BsY/Tjf6BoMflSzMEzVagASo+fVcaEP9dPSLnVGlJ5NTaFw6QUK/a2
1DGTFrh2DUSRjOb8cEFHdo77nuWm2o9Zil4YIr/R1SI0IJIRQQoCml2okoX/S33Szm/s/3loANQE
RFhfKtANWK2FeurPSPM8kuclgJD2AJPCXjUkrV23u9hKQRuOvkk62Vh7fMonSn0Pq30EVrGRh+3H
LzQX4zUPD4ztuwfNQjYJhhMt4Uq3gJ4ok4z9OxgGuvb85tipxYawxtJwUg7j8zzfHnS3bC50HOkt
lG6lmh3f+4uQDkWzjCmlTTQS5D/WWJ5q9KyDROPqw0kKUD5W99syRPhtShY1p1oZBWRQ/IbwHuBS
Z1u+yNSW2G/ldDbm+4ClUvtFuG2jM67R04RE+GgyLY6q5xugRtHbFolregF92aGWft2bXegHfQSt
iip/Pnd/umysBM4kFmgiNCyoXiYqVejOmYr9dGw+ac4F2sYqFOk2pvY6FKVXMr6olxsoj2X3Yxq1
6r6sLMPbsu4W3+XhNQifj6Dn48xWS0XREP+R4zTcyFXmn2B4sKq7rfK5UJhalvXZIQahBGntACvK
OcQiTlMbhUP76rsiSFRamaPjbRFj0VzIgYypVEsRo48/skD5T9AokZHEzRRzayxiWU1C6oaXpTQE
gJDWUk0XhSMuJYCTBsSTX1V5taTJr+qUNBp06GBUOdhDrJWRj3z/aZUBtqjCcqmgnb3TpLJWiiCO
v8qvCe5d0KteWDHSthQVvbzR3Wo4rNwEYtV9oC8xnfnNWmMfQJCab8cDRKNxzZNE3vfewoktO6Er
SZ5bgYeuGbcnPhctLIwEzsh0OCTS5o4dYrQ/KykxLiUbdBEKPFKBE6sZolkiLMG5nElIqrgsOfoP
2ZNmRxQuHbDLyln2zy8tT584NAj6QMtKz6ijJz5rqECKORakc2VmVOzgvH7gZqvJ13aGqgNOGeyI
GxV2JS3NyZx1BKvF+6GFktwObF9XvBmPZKOPgSR5jzmG4VmUqitFbMdGUrFmHsrDDz/VYTv/DTjx
cC9hz+OY2sY/p39m/+zu7XMBtA414LEn6WjrIKJI99hCorPekSpTuZj/lVHMsQJR8geTWQ6gLVG8
JMcBzydrdkIlQz3u3m+gTfrsb4ikMoKyrP1trKgk+6h1TAzvv1SEq4apNX99E24eGiHS4PEZ2+G4
agPtOegeELXe1ZajCl/w9bbPTwkOCdyKBvs+7pqf8gfVgVVZRaKMKu02t/g2ExQ1duScWM6jXsOF
hSP11HlRanJa/F8XSRWWGVoBmq0+wxD1+43xPNFOOxxzaATM1lXOgXWgc15fW3pCgXw+mSXcB5tm
ii3qb4Q76WsJpqp7kql+Ks3qALFFSgpRs18iLjso+frD5CpF+MW/7IXnxfB1J/nXwsoHA1Y3Mzpx
gCRf2B8osCN/3k7lBoXBP4KRDEDh4Jn12sSPf6IfAF1abA8bP4bDB3QT4SiXnhJjn5TUAj9aWcDn
KoVXmOElaAeazCyY4Z14JmaQS0oHPqB9OxL5qsbhpS+vK6w5ZkOZxCRCZJ00swxVLkGrmb3P8DQM
iUJjDwlUyH+MWSGS/RW+AUWjjxqJjBxuk1QIyaf9xNOF89BIdySL38bJOvXUccaV2qQrtAKSDo8j
JqtzW+/YYVf0x57DkdeY0AX9cKAHXO1nm7PjSaaBWtUq9G0zUJlTGP/C/uHLTJpF0xhjdm71F3nq
JaCdsDE7bli6rHJLYy5FTnVzJKz4kll1cJOUpsxw/phd1aQKDFx4YoAxi7Lehb+H7gkg30qOAo2u
COyZdRh2D8n3zkriZFP2XS8NJFroh1KCwCLhkEFHbFSR2+9nhE3RHzn/kPBJ81pIillZM6mmvPFl
5IzAeoYzvWRBlYZXx8jDBET1pCx6Y6S3nCJIAa+H+/wSM0hHDHA2MiG394bInLd0hDMFrpC6p003
XTqqLn0pvXXNKDzvTfvOpqHK8Elx9yXd4MY2JrARSzDUloCh2b5Y7Ydns8UWdov+jOV4jEhwDtoa
WDoNP86ahA18S8Li3rmELpfGCKuz7ZDT4pquQUHfqy8kg0aHDr+S44HZaP7gJzaGYdCraVL+2DAb
GO/37HUUcekZCpfP5Z3hI/a171hUkjuBUt6CeR36EEBttXhvBRuucAx09TWEfjlqmZw3BvKhGyAL
axA/i/vO6F2JD0XWlBBFxH2PojeDOtXX+vYo91d7JPBEHnSKnBsaLjdYAM4oF418c99SUSCT1MKY
7reFPAa+W8aqgOGAx5Ml4e2xE/OOSOaSDpA6forOgc+BL2pzPV92M3JWPIp5c7XRzUloxrXYivJa
Vm2Td5OS7ik7UsaZEMo61Cc69e8HL+/MnhLDmfzgQW49/Fa0i+tN6FNWywwb/dwK6nO80obHPhdS
dUK1MFLY0U0Dh8/+OXU4HZpMszJYRBKs5XqklBYMpdi4OnKxkiZDEjL2qzAF0tRl6H/mj2rgC/4r
Xe0wJVlaHxHfrMYv1lJSmch2/6ChIjtk3r7VTKIHLuhJGJ8eENbkBoVIRCoxOAMfq92P01qvqeCj
8x18C7XdzzeRSsMbEJn35U5ZglgwukHO4QvYVD1FB7Tq0iSGrFmIUsBglutyZq7ICD5x7bDTKZtE
KQeWbrYhoR3XtwzvpsJ31Dss+7ZczjE0y7InuAmt7IHKVZ+dTL1Qk73yodlODQUj1NKev0Bw6ugk
BN/X5r1CHi0xtjCTEIpCBvkVmFWj1pwGGC9I6Y2uV4WswZ8tSyCKVZaE9dxfVyZtkRfFdrGxLYk0
hMX2kcSp9Y0Gmqb96ZvywV3BhEyZnnbRFVK9W6E7ZXPoMhG4dGriQSKtiMtMvnXNaQL2J7M8Anwm
UAdr/kCtAO5cEx6eAXrT1zXzPgzQ5cXWi9O4z7Wma8ZvCfai/EJ+g3V75kavbzuH8m0JJEOuL0vj
2XEd1HIuD06ji4Wd9Rx4H6YI+XEPJNJzgEOe+o7aLqJZDX9C9LQIyIavT379CZ85GubtPoUdQz1Q
91tYHtLDc+PTmHpThb6IvY/OdaUkZu/uaysPgWVkS+vUPqLBi6tpvXC4seqfU9wW2iHHAa3/17jL
nD/3W+e1GCq8amgG1pG15iMRXlyTiXkUW1zUYh27NeFPWeoSVBhMRItHIYI5L8mtjWMUh4+2+T5G
isb5BSi3Y1bggl1sloVgqdZiO8r+AZ6SPDgWsSNcD8YT8oZSqbJw0HVCkhEirm/eKlRNo397wqGN
M4eF1p8elfGaITCvj/h0p2Yw7B2RhlOKZ16RXUnTGMws93dQoBRkWLF/u7PlQsPQBKXou58xEiR2
P2AYmtMcAF5tXi51wWSKzX2fxacSTe9vFHLVw7B5HkYdqBMbEsf9TzvYdVe/MHvbJkEGPWIEQmHi
kS3b98ooI7UUbcR7gPvo9ql5999ADuub63G5/iDq9dNqwzsErZKun0b5Nrriqa3mq1gYM8nA5NYt
g/xeZWhyOEUyZH5N4nrM7o/Te5yoA9vvrm6cNH1xDfvg/slKPzIggzpC5kL5RrfSVrDfmc5krNhP
ZnzGx80HbUIveGGOhMmjwWSmWMkscW+e7thgCq76EUPW6RfqGn+vppyFA54IYy70/4KEzA5OLAF5
zscrrVyuju4cYTWis86ZV/VC1oF+2s579b57fHD8WaTiToIF52CpQLIwMTJJ1kVEjYvsXA1kAYJl
ArxlXRcj0zzw6R2fq9vPi6XIErmQs9LDDERIa1/4ihhVZpjgvugIlk+CWTjo0gogfAtYJgcMGRU1
MfrKNDkRXc7ziYBayrOcqpNM6Mu2AYpUeSupCxyalZNiMT9Hq/dmwDjesNgLvrLNxyEVV0HLYdvo
FPARwEJA/ZE7HmZO9Brfd8h4r4vtrTPMGI1/gGbrW+Uk2+jhrWZa4DqiXrvb4Wy6ily6K8eq2bH6
Dt+VPsYxktJLhuGEf3Unbgm5i0YrUxhOB9vlV6dXA3eVK7DrLs1XRgZf8j00DGUC8/msklp7aI4R
CWbSEDDd9VpxTzsPjFTEC/VKUExnMKiMVzTfZibUhezk5uvff+wTPXLEXNdv6hGa3kvJaGqswvY5
e2FaeG9ixVIXI4kEGr1gyS7yERzW65W+pFGpZfLOCKV/j1mgTINxxlToHt20gbuelQ+tS1wiXTnJ
3lgtbDXI/2ZYnjxAKOtoGnF+hJ3knyJe6EX+bVvIQhShs/1SZi2AOdh83oUO8C6KfLGgHsmT7cnY
eL8+yogIZOdzw1vWTE9LMBUKYYbbvFQHWHnr0hptfg2aseVbF13iTbDd6L9sGmro5RLtXMa+obkX
bSVMpIThlQqzaxedU9LTdy8Nna5tgrYCvPwKc5wYnznL5mnB2crDJhW4rAwREUYnhtH5wpz1tJah
0Swb7fjIrgQNmLmQWNMlQltwBjisfi8TRfI+Nr8XOAxo+vpEj8oyUTESBH8XMaC52Q8IH4fzZPSK
YvIns5+yAnRsPovfLDpnrgTnd0t7+uV2Cbr59nuFymE2yZ3DrpHaTc+cG8dZ7TEXiSawgSLoYaqS
1JJNKp9K3EfH5hRr3eoVXqTvdh2qPDqdd6pyPyIbZ1uGzAiDWw7cwEpDlBgIa0/oix8XWwUE17y1
i9ZgoEswjyEArB8aGJbhlCj56hZSTQonTCdyQyPuXJpNDtjZLV3mBw/lWeIJBs1fHr7b8khR09G3
0nEobkVi9C+1HhgaH+sQ/kK3vPsqVo2xXVk5K/TygaDOC/eVZC2kGpTjBsGsBX3MPH4GqlV0w3wo
7Go07ooAdj1ZgWaptENDJRF/SBbE7gk5PnAlhWZh1GOFX7GX9tuwhC462d+uK+k/LupaC+BYcwFg
5GM7zU70WEF/TgPDxvuoUFnpXkSMDiDFXI5mG0cmahIC9RpsU6mlY+JIrXBmeN2HJaMaNu6NOuPw
LkXbHUDb0pyWJK+vWLfXR2K+Nit5zGsjgGcQobfuu2e5HahvbXya9hZr4s8Xpl0uU49fZOmG6Z2v
QcpCx82nKDXmE60xqUzNNonHlLPMpKounUIRDhZN9wXRPowoL7lEp/ligbbmcS2zfMtBxSuHNbFO
G+m7WpDgmBJh253vfPMy926CAOGL3qbBt+HzmAx6VcccPWEvp0NGHRa3xUOaWGdF9/tRrMiB+9sh
YHO2tqcnByhkoHfD+EEflLWnZgvyU/ihKlCx/OnYZtmgoiqgHZmHKrtmzhhxpg0KZwnDrS2gndi5
CM3+wQlOHYs2HZh9DFTqYoqGfG2GT8UmUK1SAJYAL1izIGfSfab4mAJP5v2AENDT3WDaUwN7IZAX
eP2twvRg5e930F+XF4dKKr13PI+tPYNkJ9MIqt2DGm63jIRa+pLpmyImUGZV8Dkk8l/RMtJibyBe
YOzGXzGX2+E2U33Oyp77smKth72LuAS1edNlS/zlkNYlWxI/CwaSQfGncGyRHlMwfasF76Hghx3h
iAxn/pHky9mwmds/JLQh6XtEhZWnhfI0jXrzvqeVCyipj77dCFGQNFjn1kcdLCu/VPWAdRb4ZqP8
PSTMykWiMlPhsKAjhNvm03E/LkCHoWz5y7+WxadBnuwlNG51VMzBdPAEW3jvdicWZZ93vLtxlnDq
sgHcw6wKh07yTbto4UcZwkft8K4PYNWm3bgp+WSWrwkAs/h4JgykXK7D4IYG02keN0fcj4YjVahZ
Ycdj4jI98Q0vf3tlYi7lhKf//C50ctrXqVi3Sbp3OK/FX4zuEQfN6uYr8KSjCzwFXrzdXHMXcQjd
BJ71/j++gDxujqgm31kKBZpkqmKu9PDVCA/ubt8hFKHlDvMbHL4oSooKq6t7clxJXJhWWQZZJcA5
ANFGUfrtbWyGsU0/GeguW1XHxcHONMOhdujgbRZxX73kuzZaG+4ZZAU+oyENEv6c5gn9RQaveKLw
yaTGKx3GvQ6ci8RB6PvvKyJxftVKFWfYBn4SU0salnwX1DXfD5CcEoOqd5T0SKMm0fVQdM3nxEf+
uTSw+N+4QL2HxIlhR9aeN9HXEVIY5ts4KKFLuVnX4a+trW3FwG2UnP+v/Xrl6SfB+wAtC28ds+pS
SVNyOOLInUsNz7YlgRjL44sczxRBLQ2KpCBFRRibJaz+FwdV40Xtbjl9D7+7+rSMUEAruff/sbBQ
FAfGObEf8X80LaAO26zEtyql9a9C+alluMK2/CnKG5Dm2vtOvTR3rXh/rB66OuapoF468orSlJKq
EE9ZKtBU1AauzaohsiCc/Ua08cSpShOzfGS09FTDC/55zjTHyLvtWxKI5qKuXwc0T4hs97hA5r9b
1trnRS9nxWoFDl4qUE+V3ZaQ9AkBj4ScjgjiueoacGcsAqN9Arwtqhb4qAyOVck5P3ElfjnuVZBu
k0pK3nkeFIAysmn2zNcbW5nVsh530BdztGQRMUbuKrpknq+W7/gnTk4F0RSWSTHDTtqhZ/0jQ8Yx
rSYByUaIrcOi0/WliiPDGHHxjxkHlgHdEmA4HAWEWNEIknYjJSs/gslpC+6IeWg9HUIO8V8sk7cl
iFIfOwm6ZE5rqj+l15UBePGBAjOmAzvMeTjgprr4PrnwvImKn4yD4LnhrQ73iGOX/kZDv3DZ00m9
0VNcN86UAOg2xRmgQUZ/+lq65xn/tn8s7XC5Xk6rIqV1cJh6ihn9pimKh4EDN0NgIUxeavsTsJDT
Jk3UD3QVAINvELfBM03bb5+vSfN64rNC2xAP3yseadTznxdD0iuVFATOUC7Xc+YMJMMWWFalwdo8
kfOkmd4QChDxPSjcxcE4X9lPHt0Ad+KEbzUF2UX7m1jUov/PAr0n+BnonZ+5/TfKOz5mHn/hVKG3
171Rowo/qYmvaXtwfr+BFsW76jcMxfPLl1/Gukbo/QPWdtsZa9+SXTP8tVyzgWRAgMV553JQbvtL
KpGFLRJWTSPzknd6xfWDQH0PIjIFf9yclNc5hNUMoLAATywjGcJKq9xA++IoIGRlyExo6LmZ7O57
lyVGbo7Ua5pzBlsFdQJRx5Zxp0LhoP1TcJP7uum+BD6h/kPaV3QMbW8zKEm7OB4Tx8CLCFRG1OF6
lzjphgTVW6AkmQ6XDn1g/RGcF4coQq91M+pRvXa0oO9SO3w5QVVEXCC0IP47T1MaE7Tv/sFDp5zO
KnWIq2d2xhLasWhpn8YLXgH+1uGp0+kVwC3mAVDxmi4xlDxQAdFamzrTaEABpBZDPiZKya/KRbxC
Ypj/9cZlHdY/4gqcS0Icu2g/DGyd+7EwY9WPyadkBCRRCwxikPP8+zfBBVHRpcAkmhmNHNc07ZxO
Re7fUNV4L7AHB6jfpecbsXmM5yiBeYF8sFcnMolzfPgn4HM1n2n+Xa44oDMd0DPKEP6GSSXbcPKT
41PMCfAni+L+N2BFGYa1pgbU7bH0o7RpRPqb6BnAI9xesB+eNOorjQG6rnEB2Q0NRa/vOqD/Y+SO
YwvsKWSpMM3YWDTxoKGkfcQduwAkuhZrsbD11IHwQBmBN8YG07qH5FojrixsgOjwoWIHC3zXQ7Em
sF5v9r9n7Zctwgxd2rA483eLZ3m0Pt3+iD1JvzYVY/yCBY0dRfGFk+LxUZP+a2bSxG3GnaBaw6PX
YZIqeMGD1Ebujojhi1SEvYtlAhLQM2KDX25CwxDbwpoZyX+jUUrZo3eychFXgIKlppGUjd09m44/
R+Q+noSDvCNMs1oD3v/NY9bT+m9HhwIXKFiojbdupqL+OjrcmMvwWn3hG7ERfjX5cclYQUpmbPg/
lV2zNpxDMKvTU8kliwB2/XrfhazwtX/euykjKaIzWFoV29uE7e6lNB0Yopj28ScRAxHsXjDE4O83
HGl+QWITQJ6WnaZ1/OhI5gpNnEHMgnDg8BgU7zVk0f1hFRsy85q6KgnLYh5VZ7CBOImtUYQB4Ii2
5+wBG/bRf0Pk/S8HnAAOWfoIdBJl3qEfEaZGuvQbUarfEWsCuFZLYYdkCtgGU6aOmb4E5fjn44Gh
kLyeQLadb+e4y79TAm0edad76MvgZM443mHtzEa7dvykgfGWS/WLoFX6Haq44HtEOP/aUyszkSKa
PSfi00O+65iTI2IF8E+QN3V5Kmp6viYxBuy3TRVNn93lzh+cn/4w0KYw+4XVwr2XIN+5U2hFYF/G
uxB2q8gOSfYUC52iRhHsgArefOOEFiZ+OfALqSfkZr0zreMzPk8Si0ZqpRbxQVxrl5aoDK+Pa/Jg
SvlLJXLt1JgKEDvsirWEkLI+Ky2mj/fWJN8YS6Cqh0cd+xQELFNUm7Eks6qHaJfKlhZLHdV/7wP4
rh/hBZfciBc1o1lkjjou/oYaDKYEAj0ACRcoDwo8m28/M5Tv199Z6ibJNhdwGxXgxR5nlDrgknMr
RM2yqNy1Tovkn7LQSiuzStm9UJnlEcqROyNeUueTCK2y5vYK9rkP5/tEsVMPZfc2PJYqe3tPso5Y
ZRPGM9kCZGzGnd6IlTcyLGpxqa4qHZ6pbzCz+FCHbgguw9zy4FUUdBA6u6bw9SGejjKiW668A8Ha
ebMmUMbPK1MGPOKKOE+BU2xH2iGJQNBYPtt8En2UBS7HPt+GTF/lOdYLFnTOrKcp5EJfqGWKnSJm
lJ2U/ClbvJ63Oda5I1wVF8m/mLHq8wL5YaXyo5UfzWs3ryqus0osRY2loyX3VTVc+ufnreO3de+G
iinMUKQJ8hrSkxwXjktCzgbc4zBseZD/R7kasrNxWkYep9alkoySsBqtOCyWpAllmIOjK5xYIwKy
IBncWxEJte65aQ6gaY30Qjpcw0DZJ1+iJXR4CXL8AT3msorl5dvi+1ZKpkrEASwM3hnIld+NC4u9
1F/XQuQFjHJnJv3z1ZkW6R9DD4HyvlhY6nZSoL046ub0rQS/+MrJ6q/Mi2LweF0kPA7JtSjRR5fa
0JbGWpSFPHZoXUw5UaatWuqs4dZd/O0bei00cjgmv/1qxU4nDoskP2dx/D3tEhn14wpcqeoIF6vr
IU8x8DmyLn35MXssjS84a5iubVhYsG0/intGFQOqBWbOCU1PD7wqrm1uH94Q57DddmLpL4/oj9Yn
bGuqQcebWkChRT0zqAdl7XGYIdvgdwzLCVzyW1hkdGINy+ByzNmjAc3WqPX2qIJdiCCZhEXyN10y
ySiL4JgPV8REVhMa/tp9fjXxp7tQ7eg3e9ohKimbioLq0ffz/K4Ni1tmZtUuYpiq+Cq37kveu29G
JSDBHE5G4xyndzhGDblLhqxyEgrf7KLV0iHPkYmR+XfYylXCXMWjiVk0HVUVVdpI+l/aLTcjOTIF
rVNBSrbjiFdl6TplNnXPDvkieLvqxxyIf2QtpJ2AdYtjTOr+dOWPuuTywSvIYbJXu5x3eH4Ft1rm
1z1t5I/KOaLJDvQ205ISBqAEJE6iorJPNCZhFM4oupprPKax7Zv3phhYHwjyCcQqBGEMT5PS0+de
M7RGVwjPgm3fUzUH+Ai4iB05jPxvFOeaWtE31T3g/ddn9irR4xsx7lCLwg8CB15QHnWYSqiWHH4i
UP6Tapoc19LoEWBCNHGGlIaOUQkAHy4Jn4QYyNXiz4bW0a6OEU37eNba/+GvhEqvCWtp7lCBVr+k
qLldfEiERsXEBWHSSemTFzkFO5QonNVm9RgRoBdQm4qOpyvVCd7L3ZHIna5lwmmOXUkEDaOqvwqJ
rTZFDlUG+/lyd1gRBrLVCaOC7G/IpF1zDeETuQoB2v0MtOk1SVUpC5UJsWE1QwwJOwJzs0JDTetq
cl/iH/oa9KZgCjFNM9KLEc7Uunj9ZSkx6fDWsScu+AH043vfNaYFqs3HV3DonqDJRC0K0whU3jK+
zqoLuOawn6PV770K0D/vkcfRqaB2YxkXFRnbIG8MeUOVfyupi/1gMJQYFnT9+4HZY7iNfRmrsZDQ
tla9qS04IUXwvxFRgIwi64sdb+vq9CEcwRnKUpTr1Mjmp2M91VL2pqus2iEV9TNjWHHLc4psdX93
25QFp7hN+LxjHGVfPfSwJ3uf9IdNZ9FiqcSjADAT5Bv0xrQwCW9+2HZFg918wXMkXRY3iy7hX3S/
15UvyETv50LenImjG43ZXY0gWwunsaZ4eOtSoAOSU7poUnkt6h406gzHKZxeNNaZ0Bxf8taxNLFH
69qOmo1myYKF4hzAVxGNbxKjQm1hivqU60o64dzv1o/aIYksV20EPWT2k7avn5AG1Ip9J9m926Mw
0nYn3EeMDrf5/pTgwTc9PEqI8CbfhFtaiu1fMj6mTDEBg75/h+YsndL2VdpGSwtKgrh9Hr+sd2LM
rRfeBaqwttrWdFy2arOs+0jm/f0WJsK9c8NST7mamG6fFexaSHOyAGz2MCZIAiANwOEZv3ekJBrE
0Gzb1wAz2z9sOeDIieIp2roLvkIp4ihV/q3C9XLAACL+mDud0TzUl756fgAgVzHGt0UoUoUoSioP
nMpVqBfMeoxoXfdZ70LCZ50GLGehTUQOWoIBn7OI8x8D0G5d3+4uIj7SCI24lxOkPEQ0T6h7kU3d
2HsUsPmYUtCUlX8sfXO9c46bUp4kwN6IckJaLKXy3V3DFQ4DlvWryA4wkS+5tW+iY2Z/leHx6SaL
9T0PncoMdoyvMOd9Ni9Do11+TlPdhyPhSsOMyrVShXInMVXQjDjtgQyLflkP/36+Fd5/UEZtxMHO
m1wRYkOMOG3Bj6df+CPsunXl1dU1FE5Ut+7Kb7Noi55IhSHbVZK+UKqLhr8AuabEGGHFnMNdkH4g
aEzOHxhO7tHRpfbGkPWFcW7BLe6kv0HYOxIRG46yXFk+DXvHUP8iGv7F/Bwk9GWXYHnXhji7WRzt
u2lMPi80RXlpW/0C63E+9vCLo885BVBNmypQQKnuY+kh7VrcohEzfXr+GUJTkVxS3K/AJbsdd9TY
BWC5Gdg52GjAQ6sYHyWiBX5O7s3rWuAq0cxiTAtow6r9voFkgsCyGp/k8Up1/78zxJj2iaYktSHG
q5k7d73UvBTSBx6kvv2Sl70EC4KNOK/+IaqvQtsei+HIynuyqyrPaKeubSX0SCnac1EjCtAes5j3
4wVPvWSTy5BVoULWF7+PdGtBG2NqJf6cUeNNZYwgfExlIIkV84GvsRdZhjMmjX3OGW3P0UXe+Ioi
yaWmiHlJ4MSlZ/KkrmgXTQ0VHkvzLe4OlshAEXdkBremsldVCVZPTJl9vObI9jmH+KnfC4xgo2Zn
mDQso4+Mjz5DL3yF5osRmQQYVBKwqm5eQvwN4IxyJGg9KYnOzNpiAIjwAeQyV9S2dAv0PeAxFGtW
dUCas92lsiVX33XcoVd4XFh4phmyPLgI/NOHT7FRhzlt8UOVkH1czqRVZyRUeHFfJFUxDCE26qdd
s/PLy1R/uKGGTnbor5jtfzceqtFPSTeARc+cZA1Syj1l2P55nsGEDzKuKiAg/tZZ9SunTB5u+jgT
40TLX3FQoxVUJ3mQ54XxFJSnk3rJX4Su4uI059vRAHkfUONFG2E9pYguH7vfIWoR3tVkWYzvhVhM
q7iqD/Ej1uDHr8P+t52aCxSL8khoil/RBoiLOjXTLXtBHafESnfsrcm5+ByAeSEg3DPBJ4knvW19
0dAGU5J+X9cdUdozAQtfxQcZ8w3mh/Mk3sfT3l5BLhc+WpkCac2D0K22u7MU4xSu+qvuK3r4EZp0
hsVNkgjshkgQl30VKt++FgrZlJthRNP0vDzGxAdA2uZuNd8OGZTRSgs/mEzhYlTxykTW/60j0nWy
D3LhWToVVJxJErM+ScjfwhxzczU7+me3wL1z73ObGWxXv6Nbz2BDdpXwJ7LDj0rqxZm1lmYlvxIE
e7nMHxpFZhKBP8Csr7BMUbHpzYpRLT2O8hwK1h6IKarqOxLPhtNBW96r/vfSfoUcDk/xj0jY2XKC
q9fgLo9VmbOgxOat4Gwk4AUa8qWJdIpinWl/XHwzfpxS4OXC2f8RtG/gqALX9DZAejCV6EITs2Mc
ypnF/yQjSB13N+MKPVwiaT9TKOhQ9GeKx871li+EUt3B1BIqf87wy1S9xmJLf5tIY9E3gnsOxqwL
nxk3SR4Z4jiKCtcl0E9sHxzDFBvVBzJKt2xMwOQgA5DYItUiQ7Mh6KsS6aV133uHJDGrXajVmjZk
i5y/I04K7IaJlvJnn/klSf6xlsJw5sqESrmAOdDevh3pYzAdBux/UrXZbwrjdDPcNC5sThcOL6Nv
400YNHS2IkuD0GuKoSiKZ7sXY5ySnUZIFY0K7dvyAvGqCHQOjyjS2uDlImT3SUoiFDX/4pHFE+nN
UP5YcegWhjYZJkOHARkrGOz8vFzA8rWnXO98i774v5JCjdu/b8eU0t2QVJ1dJqClJdWW/CdXfL+k
oOYoL5W14Is1JbSm6fogCzTrhdkF/QU2T78gveBHf37/pW8rt7uncCjj5nI2nUr5RlgAjdRajq+4
oPfnhVj+6tven63Z1kZO3aoQEHUiDJw8exiZjW9x+xXTRKcNOMF2x1yZTr/vvbZAOsf6gBoCgIud
izI0akOPdjomORuj3yQNE0TQmvk6+jycT2/jDiZEHpQtjxNK1XHWs7hca7WAFohdvj/bb3Sp+Pko
YhZmm/RFdYJvYTfL9tZv7bg8fCy+a4wfd4d5kRGUYf19+Z37+cpx5EBt9GLGhXu+q3dVXCzRRF5+
Slh/+6bVnI7nAuJ/yx8sLdnfqnxe942EZgSPM4z83bYSKgY2AknuD3U9NxLzHC+4uBZBY6E1HY/7
Lhj/xgF1xf3QHWLWZbc8Eg4QcjdE49h2KVz7ul1hhA9qWy305VHpuzl7s6AmMR0UI6oddgQUOsog
zlz0P4/j/Rzcz7jbwx0pTtoHND0fHy6FOLbIkBRk3HPmIrXd+YvT4kJQTwF2oVhUiRCWb5EapLCa
5THHt8rc96eysxHQHV9pGEfq6MNTMryCMQqw4xfIXwtatV5BpNrAT7bsmhNIHW/v0Xov/lnrBRAX
dEpudczmhx+YPPqV2KKYmDOc08TBX+nZtmU2PbqoPxhAhFw6sRGw/T/GcKCsaAoEbC22m5WG4HLk
On9RCbM/5DJFeVotp27AgzyF4RvxhpdKQ9Lt2mJMMg6/MKvo2jzw5G+J3/nJAsF9P+Mxyb/rM3KE
6UquX6bVRoSVGxj3PTafoNj51z5vlRZWNQy49RMz2MazqRlTULOdm/VkgUSCfHNFzdHD22P2wWQT
/askEl/fCFMhNGt5fZI47IXPlSQdkiE7HMbc6lRu/57YXQsAxSbgYsgW65gArDw6AU1z+5bk3Y3z
ZCxrTKjfnXOSPcpkL4vEccpxhj0UgfG6gdEk0ViQu6hnK8xFuB2mqekweKECYRDxTkB01C+i7OVm
Y05QI74kyfvVxruJNxBx5MkpXGwmeyOV/wdqRTRDKbYO/zcZVFffl0iYMjaHQHXq7VdJN89tQgKq
7IMxh1AdDUigoCAJg/7B00ZQnFX3bESHSJKbXcIgzCJYeBzN94vEKUsyriyF/kYxRjZWetQgTPes
072ITHNn6fgPA3/z0atsNGGs3tQ3WfTzK6BQFnSmpQ2x28WRx+yztHj3H7cBvBatDHqsrA3/Thkk
rKM+SpPn1O2Ug1lyC/Ft3jkFuEhW6KnWcb1xDqtrjOetZE09JNdgf9kDoBfmrHCNTOob8UqC4z/Z
pZHdEz3IqV/gKeqeI0DOWFzN5IOuDGv5ThHpVL/Ec9y6DBA+Z8+nVqfBlA+k9Te7WwRsrfHl0Bs4
gWPAmDiYfteY9sMK8T7/BI0tb4XUmgOwcOCtc1BAOdVte1h/gSMXVtkY+pA3oIvQOvTkjnkD7AME
mygjK2I/Qe7I5QqImxuYDkAXWGINrrk/+QLKsgg9MCJp4sOOR1JcmFXLEEXPadzWgdltM6hXUgbb
lDXyadZjhfoNWmifeAbI71JPF5AROhqw0ybQlL/+TEt++cjNeIqtL9e9gDODocWoAHp7Qt+4CdEy
S5oGWNiDS3kqbsVvpkYfAsRM7FHfBT/27R0GBS8Y5o4mmuMYA1Om9MkkqArv+GxBo2W4wOhrzjwX
MpJrGfKIhBgDwVtfV9uXPiNthbU3mQ4umrAzqnadDPhQlmpYCgogYn91g2bQcWlbGu6Ixni/+l9Y
SXztWzC6n0ARzLJtvoi/2OvSjgzPygp5uTp+VQgjLtthn8z64zPpyRVpbZPMFycw1o/UwmDn76Az
2V4hmwFxEUojh7OkUPrlKNbTkjEAGRbxG130u9+pxwmAhQKxd0Y2VZM/LzWJkVtaqhBTSAE6Mluu
K/3FT/oyRcexOVFiuE4rMjdlrAXcdoMKv4Kw4nfHguBwFjTHfnF7TF0DxabvV8QMnlQ2wUJQVQm8
LE7h5x9vahG1nWCZFlSKQNRdL0C8Oev5tNqyUy6BJSyDWDOche1NanoPdtsgHKPt/acGkuXEdOxS
1qlLkmwhVXga3zM9kfz0XoIhHcCYd3ci3I3Jj0OV5E878SPSZb7myfHCJMPdJwyHTuhPJh3ct0XR
TduA/+IbFI8PtlsPj5trEW2PbaJAJlMWvkhmEmmYT92gcdQYX0/ebVCwECE7AKIUnJaonSmYhpyl
OBfUF9cS/MPdVdEPOsdehDVEGg8aPvNz/cq9X17wmHceQdYe9uCNM7NiyN7ut/qwtNq89RCZSQfk
r8wiGDw0FvZlZc34DFLyJmrE5pK/sryplpfUitfjZH01FceeiSJGV8y6/XH/6fFC7Mo46YubIGSz
+tLZ7E2RQrKbWENrJPnP64CenCOIQHz68EngqBjHTREPCrclVwB2azJ6HlPQxYywHm5WKuF6OI25
iFiqAxxBqfY/q9tpAAnw8ohL28YSqnd+zFl+3k3bMG+edGyURqM0mFA4DNodjUJ7hvZsYi9JbHEu
bI8kAnqcOIQ/KY6XFLdDNq8kEXq2eK5X7Q7aymbuCJgNE40xTI9VZZS2Zyxt038HdZ62vv17E7vu
05L7UHdpjl09+HhDNR1uiYmgI+IuVuYMUuzyTa79RyVp9007CU7gTHOhkJ4tWlA/weVPbzirN0fq
VzjOLdOXdayhFYF39fRm28QG+PtSPBwLTyqXiRp8mt1+oV5/2GiGf6IhEOHm3nIUB1Jar2AD0BmH
6+JiVuUuJkyTVpH4VoGhIfaMNkHy9CjsHdxRjSmPsoutrTUUTbB6pTsDh9AvFg1/bclVTWNi7erj
MmYcKIYpWMPfuOFKdYxp2TgONDJMrCTgFMznFMizfGkZCLCGdn1RItkloHomteJOyoLaIs5TK64L
fl6p25nKRdG/UxMgjpD90waA5dLIACoZtQMW3XMTGvaXFwC0xOnieBW6faSDyv3iK/1ghhVhZKjk
1YxD15nQXP3R1CVYRofJKrRn+YWdKsW+YXiW6rscK5HCGJb95AweHKNGUH/e83Ak1ayXZl6UEE7J
EA9JKCcH7MtoPKusIm18O8kkH+syDyBzGI7ufw+5VAMyTEG0vCk8NyfhyVnCKDMfCZB8McnuKDYX
yTmTlkf/Uf88NQFy5+IGJG2nD07SzSuYXdeCyQAybpJ6ESxAaLTCuNj+OK2hNwdxgU6nGqMraStI
9ltV4zaLr7K5xl1gZjV5F8f0ED10QhgkXTriCFMfd02tFETJKxCVZifGAghXdlgk7Z80r24TQBrZ
ETF3emT/wsgkZyqiMC6iffixe1hfB/RvSDUWIN21q4iK0AIfVgpZJKxg/adM+PtjhEAWly/L0CUF
VLt+2C1eYJXcQqAYRObg9HzkTcqx7dZo8tx/Bc5eCW2jrQ/bQA4XF2I+vakVkNvkGjPxk2kVfLXI
i062yM6LYpseSemS2mZKCEpgiauq/pV+daKl/K0v0y0BQ1jwuOnTU8oLY+TGAefpMs9HfRT3lxKK
Kv4/X+Fzbd5IVButA5t8QSY0N9fXVvn2ar/caTHVuHoS+W574IdttCxddX5jP3x7u2ZOA2F5bRHU
oopkBNYguFTEfhj7jcdf7+wTi6mqZXpE4MFZ4TWgsG2jHzXSXkyZrKD/FarZQd5LRrlc7Mwjpkgj
fLrRZxxBON9pUmKk8IQtQS9JXIZk0d63vVHmMOOkk3XvlDZPHiPRDb/AG+mZeREiW1lDiUKSJPQq
WXFcaqfTzJc17Ro/eLCpT9FSzfyzxnb/MC8R9ZKLp5w5OXx4+0idoU08FzE5veCG3F8K+eM8OmLg
N5rGR2Q21pSZmkfaI7YSbwPrptY/FSrQ94p6DvyWAv/vlXAYyHYYKs4JDfI71cuBFO3YPlt2CJFa
DmUzHhu4hi6ROnjE+vQMNfkZR0WCfu3l56tHcanGjJrn7e+8iCHohcli8ykvrk0aoF4Os8NBdF3C
aI3dpXiNtk2nEN2Ys4BgaNzVaF5OGlTELanjt3iyA/SH0f285FsK0aMb1TNe8ZPgCxPyXCaHSRdG
hYmd+2G+37f7R5Dg8tZW6ApLRUCNGETJrAeMQduJsLMjFqd36rtRdSHCC1BND44NKa4BrxyFqS/0
RG6AHNSmeNgeDNunjzTBXgy8inMqi1OvTTXDv40to84a9jB2fBmIv7mlrE0d5XxS46hHt+GRTCLS
zlZvujXjushNnwV5Y/0qtK2BRGRJ9fuViXWnnQE+5SojLM1/oIA/WX1RijpFRZSYZ8L7PWTJiB63
n1x+gfG+7WdkzrMq4A8UDiwtJllUaIYHHrDnH8FkADiNb92bYtd/wIF6PPam9bIZus7VBpnRJ8jx
ZYZ5rgxyqmwotCQ5ClVKmo3PATzXmwsb/q4cq/emC9IRMv/GDFDud9G4bSYQQ9a++v0B/KtSSCV1
yEqcdbQ7ptKBxp8E6eS9U1oynriYL8Qn2uz9dnxCTI+5s8714CGRCkIvOP6bDmmyWSwRBr+a+olj
tNwHkLsajO7+H8IFlsDCVzibKIUSPMFmhrUVhbstravc2idMTfP39uT4vTKvNtdaRv3Cdux6MaX3
x6BwjcgctSRGHsBgv53AaAoMkYGyLweqTMs5mUzPSAXPF5dukKoacJHwwT2EXi/dwbmvKQJzLohN
XQIZM8STfDFmkRhUp6hJjIYrbs8DpFuJWwK6M9K5B7NNiuCU2Ql/dQ/AUukZoCiEHMn2EZFnsS8B
MRv5C5JYfI35PzOyeJZ1kA6y8FdHOI1IqC2jmy8xBficA/BFxAxwpi/kyMvOYiA5fxHT13cSsxR7
ZZMXGoV1dq9Hy26hdKjOUgz9V0GxmY6thULgB1zZHL2tiRT+fZYOfJVIePaB5yX50yAj5uPPQI0z
yQQOMEDcoJOmQvd0yS/oaQhlNvj/6j04GMFsOhfIu6kx+o46N0Y3llt+JrCFhRPEt2bVwVeJ4B5k
XCNP7Aig4gTywfaMAYgO6aoMtp2kkpr/X1vtjYDy8GpqqJw/Bhzmx+OAo5+SdZ2+rewaT7Yje9od
wQZ8WjnMdWRTQqegma4uxVokVfgrKod+v4yTy+f3gpYoqnigNueRy6x5xnLoZUACpy1doY4Jj0i1
ziNnoQ6IycAfp2OLxY9rx0R4+bzOu37MPOc7R4L8u0fmyh2GuOLhdpqt2wi3gLPhnovlwRWaGhvn
owxzXe4QnuXL9cQAiLOHAPjQoR2ptjqtoZJ74SJ+lX/K/9AQZiw7N/V1/jXI2zkFNNmH6iFj/PS4
Ze9+wLXC7Wuerwep29XIQt2qapeThzCjq+TtKJj2l1CWdJ/ZhGSCCo6Fa1o3nA2obmwZi/TOvpNY
L6a+qstRVFkD+XkLYIJYSKeA+w21PZP0wZjIi6F0dZ7OV5OJv/pP6cVhl1vRHvKp7u6V7Rfy9n7F
2LITFSoj/pB7sRJrsRCD5USDVGBoXA0t0I0U0sLq5UrYkuXyPwvNpC6CJFVx1ocfKHCYZh2uwtkP
F+kkX1hvgflyDH+M/T1KjT/AZzqJ86WqPcd1H6MV32QLhPX967oMGT22sRmcNs6kSwpKzFQS8CB/
Om10es1fjteXMhN/z213GQ2q7hiu0qkYLZiaxwIR5Y9kNdWlApEisKc3CTOZ+dn/P9k7ffqRNk8P
HFBGqUX/9EYTj19b6kPOSy0td7Q55jgAsvDW1cSmC0qMxUc2m1Zt6ae+k80KWjoqd2FkW5kqS9sY
2NGdZZejKW9KJiffmESHTPxFbPczYED7LLeu9oji1VLIyVqRjQ1CAX4e3dyt/Mgrc4DlmlR72aQq
akpUDAOVCtfT2tLQHZf5+vVga1u8PpssPmYWPzsAo7KxrgqELq0FZ8Adk9i1VjPcFca/7swuki/A
qF0EU2VgVJDV47znL9uLccajvI9EXAlbfpfNFXfaLQ4MtQ+dkvh8HhxDHJ1eAwmV/Q7DA1sQUeqU
j23harrbM32++LJI7PlWl7bc38C+/sFi7Jho3Z0PKsaUWE5vcMynLbwAtMYP+zjyr83bd7BxF8pS
OlHJ2PfHp0l4mMl1rnUtvvnwKW/2tv7AMux6YensKMoaJ48gPcla7w0+R5k7QP9reHtA8eQ8rHkf
SwsSu6xBWUjvzpTmTStcL5k5M+veMkyJS+4NRg5O+7inEHjknsXGz5d+O18Qds//4n0aiXSeRV51
U9Bwas+Dyj2L0N+bwuapdCeIG3elXwFUkSlPP4GU5EEh0d3xAcSLdNDzCGhWUzinHwipSRu8N/Sj
owax6Z/kojmQoq8yw2etIWsdmCytPYVYR0xgXJMsIueiBgMouM+yjxj+1X+r/0c1xkqdYfUgW5GU
aXA0NMMjfgQsCP4i268JzPp/+r65AZXeBmUXZQS/5Gcx6qGj2DMt7vte8qvwUMAAjrcM1yy85Zb5
MjetDNmmQ8WrKguxzCnr5Gmv0QUjbsM/zRTiSckC4HPgdm+sYGP7dYjbJKfW1stcnL0V2PE9O5dm
mXBkBanfu6bMrn79NWMV+K+i/e2vexzQYWOmhacgIdZmNYqwvdIthWltpMvhRJyIpfusTRWjstqN
ciGxNrMrXs9uhuKekhlklyn5J72ISrhGLC9jiA4ZAKtIHvTzj5Db3lhQMxlx/c73Qxst76FS196S
zsL1CUMK15c8o9MlFPSG2DRtN+t0XYxNe+dvn/ah0MYsUfGjNGZjO6HRsv3I8l+PD+gG2SiYQ71s
d/kvYnYEw8MXDY0kmsTdS0SjpnvYWs1l+nyDHBzUXRhUVqtD65T6YJ0WtyEyihUWtaTOkgMYv3sL
DuzGRO9xYu2Q4mpPS6guUeD30xSgOqPL+PXT9nC3iYL5CzZkoc14NLTu7dwoadPXxS5M4MiqB0P5
saK0v2TV+F1LpxkZsfr7QDGfxvgEokOzdOic80x8GATtKiW2QOfkSu7rEv89HIoPFY1sTdwIalNA
hRZNXvjk27A62n/zUhZe4a5GkbQeGHLIiLWcWJptDs3WfNNH4ukj8FlHGUaf/SqRqJeHV410i2W6
ZCjDyp3gLOAcVUuvVLQCGKhp7WtbxL8Pky69mizup+0NSqH1XL2Y0T2sdIbTNs9jC+o6jsLfL/P1
N++BVTfTAtXjSBmXTLliR/Nb5WRp36xTpZW1U6o8bMcY+6eK4kxI8zKQ1suVYMeCx8aTL2XT6Wpx
bUqPkedHZTbXMHCZBIo1iFol1dtV97K0DfbxaxMBAZ4+WtpwIJc7eHMZKCGZS2mUbPKONMdYk0no
65dFTUE5UqbxjiPrapSex//N/hnrpGsbJALMHbkEufukQEhyr3tHKbdrHjND6Jw//aliWFiTUsZ+
6V5DOf4ker9VXWMuTrKVwlworGodbXAveDW2cZl5sqYzLAn1+kV7f+ZEErfHJFIaKGSuE4KY/jbQ
sTkMt0ey/ZuvSLyu9dSTK2x5FtEEXk7nqfyxvFf82uGUOMfDcD5joO/5TbvhvRpdmRcqKPFdR2/9
9723kNFIqi44iWlFvxPVQWM6xeOYya3bgNlMZj8SyXDSBK18f7wbV1DYMb99SSiK9UO4A1Pwx5RD
h7QMXyi/+sJ9JIajUrgNDjGs65Kt9M9u30tFGCznNZfP+DUWj1eIDOS07sa+Msb4FZQFPtVZIpzA
1Z7kJgDKvkk/CLzFQSfzf3lG4no+yxI0G+IpZVIr0BqVTwtbkGGe8pJ99YXva3HGkqdtzJew7SVC
RjNtCc8bwzPxH4rJ+PHPwraUo9PGSFBCd4AUwkgw5e8bh3jBOmQepdXckKjnYLcLrK4S+HEWd5aA
BPVLbZCrLO55qDj+L8XcBdzP5hE3hZNle2o7GzhTMWvPBMzjiBKnUbDj/7oDrlw6kQ+S7LU+wYn4
2jo5yK42gZNYEw5uUnL/TsEFbxMtn5xDLVdAc294/PP6tOTeObor3yt8nmVY6I0Nqn41oa7raWfl
SKlBCgm/XiI64i+RZLiIIzTVLx/RbA9Tc9/PsgNNpRRVyqzS8nQ3WCVQYMZ/lVe/zC/BU8U/rf71
m13i7GjgQ7iFICR8EHwZW4HCssFkWGh+FErejqwRJKq0GH3ebhQ7cd3TPVfUTKcEXWy5ZB7ae0vJ
1xOz/8eUdN6WSN1/fJU69b2aL56aG38HqAEOQXUxED0jixOGN+RsInk8V6xgkD497sLZ+IZfEND8
cnMOHF3K5ov/NA7rxNGoll1DHmwjPbOOI+kV8EEA9n5pEIT8HhtRMHaIBQzhtmLpRUPC/nuDxZpu
Hx3H0VlIdi8lk2SznPH9lo9pVtKm8pZJqtYfnrrTknqHFiI5HTcVHgM8k/7d++RaoTivsRW2JQQn
dU4J5oBuZOKa8pMqoVfVmJ4UVjTdvNBVLPEiTH9D+sz3+4z+5/QjVpkRVChnb0q0OXwZmHskyNnk
ZWDKLv+Q6ECc+BJ87SHXOXBAsjqqpmrgk/20SYZNEAg9nULyDzNJWypWysYoE8wiWZT0YgTATW7B
CQO+Vjt+Hhw3ZhcUpB0jaKvg7zGiDKgFGjICuusYbKAj+TCvGPNl1ckvAM4NXHS9SVGRKxedG/hC
raJoy7awPyKRUQzg59rcmHE2o+xIceHqPDDapdE51dYZatb3BKp9eWeQHVSPfDVi3m6tMaytDqVS
tnr4mWng5hHM/7VTsrVSDUNN4DHhcsVIwUl+JbMfeWw48maEVkX9rW36B+rmh//XD8IxbqQRW8nA
P1v4X6YTzWTsv+rRFcskARSQrmhQPTTUcMzeQiKb7FZ3YA1wp0MdUotRVUzmqIuLs6zz6qKfJC5c
gMFmf0bdicakMHM749RtVXQDWsyiYHz5A1O/10Z8IOciYFj65p8kn82yutF+dE6LXr8DjibGidhP
4POgizSGzhJKZAPDPkmp93fTqARU62cGokjaMVQYNYqcCIfvm8usouAuDYRg39lc4lyZITJC9HAI
BdCLcvL2gS0jW198j9L/qKeL1e8gTYN2YC+hIMTZ48VkZkXwE/RtbQPNFiFg47tKefoMNV6R/I/8
/13T7uS7dam7YTBs/rrXsgmY0hQ+VP1cYzBgM06GWHemED6wOaWBUgQqQTE6RUR2KWYKNW6+7l0Y
VmxDGO1K+U+Z0waRvkYx9SWitwRCpH/7OS47aSV8rbSCTangY+5eDjE0U1Sb3raZyCQ7U+ZROuQ/
fjpxq0urrrBJgelef3oEdwKUdQSUTxoOMFjp91YNGKcldq4S9QqTKA+wJeeW9UbmnbIa3V7vilFf
xjgzbyfVcOglG0mdGwNDK68sGMEFMBtMSL1Z6DCzvOCVE6zi+f7JVOkjvRdO0jWpKSnWzrnfHCjL
WfWrrLkC+AWLYs7D+eG1ZxJ/p4NWZSZzRSVExpH0vqQSlJxxyHdHMwV50neYSUJ5KssmdUsE7RNu
jMWeMTYWm0+Gw/lZDT0BTh5FTB2LXV3axehosCpdKKsuPg4CS5VqSaZzbQH0QraKIhG9wCfPyb5g
QOOB/L3RodbCiRZsQdMOkE/Od1gr/IqQPEPKifDVUpUx/PSK3E+ET0aPO6oz68y9Tb8I39nTbYws
+7PhwIRKITuC0nkJknaoKvNWPPTMcTLd7d3iQoLaor2taJQ/gkZlfIP98kj9hx1ABZgZMfZ4hoqw
A3+6XzxGEccR3bMVwoSHfxN83RrnjjhJfKxNSpGivHrRn6vABKlOu/fajA1G/qndXpgk1/Hl/6Jy
cgUFHJsxuS/vqPBJ8U0vjxHkDRB781CdvThoEf3xRaSWcC0ToXXMVo8kBlO4F3SLia7UMp1Wd8ez
nSk/qnH/mc0kgBIruphFH4ukKrLqIxT/cSTJ5//DJhhtcbA5KE30hVqOiq3sbzbwimu0AltvJ4se
RFNM/W6A3ikLaQJwWAvShoj+mWYK4wlTgUBg/+LqtvBBVNuq9iKG9t5bZZ7M1YL76Kk69MLcIDYY
mtoLfSEoYEmkA5DNa8b38nSyRvbZtngDDVHng6O1QJE9IcSkmPT+iExlODOZUJJYJb7ly5gAytT3
IYQGXh6XVK13kVBm08uE5GvsJ8hJQ5TqZrvJcNCzcjlNAqJz4jwrtD7kkLL8YLATzC9lM8vojzM6
iKAFRrwJ/xvYyyb5gh8giZdEYomn2Ovb0fdFdXBTVrsMXAVBMhE644wiWt8IxYpVz1BNVteLmpDr
NuP1Bi4sbo7UDKR6GLQ2+a82sFDsfLEFGCV74PCIfqurUipXN2hbWU0LoIDGWjwFUiYIDBQaJA6M
01pRPEhPjU6bIGh/hmjYeSP3rEFXm1yad+13/dICj13PwBI+04rbZEw6M6bD29BM73FU5k24h8iu
jP4DWXeHU4dn1wENrqLZXXxWmBYaHqZWfmcxKwmYN5nZlM1E09xDPvv8kBeg9ATURVFvEqMBlfcA
jkWY+DJ3MsD6KyD22QNScyWKfrDQfVgJcd9a/WikBxSnc+8RPS/LwRzdhsDqctm9TEsl0nxeYtHB
EpXhou89Mv07BppPUnUoow1HvmW8gvaAIlCc5RPyQmakBgBjrVu86iKkliTbzIobnL72M0AA/iAf
n+1NEMFdzBGR3YoMERUdaUc2u5NWvHdSCMrIfJSc/KLLHulHUJKRbimrTFGhxlIcP3mr93E6R0MT
iCyknUABmd3soE9m/drR0YzB1Ao2gA7ZDA2jO8Wh/0UkKT740KjXDPTjtrORrl5xnhUnKnhLSKp4
y15+k+D0oNbVlJIwd8ayJtdmYLaUysVT0wUkMgcCD9o4XasgVNMcHlumdPaXOB4i7+uTxmO+aOiI
g8fWthV8dIZ4VHVSzIb0KQJP17nipOzEF4XZxr0srHnrbnu9GYvkyUQCIblWo2qtEWRRo30+NZAB
t3WXfxuPNYLxEmBNEj9pOFZ8cg/VkA0kfx5cwA4HFYJ2ZnNl7zUXr4lI5pSB/JXwbxmdueSlmC8r
SroF5OIiIvneWJ0iNqMEsEwNIlyByp2bkGAwqGQU0axUe8bSu3SOMb0gczrfHT+5gVJldnItj2ML
gR/n+TfmtOLg0Dv4Ub128qVVhzWs8ZMZsNGklZtjD850/DffEjqektba5dgbDvU17hqlgWGHJC05
fq2VRzeGbKeSi/n3RpNw7syMqUMV3lwjD9fh+oSv2IaUXcZJQGbDC3prSHh2Ab+hnmvbWMnQ46k1
uHtQvZaCPY9jybXBu8EddaVpvbF4PgTkmQZ5qK9UC0ifntQ0Zol5KuilEr9zsliNTjY4vGkwsU66
Qfr4OLWnKUcH6dor4/lAh+QW+e+oxWshmuxPwjvr0wky9zJSTIJtrP1W5i740JYXblB9PPOppHKG
F86AMiR+krw1mbHKdSLloaLjh5+BZBa/lrVmMEdw3SwvwL56U7qJosn/6b/rWKtP/y44T/Sc+QSe
mjUYe0DuzbJV6fLoXhs1560+jvQ4Z4NZUlOEAK4j7lS2Q+JcwBGMvSrwCUw8gmfVVmZh4195iCbu
SivYbdW2u2iv2GIyhzGs55lD5jszqNv3lJnL7sDVfY83qnuELKit9Hkf70BJM/WuOvmLAkCpf0+s
AZvR0YVfvHo2CcHyKdoW1fXrCCUtIDd3SykgdBwn0GzcauiG5PQAmgUNUStcucp1FRKhWgG02/zU
jMuesa8P7gdE7YmdKLD0Zv21XyyCS7RF2rQsmWhQ6i4+Fsl4HhTHLRtTDig8c+KAhbSd6ZTbfIWS
lMsBYuyNmvl+alj6ZkPHvPk300Ft6WIPQaEYOv1Gg7RtrekQJfORMGqKATNFAzoUZmpPLW6IEbPM
4M9V2OZE6np2ahuWHv+Z43HhcLlWIvd/P4DqPUrSz4/jHarUunkqoyz+qC5sazchZhOldRVdWdBV
6LKylivg5peFqwSQ4lLT0PPfzsyeA3RILW0+P2LeCte30JAwxf4748jFL2oK7vXw60Ncuj7SiK09
/6WRj0zqmJsu/Uh0PrDi/48TSJXZtLp0TKHXEfSXfc5EJ4Qw2dOLccZrekgjVYh+VB3Th8YiBtvP
KDW7TgVhWO66Bg4nh3HI1hJVJBC8ZwzcaN+r5Gs7DIpO1abLXYYHVMfM5YesT6Jnu3kHd1tb8z6r
SimX+xCUBpY3ddhtnmUIPqOuFaRrPedBSZ9lhqA/WjiEAj+FMcLw98WqQJ1DKG/5MfUbJ3Fn+jhK
ycgj/t6pmsvQfCmdYCpdbG0QvgmjO4/hmiJTig7E6pBuYs3SZkXE1TcLv4hC2GEyWmcFKM2fKwF6
SRuf6xZeaCJJZLOjrLB3Y16LA9xio/ozC7DJeGpLKCwzk6C7Rf9alUiNmi9cPSJYjeGmDg1kxAJG
IxcTFokWJ6eOb9p74IY8rnu3gT3Jo01faogiYBOJKTUpWN2nLmXLxgHDVWsEheieKADv71Hr+UwM
e45ea5Cke991RY9XMrCN1WPB4kGJ/Z3KqSFSvpMugZZQjEhK/qO/5XG96ZqvKHhrmCzfbIjpNt2s
MV7Og+YOqYew+m7PO/j9i5yKfTXPFX/l8Un3O6RDpliLXT2tKMJx6WYTBJmQy7ChxRlryh672GcI
godw3V8v6pLBz/x5lVH735KCQhVuZKnOV6NlCnjYun8+Rpu3i83N+B3CQYD379oPSVJju4vJE9V9
zt5MoCvjb7qsQgtg37KQxkhbI1/4OyNRfsj1HlzBpXod1GXszX9aXZXWZNhUvuJvGaNUeTnKpmqP
WzNJ4ukH58aEEswR8ENrVXPFkD1KNcKLKTCiGJvJTzFdl9/2DQLoMAurn86iNo4/CRgvpeS2cKI6
fzKchmXVe5jvj+CNNPDX9cqWSohu0dXdswk7qUt2SHtBLeQODw7zt91VjdzNj2/V1UXgddKQ/REC
uthCnzB7BOuVfmaUDxYM1bJUEcP194SUJVa+ovhqpgamXgmc+ydEPI1j2hTMKLcreCxGPTrn0NVQ
5IEVbyW78JCP1k9a0GL49p2VwkC7kq6//bDQrU9ILGvXt6iUIjCJlGvNvdIoehb+PBkvzRO8gU+4
RQ0JVoBSBpu581VCGuJpLyrLqgSKUgp9+DsVSw+vr2f/IjrCKhZbMNYoo7uGFe7rg077kABIscNs
HY2AiJg3NeyM/eyH/CLXG8ERpdyl/IhRFT5mwviHqfB394HspYzJ2BEAEWDt984k9bEFGisna/yd
lW3CuyozgHkYy93t8R/azwN3rGycWCGOwTwwSgbHXP0UUU+zOOpnBpW/vu5ZC9upW+gUEolB6jZ+
cSG7rJpFNqPK3IT2kBR7Xdi1Cc4sifnFtaCilPlKWkCt8tH8fkrIKY4koP9az2whEHP4XfiDnGpN
pzGQY6sjE9Jrp/19v4mwrsRQ2gd5fXLwhbe+4jXbwB8QmjQ/A2n5dlb7aye/krtEOvgVUdkSR4dY
ZbQvz8UFk5YnZAcFGUdWnX13m/1a/8cmqKHkfKXPVGLRtxLUw6XlcYrxAWrambDVvnQFlEF6LMXe
ACtcmiqT1K/pFyZe2cFZpmhPzWPUzZ4KsTor1y4wTpGcZFvgvO48rAQ0CISAYZkWMDyoS85mXiMO
zuLAom+sh0NIDSxBCK0b7FZj0596URPuvlJvXrQpyR9N9/cJb9tFasXIAuAq6d3EfpqAXCyRQ0n2
i0n48dLbuF3T+UbhR8MdHb5PEZDwS8WuZVarOISavUrcn6yOqd5nUFQWT1klhZZ7Yfwx044M6C1b
IQKgAFA4w+szWsi9Fpl+Lc1mX6xk7uod0YGTUw+yuQKFSdR3hiV+PpsiwXPSlTyEJAu2kR8WFnCT
UwoR/Ks4+SnUv/e3evihPMbYUFTvuONfEKZGmPTSfnblZdFcJ7egjJOw9vpyCCnweu/+c+RDSqN2
5hy3wkAU+4g2Ew0983Bo3VjmoIusiN6WzBqZZv2hHLsesKGDqL7sGREklcI/MDCWsGwZKayQRGS8
hTjBugJ7A8rVyx8cW5izLrjmep63zKZYrGWNnHkUEbr2KR+qWqyl7MKY1Yf54P1ap3e+OHAIm9tG
rWKQ8DlHbbMeUt7uOaj2tS2RM/kVsXb4Rr2AMEp7Jolv4RTsNYbJnkOJ/GTl63O3O9sOwLNGl3OJ
mKU+dJI5EYNp+rh46OjyCEMX5r+27vVP+VMJJdVR7l4SNOfSwpPSIqqUAu+Kdv34o05SNf4muo3K
/0Vnh6+N74b6F/qajGCQKOMCiIcF/6G9gmgiZ+iFbDwxRQFgd4NhTcKiRPWnohQAZhoZdrT41R/a
5HJJwU92+FDC8+5a1iIyZvgC+xrSEol4ZQml+NxruO0ZbCMC+bHNJzDS1h1GRJ3cnbBUULEGKsRO
sLBsh+iWr6XVfsDXjjbrQxh9cNAbOfs2mTySCyHNlyutdmMxTJBh/EWlSB+As2PKWmO1cc+ZBxLQ
zEyyCkn9cKuxQsox27uiI5zuIF6FHA64QZENoBDXen8j5B1ulChNdjF3D3bmPhyECrp7gQlOASoh
rap32CNGf6o2tYuilFwS41QAkCXJCqZq2hWoYns7pRlfdrMxg5v6pqbm0fK5Escc6K4hLeEANeuO
eeoR6cn12L66WEyNXwUoAkj6hp3ytDqHQdBv7lTesI6YpCgYy1GzAR9S2C4dG4idhv7Ny8Pdk4PW
I5dxMxthhAFY9ZC32QmSoRxR4snhboYYBS9UpPVa142MTM0chLsvmuuA+9prR7i2naXjqdpO8w5v
HICgiwNeJgFUYWIEm/pMrHD4kg4BQFlex0WuqJUC2pg+PJdFkhWz5kJhozFYqAAMaC8CheZXEK50
e/GK5r1P7lGUgWgaloaP0FtgqJ7zWuEyjGhvZIVNFKSeD8C7Pe8uv3HnJrt3MFkzkwYwO1cm0P77
rK/GccUHrva07GFwgaO+2YCNXN9FJyNB1r6bNMpLkmaYlpzxwDAkJ8M328wCwGIEPFOHV0X91Dnj
0XCmhvONYQPkldn/ow62OyFMVHwagY7WxKH6SEtYRlIUWMBdpbSZO2uxIM5v4vefFXOkQXotuBs0
hcIioyrM8RKTFVk6sWbHro46eX+cGuCqPX1a0lWmZBOWTkBXhR4HlzmekHPh7iF2J7dezeo9PGr1
hW93al5iaoEocqfGQl/hJVrthVeR9QBbJ8Ak1wFBsy99QsvyPPoq8fthlltRYwluCJ8ljz4wj5GJ
Ff4e38teJosppkPyr9zoJaoC1s0SuxjhKGSPVweRtJFeIKQ7gxWlLtjfV4IqSvvE4s1KCBZjQQww
gMwbUfmEk5aRBI0vq3e6G1HIqVGy8FVGLTHkDyILNtVo6WLIuf16k52k0kYLppLk+AmLcUucONBu
l5ftpn3KkA50WgY8Apw1uEgXN7cR42ymJc9zXcGF/ixyV1hvuphCo7curIOio9l9L6hbDBN6PXzU
mdLpM24fuHiHjIwem0AFzZiLOBU4mLDebqCYBfH7TdTUIsGZWSP9asY9uhHG5b3b3yTYnyKzHNLa
Vmu/y0gz5HHaEVGmqW14q44HKSdw4wgn+0obUetXOG4g2+kjS0gIer9fqkwNlTXrdLVhEMg0gYlz
q3fjPou4lYPzjiPYqkLRqfMDL2RoPj/3cXwIpyUOW1iBq04lPFTdt7+sgRl70hsTZrjvGIdjhEK2
rPSx8FAEvEOz3W8Y2Jr7qiF+nvHLpkWHqx1aCSeCWb6uh4/8umSBgUnrIB03ZPD03UtgUvzwlQfU
lyj4rjnGfLArxeLJKsRyd9+/EPJe1yqJ6/mfah650TtNJsTQdwGE4SwH2BMbvwJAF64r84hJiNNf
+Z5EDmkDmu7B4zYaR74nD8txf+qq6Z1mqgDu3btdOH8zcEDfWFPzrSWaY6THITR8Etl+vLYZO/ry
t8MyKBeTLbmyjDVijuxhPWxUsn/Y0kwX2o+6VIVFit41qh5L9vCOgwZlHXJcZSku8d5tINHqUWPE
RcTXuacQmuX192RIFB4V+xjm3O+H/egyh4HkAMIDxHC41u67XBePjd/CgDZouVmKNSsg3kOQtbZu
hpSddokJVGYGrALCd6/4QZj6h2fVANJWlf8GST0yC1U+KiUI8HC4nEj77iwBqvOnL1XKP6LPUIG7
jkwSJnZj9iYFgEavc9UmxoorKAljgyjD+KNrFExe0PcwEBtXCzNxukziDogeEETOhFfPqja97srZ
04Z7xV2fPGse1eJhNpqkkapp+A15xvBSWVh2LndQFHkyqSZjjDH4tMB8brKLKokF7mzIWK3P8hJn
QBGObPsih+VXm4RLOxM3Efb0UHADLwmCFr3tanBjsKLargXIXrNGv9ZG3eCVwxtNYZIoqYRNzBQz
ZT7lXDcbEFBxUI4mfWUgKD0Ks0I6r5B/b4BOkLiYmAavoViVJ6MRwKTP6yeuLAn4Bi7eCVmdfBvC
N2PG7ggGR0ldM9ADws5WEoJgebjDiYtZdkvV9/Kef/o3enMQ8NGFaswR3CpHU4akZpl7R06vYFNM
xlKEVBNcXrciPcnYJyrNnykbP9ykYw41mpMLACsEoefQklcwZ0jRlOc4QFGLHYpOKdaVvD2fmOVD
A+8Uz5hAE/14U1Q8lKTixbUKMank0avO6CrZ/6zV1U1eYK4NBoFlJj4HW2i0rLnmpl7BPEVKdt4f
v6ukiA1Ka6JgxChFUWQUBKNru2XYoKB1zkL0XkR2szsynaJ+8e97QzKKB6oEdSuyHfH5OY0p1hp1
iMZ6AsSz1umamJfXiSnZeb1JIyp5USk7BUeD0RvHvDt2C0XZ9S9glanq9Z7hqaJMryJPOky7nwK+
0PfXIB/oiXzEhJSIN75m3OjZPpUgM6bxrbCFAwZU+pZcXo/r54/hMPHW1zgVpyVfLPy+2vzTa7cA
FcknNFuqiVis20hgBQo5XCUNw6TnMIWWu8ARCO+QH47f/eC1UtSj1RPB1DUlunVtE+0tlSUkcM0S
+CkgmUX0QNEfSSap5ADOHqagiPSIX8wHTFoZ5EGZEq4xLNoGxFGGX2hG+6yszcNpTnBYTTw1FENw
n5XNAr1KDgkK23SGg7DcCOkk4riKibLu0Mbr91ehp12m+L3KPBtOxBF2QEGoab8oWqOdga9ilks4
PLs4x3uMACp4N4MnpPWGqZ5a9eTytT58f+xl/ZwF3TpdyQdFl/y9COGnqO5ipdfT5Uq5Q0q7LFwT
thTMvMlehrL2WWafOtsAzB6a6u8catFQmmscyjp/Ko633x8SSImEni0vmHsSCqmLGAElQGNt2Xog
Kt/akAlHJ5+ZavXqvCO/X5qe4yxwk/N6XxoqhQQCAD/eVwBcCcq4JjLtDBI6E8vBuDygwqEliCAN
RTd/jLRsolEORe3By5gNCmh7wt/2EMCfNOEf2Etb9QChsVVfhGB+ZdhOZOufVzdlQI13y8+4lmcH
6L6zsCjv8xtkl9EUzPojkm7j5mDkSj9qCbPW0IIDxjoONOdMTRGHGw1ugIiwwZQHG5Wqiv7jdviJ
CwpTBiPkAkIzGVI6RKMyjVMEZxRl63yfVW1mgyjCGgTyDd98MW1xx3x68JtDiaSRLQhljFkNwcFu
mdZfDifRQsrACFftcmOY1m01dHolsyAEbiBbXfmMlQy35UgjLMPreXoxBKCz0rJDn6KT1CHEES01
f95P/7nutmlr/hIfqmYrcU02IeVNjKyYTh4zfm9Czp2DGpzW3BpBFVLSpbinKOCZ+hBulzC3tHW9
8e4c1lDbaV0WSfaFkblyeQ4FuG+WmCJT1qFRNhzbyfCdtFs5r52FgCqzTbWiS4qFR2tIjjXnT1Lh
MzA57dgm7qEQ9rxdH6qwCpIfYdccKQEpJa7zcvvKBnqtouFoW11uoBkCI55GkOWMRCoP7pvx1e9C
VAZiWeeNevrMXQveZxcwyRNE5JrwGVaysqO/W0fcI1c1CjmKclIQeEg7heG/JNMQ6wt4wvGOPLQL
kjrVQCc4SVLRuIpiMnnzzZGkOQlofAZp4U5nqmcfCX/CUaALkHKbRLjuA7ITyE0SRTa8F5mrHV2o
BM//bM9MoKYdiJtI8kp+jniLOxLlLtHEcY7Ihag5WCNUTG79pgbbTuPuevcxw5f9nfYX7+d7eIyD
ryqHCqT41vpWxihfapofPnyI+SN+8baV8LeQGA1WDETmm81GV3Fea5oHxktwW96HON0liOcC+OiE
B100hS0dq51m5zrUCvbVZo+wFfzauuURl8jbuAaZPpdoq++UCm8T09OIIpP2obpd2CfyTAn2+S6Q
UZZv2TizlJy5x7ljO6dB9+DzeMyVNY0iQwYRFUKZOrTQINPGH0vtp6tfzCaH2I5h3a4gZ/7QBwf9
B8pQljMU2lRTwVotebgNsVHy4l+DXM2OYHMaa48/LB/0ik21KVa/yiEFx7RhyxSH3KpiQTosk6Jw
XUk6ibyyaeC/1ERZEZaeKTVQuUlc2qhZJm0EAAJprCWZhBzozD5bNRls6OvkREJaEPgmjbwYlteg
2zoysYaJ8Vw9Fa9F97CIojPRN4lIdtTDO6m1Z33cygp9IQTVYgxX4Mrv0Mvu2frQ7dZC0cyk9Sc2
SRKIqwwmrdGy4tjMCPJdP7aOvr1+BmLBD1uO4XanPJX0ijHi83xgD4ymU7tG0jE9ae2tmeADMNAt
W7meQvl1M6U5jHebaOsbnhgHnetlnnlUekSM/3iF/TMQag5OPeUP6zAkTJIP8QHY5P+LjCn/KR+9
wwcLrZ74d0/0Vn7rlLepH0S4QArU1uWeQrXNdmLyboDd0XAeHMhP84lVyP0D06sY5gRs5hxKQO9P
4O3C64/nE0fSM01DuQ7/vSMovoeIAyG2gLu/rbx09oyMcde5OqoKdicSC0u9gFFDgr6L0i9rhM0/
RzZ8hcskW7Xhk/UQchX/HurYPbcgIqlCk+QFLKbvnNCI0ankb/3GsphsRwE60qqu8rCDcopdh+Cl
Wd6D21DpEu3K2jA0Bu/2LK1feaXJ7C8FseErvzz9x0/i02DVzz6/enFn5rOXQgzLGDw+vDny8Eff
hqSqzIeq46TfUfHPLT9m/x82VfEnWS22KGfSKpbxQEsLugn7dzOYDPz0MnKQ8dyIdwm76XqmHij6
bz5zZMSQORKfuv91NJathHhYnDEL8fGow0kxNtNnQJvadMGdBtZX2JmLSQejOn9NUAYOkyj0UUy3
z7IOAfpImcZ3m/4EkCXmxpLb6jOCdwMVY91GBKY9VUtoYMezaan6LIiSPBP+SbypwHLe5NNEnOnZ
XPjMc3K2vpgbscXM4G9kTfZEiDV/lGY1bfJlyqcbruobVMR4M6eNXbRZteyh/sAMX+UDF7sLrioV
aX4SCU+Xr6QGq3zs3A0w1ivxBtOJBVvO3933WULtgIy+4McudVGWZzrBa5rSqkf/wjvb3GahUMZb
7cWFbaott0n5Nbd0xqh2COs79h6PIKb4ky93INeH1l2xetaOICPS94cotc3UHusUwRE5DekTRdiz
7JU/YemoFp11WgguR0aiqsGWeFHrBRN/pylUDo95iWJ3XuUc5tmbAndjj4FwP+b/3G69270hqcKL
VArznsiHUd//sB4dtou2EtfMbXNcEU4Zc3ewzixd3seGxdGl6jPKyo8WCocML5FbO9ZuiveR1fQB
90mlLiQhLZIYhJB12ZKIeCDJA5sMtwzHipK48OSAhtAO1V1av6PHrN4Ewn4mFIhVJjkPM1bRTKtW
cVnse2lEyzO429ygsZEk9roJlGAAZ5CsJ6NQ7vdbdElVL+YxrQpIds4eYcL+Pf9XxtiXnmXEySu1
4OnDVBtlz14lMZ03SD7Nk5ucDbYdeyrHfPVtw96UpMGgusN8QS9Mmyq1FdvXcQvnmIJhSlefwVvA
QNNyS/b+Qg+VI9CDIwJGbnugP7IFi8snubZCQDFGCSQvYWzfwdeN4cVlQQjw8kYNwybzmxytpkaa
Ia+QMWv1qItX9pMcnBJJxPWgK54UMEy0mlQFZbcBJOx3APVPD4XWcj8U7ZyDRhuV+6on9/s4BhIg
VeVgJ4vpCVatovbYBSPi297tN4j3mZXhyBTGzSLNpK68cdc6ZHnG77RKq+8yb+B9c6dCZaYSaMVz
+hC4I5wXVBJtJG1k6qtWKYmZjqVyD96TrO0MShrwrpZb8F/8Tdodw5hsUkWm14a+6YeZ/v/tt7td
18wcmahnxj9yoJC4jmCC79AgFZAykvC1YQqY/CULKDT29zPslsM8Ng9rs+ar7OoOV5QRsVxE7b31
aCPoVpI+nE2km7G0mDSne7PPRSOJiyAoK47n+858sNUWq9x1YjTLWaO+ve4wOuonPLTv0W34G6pu
bwEmD4E6r2+pDNugln2dMkhf+DSDdjw2mL4QF7meith3F83PqUyjKSw4VfdW6XpqGuMELbI3AFBB
zJQQcrypz4dMafRMrzE01XbeRAkpM8ito+s5kBdAtPoeOtfVkanotWAivrU6SkHLV8Hy/B0qdXhT
gd9Ac2WT00F8TaCUaLtV2QPys6aQhD3jTwX2O1KpMbdlRf/DODZSMeTEAAeErJ+prP97hG1njYiM
SWwrNxhxocl2q+ku1G+6q1mYv+gQhpdGT1udLDrbZApC1ytlNAauVyb9uyOqzT7Gyrb+ra5iW8Pi
zaees6EtbTPgYxskWLVMYGESB4WqGkox/0LA27IWxpqhljDD6pPw38GezoWl9W99OzvGb0/o9AdD
P5znFAKkRSLbtZnOsIfqNawSpRpsLuVL8v/K5braugvSYwXZVV8ufXDR4XO9tXkEdAh4cSa8wmpe
GxwRZsChLO57cW+mm3/kOJL+BOJeUnyTgfUSSaX2SOHBJ4dO606HUlTY7g8S/Tr95uE6Gf88JKPg
NjB2cTD1p+eJQRLuSK7Nw8Frfn6jevJ8nxINouZRmqwQBAqdRTq98+aPDdhFJr69TIplRty3jxRW
IMtUk6ucjpVszmq4HjnT9rc3vEjhUryaR6L11sGZGPO7jYR1tnyCLwJTJprzh0QmQFAtzOnACS6h
IQRTfen4BXpUPPR2tBFgEWp2Tc4c3GMwHajSXKCPM+Lrqpz62A3jlELrI1CrVXqS80Xp/9UyCA7G
fg2CxnZh5aTNxYp0SAue2lM0AdRuAUfR/j+H91DzwA7bi6Ul65KUAjPtRzDoRfrUhPy66ZazthTm
9NMArecHd371ap+dpEV/ViWcjS94BGtwLpkCt9p14pd9suEa48ghjTUCW6M4dab7Zf+aTwf54pbc
sQgHyxtouc7uWmRWCJaJISXm2J59HUTR5YaZE3WVSlV/7oateLfjcVPu0CZsvgkSodRCTpbyjROH
kIIbfJUHhribtvRpwsKCxNH1TkXs+2NjdF1wYflXnmB/l0OsNB/M4PBJwiUhIXh06OctHhmhdnvi
Rwi2WqemqDijv0RxL6riGwVdEvZb2voyWVdPmR9U3X+rqDfg35xnmnxRzuRLTwAL1Bkub5RGfn7n
2q2L9jNfHaWkAaojqf85EU3sacKn6AfBSwwT1sisOdV8csAR60d8uBVPGYp7b1JYvgOCVroxd4Jy
JfbZHhxxF+qLR/8EOEdFttkAw2tDtKgPbS4rxlFTK1jP7ZRZoLXG+S72qWDf/7CcGtXQpg5oQH37
8lc4Ik3tnVzf+WLjirfrFpEGgi/y4TnekMB8sK7XciumySN+eQhUwBTXGiW+HKeymzlPY/nC4eqX
5Cm7cRoP1rT4vuPzOBBaxSOa5+MBOZrhQNJbRF9Bg4csyqPqxLaasYyfJHzBPRlAmLsMMhvauGZ4
kciOZ0BJOSn4jRBn3vQZ8h7CxYidhsJpB7b63q3+y1HnSXXCHhyR+OWyhAnTRTR04fmy1p5uzDDP
sgPXhn0xuQlziYtrv/Iqt9vELbK2NkMSrWaeqFll4aFoC+c94rArXmQGlFg0ardmKBavJonl180/
YAUB0VtsXKr0kKDOnrGkcUUdcGO6Ae5BXpAk8nMWOcxtom7IQB+4xzYdhXhLsXGZcRySjKesP48q
fEbe1uQj8/KvZJJN/RyRguCiAPHb2CnjsZZLcfCKQCfPT/ktMkk9b/6OY1Z5QzWD92LNhntK+62a
qHhOiEfkivqsrlpyNPf1++4km9TGfpnzAL/Ypox/pBSJJwH/1rokbBdkj6ThZ1qN4gOmZBlNGQQI
23LaFg4Oqo6uCuPTAeyeZclepFIv19oFuY+OuUZW3Wygt0xKcVfHOVmCmW1Isq5ELSjSwJN5P0kx
vq/df6Z7+vuesAxndrsT3pAggDAWTjxYw7ql6srD0hA/Uk7wYANhp+sR/mbB0KH6YUX7SgbtDSZD
iboy/ixe9Qs2asU9UKde+x0nAe8f51nt3AvXrBB9K0bw+/1Cuhuv3YjVoVrNtTNgHhMQpmedTxKp
KN2R53ZjgYnkmLAclHEG9o0B7zkWi0/PAVTp2qqPVUuo5Li9qGin6q7qWEkwGyMMYn/xKh09v3lY
e7RBBfghH2mzD2P9zdTHt1yBY0p4Zd0Lu5g3XffxQGEtfeIkzzH5jv6/JvaylIgFsBVTB5WTzENi
Bwql5jXoqXTD5Q6KzVs8gcA4UQYUADPpVEbNOskseqf+EYWY7//yEZC4urK3U8COZ+gSR8wxjoJZ
mFB8tMvIC3sT8wN8eZnRR/9MB99IjP6KOXsUwnwXy8KtkznbzE1bBgpt0O8oYJjlaDXm5NMdopi/
ZiJg6OF3Lw05xktXIQhomTS70vCVkqdak/ryYdOk1shRTS8wB+awDAXs9CGbyQKLxiQJbgVbTFhJ
o+q3Fu1jV0dgJsOdsZ4WRqMNMAlLQmbDXU/GApBwEPdLfDhmZ9SB0nhEtmqzEQfv550PW8Dny2gq
s15Hb+4fBqn0aWqgx7M1Pbm/spD7lxbaW2lNBZ1Aw0xOImfGjaTnUKBw5izFqmxpq+4Jnw8YaOD2
41m6D10GvYZkap49rUPLEaXvGbep0UzZ8QRnCiF42oiCEOazMAPDazcXARaCXzqBOcjeCv5sf4VW
nXuMkzjuUkifd9Yd5j86aI4Dp5WA59yDiQebho3t9MaA5iFVU0bDWp8dq89LSrImFml5jEMikf6h
EefSkwmOeFYj0TEDmhdxMRfrureuceu4UCc+krymY+w2xLrYwapmKngRQqL30syDfR9A3vKQts0O
1PyS0ZffkeI4bcbKUz796Ex+UrVjxUwGIVXIR92cYlhSnqxp5hXUpHuTDLTc2HYobANJCbrBZJUa
VMf5lyxGYHrIYd79oqMW4wAM3eyqFKaKwfAYG0h5F/m2p7e0ZJDjC2OZZ5O2HtxZlgBm+DH4GwgA
Jig2vAIDjm3p87jZg5YMC4wPHubOypsDR6NQmhuQl2Kx3fZlvf6g7JQYd99I0eQI8S0zO9xbdrfi
zwa0m31vk6Zs0Xvi3RjfSsMIkKgTbro+NNOj3w5p3BC/V5QKm0Mmhz+bglW01lFsXaxH0e0i0k18
p16kYRLjaASe5VcJ4zWHK8dBEU56BJFyWBhmTQwQyeVpkW76P+L9/1j6LacdwmZGXp7qXRsXnnb6
Pwv6uwDKzdFrPENTR2V781LOHGPzP0r7nvzaLhUJGclrOVBxvMxY7WXl2hVUbhwMPnlebuoXsX5l
LSDq6l6sJvh4mCa5J8hhovMbJVhW/XFZUV9DAioqrJLGY6tpVdqp3SWwvceub9S2lUGNzzV9RUxU
Btd4f8UdTBOhVmynVH5cHy5BCkmQrpvE07mCxiYKnwabM+UgHT5mYNPvmaUisfYJVjx09RoB5hE+
95UwOaM/z8oe7j2UnGVBDg2JvFbq0Oq/lVSDCEwQ+51f2tJGOjRms9j1XGF7LbaEq7Ix2k4DSZTc
MGDeJQPOanPu8rte1VQSqmyuVGu8CRJ7YsxKzl2+JmBBc6gbYd1ZsqObJwCPzQnrOK986rGinL3d
b751ykUZiFOFzdu3e3ex4Aw0j56BFRG0UIBQ2QqgNaUu5Z0MoB9cAmkj9CvNyEs4iRZcXlzNm8rr
b12hn5a2ZgmmcX0DFEZBwXVnN373SuvazaOSlz8MiHBFRBlY/ie7u6hScaVle0s174XYok3jErRk
LenLpeRrpHUvMn4psNmY7fma1tssSWWI1yiWrRQF9/u2chJzTWjyTdFJr62t/k6XHsYEsFJ4oQ+c
22NT/gGgU80ui0rhCjqWVYUhW48wPNspzqrQOyLFgqUyI3pNtQJu73uYeqGfujuylv+wCDt9JSdC
MRejH9vXyR3ypE9dL1OQtzPk3PhkZ5/HqsFsZYi9rWokTn2oSddfjOOHINNPhsryVQ0GIJIB1HA/
Wv/PJmVj0pt+W/g8K28rXIIg/Uam4ksuruqWl6eL3+5YdcdjrPpyoD66emdSgxnHwoYl9SGZoTBU
+sd8H1G7l/wIaPIeIK1Bp4DNIoFe/xW28w/0mTiStNJQFHF/HwaVhNtnGptFx5bc/bK5PH/bg/2W
y7JAL+GF6vZ1dBWb3yS/+VdmBaU0lEMFfFePQjOIk1AZ6WXCHhP7K477SA/yoSPElDcsfYN6OG8f
sWWbVQ7YIVIgyVlXt8/tQrVqGpy3JZYoJ9eYlCse3/VgS2X5FTzVd4VVVRZb8Z2lZND1J34bJSsi
OlRNIFxGo/RslLBBQqBY6oYcte7Z1RL8SyRAWfRD0N5BIyVypUMBLAgboJsF7tsihDeNghyBcUHv
schZWKWhwsfqkd9Hir8J35bx3jbeXA08Lc3UjRpz+gkmWT6mgVtXrBSLiUgolNCEo6LvcQDvmUyr
IUvYrFQUDH0J6MCuwomZ/tDKPN/fO7c0dWu6styQHJaEpDJl5ojAxxKK/SfVkIBaPt+Kr0ec/esd
VBTxe624YrkWvLExaRNtI+KsygciNR4+oIMNARABNnWsx7LQgzzRISReymh0JqqbSWDCpsfmm9CU
4Fw28Pxyl4047kmqXuMA/6jF0hK/Xc+5Vvd2O64XFwC5FY9ca2Y2+Q7fNdyCzGfShpKC/eHc/dp1
qx3jFqfbsaZAYG2l58AFfQU9sRoI1yolRiCv11lwtyj3mSQZPQwYsGs85ByenIBUYQ1RmrLuILfB
Ap5VGiflViVyFS/gBSJX1tAG4zbJ4cMvu0GzIUW8YFk0jc21RP++h78M6tUD8VbJs/VsdH9vqfTD
EzPzIy8OkZdzCz6ChpyOpkFUOsdrHiQ/JqfSswPgiP5PiNXk7axuoU0OSFdzDcGlM3RedT0CXVXn
kUi6NUUOBCCYD+JrpPkAT9C+7+gnxuXo8uhbqL59TrchchQzuZsTsjjfVNN+AsfwLxlDVLaZF7+u
jYmtvesB7sqRFNXNGn+WjUBFRhFOgL8CCq7+oNdFhPJsNtKPUr0j5fWwDMCCoKOmvN5/gClopvW+
oTl/vwuk1ZF8Fva4r/ZSHj8B86nqknHvEgyr8YyIr21g20LOBNZum97Bj2YGifbH6tdWQt/gIuFz
w60WCnkb2ehjgsk2QKJC20Sc4eJ19upGRoTRNOhWupeDe9S9gsplUhSIWJN+GCiYdNH/WUzrUJxD
d65sq1hqUdJPXRpEsuRffw4RzXeug4DCGeSuJxEp9n9krECUDp8xGu4PXj6N53Z3J2J2c96AMAIH
JVkSe/DEMIRqm0h/S5L3iOVDrscocrBwO1XBgfGAZZFdmsbYI8W+ZbiCjcjo6M6/dKWPdOQEMave
ZYlzic9js7NvQmSHnJK4kiqTfhW0EnUDY8QCtggU3BZcOyDvF71Lo2YufybDjZbi/cn7jbfjMSOM
1APbGhj0N1ffXkHy9w/FoLTbnD46Mnhh4qZIxouRhXcp+FeGKEizVqodQo5jCZgJf+G/6PIljHrj
C7RtHs7/RfGzIjwz/Ixn0nsb3AFQgrV12/5kH+5te4joALReglmzFPCwkm7guFPVV7l7Wxs+PO8R
WWQlBKzDH4XthM7/2yrU48j+6sFqBsDhCGvR0on/TgnvhpjvIHHBT9wSoVSd4sjzdMs5OsV54rgz
vxszaIysp5Z/k0vWqQXRyfR9n31OgavfHUVCAtl/v4XLpsscAWluFNIgjYu5nfVPQiWrkdv30Jqz
zDHgnr4qKJXqil+9McvI/0TyRFDffFb8IjvkfnRcSntkVgtE2dkem6WljaBfT1lCPwi93iHqKVBf
wkp4e4G4nVqfE4cfmn9VZSFf/YfRIQim0Acy+lRKdaE8mmMdRawdXqHd2s3EMw0HgMwWgWMOoGGd
Bu/idE45Ee/oRp7TQzc7Qsab5d5PAKGHEaXSIj0I7DZmoxvTaOx2Qzbddv44+5UTEQrUtvY7EYBV
9sHrIKDzW/tqjNjeborUyV3xlj1RKsCx17x5cRN+IF4lkzuIMrukKnPejvnNA9UMWDObNTncp2OZ
8Bm0zLv7jWACmiUoaPABgl1Q65HO6tXGLYpAvtzIwQF4Aj38990oxAbVAHOcnN3y7NwW9TONLpuI
WBTKWjGt8ZfSzerGrV1rtjEfeiejLujJeaPQhFrMGVMR8HwI6mZYGgPbeJXfpE3yv5oJsU3jGbr+
8X3gKKAKrzH1g77W78p1JsLd4kbj3F2MOSmXO03kgSl4DRWk7fCIUB3Y66Jb9VQTS8eY4xKQxP/1
oeKT/oWa7j3jBKAtZ1wonTnKpiP2lmWGylbJyIbeDq6/eYhIKrAKeP8MgNY2Yg3/V4Gey99d8XUe
g8rTYNB6iEfkQY4vjV9vbt3iT8SK+/Vh1gfaJ9HjUnB5BRBLt6GMb1k1CBSaI8U12ZDJ4RsOwevu
krEnCHF1acfqCriGJJmYAipAH3uOwr09wSg1sPchI1pZu5F/q9TrBNcZaljoCyTQk4ms/Syrw9Q6
CpnVje4Oe8QoRNRVFzMTFOToyoeyMneF+psFudtyDCphzu6YX3WWC4veLo6Mhs7sVE5eDYLXJz7S
cgr1WDXXP8yo8+gbBOGZT4GuDvveHNhjYqeoTsbZKbMIJebVRZj4csnbDYnXg7cINaGXJcjzHrfT
vb6r3pPtbpvKoASlvbKiuye/8ZG/lOpHXKNUPVfKYCJw8P6EVBjwg/fHxUL3c+CiQ3dtzhK6kTQU
/tGsficv4m/fUKQUOTmg2QI+Ctk7P8i3EIJAsjNsJuhurUWTTRjmli4fDzLkmmT0GViy1/uj0op+
StTihaEBQdaHZJpKdFizBX0k/4gVWDEHTTFiipE9uSrOFNiYY7UXE0X33ukWQdV9TMe6vg7R22mg
WkJsGsi/Ex+13obo9k56ZjqLQd0Ua1oUVyFmztTuZDrb3LDr+2hzByL9eozqDrHNZYy8kCGF/5oH
KWJ+zmYSGLcvukiICODjQYE9WuxM9fNeRbmYJUoaG3n/hH+qtC96qReDt2+4X2VhxcFZyrQLVfXo
VQY+1NTXkvuMQk8NhyYctmYsWxRnVJ+tajfO1n/c0qSZXRserftWYQKWx4ZHXLAaKWzPMw4s7AUH
z0P7UKu3tpyZTuuHNkmkJE5aO2t2ae1rWOg3+XuXECRFYVL4eFXy/H3msMepxRdO6f/O0u64sA7u
jji/+4S4TWzOxTo8PIVAYhSy0/EbFIGIky2D3UqKlgHS8Z5R8VEuDzVBbfxBFBj7qK1F7uZ5pqto
Yxy5J6DKav4mwWsZUlSTNpUkXjaQBy2WAYnDSPr33XvY71MfHQlC6zpitfKPT07fSAOS7TOGqWow
rSbziI/Gq1VXwI0Yr93yThPXQk9LlwchdcnCFHK/ALLsjzkXFwoCgIqzRisbjTrVbCAvCwNfFtc+
FOHlKtQF7c3+eFFR850kyAbYUaMEUmV9HGV02YuvJO0CilWIs/dvODRpZcSuishD1/FiJhN7FsZD
P1jXUzZ+2RUwIueHGyfI2wzgutVMpoP2IuCvGs8sBWU9hufyD6s4FjWwkDZLW+3QLpfrys5UMcZR
Gk0PTLqfMnu6r60XeWacDXYsBbta2EN6pWeMK+FaZajajtbS5fJZw7PCDNADrcTc1FZQYrWvgDWJ
Fo6udh4BBr6tHmrKsbffcS47eGQ/Z4axEHvezqm/rgmfunWwQyEfb01Onp1eEKHDwNQLMPR297qT
pzh032jkAmVJl78n8x6TTBaUG1OsuadmE+wKm2V3QwddVU/nZQhu2sfaY8iS9rEMUw6Vwb59RbMA
tNKgqNpHvjjVr2aC23nRS6SWsFSKqiU70KCbVzqq3XocTSybaeu0NAC4gqb903KG/PYBwylsp9wS
fwKsMGjssOGLyZtzvQZtmQOYmM0wpMZMx2dy6Ab1bn+q515kMOPosCbX1lILb325lXZjZEVB85gY
yppNzoMPIV9uSJ29Wi5K2mrC2utmYDwR1cXSRbdiSVUjem3GASnXM/l27Kw7CPWp5d22hzgQe7bs
CjAz/zFZWuwtjYz3EWr3cRXM/FJXpNJnBV/6+sa61KOwq1z3VF4h8OzT6nhCupl9Gt9jgWsyMRDL
KNv+Sbnqdgg9jZo4cqB006bHy5GJtikqpAYJ+PEJPX8a0VhBbtkRkAjidZMoH4+cXi/Xdz5c5Yrv
wOG2PSJhad8cyzQeySqUnqpH0PrHCRjdnAS6wLJH0xQ+VD8OLE8jxhaSuHn5mgFlsyrIKKk2/kLs
io/c/Rhw8OEwyqX3yp3L5D4OnDX66lBamHK3oJynQF8A94f8UzBSAjl8jMuyeBlLIH0tytQfyxwt
R+Cpvl+roVIuzQrag0vZkLVtUH/8pxoccNxS1uw2qhu6QROR9KoPv0Wp1jItl0PQMpEQ21Tm2+Yz
6qFZ5Oz6Cw1Nfc6azbIJ+Yji4bytVombYYna4Pt7vbMV9KYQvJYqZg42hGzjjU1RHKvPdNcZ3DIz
1BlzXqfMErbTXO12ZpPKl72dan/p2FBbUcOxTVmf/xKNQM2yk19GY7dfhewdoU31xH4GwNVK2DKY
xKIKnM9MEGI/lzWlqJ5UWdnovVtnAWWEydlVHbmVme96nPB+pKM4kBwdxfHe2WUzvEwYN8jwuahl
FJ561HGWQW9f4AOJVVpSMu44+r3mlI8myps7rehCj8E4zcgaWyGrWEqFlzgcyBH9nmUiv5vxSqoU
hJBDdYcOkj/eHVr/TN1re78TGre6ocEhRQ+V2olGpMXxOKxb678OuA5hDBDgXJTMu9yhlJLT33QW
OlxBWLiwpUcxPEW7nWwz9YOv5L6OF2fm5X2e0Qv/qgHVpKsc9bl7ujqgvvO3lLDKwWPlFR0lm+Vu
tEkH4qgBAqWEzZlRateI8U7aUdeJ4xG1/k5QklxonMjmWjE6Oex2dRVa1e8VElBFQZ45KPviG826
KarmWsQP0V6nxOmsK23pir3Pt3Lx+L3fw4rGVgV8FPE36LDu2uxVqHiA9uNjTkMUZ7F/JKHJ5ofR
lfUhoPVKlVIpV4AxnfnUzjCB+ESSrV4QRun1iu+zZ4grotUp2sp4zD4AlRsyjNZX7AsaCIQ4VkFU
pzBu01h/Ekw5v3+acM6K/yqIpDGQm/v42P/oDbExQqgUBsIhuUisHgB1Sk5NdM1X00oEeBdSgrFG
v4bD3QN3McramVN9WqSiPYFTpUo+v7flyN5ZkDRXq0dnxz1G5BtbuDZ03yJff1PcrLdbeUYe7UtS
c1DPjH6N+mFO9F5jDNPvJU0yladMoJDMNGzJNUAyvU47+s8lslMIyGLCViJb24Xo9wQABz9bbssy
MdIic+SU69xJTGGd4LXZMlJTQZCUqu103XKSaemyG/k0r03iRcmTAGJXRSV8z+bv6F3qX1VnMdRe
2Hps2ZT7qO/9iZlmC+SYBcWvP9Xe5V4zyuRuGbhzpdcmFTf6fUJbAaV4VRFiOYhNodiolIQFs6IF
VrHFtkg/vxglmbv2LhazrNOAmYFZ/gaAGiIq3yay93iKuHhzBUisT/e3zlS+iX2HNgFn/i5Dnz9F
DnrsCjct4Wuw7QeSulnzfrQRJW3mb9l/3dTy926Fh1n89zWunAN05uy/bqfskgPqbEgpMQV4EpmQ
Q0KJfJalGTvmQt4o+OQctF65gOLb1RBH5vCc0CmgIDHJkyJVeLX6q+G403FFoMxyFNwKMi7ALmBY
O3Ykbwe/rdra7eEDieDExq8gjCuxyhJeqJnztPyqxZyO+Hh2wDGXnxX6eoJrYPRne+X1VR+UmxGK
M/ZkYYueISx+72y5gyVdoiIIiZGXeP1LmXiSxlhqiwBMy5LXNtVmZY8nE3zB344yTZ1TCnKkL3LO
IeyOHGb2cUQJOmo3fxnhKhSkwhXqhEDgPX3azFJSN0a0Que5UfWtfyKuN40GLHohZ7ShWZyAY1Sp
PLa+Ol/OeCxdxjYRK5rkxDrSdPi7OEiTseKaIsgPe8n4A11rq4qoRcfGPchzn+7ehMGbHUlGKEAH
XgzVH8//tmieazotGYLFcXz67RL4ruzQmuEtZaLMqJ2QOL9pi2wVIJrvlp3XrEsAO68IIxYhr84S
8Y0R6OMppYaEWrLhmR7vMKXlKzO285AKzS1tAhUku86dbCuRan8cOsQ64yhAXaGNc1k0CxybdOTS
owJa8pIvNHjtOTYPQYA5dBC0qs2fSiCK0aFT37bOVGwXWPxkLx4zOCxGSqzBD5MXdeUS/2zshN2H
OcOuWFG20z+2dAxV9Va547an1bI/tTBBwSnChBLyufwFm0zey3cbRapvs13w2U0Rf3JXHQ1kfEyD
lRpSLVATAUyMh1pWIpAOaAWIuePf+Y2EOIcxby8+vuJZGKe0Yd14pHfMfsvdWZIzG6/lQ3cK/5SH
sLrZKnLdEhrvnSDGFY1ORgxMlT1pHObCRJupMroTyh1Nb6REw9TjD79om9mWWzgqVuNTGAr8cyLH
BMuV78jhH8yLmkpoGRgS8yAXZK708x2RZ59PStE9TMnS6GycmjCKwjL72OYukOCA4l/cHtNmoVwL
gqn8qPdexI2QMBJqANqZPmwK7nzr0PmwesGE3ND+yVQnovkgVJqCjdsYfafXhlQIjCtzQ46IqHR1
EtBTVvid7XrukQLPRW+3xVb7ecS0O7Zv3yXlu35ETDoMbB5Zxhb5lXYuJmWZOV+sRqx6tDyuEqDk
DwWn6J0EfoOCWo9zRpOtSF+dVy3benNbPxOBm+6rkRQcaC2y8BZ+E39aqcm8o2qh6QqqAzyGJX/T
LFGj6G1AHPW1w2adA5QPubaDQe+vdBSkwvg9iPfXr1CReT6qHte4GsH+YrUaP5LMshlQpfefZKTa
jxuNkY7VdC0iF6A52r5U4DOOxGpwY34Uelagp7wpkInP3krAos4PBPStGq166h9ZzOFW3ObbsZN8
0DUkG3bAzXN0qkFkERwDMPwjx9uvj+slEGISRMA/wjg7eReVGK/4ZLT1j0CmHqdV6Ef5aD9E1sOz
PJ5POW4SR5I5OFgqDV0qBqTb6n3EABLWAojDHzitOTUsaCFgP8Ve94oKnRCFMBdelxpOC6jDHVUo
xa31DV015+nN1MtVQxKIAixIi0q6Sl+gjMQbGvBT2VlR+vBuyO2sZHgq5no7RPiH+kMfwUoydXF7
RXXYArJi/cJcr1HZBb0+4EWpV4xHqAmz0CrALVXrM4W/95trvaFtURda7XW+86PG/3Rf0lIGGckj
fpr6UI+eZaabb9haPe52eo/S7ZBb2pgsfrDYU8Alh5kSWXJssV/hwsf2viZbwSG8ZSO1FXXmoXIb
UogVnJHihbmejrlWzvHoSdLjcOX9KuaIz+rf28V63oBQaB/KVD+pIaKr4X8X6ONqPOOIKJsVe5AT
9RWo50slrrtt8zpPeqCo4+sjmN9p8Ia2ksLCTr7XZN/eycXyuBoiVQ55oOl04tFdNdOkmO5BF1Qg
eqZH/JdZJ+glTM6vDkfh2U75xiy84w+8vBRDz48k2GK/jXcdss0cDxdk359GcXIISzmoJLMnQOwG
TEn65T3i4eQ6EAf8Ogy52MhYt5dXEkN7I76QUhPCEvUa3fYvz2oyxpO6j1In+56d2EkLNWl+kgBg
mUyDZ0WSqhqBmtNC55OGJiXWpRUdiTXHs54pIMYvp5SjSM+EOpPHFP5KlJumw9F1LZsLE8+IIAuM
HGLBQiubFBBrZ9p96zRAFFC2gBm62xPRvq50qZ2NUToTcrQDbs+HpXSDmUD/2mHkcb7qG0EpW3ew
9+SWmat8tt47ANNmaP3Eq44b6xtuLfcoOjXW+Z6B98ImCLoGGAUNwvQCYM8bdPWxYvtfXyzRDkup
y4RZ2Sh8L+gYCC/wRpvby+bpTpG83MyyAa6FVHM6Srjw+RElOX0aB/LcI6bo02otgr/WEkEN/G/g
7ePaimQskh+FAvQmo7xpt25p0kTFPZOhtlTF3gS8INoUnHIMvAeaQwmZamgNiABKF1Qmjv0gY/k0
t0NZqPUp81mqspc7MzNKpYW+DUi4vJt9U2PkAwIajS/Yh6mIzx5B0hn+1AOkTiKoFF7NPRKEYQe0
HSrAOiToreWcL2h+TFkzGnhYXAKMwqRsAF6xPlhjXJCzRlBCRsbDPf9py5YupnRlDPsrVdkD5PQX
Vx4lN2yMQ3whC/Vdd8XCmDq9ETu6ENi8ibBODkZaqVfPvMqKsPt9Ps8VvcWfWf2yfIY4DzADbx7M
XXdMdqChoMaqDoQP2mZdDZYeXXiAo707Z3SmwmSrZbrF02+vS8bGHyl217B1x5uBk1e5b2PoMBVa
VRAusEkYoYDDcN0gS6y1ttTjdwiz0n+g1//XAx06muVVK78N2Qwn8JBFPv0iaPJR9bm65jJzFL8b
ue0iO/TK2AeFstDH+Rck9D9RJhWXTvDKgLzx8VB1GblOtwMS7eViw2ZRTSMGwxOifzpm+CstL6eu
EP06kr7tqwuLFr5U2UoQm9JBtXuG3f20GQgobGRWs4XCgy9EjiCp7eQZvdhVecf/YCrIiGYwHbhx
iUqOGGM1Zt6HG9OnR7f4Z4JkGqYUfG7XDd/F0ps9g1Tlu6UpZOoYHvD5HbvIZw+CDjyIEhVELa98
MNoomTHJvJq4kWVN/qRXy7AoCZ0t3XULe7ufyZjYhfszKGmDOFZ0vNWYMBisjIXMdHcr5vQx0S20
3PNmIY+UdH9bADFp0nB+5rrsFgrlXsakz0NubfT+8XVb10NZVYMVFsK5BBvY2jmQJgM2PKG3WKgL
yCGC5FfHVP7FtMsmRE6kUSTSy6k9VrUBr0lcplRPpVhifdWTLRTSCKqg6QYzEilo5r7jx8Pbye2Q
B3bitHr8q5pvaHm0OEVBqMKOFQkqGmGw1TOBfmXxNdfnOuvp69udbNa8/NJ0XrYFRy3aqYg6Cylu
eUbi4iwkXfr9XStESzmXi8YBOUu1PTnInsf1e8Q4WbrsT6DCJL/R2i766wtjnEiPvwJMmf3wyGqt
PFd6/b5cXgeNP8VLUcv2UTjkynucwec1NWVDHQeMW9acYaDUQAFzI5rFcQ71snwXY7pajnB02uNZ
EgT6HH6OkroBt/6GFmgCfHFYHyzThDkLJy0bDeTeo9dR7s0wHmXF614BSWdrfCE+u0Qfe32Tq1vL
l5GDtZ0x5uLkwOWpB8mGBUDLKwkC8/O4DrJKvHrw65JzsTjJS6KZi7PJCsrewBGS49a4yw41Tsz2
50SHfALO2h4mpzlJVUpjf8rNO7PvP8nlsFMawoscppiNLTdm4BMqJJvsS3nq4OurjwJ6TVARqKyk
9gY8+ooOc9DPYppJSi3kY0VY+yc+q1dYxv90YhjSSKT/xVvqUN5Gx0Jpck7nANxFZBKL3RT6Hr7L
8zEUmx3T11AXRC21690HZxjUqL1Pc5/L8uXN9ripXPhVaeMnaY+NbvoQ0woTvAUpTBCljGWyFChK
V91/lgFwh1REP5CIzTYfLWdUmsgaVzvd2fcfm6LtxfffF8AdEK8U3uR+IEvV7DojRTD9b9Klnpuw
FWNsGTOkdAtuF2hcQ/Z38vAEWdFh0DViBOfwb/rZN7ghbg7tY/j6jIFUm10ZqfskWwZsbAd9rdpA
BELTGxrE7IWEBxQm31NQtaAKVq9sBqw9ylk+JkfhxUCa0NpGckwFb7GDWgFoOShskDywute2LO/R
UixaNqACfjd19dUIlA1Bv8wxA56/ktAJBdjFGVbN5D0xDan6S0GR1c7SJeUt5lnjqWdPdy3F9U0C
EWg/SstUCOARYH5OI1f4EA+fvwAmkf+uyBbY4cbbp58PmmEslXlBQ7NihxiqLmbiu1R2qdTaguwb
nQt3tF5RRbcDw+fI3x8kx23r66rSpVzcQiAoIqTM/FgHg1DvqJCW4H9teIi2R4b1Pi4UjOwKMvfb
4ntsfUXDFHxOSy2mbVnjjwuGpINaLVL6HHA5BIu06l8/wV3qnZ7Pp/Xv3v6U3dsikirLIrbUwFtf
1vvw5OvouE7+9DKhnvi6g0fTUlbPPERWui1sVKZgZkN7v/SVB+haGQH+6EWEK8dFtWoztevqgauS
jl6JabDq9uilo3nejop9zCm/ELX+IET0yW/ehIBu8Q8DZvRWH/z4rCPAy9ukRsErCcZdQlPPF98E
v1Df8WNGd229GYCTnGg10X7puQbVCMiBgg9CjoSeWHNE1+rgnvENJiW/IVzCkKmYB6pHx4ykGfko
9JlhUDPNZWzBnU36+vnMoQXmTB6M1kaeY/t+ZEZRW+6XS+qF4UDsHh0xNRKLRj+pcnpyTqsKckKx
3iki3+Tof/+jgecSBco7MIJo0qtdh9VYJz443N2dipZe0mEJ9zZuOaVK8zbp/SHgYMK71MYxQxOb
927MUXNM1BDEoFJBqiXn40qisVepNayjfWecZa2DWo2Fqe4+e75KScRb7629xPvRz2MbzIYWfAPO
G/SQ0tyT53guisgiKlgp4XSep/5JE+xqOgq0KuFnbRmr9LwOYEvRjQkLre0qgHOdv7gC9i+lt2to
uPGHZguoGK0xPj6RCIWCScM/ehThHZXsG7D72w44UBz8mn9+eSxlh9twIp1MJEvBo26HG1eEhdTF
yUhny1RLEbUWpNDg+YxeUOyVca420xNgjbDGyLi4Jk4R+t+pYfeKk0hfhCvxDkcUxh4wVWY/mjVe
z0lDMtX84vurkM38eoNCYGtlsdfq43SMgbePeACOFMbG0gCHysHpMvzBcuKYyIcmyKobTNMnYA/y
3HpvmX5nx4OzkVD5NI/jFRYhkqQi2BXwD0MryARJ0T4dNz/SU51v5T/E9mN/UKR4oAC1L34gbbY6
zHC6Vq0jl3FfZa+uifCZaJlHVSEMhQ0I5KN2KGErLNch0AcEy1PgbMFz2VfT4Q8oSbhD2euYuryD
Eb0P+a50YHXlsGuMVeibe22i+NH57UGbfd8fR7pskKSj8LQ2iw82hoBapUQWjt7X5TTD6qdjkxPN
UTF+JlVPodSTRiTyzIgnJHCr+v7PBFrPAoX+p5ROotg0/tcpDSXoD2XNCOw3Co8Lu+ykfhSZXTjX
MKA7TaRzGVd8sDAsu17arOqqsARGkHmcyQK/ekulHsUDNrF7HFq0XBhyfBFpUyT3zu7WpVcxwTdo
mS7CClmy9uueRnTJ5z3VkZbOpbjy+9K8Ua1FhtDr6sd6N7dU4tVhIK5GmJMxhaEd70oetW+g0mQ6
NMk1LT28/YnOQe1D7CyWuZM4YWt8kjA8xUm77Szd18dDL7iTvD4/7Nejx8B6/dv5KxkC03fz6zF9
hnSlIf0WKfEgC7EgyCObV+Vs6ETyWDo6QWfYJBnC2vYEHn+yrO4Ij4S99pInoHvN6wnP7uJc4lGe
s1prp3vPM9F4VeQbV4xwBUhP8qhQXOjj+cDYyaMe0V2QOFy0RGbadBs6rg6tuDiQIzklGPnnIFTJ
2juvDtW9KmzNPtA4sczzP/SNuNb39wi5NS7FXwXRj4gijGOkP7mI1TRAly/77YyOhv/o3L/IfVHA
+l8EjtV/f2szwEOrCllXI6s6g9IHEqwxcGdn6gNtV72/+cZ6X3un1tSSIv773nRDsfcqlt/X5ZXG
6y7yYBlnaKcyYkpBFNBj8dViXTcze5DyX72FFkihRLM9Nosl7NhfY5bA+qDE3DT1WpinILsRqn0Y
30AI1nT7NpR8Jo8gKlajaAMqsKbPmrdDr4v3DVNfH+BqjGJKDi32SUR1gZN6d5AoSdfRW8mmK3Rm
VoIxGnzUdgbbA4LtpB+iUSlVc0GI13oZU+/xvFKDiq1/74E74Q4xUswEPu3WxMV7WY3etZczQvVq
0V0UaWPLzYy5+QnSZEnqNXVZPh38DGS/IfTZFpsAZ/Q095w5vIRjsSSdD6gV3UhuU1KlgoT74sL9
U6kLrqD6Ma7ymluUDtlSFqFB+oqrHq32lLhIOHqlkRmy84I9sXP0lBzqeoOIEoX9AIhL/+QuUUmy
o9x46bGER9BADOcpoOQWuqMvK+2KDmqa6K34HiVMI0ApVH6nLnXuLDFJKZ3UVQlBgYLdXnQLE+Xc
X4LkZ0TgYt5gLdS/gKmArpYC+Ntc4oKGZmRNr/UtuBHndeLh+BI8lceucgBaKVvceTYrn9g17l39
sec8nPGIfOjlNLMGrvW3VHMGDXeRE8kGIO8Cxcyka5kNcxaaIP/b8redNzJgm8upzr7IEd6n3/EV
K6blip68hubJi77DTIqHgurM2c+AWfLkCujnmjSmjOJYJdEECc08vUnqasvheML54bWK4bnMKFNW
zLYb3KjwGgmDxLQ8L+aEU7H3MUJhGOHqdFPl/v5T1+KRa0Q9blY1R3q5OQDtfiXZjDnuRSNqt3B+
oYLlZ8SflGHxUnjsfdDy5NfmLsAUycLVqe9SPX0T2YVwD3LMR/g5IZ0/1N/XcwUSVDqPKPDrIONQ
M3UBG9vfmThAQP/yFWgHau0y4+/q9kILsW+TSian2KpXCREn7WFOCz+Mff/N+oGiDvOTNWOXTOEk
MPrLuWc4QWZwwSgvAynSU5d506ZHPoW5vQ1drjW+MkzPGuG2pko2q71BwT0Qj1TQgX9F8XE1/lHG
975SkVMyiJ7oINeqF33u9yS5hXqgqHpCigEpK+SNipUaLuVf1r7VXcayJhlJy/D0XWYys90ekMaA
LeAkPz08x48+YqG264L3v1B+o15Z1kgps6J/ehVGw3qADMqfpUa/5/ePAToRfTvabdFLZdvVI9Di
pKKPuJx+ATD176spJhJP4YLQaTdq5z+zt2DUr2XuYAof7ya/B64dw5gKh8jFniFJ0sdMjwkN1mA8
RrOtBXUX+jc0ptxi/YOz6YTuVlOE4Sz27SIeZGkevOhWtvYw8pHZt4whhRymQdKo6EpiWPZTFiGl
x/s5DYqfnQ1k2Zw53MjW8gD/s9w1wNmUE1spzMyuzceGH2zIhEYdL1Zeop9jJh3Ft6fCYcAGu5kv
oIMO4rYIXYpohVFnw9DLfF05WDq3wND9U6ZMOm6cJP9bJ3KvgEQKK6KQt4TeactWbngHsXXqxQeJ
gx0OMH9mmxsC694KzZgDkesE68WgzMGxL+bVq40QLqOIXDSis9mzD9LDZTbWQ21KrHOBXdkorgeZ
KMDLkv7Q3sxHuqq02DpehT4Ka6Vy39EIdN/Y+fmDWViyBMsC50jEYKEqNt34ml+zSF9JwP80xe7m
p1NA3Z5Zb3iIl+Nk5/jz0H2IRlPJK67a2s9KYvH8fJ+R4QUAFHSyCul/l6aMb1FHPELCpzDiLtG6
dALUu+u3l1cFvJv6RA4G9qKqHx5S8wEWHnUGguPhrtrTLwenmKAyDQuouXkshqLKQfFAgzluRhpY
5Uj/aA7ERJsIdU2Xb4IQM2mhZNxLhXI7eP6URAMxmaV0uoah+lJuWFYWGht6Zb1x55VyjCdJomyl
13PqVhqjfPckn1ZGXUumLTxYFH+yh+KUVLfOASUhaGz9DhR2shjoaalclIG7x53wpR0f8joE++xr
Y8sEyKp3gGErFhMuS5EhjoZ71MZhwmTR4AiKdBhlMp+GajY1HdBWI70eb53ZAXIa+0r6kpdw8XKe
GzeLVGEZGeIqXQXUH7OmQNTfiIdPyZ98GCsHHnChlJRayNj9Cup/NZrcs8quWVgYKq9pT5YOnOeP
NWlu6mVPIMT0xEV+zVRET2E8wnbWK9nHdd+Ho/ubRTBOaR2JLWYcvB5rhYzY0r4JVa5k5q9/3Acw
t0ZGxMCzmJDu/0I3p7gVsjanur5GnJKpVVdsCHevt0wXOiBFckszX97E74tnkpKm9xqX7ZC1bhfv
4afUQ3ekgBO1aywyVl504Z/d5l6YuRliGXFBwWNJ+g16YPU/MiNAKxENETE27j0G2YOJkyvDUx8B
MU6RDxzCX9o93lo/yWDqKcRRMrUKYLmB0m1P8e2qkgCtNmSrhgXi2nyd+RX89kw2Q8mq62rN6Bdx
hrxTMWfaHirC/nsVvvuiPKQKR2HCqQM2+Dkr6zme76elBi9FZvcDRqBEJCBKpdGl0wfa1oEG2jYL
INlqluJwgOHJJKMfQR8DfXh8ZT28oMrSFvkAHo8pkQxDMrGhzJFfWGwSBbxd0pd/RaIrneqhNrX3
falZvBqMhQPag4XG824DiX3YIzqVT/G7UN5Wtazx80v8RhR/8LqrD2YjK4DvxYPvIw/6x6uFFo3S
XQH8PIp+4vmMlTjwL3BCDt1nlX/bKschvCWhZD5zHouRUwKG6U3bSK+FtMyXu63/LMtfgNi0DicQ
RNAdEQh8HIkrDRHMQz7fxu99UAYy7uHHrvu5EbC0RtMApHi0ZnmI0p4f6mbwymbKLt2VQAPWaptq
zzKnufOHmS/WgJ2BG125mwtwsJqPifUG8Db3hdRsClPsj/U5zhy1G6QVYul+8ah/kiJyBda0P6lP
IjHxShEfu5m73HmOmyUXzYaTNZrzejx6Jt6wA2xexDQLNoiHXBr4eVmQ/jVLFBI/zP35btS9hwpF
oOLsrELrJT2BfCAOK/4kDQl5YVxAeOE+73mqb94DR30fWHvK3J4FACFS42dieDvkBqzMHO2dl/K+
lpcVY4mZSL1lTNArFA1jJYEVtS/a2x63JQtszjjhehCnmCZDuWVlc+AdjjMtCWyBmrx0+TR+EbSh
FQ+8yMaly2Agbf9yU8ckA/M8jXIRJT0/T1Ys57HmL/DPDVnCvPtP4aLzXCZUiuoEy6F3H2yIHt2x
kTglhb3J94I+DD1/tldmk8KW9XJTCZ7v6x0HCBKBaswDW7p52TZODMV835YHblqP0up1syteJymI
nj4mtRY+z1Btb9zFDeZB+7FBclvPnufTzFjSpmKKeT/MIpo9GGz/2hzbTtqGfGatIsMiNq8kRypM
axDiv38tgfoOC+1QxshKsLyt96fnGA5Nw60zuIlNaHkDIjFmYaTJCIbmqtuoPb2WuU3XlWY0XzRS
JFjBYlDhHhxblabUp0v0R6EclKsLhtenb5VhM1sdWTBh9/+vpomxQpHw/aIaXgSmmlHo1W/ehYUj
tSQpcgSLkzCl/T46RpGFE17jdT+byw/cEf6TPAQHsoJecttUar2JW2XIJA9ARO6esTJCRUCFWotu
1aTEXtl/+rRbuhIrBkHimNYrW79oHSE3olaYJ0t7oQ3tisDSyDZEjHvHZeInqr7ZooihpONLxS7W
4Sc53pb780+IGceKkxAaS0iAd8ABoljUegwYpxx05ZTDtouA7UqchnXy4BxY6nFLIAjag4GeOgGy
Ah1ZXuD7NOI8AOEclq97U9t5KXn3Y4+Hkb2qmI9gDdK4Llg/xPK1ZZlV9mGNUPUVi4gQL7ug3ZoQ
/b9JGfdyoX+nCYy9M4BNoWFupaq1RQGIJ8ecLD2nCsfNBBnLvqWWFksP2Z0qNm9zkTGtZdJMthkg
J7EobRqMNQtd5cYxVgtQNnNQ8AYEApX0I0DtrIbDWE6zu826VblPwUUrjkcq1FIeY9dZMQk9V2PD
uYn9LGI5bDdcz3FX7tOVHuN8rnQbDBbdbwaewxAJVYOfYkEokH5hJtPVCKz1kb9CpKZU65ucYFha
/hchEPV8xmcX22Ig3BzpSknWqDLUr9HVpSTYw0G27I2tyHPMQsKkxjd3fMDK5VFOF8K66GzuPfNf
UL0dFoLNThYyUSif2SQIusqaoTx3bpJkJ1NriAMLBQKZ2hTjiNxnk7ZChOmuitngljBLG/I48zLC
/zVdMzzhx0jlkPUw11yqipqmD9SlX0CprMqSHq+SU3qgOzE0FtyyXeEzlm/WlmK8+6W+DNUggYqc
mbJ6EQzBG4k5iVIXgHGEDX1UXt8TD9A+pBsE36mqV6KywMdk1T5hMgfxJmrhHltLFYlqnK75f2LM
3Lj6OFP+k2rbPJnJH+7ikMZN/IsdGOisNNMaCq5M9VjbcrBgE7f7btslzVpCbbNsCuCMXkK3ezH2
vB6SunXJDWFQ7zgtrgaFsnUrtwOspWdZ9g/DqJYbeoBZe+LxAp/MFigfMqsOFCjMY94PRU9jS1Pr
4qRelFrUTOu/xg90kaIvvLewCjVImAuropOiDwlh9J5kGK2Sh5f7QGZ4OkCtebHMM8T8+hxJlxgh
5oAn0G6NYdIYWpLEw6V1Nw0miK+gBDjaKNKqF0e9wQIeULRy+N6nVMfRewqR2u9QvWzon7e8B9uG
dIxLKj8Ee47E6RAw1v8BnboIunVLA3O7ghXoFThc2c9tggJELc6jqRnBuUALnfqLLF2kUMs+iY+6
eMJhZOdfNsFjDjH0dmcwrv3lsL/VXWCoRlbt09iBNLxBt+OWgSJ2dwosbGqAQGFOi5VEvYsI8mVw
vqVGcZQAemw1JKPSxj/GfbfGilaReTcRDVWqE9BxB3jQ2pOX1cvnFfALxsELlI3en9A1t7XiRp93
U7Gdcy37qpINgFqb4iDAs5iQqQkxsx0qZAYydArMrBMVwqivEMy6/TEbHhF67BR4mzcGx0bkSdXg
Tv1V6rFu47QVVtwl8s8PtDSz95gqXhXavqO+Fwb9DEu58inmI4iUf5T9s6y2QmXzALzHr6yGkPTT
IgZ04cd3ywIQ3u+Hf+qw1EDcJ0pZC43wHo+lXK3spgoRvHmR7LMu99pE4f40NOHkiX+hUPnHIFMR
IM+tyGhEcimYvMYJhCjldUJ/g4Ff7a1WGLULZqRNg2XF1mBhuYC/Dk8w6aUZTbO/hT/e6VBVnthN
jGCdC/B2mzRjp4Mv0nBsf0MoTQuOlSWkS7xVjnfZ/Q4mKzUIV70Y60wjoN1rQt75/9PpanR2OOTW
xo9dD+keAMn3VmSx1m0fcwX40ZPvh8oaLEhuCgjYVaOm1eME/DX57tfpbYaXB49lvfbsZqlinoFg
O0fBlQMfxTDFdGDKj0JBP6XheNQBuTI59qprkVZROe+hUb2CF6SGypk0+f5svFLDqdxSZB67v/gc
o3rTfGijrW4obLNxfV4gdMvSNJrt2fpq3VSBBbU4RahQN24BXSzV7c0kODoa+bgl6E8VIFardwVn
miqdkz+53Rtk94Jx+liAJeFRwEP90+4UXq+D+timP4CRKjOxACEvybFcZZF4pR/1wOXPSD0rlqLM
Koi9Wokj3W+MSii73d2/BYCw2fNbb1/+JYp6dBc1GDi+5cDpnFERgGC8vByhJuaGls7TDvVyi7kL
WiOjh+JOERbTa++OXRiWGFUGFimoQGtXBTvn9wKC1aRmjWvVFhl11gb7KVNclFSPV0XU9ZhNeySB
aD3yDNudcqR/vz04o97+7aFKFq4SErBrNa9vTlL7noj9Rg8yOXDy01RXbefnqqQIkiQhgPIB6yn9
7bFes1A+bG9KtaGi1ImKZqCtNuGAL8w3l5szUGWmeDPgxleIME9dPKzSPDiugghf2ildQaqPgoX4
I4iOGQKVszR33ba01l+fFeS71XcBqWqgweSRrGuX69QRYDhnZSjRvpNg27YeHTrXrEX8+wpGus2B
e1nr85WIQk2DICkpcQc0MM54cAI1dLIibMDtvB78CSkTm29CJn8HThUP5FFDEpTh+3v36kMBIit7
XmPtSsiG0k+ibSSTTW0noN5AqQEwpJagXaIohc+kL9fcr3gPbfX4dglg2FlHI8VVJdXhluQis9Uv
aEKAQvpifBGVFBg/ge7xHWwVvV5IlplCNSJdgal856kEiratCYm4HNZJUbWlJEebD11WhQYBGnPF
liwSVi8dWBs6RCB1nDu3myx9mEXWIAenb7nYouyWx/TaDD36K+GuLFIsf4agthO9KLQhTGsQ9esX
4/2goCLhhhPU/sKj5hPMVzuyby+M4fhRSxhD09VexxC+I5HaJ1Kxm1sZc89Y0b3Xzpa4RZUTHfrR
WKxX4jL9uZSBbnSFB2oEfkytN9ABFSGevhTXsIafWRaNSWHXk8XkuzWC0rINIA9XzLrVW+5iH/W3
LEIDh4f5G2qACsOFNM3KuVqUjBxgIDt2zQz0iSTdTYdETqF6MxWUSsRzeX1mO5esQk18tzDeWSNj
3M7gooITU6XUUsbqN/vRy4QG8dRiSus4p4/kGoiH8DMnHgfnoNwiyisxkNR8Dp6Hrg/asJcubtoE
gBsfPrXi5BUxP5mmYHmP2aBZsdEPzrV+Xxq/cPGg7OsZndhNQRH8M6u091r3xHszOH83lFi4PV0b
wYn1trbCSakjhdjJZzw6BP6mRorXB7VfroHMeXDGp35rLNyyB+JoGkMKcB9w8SL0e6/Uo9ZKpAXf
4vcCJCScAe6IkBzovkW14nNhFolmJ9T+5DeCy5Jh+qfSTPUdIySigByzoQOEm2c7ehBEVfXWKMZm
WxUWGDFBqw9wb0l+SKFKd2amrQgNu3vFB8kRZcfczSYbZ158P480Zn0nQTP3HpKnN2geb91F8+71
scvGHZVpdJm9rUJqOwy03CKMztUORlEuTKw64e2B2tKCWF/gk2PpQpyGKiVUQBVwxo/v/Edzmudo
1HfZkT34wq1Vtc5tl0q983KUfv6HH9tz8PZUdAWqa18Mg3KVfW3La0l6r2Nv5TbYcG2+oHFa5rYZ
Xp/FLwux/XK8mCY2vlmU0ZbEiI8/Dt3pHsfCQWl+MQnanCRxQY/4J9xDU7nNtWwnFzIDZJjPPGnp
kTpEVeICb/kgtdaLrbxUwCeqjQQEGFqZZZttPJRQm4JQzxw3OT4xGZ7FwLIooFKQN/Kv2fBFBI31
kTEigvWm9+MQdH5sOpHjkCWcFiJ3bYP2p3LIzVQYb6wVqQ6JYZD3FZADWlq784Z7pAXmmqonY0E+
d0qAM9it2ujAkRp99ONKS9BHuTh6wymaQnUIhYaPSpbsxxfdIYLNJ07jo2+iCOcppplKr2U+MZQz
ZHg39MN1DI6uPtV+5d1LVK4ZOSwmvfH+69rYd7UieUuu0OKV9g/QMO1VmDjrz/ltrewgXf6naxjE
029LfAeidcmMv2OL86oPjNkONgeyJ0AS47m9BeM6Mkjw02eKNz2WCHMbq3DjTtsR9ESS8+G6sQTo
/n6z2PngGB1SaZIxOjM/4gH9CmiY+YKcRdzJ10r9HhkR3uw+k+UJ/23FyCRpQMGCX1JQYaU2CiNa
I/AjA6EHcy1HI5FRol7IuO+X8UiYiFk2qkkDtst05wreTDWlhbUx/D4/VDT8+mtZTbAgEFW4CAsZ
Mvi+n75+XpCWQmHkXpzEnWX9NlivY6Xrthtu7pz6P3Z2lnlNWgI2+nAUVKHAjnauvSrMLTZT5Nfs
BrbA9Sr0xeChO4TpJV7nr8reGNbe7NaRjFA7pZ5czm+ORlE8zthLRCyYP9ML9BItQSrtOv7+b8Vt
TFlD9JzL0c4s39WRsdzkYcfJGNOYDhzoynIJlpbpSgBz6YZ0aVT9VM85y0sXa3iisVFulKFkqyQA
8x92K73iPRexKFUT/wSfec/r1hC+VAM8Kixo5FYne7YXzRPFcFlchJCgQHyjxJsmtD0AKQ0OcQAB
tkg7jc8gv9Swph71vi8zY4CAQWqzwseJJM7PjFQbzBcDLdXDyxOByKDWXoGACKHEt8NYGthVH/Vf
2owxtR6gjSVF1yH2FIe2wnGA+zy1QFmHdVWpHMT2WAnJtJ91xrIa0THBUxZk4Jh+Emt+GJ01D6tE
1V9YyFZIVGFwmOCkEAMt/qdFxwcMY6d3dwT4PWl3YCrbHiuMLoTLuHWU8ktugwRL+H0Hji/DibzR
DnM5Twnac33LCcCakQw8w17sN6fc0DPkSnY2AuNON+E2E9lw7erQFKbDicQzNKCtkfd/J2MfFJKH
FMlKXWmCIReQUy9hSyYTiav0TocG6Cfp+l1LaMryJbPRIthApvOenNU+ZbBEqpTOxJrPzPARRqlE
xaBo8ukRAGP9iw7Egk+9OZEKIA7sZOpKNS7biq+kfQfvSZxitrVo2XHBVCQirevzcQgJg+oN1sZz
5Ty5hsYx7Ir4px8HaDYSk77eP0COe2u2naw0vhkOlYZppo9kCe0P+ivJg2ud/wsByVjv6q55ank+
oix1r1rjysePcZR350BsX6/K6enHx8akHdV+zdhBAQeQxM9dYNao8J4exWy3U7Gu8vy16fTeOmP3
ZVBUtYK/DHhu+ZILhSGGJ4MEyHpvwazSosXS+b9Ehs3+UJFY/k88g7JSab+NzCmmlxuxLtTL0HOd
uhnXA+ezw8PkTrspA2QayG5Z+wxcGaUZ16ihzOKoyAhcZkBLqWlvbuqJdd8z/qviktYJpPDm+5r1
NBj1CZ5SmM2r1rUIoG1KGFZiDHpTI/CRUpksl0V9AR3qBnb+me+MC6EOnWuH43dolCJ2aBxv8Rv6
naqDo9hoUrVCXSoiDbjmUgO3lf8toHhVpMjz+2e9rS3N0AEukYoVJqRhlt5svSSfcFnzU5E07ort
uT/dyCZ2rEQqo744+/bTjlS3gGgvM21nn4DNHdU6LPw2C4BMb7ti9lY2whN3qcy/i+43/mJLRgnm
nLwKtO5l5CIC5/tdVNdMaWtwkemdcjs7lOb46xxxzic7fQzx1dGJiTfhUQEXP7eEjQAN7kZwCmg1
VaLeaF8WNGN5DBG9ZatNI6kAo6f/hrHtL4UamSwiRqaDOLoGoP+RQVurHHt+h2zXK8H2m2IaTVpi
Qpd3vFRqInQM8+9i6z8BvlxNB28Om77EVeh2v2nphNxoCbwIWXMmpqxKjr2usB34sz8tPkkIS8J8
HmrjtRZcj5jtCvd30cmDwwU4k+G/ZETNsUHbDM4NJbecBidRO/RFVWAvsSRWeuIXtjXj56SfmVP4
6GMiGrtijaIreAgwbWrZaX8S2+1TgukhdTvFOEhYwf/g9KnsFt1zx9Zg6/5CTR5bext+McDsXPaR
eiNkqd+b8sOqAbD1/9oUdeCKvoA8hhh5FNLZc6P5WzTyYdEfjhsqlOdIk7/iaSjg4o/MvsDT+PPy
vNFErMnwgHix5hHfwjKKwyiykwne5BWJmBhpyVlpQYZPGy500edmrhqeq8qNNVbvCE7leCEbqwn4
lA72eB7ykdj6oX/TQJ1G156CqmjfUYC1wveqb7OXHpXqRFBp+ZMiZMbeu3H4Y3zHC0qpPKSCowWw
dUyaqOsDm2zFAx/mDMDuiaZvQzpvHm89VnKnzl5jI6O9OBQsOHnt5Ok2iZZwin6nc4LVQ/1DhUhq
/cb1I+PJE1PZhe2uDP7aoCI0ZqENYBPFZAfgw6eOtMTU/NULRXVnDvdbhEl8iRUVBJU3OcPg2Nul
XBTLmS+BKYoSOqwnmzeiQXSnOGz3oOa8PzAy+JkfwU0cB2plyhQ8WfdOp7wOfGrNGPhFzncnnZwR
OF6Nt64bX6R1e/P4BT33n7vHPCt5lpB3KitMKup6okcvEhO+2A1b3hdaly7ePuFy18iU4OrbXIQC
iEopKlJOSKrJCqXOzyVrkI0rBohTYN/Bk2ISJdgt56kBdgf0gJU0Qa05CiroSvBF0XhUIw/QtZ1b
PdIrlLpc1cdnEFDLyTAb+zsdQnZxYGuztK1GeThG23+cfzi0zS6fdCvFqT6WtzWhEd8+ig5Axglr
2sot2jcbF42wwn/wk0RR8VrjsjNgf4t28YX+Yky6gzLbB2HEsneNJpcebi8E2ArkOIkp6rfOhfMF
+tDdFOcuGIh4YX+P0CwByDxFEzqyEwMx6GkCmQ8MgLhVIvDODeNmgxVpkYVelqlfmvDtChE3C3sB
hqryir0qL5YOPQftOCcrHWPPhjS+08PffrHPo6ipgUL7qGKoRjxlGXEOX7BKhrW8GcK6UeYPulZn
ijsngst2kttG5bTJhlbN6zPpTy+XtuYD1y//8Tix1jUEZMx59WK14F62oDMLugVyrBh9CoOp7fzC
f+T1KrmqCREM3UeDJWVFh8iljJKwcdzvKIvylKG0jO/75D5+p31w4i0zfs97a7vChWcqpT7ZuKtq
Oydanhnzq5+YKzuw/s0NDZ5yuKh/NVm0HLBwwJrsObsGWwRVdbOMHo+J6kcAFeW0OlqeVyajlOHa
tZ+TSxEsmwucuFAcmMQb94ZJFFKxOsSZfQ37dVck5sEMAuQuMhSRpsorGQ6Ml94eEuaqFRwzN71P
AEoArgd8gLn6OFrvtRXMP1N1gHwQRnq8HWLBjWvhQAZLYGZ5m2byhj6OsRBXx4yyRI6QhMisrrj3
Q1ZAbN7H0cB5U/uU0Aro1syaVO92f53Ffu1fQ/gIPC3kXXRW9U8neN33AnJiCaoDxcN9iHVLkK8+
f3s9TXcRfR8nL7yFAgvzjCkokPl8KnwIIriQVvuVzttMwSD4M1+zm4iBSTGaUbN8WxpcUwOPKqxR
Xv1IZQyl/mOXOhimejzOHSMe3ux71XzUbiVwKy7B0UXyKCbADCnXiAcVlJcgYJqBDv4mLMOzjON5
9BoEGokel1eXERgZJYm+qz82CiTPqH+cHGArFy0ztUTbm8zhTXqLrOJKvpSRIX21kI54gyDo+UJh
4+0uFKH9vcwyz3PGMLdUrCM/NIyWRcvHV6bKF+gqJZ8YlxvPIf12ISikK47ieSld7dHOPrMeCWbD
ofBqAp828D4R3L40XdzQ28ZGbLvnQ3vwiKBz7bEtmAEvlLPAyzPbLDk5L5FJ0PuXxTIHuLy7x9jK
J6RsfAIm+NBGot30YWuNqx8Yv9mBYw4fE2G7/l5kMgFoXjHQud+FwOiTxHLVe2XSL5MNLFZFW1mc
qUa7t2Kqxe0ZnodhXVibrrEW6j+7/oTwxOQ4eswCpHEaSYowGg4w1qLOWbwuwq8CEdmFWWHCAJux
t5al5PBc9N0xrG4uJukzj5ZXIwNAEc6OorJ3BbcdGQBcp24xGt4Joq2m3XifiT5vePBMUMoQ6NXo
T9fHa32S8Me261WtkIlbJ0WoiLC0pduQlVt56/isgCED7Bl0zBrn186tYiHEYaiYhg7URGZDHMs4
PF8UgZ3cqVRrMcgIuXAKp0D19KRZWUyYQeNyWu+gwBrm4wxpm5+/mhtVzoXsDR3vaFeUjOfCMLea
IHjW48bN+MjuVNca3JO83LVqYEp6zNjcFlqQUBaNRTUIqsjDYFTxXr7KbAUFej/mdN72OEybvbx2
vFQhGptmdHb0iToA0Z1+Yf7HIN+Bt7qEA9NIjOhe65PkKipZQ7P1JXWsJZwzdNRxaw6PMYYS2iR1
QVYNxXV3adQa4MCtmouDWGRzJcYu3W/F4/5Rr0oW6LlXDjZsHFtas/MgBpcm4Kj0O0OJ9yNtVqhn
7FmGej4G1kIc5RfEIx7i97ioaWmYX8sDiEEpPQVnACv0Y7ssuyGoqhcIUyjA5Rex0sCZs1wDxUpm
YoMP7kQVZ/BWM6CNlOkJYQExdmTPtIdRLJE4BMbThHMLW4C8ur6qkh5zRHqddAL+5fGPsbRQZLsP
FVDbPhrpDjnd7UN0W4Rb7Z5c/1cBx1VQBHxiUuIhk6x6hRYBy+u+ZvyZ9GJnyjmn1duY/+xSKOAd
RrrzjPyAwYOAZhXbhYHu4TYTmdjgWBcSXGBOjV4VzuIPuqeuSJUITmWUdh9V/wIQdAApljnpVpX8
c871H0oRUr5rVqtKs+kOnFFJIgPSkZUez3ItLUFPn7esQnxmrcJqHmT5ql/9N7OOhwGrItI1L2i6
+YoFAikEyiBgqxPuW/eshmtOW1DlHFvCibiKKhjPl7JOByb8OqJkhZfSkUd1tDmRMUn9Gk7LUKe0
PNoa6qRVh6xFZf+WJ7mvtgD2LqFEnSJWjeZ3Qlqk5bY4r+0twy3lgJghD3UcnoAJ1IGmPUfxkU8F
PN1z1f6doLK+U8ZSzfqNleiLmJfj1eVqdNnsFYK1xLliH0Ih3IFascy4525PK9B7dSbqDqXXYN7Q
yQcQcdTdgJWA6pMQzQ+xcBYze+zu5uWdamB1OnnBWxswy7Ij2jeUQq5GOzeCKKiostmQeg4Jw+Pf
+zZ1XZw1iCQWhW+vLaVRNjPzBsK/iY/CxnWqCUjFQa+B8+b/9kpvv/y0TuhagGTgIRltqh4uHzG6
icOnQoVzFiQR0tjmCm8FfDnAFXNxPUbH3FjbLaKkzvxe9zAYQI7oRf/auoc8YOEvYQ67U3kgFda1
dJEHj1rzwgHXgwwwSyX8CCN3BmPyI+O9uhT7FhGICIVk7ZGUEGhWvg0yMbHanBOOaER/MGbSiOkF
MHIer/u+Q5j495jmJZyGui5UDHcUZtoig5bOsb7wYjF75AGWbrpupcYp9DA8V9W088Nua+wcbsFb
8LcqGeKbIaJrq74gJ13TkZGAoLoDyhZ6m8waV1Xy3g/EBfZKDWqxGKA8BNZq+G4fSf03yJlmigdA
18OY3ofef+OT4oDi1OfhzkmxTjYcOa4+zW5gJGALJjQX5mzPQP+7b95n8lz41lPDGvVXbHyNRJ+U
pEa9XETH57ia5YeJwA0iwCDJhU2IqxLagQ0KbhBCWpqOXUBoI9L8O2wTrQKFCTs/NKLKE9i2TxEP
/CBy03Nx274/Foir/RDkeibOaeTQKck4q+nDx8gOrMCJfg/oZFVmmZaaEKkD4rn6DPmnDNIDY2BS
HA/3RmyQoI8FtwSzwtnld8SJ7UiUd4/wHkjorPNfx6NRankOtEqhKuebw1c42w/YXF6B3KcTy74M
C/HA7/9zvLBTzwl74ZUSgTnt015z94bU3RCtnSVbmBBLEiUV72snyLKV3zn9pjDArRePP/j2Z+55
EyXVAcwraLkqTWWvzKnevBQHTn7RBrFx28n67XmSIs11ljX7l5KpxiOXZ15IE+JnDdgDM/6nkus1
NCMdLLHtAx8+qu3uIgETDODrbifOJm0WxPxp+sAE4PpCBIpH3cRyc1VbVLvb6qhFRTcrFvg1pEln
VZBGWgiTJdTaY7RrIItS5K5gfG3z7VL93AMfx3r6TDbCn3Fw0Y+sBXXg5FLEKWSjz3KGbSOF9rwp
30MXrwxG5/6bUgSy+FhJWoH6moo+RM/A8FMvHHnI4sQZgZISCmPRtj1o7JrcVWUiv3eFZxcGDLEv
fe11R4gacsiVFSoR8p1MDtKe2dbyX2UkPQv36feiFI3VFbCmP46WPnsoHIl8QSifP1Dq1BeCdCa2
vXf09oL74X4Zz53M5hfV77kVGz8SdwtLmvhK8RNbjF8IvPRviVgkU0SoquA+3qFsyPfWXZ8e2x44
o8rFLwp654YrdqkNsU1hlyNeGbFAdlJbfp6EBXfzKBmjNX7ubAt2Hyhl78YkVNfoOAHO13D6rXv3
ctpSAiT2osGjtQGjdQpGv6SIfa57n/uCdHiWRbmyzVlloo3tf8/bS9sw1x0qzCA0kNA4y06ZUtZ0
fn/iJEnzrfnPEuNaXfBiOvktVoRIYBOTGp2AhJqQtEJhON0HODSmpfWdIBzseCRvA3uwNkTNqGBv
duhO0zO9ElZQ3hsKZlqsgzcyJ+175kLHuUFx06l9tNSkj8QNirXBmyutgPo9/24Nn2bX447ZZX0f
QZzgj9rtGGWCKcW8XgUT+gDew8Kn+wqSLCrlZeggtuOHjAjoQlSnRvgB3OgK0QDAyGfcIW2dnIS3
L+Hzqe7c60vae64mASfqn3pIwuqWsTnCsC9zLcM8spkonQcYz4Tp5UXbzZ95TK3h7DWnpe4No17J
GnuoHGw89CY88ccOkAainJqOOb9cMHXr9WpRCbP1lcIInuBWjH3wfYK/tE3ZSUWJgklri3uQCyA0
qfy7Xj65PVK8DJ0Q4qagqZ90ZlY5Gr1AxDktsJmIb+iPNXrCTE4PlmfjRIPwTMZrcvoR7Vfu61HF
pb2kTBWgiASpbYXecs5O4GsPMwFTfbpOB7wE1ZJ5MYzCLTh1YfTylyioeBs1lWEaih6JzhYRTwQI
BTxiF0hB1qyQIM9SuqaWzwiz9Xy0elq7/qg7nK3BBMr2yvTblrtxMftxhC1bLsDB9++BZYf8962H
/J7rGWgMy8R+6NYgrmNem5rMe5oBdgKVQc8d4YMqw3DzEtYWO9pX8BjlIvtqiY9bDatKfJMqxj9a
mXAM5TV3IsRlHPnPPUifQOoizIFc8BJrlyqyVvMLrSTWh2W/J5E8r7vb8+FYvVEy0krcoOPFUIzQ
153JmyLLIzfDgHiPxHI00jeVTVZ6A9DDE4LhsP9rZLyzBpVDqWOt4msWP3azfn4SQL69yQWQ+NrN
UN28fyZWltvAj5VaqggNtk6TyKwdvdHBQl5iQqEEa5iPybCsgyQi+4yFLWbradmoe/yJ5Jt084ln
Ub4FVwd2BNBNwrnwiB2809eOJG8Cd6chvPOJEiZxmSfYc4CHOvYKjvWBMswNwlQ9yLk1P8n8xaxa
vBMnqV7BhsF2Vef4AJnagLhEfZu8laHFyXliF99JVrIdTLU3OZJYFYDXgcUP2Bm1UP60XwahNQ3U
bDyMWXhHv3T2YG+FmkMXvDPmuWM6IRDeEYzraVtxvkPYttKtVWiRjUVBg6A8mVlZ9OQ3/aof8u4I
8ZcVdigh9wr8c7oYJudyud9htwKEwfu6qM/lxQbhcuMK0WYdkY7zX392FX4n84l1LpIqOnjQ8N25
aHeyPCvHeIyDBsyNcawO/Y13ySSwAIFq3kezVjblpGgPUJOMSWROZHg9TTbXYZk09C8E/fHVfaju
wRRwBTo2SHNZYhcp/XzV5wPCji2PZc2wL58vXn77I7HAom+fPZZet+QJTI0BCCBX+CxZ4cpDICSf
5kwHlJ5+BIp5cMHKWuuFovrb6E7vHUq0UPnQs4Qt8Zyw0XlCwWExhOqiev9QpO0QDIqusLAUhIyD
TOSdch7Bnw0lOZB9E+2XTLOroBuZo/31KfeAbjRyzkbSH8A9frvAKMvIeScm7VM3tVJEMdW1ufuk
ouZExsm4FqENCY+OXmla0QAmEmAr2DZ/5pGFsRdqc1dJqfsFPPYW/ioZdzsjk0n+z6RmmLEwqphj
AONP5pkLDAltxE5Ypw+GX3W3rZTWpCVHjtPqOHWsMQylkHF5TFUn++QnzlGGfhWtmYN9jxEoNCTh
BKScmJ8L0BlJpItC2fOKMpW8f/xvc5nfA5Ho8b0cElUORKTJDwTEjooThJMs3ey5ogB95jPsZPGP
2h7mZjIC1ySMAggjd1fihIFO/tqghgNoL/+x0KUyOqS6GBJ9aZqCOJxPLv6YnO4tm7hvcNXFUvhb
uCE2bQhKNCG9Mv20n/CwQmDKieXSM+WAxfED8Tbpn8FZp1WjtHiUXwnQn/R4W2v8eVEE8ZGnp3KY
wpDo+XBpvlUxUV8eIwd5IFDgGtbBd0tBWwtQAyKatRVHaXubjgUm/9awCU16OezE2XbSVxUVTeAe
0w/i02wHoBGgE2LAIj2JJsSrXskzsV6xROtLPLImRwfpcR+/XTDTQnu6RztTJNd3IgZqDZu50xIr
mLiL+yjdOLphCCkM5gY1+iz1RwymFymsVJUV1T6mB2BYEAXMahAk3NPCiDFeW023nXVEKM3DDnvE
bK6pv4bpp49ZQjjiY3XOg0hyQdbhNYmHnOd4vTaUodb86MJfPvsPYl+yHrq0UrSkkxkB8jBTPte+
k4hVHW2b0hjrJesC5vDA6MMFnkMyEz/i5OZtiawQnc/eioJhqYdDlePfB8cJBnvxwLE+Slu68ONj
uVHUZAbCWyuAf2jG/yUym7a66+r5m7N41N8PDUh1enm+Qrf/TGFxxsSHI9mULzXKLW1uK+pPazWp
9FNTwHsOJE/y8r6Lx2f3bSLYfgJgH8bFXZXD2F0buEKTfbvk4gc1fXT43Z1ybZOnDJp5lbtvebdQ
Bqoi3wG0RLo82FFxFfzvdmmcv8+nwAjiCI2UmBoxuNUMokt2l36Hh3HRMaLsEVjT+bsAMNWVEgze
b3uuAsFzsRE8ClJIbjuhV1mKu+jtXSvotINq5rycrCYc9hA0bu2EOb0HmsnnPycKq0gMXX1Zc8nW
Xj028tigz8XVXjepNUQyBXnPdHa5chOfFkVeTp4A5smczB0NpQb46yQWkAZXs0dxQkloMrI8wn3t
rsEmzt4o7UhTzONPqW9DwX9IjryFbZlj3W7rQjIBqv8H+9zk2RXgAL5MjvqGL+NzC9tyqNm2ERz0
idHJOoe/WFfZAbS9nNnCKyaUCRMjxNHTPz5/gaTqXnqP66O9oHtag/4mSti9OzcTnYEFWVi3VqxH
ynfzN5UEqwgNccbXXUnGTZc6Vr1SBWAdzJ85Lq2xVEzDkhZdz3mC801r8/ATB8RcntGNGZG5PUkc
9EuFb/Yic+Kn/zj5Yi4lrLtUXVK5NNHTiwRYdWjYDN3BHOexYaUjlKpKPPL/CH+gAEnjRZ6Uhu4x
Zrtw1vNrLsmGL47FLgZTVX9lBM6TOfQxlChjB4fLGO+9MzTqTM4y4YecbUPY6k0sFfOODKiSR7Qm
+0IIg0mPMWuHzxxHeha8D3ZELulZnLoQJtB1agdCekBJItR59RxbxwvJYiN8ZZyhY1RL1R+Plojy
QSTQs/zV6Z6zVrElmJ8DctLiTVbSAmCWivj5/jvH+hjjtyyB1TiF1s+sjlIP/d6QlacnbYmJpKSH
31mu9n62U3Og8C0mOQKu2k4dV0LsQ6vIkQ3vcnzq8yWcNk4IfEb80m38RtynxDbM9I6sO0O/xOA0
zF2zDkwdzyqi+aJ6yotpScuFDMfylrr3kAyUn3Dyf69xe8nAJ6jApgMwmx8OkyQF+kmJ6DFZVmKd
UyLr40KpluE+SUFoqeRfEs7S0wgyEZpurdpN+A3sECZPO3B7EpTGj0/xmYHXVRMIVjzf3SQgnkzH
EuwW4TZOR/AQYllK5zJS9tfxIPSMCqCT26y0CkL/rUpbUEcemt3YmxnB7agELFbG7D+/X+A59NJR
3RLbyok2TmX/QltEK37UAgao2xwWggZLdtFMEBPDIF3GyN8Yw/tX7CbOGPjGpXtxxTPaHDDCx5K/
ttYLUSZgDpzyoO4ePUIuoeBQ/fUhD8UW62kv0D8fIxFF/Js7tcFgSKw3qkUi+0HVKS1mMS4MKfgx
8M+ryXBUQcmpUX/e07GMa9AYFmxPKrJX7xWviH79gx3qYh9gQtwM+lMBJDW+m3LN2za8uJYaftwo
5Nk/r6IrEHXq01+gvzRhWt0OTLxkjoLVs3tKqxcDQmF7tituSJFqBg5QRs41NMkiC2HjzFJNhOah
7By5muKfigawqjIgJtOaHzPPnY4gw8ZuCzufa2b8lC+fnobcpvEYnpvRFc5l9hcq8QXNwGbNLHzV
BZZcd40PnpQ45/gGqUOV+0NRmxnsByZBxdIvLVZUAsyKVAGKRrBfONsgWV8Rg4GU3gQHhZHA0KBf
nL8gVew1cK0A43sSSzbi5/U8C5PSBv3iOCx3x5HhvwpI+7/Iw0CvrRNRN6Y5LYDs083S5zYBN1pO
0fGg3h5yjK3UamYRFxAuiUZyK1EPMIiJDq7AwhVy2iQofvgWTpDnKourcJULPyfvfbAEyjJ/zDkv
7LoqdHnZEStQrzmPQZ1vqAXtJuD0e1KHt2xQ+Sa4as0XDJjhPot2hj3nmaG8y00oTIYPrcuxW99o
T+jPDJRWj/aWR7mxPvwT+35/7KEbG7Oe/UdiVdO0JUCFM4vZeDjYaqfqX59e3II1JVjp+h9WA29u
mYJo7Lx+ZSQynY4b/vVKeuzlY+xNV86YXX0BR74yFO5ulsPGYEBysiq/jOevdGPfhCQniGOqlE1r
EAwgXtZJAsh26/ijZKu9FHKX5crNTdhX8Ac7o0/HGqDshQYtsc9UeTRm205xiIw+l5OLPVmxVE8a
j/UoaLY6IsH4PNlRsdIiCI65YYta/pMvHMTXL6jpWSlEsJa4uuAEw8ZlCag0m5UicJDleT0kxkMN
7aRY/eYV6eB2YSzwNXR8NGYfkvrLYpRRXIEjXGdj2WWmMXgR6GzJIZrdcWdKAKV5kufEKVy359BZ
Tg/x0cpt+0vnkap2RuFPuKY0zdn1Csl1z46liHo9EgGfU2nyXWgbZsv2g7mFLjaMYk6JS5B/nOuI
LA9dNhvyd6HIafXuuc/dJbvSy7LbiNg+2xOCCf2775pRwM9nI1cSdTget9XzmWbiNU8+IBb7RTZR
P1dRL5qefqvv5NZX3CFNOQoFdCciwnRsfqPBaXrIGs16ymiyS0j265qsRnNKP2oSBvHUCbHcORYb
cnTUdi2z8jzObRDgAAraK9PmobDhZqVTr7woZg9ScjPWUroY8dca3E1k4ECSeybsPY40ekYLGX5P
UoDK4YX1MegXIhfp8ncR/WepyUXeb9vAinZpS7DE0ZMfyQMWzLeHdBzxACbldQXRnvQtYgS8unzd
rIEF8yUsjZil7i9dF3UzIg5WUTAWdh3vAzW9I/Xe00lI1nIZOsqsRR9DUm/83amI+GA1XQ8HbD5m
yoesvY8EWxM/0A856p9rw+iWw8u98S6blbB6dePIpnqffuj80WW2SneVG93SGdTTYeAV2u0pS7I7
5tlOhyPj3eEjUxgeKjdOfq92uqrUukfqe5Wkk1RWotcCgd3wTob4IIYAub4fKXstwvlNF9khBpFT
gz22XGefpJO7q8tmkjzTgDSjQkMTgz418tDfWMiS4S55YSCjcTmLQE9xRPCLc4PRHeTpxsxGxOX4
Y1p1VdeHKE/kuifVfeFcoYy9rco20qijG3OSb0JY5l7UWraCyH3N1HOnCpd7AlXcZKEdGL7wqHVa
ucKgNtv9QVJ5M10iYbc3ExM3Q30cJHN31l/F/DVl8+kYnYOwaDzXoxT1es6bNDay2dtkTpx9jHNp
pKCjSdkT4kXnNWX+6usbPg9ZoI0k/FgJAs9sM6QAGhnGvUhF+bJ1QTkGZZZZTM6q3pjpFFiE2D62
3VDh78H1z+VpWunA4bMhNO8SyDVCZWnyFDvpoT5OT6OWxmMD5q2AGQsKAm8BH/nfQg1aSOOoYL3T
WU+0CIXmzYVBK9JPQZI6Km85H/WzvvWqcNWX8zjXDbW/1mR/r0ARh98tTarSKCJf6ybDZpFNsjdY
MEL2j9xsZDD3qmGrpbQJ7VdSzZq9tP0Di0BS77yo7V+zJa6rVv+fxyr8CtUv6Kww7OhcsbpxBlab
6otbLdf8GXEl/MaGvdUqNaZf6y+qQswoqO5Y1q4kcijXsl/uUS0pzDe+PxkQsYLQrKB0jdTnom4g
LPA0K4gQ3hPvjlv1/t512ZxbCJXN411sRveN+t0E2eXbrSELnRqWHtlGJaki84nt5qVMCYADISp5
lb9oMh+Mc7p4kCOiZ/0V8SmX3PADGAVUpzCRoDyQyzRLIipOv1TuSiajV+ICTpO07XLzq5KD/FmZ
wdWry0mc7ejB3wiVz7lk8TIPRINKE9pWgckacdXfJUXf4hLrQVs9HWomcrHNRY0BUMkmYmf3mwJL
S4EBOIrK7zyu0hB/PjZxZ5+TODxTblll6d/jKIrimRO07w39min42kwZoZTC6S9SXoZkLK7pmGxO
wY0O6/t0Ii8+ocBY7IKNZFO8A8Vaw/Yi373zE15Maag2YXM5I7OhrcEjccYSj8u3q+MjOMF84x0Z
e33Djtne0o6JCV2GSj6qMgRf+v9Y++3pIEYsuBLGgQwk6YUh2IgjzptA1YtFFZXuYxm9wiBmdHgB
uRXcvG/m5tnd0burbYVQKAuQvD0bxPkHPxyuzYB/sbA4UMgYV0Dw5tVoEhc2YKwdA3MtMj3o0yNg
5jwb+fBwudY+MsLadapbZGlXhpbAfSEvc3P4n86CpBrnLGeAcu7ZSPBHTH02T4VTjCdXwduV758e
zEhT8Zx00W7fXoxHTfwxsjEyqY4xeVibS2qto9ROlHq4iK4PWQhCkReapD+AocS0bA9z0xwoJPCM
A7r9vxlaI3MqGAe+L8hs7Of0RXwRg+Ei6OJBqi318ZBe+A7lfnhGJ+lZh4dxsUA+dyT3UWCvtep5
OVSMgyKL3VVNV/XGWJt44gRlzg6J0wppYV98MHkEXgtDH9t6h/+Stq1iiEMIvR4ckVQ9oMqiLmlJ
aOBgcUtLT/opKZPZzSRLJcbToNWITTGB1FXh9tXmaRgGUXdlNgV2+BtSowNmaA/J5f1jY9fk5epD
gTjd8FsdwtfdUcyFGAGqUIkmG5MoUbO3esIDEdccaZGgGU3Sw+Oo4faA3lPOL0AkfjnPe7WZiQkV
Pf5xdO/+rXyhjsAq8t+7xUrfSZNc9hm9JzjFWE9iaHfAwB1ks+pgzIYmoCRO8jnoxYO6kX8cxUuz
FYze+Fwg/odzfK9q6D6FMG6VNhxmPsCGPlpFmmkF9BNte2gOh1EvydhFQ/zqdRWBgACA9zC0PEDW
me0yizciTl9O4/e7OgFwMo6jwknK4dP2lb6/k56tzvWbcznkbY7QhMDxHX1Olscet/46+Jr73tbD
bwhuJlHakbk5YlQIwC/JtieLplRVwl6reL6/gXtS4siCeKiGnXxZ6HC2sy6OJBzjgQtTkhPSPahL
QDy7pPaya5g8CcpXV4TaRfLr42lmKsb1ZAEDayjE30rUpkRRjmtVJEkX8jl+Y5z8YiXeQIkSY/Ek
BdqtCGUdo5iyb2KNvtplKjd1wmdmx+QSuVz9q43m7K30Sg3wcdmHknq8Lk6pXY/pNfCFUN/vk/Ux
nSF72zyW3FxzD1Ot7dwLi2nK5kNWdUri7PKpZYPIa+brMOSD5via7Sxln3CSp+HEMzkeWdjw/R8A
4/Pfc/HHO1NbazLmQS7mYSOeoPmJNIc25IRUzL5jJGm7uTm7V8U7r71RtGNi6BDh1fyyEopLBYGr
kzwoqjcuZ5wYn4FlG+tWoNimNK3SfQpe0/5IHv8iGs6nWPqzLKrchy0MnBXlFaX293QfftmLUbuu
Xrkjntsq/apO+spRhv/DGUTHW91jcMp8T6WpXSzyFwoTk4r7u/lOgH1Vzj1l8L2eTit2NNqm5RO/
k1HZzFyqOdZg1LFzSKpqj/sPqoKDceGRSLK2kW1NtbOfHHyYgysxa6JH4GOhLLMKSxniBqYkVGWY
SIpOGtQWGSci3bnKSOTUFjyN+Hib9PYPD5J7oMznrAtyKYwenr+IHts4q76JRZ5L0U87Z+G2zwyt
iCtECC++ApfIKIpOxoMfMt09xo/3NfORuETRsepKRKKx4fTqfysq+xNckeZqpEZcIfoJhgdlXieM
bUdnDcp1Czu459AGZIf/3bNwi0smVOSdSzBi4hwgj5quXDvNr0oQ3VrOkvoF5Q/kVMP5hjhoSOBL
5Fv7M0czUeC7lIXlajaGewbVm5NlZeMrcvUoKf786l1a3vOhrfAUjqkl95mys4b1c9MclyVxiam/
ijsQk/SUDWOJQyAIHO3EMm5nST4jGhPiRgIHHRn6qDWXT44QhmmfnLbbXJ421C8+251Rj9FXUy9a
ufAknnNvVTRGbD4uFXHYX9G1MltLBv+uWAaJDSVo+2BY+QrQop38w4nQ1kq9p6alkSnRq8Y7xhtN
cCFffuimGqmn86K9TeD+H8fOMp5z3vEp1oMavukpKur6dYD6NqF/rjFkR/0V8+y39v2/KxNBHG0T
WGRPgBch7KxnLDiA18Cl0ddSI5qLS35DZz4lvCu1VXswMIa0O3oc5jmlG0zOthNiEa5ZELVguvQL
sL1GG8JS5IdTlD0zROYcoigbB6/GwWQ1P2AMXKatkz5ZpLzMGhiI95C0iGSSmbt0lPrpeGe2iWeJ
qysubkMPtN2bQ4fbymuG7KFv2O8thXhG0nVncM6fjgn4/+h5L8fja6YoD2Y0JpjtCE3DT6OtHs8s
f+Tv0xO0p65+0uIvOGEMWWp0Y/RQXEDLY791b83isLbkPrkWk7i+DnutC4GkZZsm3r1CZtG5vWt8
GmbbSElzCc3Kcmox4qemWUWt2mp/F9VwPoPPKGRyhTKsVQT9uFTd4p7PJfRpozxCdHcAaXmy/Ysc
n9rUrMgy+J9UINF69+ijsVfiBUa8UrZpEWZXJrf8z9I6H41G5sQMREhDGXWXUStTjKjDWH9817xb
AsXX2VdCs9egbSOmBdMeh2ckzlyhSe6/yI5R59xUtQPnIYoUR50PMB75YamcOPy9HWW/DVID4ype
EQOtZBWN4anqp5queW8HCnJLGztsMzEt02ajtyIVZX7WFZ/QnhqPUA6EuiCyXMqEodhs+jn+Gcg1
V6ufbk4V2R2QQkLc+WpKfNWVq6NzH+Az3KefTF0QNwVILpYJ8fp9LfWTFWZZ6WDILtEE/qdKLMPK
LaQzI3sNBiGsyibqDD7834/Sw1E/aPzMDhMhflh1O9Fywa39+pNoy0Y0uW1uhsRWkHrAHT7gSNno
vASw12iZ1nc9mx5kCTohMW1zNJKfNmz3Uy7yFRrZtzFF4RzDn5FAqNBUYkYqverygSTAkyGGLwQM
VdrbuIhc7k7BYv2t01rzVZpG0VXC7oULcAsf/t7xLBnBhTC7vVrGratKkOLXr+LVo9f/H1bR63DK
5PQKjsQnyzedaALU9lbkE1HLKMYZJ82wB53/09bhDFA7B+Hmo2X2KwuOoiGQ70vH+kij0z3p5TD6
4vBh+J+PwzP2G/RKvtt1Rw2qnKTDjyEMZeoxlWibccEUIzz9kDrh7m7tbnrcrHixt6sLg07VOvUe
GjFk1qNo89WNKturCb99D97KP0I8FH1HvNrDH3xu3Rpjt+Vrx7MAoC/E/Geu7FlUSBum5KStsyzS
nx0u+SHn7jFlwDN9t0hYre0WQg6k1C1Mvt0k1/hASdUdaUJ82HyW3h8cBbmnEjb4Fg71HbGXfglb
tW/9jzjWO7O6VFQapHPvlgpTzsNdViEXU8mJDNAiWM6WRPxNJ0uHAy3HzBI1vnw6IdOfv5z8MEB7
FAXGfBMHlYsOLYRrLjCOv4BVMsW/cC8fhCVGQsw1RgU1SptM/2IE9pcJi2CcCrK1hI4NZ0+T8ptC
iqVhL9BVmpN6vDYTt7jT+BoCPCg1Ust5GyyOYQRoy2c7kGv4ZJsm3KxaBFeUtRFzB3txjIj88SR1
xTsKrFe9b3uAZH4SFNWxagxCk0qDSVXjAMoqtugOCI7ktCtFytQDf6mJCdyV+HBbKsiyIliZiIbG
Lwbd0JM89xXgAyHJxfdNTkJ2auRdEAa7JvLs77Z7ULVbbLMpzxJjafBj4QVsTtUrNL/W6K4tqi+w
NdFd142DFOSD6wFx49TIGdQXLMBo04ceGzXvrjJSDbEaGQ2jqUoPfJqUXANpgVvPl46JVCMsn+ci
SyQNSH6hpiV9S3rnffOXW5aEAJaLcAR2wEYi+QLtTvZ5P0DWROCsGoxGyUFJiIDSHUcahyrApgqQ
gIKMsWek8IxzJLxeFUsEO2nM7p/hBmHWgNuSwXWfcDZt4zUYhBepBogwBQxxxs44PWhu744Oy+nD
WL6vDFCac/h1E8BTsMr+3QSzJS921N16dCMxNRXyBtub+tQrmD7jxxbJp1Z4B1418UJPP76pHFvI
d2GK1LlfzITtqxOR0tBqVBg4/euNCX2RwWwKNr6VYlmw+H+x1Y7BoX3O4GlS/UGw6xs8WffMrwg2
GNQPt17oY48DunqvKeG8UQAXaabCKcRkAsjdxgT5tb5x/CnLzDuFQe0219FomZwzL3xrSiEge5ZX
tUqO2IpMRCMoC9O+2BvvfYjDspV+HD+cXUY/+2VoqUCfZffpTNjiyXzYLHbI4ORu9oR+sQEW4EvV
RQJpramZwi2ZqlyIWfz+I0bT7q9bVzOeB5b8ogl9PwuD7m1SYAI13dgeTsixOHcUnygDpGWz0s9e
gIU134RKxyebOL3wGVJcgHUAzXAfPUorGNqbJNXeOnWZmmLbrIS9GG3UujeuBRcJBJR1NIWGvUmz
cbppICHKJ0CWkie+XTDFvmujPdwvQFQMQPZkklmmxneMbN6dr1PChIiVU37p1ElF+faGEUa9Hjzx
uWifYONdcN76jNkl7fvfreb6wKdEV9xvCT2SA9YHMTVFe9xLVQ2QxM89L9adgalRSXtMRrMlwP9H
R74DbiyOckHkCRTSRozXy4EYZ1t7FZDdGXMQLqqur5os6B2KDj41mtmnJmCjVtvZ8fWngtdHN2KX
4YbcCtTvIrbXM3NsxN3XzJXNgHraqUOBkE8dfKh6U34oupi0KPTFCjZT11ObBi2pD/VriwvW7is0
t9HhzxZYddGxf+zMV9IWMPmQ6NoIYD5aQIcNg3oZhX2HcUeAp0WBgn16A1vgftCJ02C4ykdOzeRF
LPiR1l57+x97SCPyvWBBuQTZCe51leCtpKtmnKeac9VvaHRZvpT6eVZg3KbjZQt+x49WzTQQ/ezK
RRQNzKTJf74rvFtsNeV9DDk1hG0drFxAsktvJA67MtJAW49VRFc+0gzgJvdTVT7TpLI4K5vg+NFb
P6s5aRIli5zMxhHGU4OWrdl8jEJ4yrXInMN3yFzE9jIBZx4yVgHhf333VCEulBpYSJD3RNL/Yqry
2GSkxJoPqT7Bfj2PMGRFWzb3QzoXLT20RU5Zda6K3WV95AJTDA6oUvHZNdJPcL9u6Ustesj37GNn
TiM1f7Jg2ndOI+yevP9uJh/jVfdfH/mW7a39MmdJT7u+732de/SE9IA2rOusHucnkwaVviA2rIrU
kzIqiZx0BiH/SgQjqpUt1svKzk2oPHP7+uEczSLTBMpRzrKW6e+KvrvBxctqXt4hpT6nQKacqz2v
CT8rju437kZIsH25n+BZkt7+mkCbPK+CL8qSspVXhbwZnW3Tjnm8/X7bazhARQCTuWh2mDApeb5y
gfRu17hxnv09iWUHr6UndHXcbXpskJJ+J9Esne5hRLT7JLAHnFfXbS85JNCxy/CiC9Yv2xapXVeh
zgnWdB09KWowKtd4Ri5GOFM27ubcmWN/HDysgUQJpQAMZsfZ1bDxqMm1DVA7njw3wPUinEtmJbmQ
gLoo3mUditfXVuSM3UzKVa5OpznjMdCsG6nfErc61pguqwevOC0HGTV0Ml2znX5zLlhGBLH4F3O1
jXQy02vMFZ/JpdJDlLtPEp5tbCrfB9B7PHAEMDDZ+o7GxwZy5pj0OSg9/gdUTiONQ66+Q0V9BOAe
jWWCdhtQAz6otw0pDV8uMlRrZjAGyK5BBtX3yXQNTuVBhAby1d/Oims+wzmYX9XmvJ16VFuf8QsO
60x+1z3GXhRqQw/FBCxyFiQFgK/2FCU2we6hUYAmwwOzNXQTR39M5Uin9hUk53U361fKSU+af5V7
WVq1NLdCsjTx5JR2toY3Pf0LFSA6lDhHLjf4rq5VBWSLIkYzyDPOPRlfCDRb43CnP9fZu6cYOwk0
z1+Z/0piqHfBXOvhVhPQtyqPI0ykXOqKNnAERQp3wInjrI9/4TZT6rrvVbGPu4vl0c6i+G3v5TaG
ZpbTfFZbJ3HqvOa5Kq+IbS/Q1ytRtLfP8kPQ1gk2wmEEMOTCFKGfiQjGmKuOBdJMWNEyt0hfabcO
81Xoi5iPYs8B3M7f21ntPV6nFN7Xu/OQXHuPJXVVi7TJAUKVl2r53FoEd9OIstzR50O1E9EYgXrZ
+NchTrpsFy2BE31LtHND1HqzaAGJnPLYTEZRJGxY07nuoBoMDDmCZwMy47CsPFu+oK2lQiZszewT
Z/U1aDce2vr4i1pb1aKHvyrMEwSg3a2kZMADSYrnbg5hh1X8EYxwjoMj1cM8J4X2f7gLz5blTXFH
K9QDJmovstm20XuIFPCmLO9I5OiEvaIgOkyMLycf3FeVbFcstVULmZE6+qw1LnMiMQTVIS+/t0L1
B7tDvu/byMUPnolzDA1eudIk77jPPpdETiO7dE3dt0dVle0ihMeC0dSAdEAzieryWgGcF5DZscCB
nbhXXFjd/Ny2dXOPdnt2UMkGZeCxyrAyZF/PFf084bnfKeUO4lnKDXxCHbEJoiGyHIphyy+Px4D9
0hUXu1dJbdAdiqYcj+4IDz9+PCb99WRfcQ+qzqj9oViAbFbSq+Nw23TdMJkOWn9BQD0Ph81ny1jk
hb8S9tgQsYpClFQlhT1oyxDI3fmHWntFQgP6sdlNCAszfP0XrMBQ3QiocnROFHzI0kQDUYq6kxi3
OA0kmKWx2N+LhjjxGmuCEQSTXhNdsQmSdi8WnUFv4Wgq0ZZBH+eOFa4MxAWpreSR+XF0RmMvmWKj
7oGLAQ8Gct3/VqNYcf/iCFip2Lvw/KN+6Nprx8w2a6aXUB1AlUx1ocxwMwNWen3tnvJNuI3QrP90
hMuFwE5pWz7Hem58TgPwF7xqKUs2qDD2Rl5Fl8DanCgf4uv+WDQjH3rMN7t2ZX8AB/yYHNJRiZVa
0+L0gIxZF9YiL4p61YtjmLSVg9x5cwN7EMdxmY5VZI6igXYI00xDWF0Fja7s5mFIsOD2hXkIuVzo
HB1HWQtWh3ia2FwXkkkj0YqI3BjfhKBjcmbYzoHbD5tESbWl8RqQS388ScuomYsHaPfq+LUCPeiK
I/+Xgq8HtPm7Cm1NKIXSn91l3adhS0JHBUdPON0GgrCzuAZypcROHrU09sPdECtyRAYByrgem0Bz
Xdk8Ls35GT3kvgrBfFi4dpMvfKYmRi8GwF6UNo9CABpuwwjjR1DO92mTpnWFT3RdYPbfE0CPnh1b
lgnMUGEx/BI1Lftd0oOItCD/BV83x/RBgMziZgv55ftCmWe7cv11BIFaxxtRTA77MBghCYZ54rq6
tJ8qb/pCE5hwBZ4e732oQN+cFuYZbzrpbiNaLlAAF2frJKQoVNCRstGtGUdjPEcnh+8efGjkTvPl
Xa/2quq8yPigDz1HV8qIMmo5kf50aU7rKZfHv5K0oDxMMseiIp8eAJh3SZqlaoYiUPa+NeQCsky/
Zt3LdDUzNVkh5oJ0Ie6gooiXQVI6OgCOqzpqGgstYt8+ttrqFZ9QMrmB+BcAknzSSxlFLhrAOjGy
0RFy+tTj0HsABOeVSbbTnd6UDn56M7mAnrjKRi2tzscFEgS34ge1gT12hpWTtvCNRa6MNQNaDnYs
Ffu/NL9vWvJIxAUJe5Aullx9Im21PcVuBZCOlPKQoRnX0q0bmB1YFALgtV1MudpCLPY/wVruK3B/
L/p1wj29OdUzrmh9b0ImLq9GQ4ZjUskgUk/YDFPoukV66NWW4oKm8PdpRmBfY/GTYVFVPzhk059C
wyDduflJ53hYHUbyhnBkc3pWbHavLP71UL9lpsWKwM//U0kfPOc39uW3WRJfeS/7CYh8LhIl2/Cp
xM2VPJoOxwKdUKHyJughyKqaVxMFUMCcdeaSHhdZOpyhZsl9ijJR3U0GD52kYnrwR3qoyU2bGe1h
1DWwhaFnBlGDw4EjjNP45zEb91DmUyRX9K8A3zfaGCYWrZ1ytkzNKA6mFufV0828jk9P6+vInUib
32bzyp33/ZnaZ44tzCkYLsosGtKrs3RQS7S6y711+K6wt1O7chUg920UTD9UPKR818uiHVpcTzdz
ZLrIhdRIOHAPRwtKgnUA/fgaULVpUHO3AzuL2mqeYkYQ6S8204bTdN+vU5OpQN0GSvIDDS6LHjnr
T8TJrSK+IxEkT5k6FmigfSjsqlq0PY6/5IHBb5eEctxAUWx9zXrfnuMJOjLLEQcFPuZfUrnLLTYn
0eqb9Yf5du4s6IiBuQGYf/LGBCyBUuBTchXHh18ZBIY264U1XyCqxHoVW2qdplMxJK+ZO0jOey0n
H7gdOW3c/w2msqrp6GpDnXo5pkxMbMhs77gmX9USqSvangj3vv88hvUlvhehskD26OUoOOckuon+
cml1awX43OiJsgwNgAk0Tmdc9jYzs5HECG4c38GLOvLSsepRw8wUzT2Qjzys98RF9pW79ES+aUto
ntUdpmbsblLiFJvBZqx2YVpXRx4LU+357OM4A3ZeQzhdNQmUns+4Tgymh0m8Up+nKNyj3Y6FjBcm
TfpXkzAdo0wP2gSQVxWy73OuRz5iNItSnxGPxJJ+Jl9A9KrbhP1eO+JBFUrsX7OdYq0Uq6TX/PyM
9JC2WTCVgaJ4y7S1EdyRNIGPzEtowDxKFeD4iWwE0x7TbXu7+gk4Icep3niGEhjv1aXyz6sAeE17
EnOiM95a+F9qXydsQ3k1gsWK/YxN4/FlsZYbvwN5dk4+vU84C2XzCtxLnddownqwS2dTqGeL1xA7
bmCMMG5yQ0cVHVNei671Hoz93i4uf0/wpN8DjBP3LAjO00wnBr0AP8Byy8RDy/paf3qjMV7wMntX
V/CsRVhG7Cis7vUFs2cK039E+NPmsz6kPQjeeFrdHsDjaA//QlqXdtyl5GWTwLaWQvNP6Ut+zA7x
5Gs8BCg7nPk7f6xAaEWjYvvNakK4H5V3cunk1UGs6+Y+nX54RD5Upx/YJRo/QCnnALjK2kvmpZu0
A+hcvWHONHiAUtPpsgWkzDumHzRkuzWfZeJTsjzwAxr4wo6PRtvJyy9awmd3RKet3i+SxgPyuNOa
IMaVKnDd6DAs7njuHx7faLMoEHSbQVMNf9dhoDhxzS4/wCh/ya1zfqeRHn//ziMjkyrmoR8aPWnP
kkJw0wSa6fGBrAQXLgwVejlyjuaqZVjkXcZjKhwkk/jh0ALrl2RbnZUUXseAmREG/tJBK69cWKlc
1GZq13BgafSoSXOXP4VxOE9sY3/C5upyDyiYsl1Ek8senwJpPZn4ObnO69BKTp+MDRRW6LeSp1wa
Wns38L/hkTbNJV6lNDXP+C2fsI8h+uzCmq0FP/jX5h/C3HhdBsjg3hu+X44IjZ36bZhdU5GJbMfo
39cHGUkzlz1L5RTNQqaB69c9ogGekCi0rPThhvj6ChzXhCWsNQr4LRhx8IVeQubOA5gA6MSVX6Cz
HRykaof+oWNCSb3CGxkMBm+GPerQqv22EaHxBZrzFouIjSDAnySadfkpnp3u1bMd1Mo3VSDwLHIM
ZmZRkQ9QH7UA4BkX6ZLO57YlUGIDDZ3CmKs2Hgj7VhDE/ceK5VHbQeK6g2wJIq+M7c8nPCu7MChc
omkUtMa3hZNGXLkp3JDJG7fXzO4MMPjKqBa4MHkQRkDzlvqFNCpsg1H9+YIulcQrKgpohKt35hOK
RBgvkeGREvWonimVQr0+5lXIJfxxH8pn3N97R+epdp7U5Ue71G6H5tFS90+4qD2sx/d5r1lVqaWI
jwlOOQeYG59nuzccwOOGOMcQdgPrCyG1QBa6IA0WKEglOsZtVlvcZvxfZrWVM9rp41CMif2o0EfD
2gLSwes0MY1KC5ZyONoaSkpVIGolsQ3wHLW8OFWS2Y9xgmB4Y+lSY2680ElHuAZWb4a66oxpmba0
a9tIZbkGPIdjT0d8ymg4ru39sKe29hMdKc3C5xoTLe0D6bvlMVCSpXPEYdkBOsxfkHYbTSnhQp9s
0JRPWdxrFt7JtK4HhvsP43eS9yipDuOk+mroSbfOdyHaYw69X2EmXEOzE/GSEpPm+a84VkfcsKM5
pGpSa4wnp76WW0UMPYG5Y9n2LsXsrYY82gyAQTU0+BS1NxjPtwO5bpXxP8ZtxCjTLv6lbGpFBpv0
hxr6HD+K0fXx30wHj6pTTitsXiuiH31x9kqA+AjJYIhtVX5w5vv4laFrVE5OzLzH5GPaN/pjapiW
QQuPszqe6q/nJh48GCXPadjCgtM8SdTYCeG3sDwGLG0V+iYC2L7E6pI7N/2KGp7+8chgwRtWyp2W
SvQ7BvFyB+xCHJrHbqRrNJhPw5eGCadzK/GpYkOQYbFHAgA9+BA7YMVgdeFewIj4tfBhthT8Hn3M
zxBshQQG7WplOEi4e8IN67MDDHk+0Zi7uQc7/x4cNzIgq0Bm5g87bT7C0GG6yR/CQu7zDRCMBqsE
0FGfpk5tolGr+KSGt7AXehl/ACMYgKlSOW0S9G1XvMU+0ptd+FFkZ2SnRGiO4hcMKDquzsF97ub2
Z3MBqrEidrKqVcdlASQoitVJJ5hsXKRnL88gg5gTcNOybpnJE2F4Mnu1dw2EWu3FgR9DT0BKm11h
6/kYG3k5auY3pPkvsvzmlt6n2HnkXFZRxO5AUGK6sh97OypuzciNQE7uVKde2KatIWuzZp60bKyk
fba1CgvX78llEHqPKS9EDz+WXpTaG1/P71iNiunSZEqius9iKwj31BvlX9v1pLNp7mutqS+KjjSE
Tg3Q2I6HG/BXc49PtS971xrEJnqrgeMZT7lkrWLQEqs2ByWNPcEp+wW2EXNQTaTujJGFRnq5smP9
AwuuLzeZioFlGdQHkg+znKFNq+Khx13Ezz9RjBO39qkzxyfi37o4eILsnx913waHOzM7Wo+bA09I
7gqo46e3SkUK6VoY298GFHFAelH4dRqMGwFZ7eMw3Xw/sKf/sfgHBNm74bXrSnjj7Jmt5z/ZQgrF
i07f8XVOcaEwdtmqO1U5E4dFmFRaQwgbxRTlH6V7xtLtmCRuiogiO/+nqcN2d14gNod4k2LhQS5N
vo48cjDGZNWToe6CsGSALqSpVY868bj3PKQ4gPh41IXdFJR4KLOhE5/Jxb1QJMroLiplDOPKbRy2
xiuZpWOfPGD7GoQfJl0uIXXmZiN249EWorNO4rPbpe6VVSm5n+GZHeFA27bh0i+SQXV8J4mNowxs
vUfsMrRAXpCEYsuuspjclZNh9p7GYoCFKZQgQ08ElSnj0d7kGpadVSf0VRVQ9obEWaK7ZqX+zyYX
ycfvtSRgeeR5E27wcM+um0b11a+u4/0cWNfJCgPUrO8tlHgLfQ7LvrTnwz+rI1JAMti6vKnFAKgx
oX7XwD9mjBTgSN2q86yRIlR7/iWRZ6mRO1czWnjBWqLFV+RlH61g07yVT+jdb9Csgy4T8eYDtzbx
SLCe62uJ8SyyuY3TRu1NNZLctEq1OUj3odvXTe3gnrvGeRJ4kcY13LwOULHbIQJURJVkW9ftUyFg
s1Yk25tImJm/+b2LwobzwvFkkaF5+npIK/gxq3UAlP44QAxhgIL2ZNtwmixHrnlUU2Xqylw3Pl3+
ibt6bNOJk3+UH6F0BLz82F7YOLbGoKegHNvfHgLC8zim+lqGNAJM0hrlf4PjcmaS9ARSiVEScAY8
fX+BUVQbnKm4cQMn0ZhreOINtwaoabZM1mi7EI9h6vc5zBWPIZa8vFGDv3Te7C+MC/BjyRaR2qeO
fcpEMfoFOwDSUJ6dKWFLg3VOwfG+UGwUwZZylcN44c8o+QHe+JULougHnt7yqWeOYXOtYid9Uwbe
RtSwHEpFRfxE4GKaWOozaOl3xUrQR4GeyLNW9E0qDKDEA3XA0QbSyK20W8aWGXUGUHVFAoqNAYtD
3iswuobvd3CwsHRkvt68RS3PuhtBz+gDonCgwfmdO7ixUSgjlI0B6cxthXUuNwPZGUzYR8nfLV2z
db7TP1O/aVZ4CnciTokNXrN4Dfuxcjk7uma2jorH8q4P1c9sk2KT0ryNMtmgoOleHEQLXpVXcpcc
PyM3HtsynrEW7QNWLhNxolCjf2HZJpC7lLuHPfb+XJ7IinzzfTmXt92Qjo5VJN6JDmma4KVEfRoA
zggCUR5FyhTqtyGg3feVQ4yqSw4ma8j6MaK7cn4yI7gJKj0O78+VUJ7kHvUwApY7ANyWMAFOvzwf
EyfVWDwSYKEOwVpfNo+W5e9EYfBhbBrfHfpQpIlM6R5AJmYfpZTqM3zGEGgxkab4tBWh7Izp4B6I
+Gs4t4byRY8dVcCGTAtXRHtDqJU3Itg9rHr7ACcQ7d3JSIhQ0rsr+hwH2RgSxG/1LNO7ibL9yFGy
p4Gdla/jFujyiu0LAHyOTAmrpIW4QfU13XAaLZN77KNz9xX5HaDlx9dr4/e0FMqMNufz+9aTpYyJ
eEIAQZ0/Q6X8EQC6xAC1WVEgJ770+zlrL6xMvmnbVbm5rnUtf6wMSjxzWDHaaG/pn05i4uuMDGWq
ViFR+0QE7+C4Kgg/LZpjgldJFlE9EnjCmYd83BV17gIZrAWQzIckDGsQb4ElHd73A5oxLxQu4jx2
927jJtRuUcLemg2rigxKSLjz2ALAJUDqnL6r1Vj40v8xwzxWA/5czzkWChqRnYyEQMsRXYoF4pAW
XZTY0ouYeGh9Ao7tY+DZ/qATcmygCLudA+KuUzhWnQpu71edS8I2gYhwUjgAstfxwToafNnAvwjr
aDwdBA0IYrKi/tHUttwQeX1lCQnVoj0NDDnmF9d67QUXVU/vU9TwxUUDZA0herljpwsdv1TAFPAy
ENoF9G3s0abD/bSeu9Un1I7+8fDTM5Nm5y/ZyWUCN4QGD2rognv38AtPNUAQRFBaSGvLmhwB75zm
uBKW09BrLEq/wMGbp6In0JW5wbBaYr7BSbYcPgTEItQ4ILAcbr6LGGTqc7v8KvQ9SoZTnpZ9t3G+
+iLl968+q+khHMr1miCZBpeM/omnYBup3YtoKISAXKnHhzsCTxXOqjN5T/S3AsIExMYFt7eKfxlS
1CES/QXqgvJInctscZFZaG0jv4olYiuClufdsQkH5XZjg8KD0+qdJoVF5mTa8n1iNx1D6te3SECt
VDWFWpJW9vEP5/SreiXunUdFugVbo+zVQ0X16FYS+UL7dO5JINlfUWwAgukS0herpy1kttSsTFiQ
KfTvwUzQFQCtchSvGFtKa5ou0bPkBDeJg5RdGU8zC6U4WBJn+4aMAZg1SiPX6aNvZgXGguHEmt/y
8suKj9U3IEd5injHvlamPgGNeA0hR1rOTWf3SSxto5DEyBlXcs7LvW3ByB1erDXVAJ3smOoakD0z
7ltFdkFP5BvdOaz2N1y8w7F2LkEeShe4bW2M7daZMJEJGQaERPxiwG5zDhfHnFR/lmCyaQa/Bz4Q
YkeEVyQkSGA/5aIlPo+NB9vFmgj06lSVBga92+ZLS0GLqOdg4FM5i1USjQqTcZ7EFmYCsSriYJQq
xfJInWhZhWVlLKCbKUCfGoIxSQBEr57Z6Y6PC6H1y7jOIKzHlhr0ZAv/jJ+Gj/yb8bwKGF+vhOJt
3Mtv9+QeL4ZRDAlXKquHdossYWNmY5AVxmUd64p7rGoe4bvIhHypGD8cK3gzQ4YbpfIQDdcHjgNi
mMeqV4/i0PHmCU1SVQ6oMNhgs6hZtqy7W7yVbjmp5wTgnPI8pcs/CUCWbRzt1tdyJeZR1wvJyU4I
ChDhPwxktmO7ltGljEoYP7rmDmKQBokyr5s3N5cvrRreCTlD7faBCyXT+vNe9X3m/oNOFGfKpLWI
5VVW7skDOXJgI4pQ7V2nIURmZZ7HOSJd+jH45i00IGW4Vq7wlxl6UrvqulK/xIT/eiQfXr1Hd7da
h68LUfHhuwe5Am3pdCwpdLE23wwdxAx8AijkyBP9JcVZ9S2aChA+HisbCIvHxgY3uR9GPC6pEN7E
pJ1vCasyv5BmF/AoadsVoZGLyEQY1NAoszR8FXbbaHn7TzcDdos2yKpRS9l1ecopKiWBVE75Q7oI
y+Dr0lP/6MgwduGZVr3BBCBZrZtXnsLEscFRJjS1fpm3JsIkpgMfG72SJ+/1Y3IKK32uxYBl8Vdx
8Q5lB4BMOwoEWBTQ9CJ6qEKVPNNS6bR+lsBYqjLwnPKfrlT34O6PiXY1bNo2dPFuTmMcSUY7ymnu
VqOLIMhPKSFYUQxrozwZ6pBfGuMMgmlrlcvbg7g6z08tU1i/CvXvwJco/j2EW7RYrQY/9UicCKpn
AWb4GetmxwuweDuU3C3sI1Lm6rC+GFQC6uHisLB2rI9xCdTA2oNhqHuRXy4TATIPDveCUgUIiSJw
Dbmn25MRCbO9tIx8klSkxs7VJTVkYsIpoVo7Tyw6nAykJSOi/IkR3TzEDr7jg5hsdQzA0/dOXSXu
nzz+vXtWw86xVDrXApLPT9mo52hNXpWED8Bes/1diQyWfGHvSK1NRTp0Db6WiHxYc+7pREj9morc
HWB2Bgbd9gbeLV9a14ir5Now8/0e9fhzFubgz6T2FRSDpjrXRvadEYRiLlN/u+2D6jKQW76i+uFm
GfdeSyhaqbUqJjAmPi64/dlxhvr7aTsj+kRYrrP/D9PIOOABQpifJdWO6MAqeK1g4L3GQsqx3Teh
DukOSM1HTMYvW3mS4frmpUji90rPAQOOvh+5mixPL6/SEBj/ssJUoFPWTPGzd1D1N4f8Gb5b4KRG
4a4nuDB1Pgd0+RMhiObdntC5b++7zkVwkDoBOkmxnROCE/PLtlnsavkAN9LkD1A9m5Doa12cLj/L
c2lIwhIr0zBCgebLr/pl8QHog5gyAmIbY5E+r7JHFLE4WO99M/C8iBkBiYFm5E4dQJb7AyXRxrz3
cV9w4lxi50lSKjnEjIH1+NdXqC1/1asbCWfErOF6ZqMuP5vQAs+IRhoxSanMQ1qka/NHFRTB2F87
GpMbBXNjFQUTi0GbsqBYS5t4Li+6O2O35paXItgZFS2CAO2sCVrUvpZom6EoUHx/PHgjLOaGHPSR
nFT/vP+fTXqY0gFthaLY+V3a4bbhwPV8Qdbnn1DNPAtbgmQFpfnSD1vetQfFZ69snzNSXMz88jVQ
7ZODvhKZuohG/s3TWZUtJMaTgvgD69nIDXKlRox1PgDHN3Zx+xTw4AHvI7bemrJeBD3QGSLDrZxe
ClAqAuqiPgSJR5ncVCAZOOHMH5XJECqd75nKeedx8SKsDz2z07ElbAkXjlUFMgWIySnIr59Jg6jy
3Y7K/DDlgw8n3nJKGpv841l2pR0AnJxwF0N5WaTNTvu3Jk78+bC/ycffGHz7RCxJx4Xyt1avZuKE
7ueYN4i9HpBxp3KT4RHN2GUkQ8QsUFX0EnTNeg1riquIMtA74toxcOcuDEEO6HO04SU/JvMaoCsQ
OP1FAOG0f7QxV1GVkvD7AkInxSrnna9uTXOAAvFmM4XwTouPLTgtfubavZpqD6DrZanXAcaYg+PW
n7D6+69gwVN55qQbT+yHrozKI3hgnd5czzk5q+Z40Am08syULkM4KZ0mFjHL+ZGGNxU2Ckb0KEiI
6yromORcWuLMOVuF31A2milHBenhTwqn+KXC0Z9nKrs+o7C8vqAMV/pz6to/wRZ3wPhGmObN1+Zc
0xhF8nbz1mgOnE/tboItxUc2vuk1FPT+0SxSiPtnTB0QnQSMyrXsmPpZ/W3hpM6CI1iKiQBr1KuN
LnhuOGcr/F43T3mxC/SZXlGuAFSrRbwC9HyMGNfEV2ZeKp+qwz6Cy8tLjJ1GRa4a4IbTS3wmT+IX
/BT3IRTXWYL+Sn8nRcaYLApfdZ3vfoO5xS6ZnAxXsAh75GlMpLLn1N2fABvCrK+j7YISgFpmUzkh
upS+Bw1NgG2mjG0A2q34XILDO2fZu8OXJ0tlPDolBsaTGaVZGnR4K67bBatrRyov8OY+RbBz+AJ6
YPjzkbX5C9a4UTDO8dctTca6RTr4uo1ovkSlUtHUQBrIxJY7SwQU8Cj8Y1WAOHeJl6zgLFn51jxA
kAHvxxZCVSizbWoNvYl6qSomi/QJSsgHbns7Yg4inqMg26KuShLxoj8UN2816vYBqNTQFFz+r18N
F1CmHvyYvUm49odi/Kxs9c28+apjbOjGsizwiheFOJvasyf4IvhYlGcmLkW9iahMnl1nP9onMETa
5l+yzuY7WKXN42ENSm3Rbqp8pu9ZjdaL85pi8icDm+0eUnuXQAaoJ/A9f4aKvRAnvbPeVl+uS2jQ
xviBIbQPzGEwaGUT28bvUszTbareiYgaHfnnK1gvKMBNi0o4OeqLSslcAVxWZR6r7ulRB5KTxYCA
SXB7FnbzcwUl1ZxydEQOtFEpBWd2d01tSJvTFQEpjvvGR+kDQe4wjcgB/tvrIZAbEckdxQpyzNKY
ViBnNoIY/2Kv9tetiDJIFWnYlFYxiAhzWvNm10W1EHMNUS5Tr+6E7aoXa4jlhmzKH+lzMNlWAHyW
Ap5NSgqu3QF7sGeNstcVmJRDjQNuaYIV7tVOBuRuTkL+l/ZZwrnaNumGssBNC9gnDRgdumt4Tw3f
fUd0mSPxvFGd28MGNSvw7FOCLneey/v18NckMJ78BarwilZn6Umb9dSnxenMg8D98qUwwJoblDIM
fe+TLKtUwqiv9PK1RblMA1WhwBQUa4e503RD2p1DfLaOLHyUBzDFHv0UFcA3jVRatny/kmS2HXM8
QlhvAlLLWhut2mGXaNVDpqCg/hA19ks+DqKUetEWDAgWz73cgdEPHk1/h0mw32xrICDQNKosMS/3
JLSTvedzZz/KKAJE+CLS0HoIgAU1Uum2Mz9ida3X53sC8lK9A5gywqcg5UClfAJ6EkV+yAkxjtIl
DOQMz0TgjfzgL2z1PAXaMSmwG/F0XnJtEg6DrCVrqwU4nKrNtWGTDo+a1kzXPNdfhFtGosz4klA3
Nyp8pBNoVA8cZueuCcSblcJZEd9eC1nuRqMOBtVbYb7YNM3Q6blqcf5/kdVHjaSd12gnDowKX1dA
YSJXNP9QC+WzbHDxL0CALTnKbE+xWY84uLWyWQsrWFORariBUjoYvyKfF81wAdS6MM8URq9t6k3g
KWdjDAhTr+uVnaztU9RbwhxhRwryecwsSx71bbLNTMucTpaj2eEjV6uSWYQuZKIv6iqddKxRoCNZ
bEX3OZfBotExs+ZcB2AoVSBJD/L2G56+KF5IuDUP8rVcuZQjmF0yihS3WaxGDeRToDNwP4nIR1rO
Is6YvgbOrfwg2d76rQpiDJKMO8dbQxbzVrtWLavrKcUvAKTCQv/vd2zz5oYlMlZrmogJgoZKnZ9q
aRKiYvyfJLhMLllrPGkLGbFd/eN9J+OC7RQY0HafszXvgIainnRkn/enyEzqz6iO0F3gaPMn8iol
E3ncdRy8LkI6TUtO1h/odYvnWNjjMaKFp/p4pOIEpRiIbktecoZDqF52qOg5suo/0OHwERadbR26
NRMcmucWfzJyOuZBsVR5pIsQWo09WOdYowQYO0wChC5ul3V0GgbDRH13mPynw7EzelLogCG8wxKr
/IBrJ3xc8J6WTN+j1PGJQgAjn9sRNKq7qQfBECvnegT2Z09pLAoD0pRecxzZ9qo5g6rGHmUzhZl1
CH5zHoxL6NRM6BXLtS+6tVwoMUHwvEt4i5Kj3abSQbmv9pYjAKOqs7ZnZSixzZOIjDNH1ty7KbkH
aCtz4EdOORdbwSL2VF6h8r9SheepzQJPxVPQJ4pFePdwvJMVgNVqKRbXyNDv7b3cNH/8MI+jehSw
kWAw7Nrb9BSJqMJnovWuZKTIBd49lAxVCuDYYBPxKVBwAjgVRCS29fbht/rDWH6ocerYZ1gMA0+w
FIO39Op7Iw/MOqlxPF/TOK+/rqUY+LqBvSGnD444/nEvx+YCskZdUah1GoZrXaHkQVfVfYoQRZ5i
scDUgLIDUZJ8/ygoPtuy6Ze3nNzHtmX8sElgDDjIC+i4P0kG0glTGI1jNLg9/Ui4G7xY4vgf+kqK
nEhlJizT5uziFvLvIOo15yueoLEiUvdG1bZRPR5Xf2dy5eylUOXmcQ1cLg70moSBCuBwL4ffrjS5
xiyrs7ctBsAcy2QAMqXaIBNRUsdR/a4MPd5b1xICSWyBHZzqEwSw3QtUNZvx5pWhNgOXsbSNHIf4
+w+T/fSIEgGi9Y1R6YeaKGnTQkIBmvTyct4SDwOSB9kktpp82UEJIMKXV4Tasvz6N8nr/hWasyR7
l/aaLNGO2oTDnp76B5JCO1/+p0tK7uLUS8dNdrESbHdVqcJvtPr4aOjHbd1H4MNGWxK8W/whzJYM
+HjE/QqjOE27ZBLPooGmn2dNETocuVepwOJghhruBGyIjb0tUQVsOINShQXE0VPdgiY+e2YSV/ZW
KDyuedZIyVfF6bmFyje0ToH2hIfAMHUwncvJffkgil7LnNrvyAD31zCADct0xghJ9SC8dXKyN88g
jGcJmZ4EOba92/mfv8PyoDXuEKV0dNqmeX4W6zCv5D2zQC/9i5CyMDUFCcqge9G9MreVcmhvb/xV
i2C5B/gm91st+Gvbqjo1ELKK9xSHzmenrS5EXMO/jWb9IGu8TCeaeyREkkUBkG2fgCjIni3pUUpo
dm9WR7amTsJxqTVdlEA+JQDzs10dYmrCG1fvsLZY9h2faJ1Kjow6tearFuhRlm4mcDyOixddeDFQ
mKEzlRgt/kBwVP0PACXVjx1v3d+DC1OSwb0qOTp+Le0gz8vi0XouiAjbiVTu3UVcIGDK9xrMALdS
231+fc/M7pgN7UFpUOCHy5RZCVfRbjF0F4mnmaGEpl35TRa9ejS6jYhzpKfi1clSgbXv09OoJz+x
6tye4dwSWg+ZMtMR1ecva0fRtQIShEpBC4FL9FElX02nAqzbQew8adrnch4er7uVHjNrhVZOq1On
dYsK9qOG6sAkLqNrhELXGnW3G7Q/IAaYgsRn5w7U/9IXbTXRKN20k94uRMmrfcBpIYhEwNt7K9FE
hDEnG/pe5XAw5HvhVwUJa8vbp2aWj80wxVFhifd+9BhkQYaLsrPM/8eP2fuIb1kqa0/DgrNYW4Wm
JmbJXed99WKXo6DMRG8q32eMDkjpdB0KkEYnRFUdKCBHe+TmzBOF+uhQhsWUC/A3kZh2zIuc6Buv
j5qQBSBGoMKsETqjETPm8QDKNkiKxi5m8tcGuHS0a8ySSKXvpB/YaRMz2Tx4GCC6CBYZH8JvOOOl
14htveTJUyHF79/SqDZs7rRwxD9CMJ251cj+ZqvpPGWlwY/HrYSaXulj+PdyuPpq7myetXjgo6DG
mCecP35M7Ep10HUweSPxqrYk005euyQ4Ubj/njzadi8KR3aYWlnIiLU6mXvlgsIlz+WNkNivHSNo
qSrI17Dbqsl3O7JQMiuwrmLQy4enHcfjojMMZCRkh/Qakau41bKhMWuONDCALTgPPYK/t483IU9G
HgV4cu/bG588xRaj1Rm5htJHB6SilsYEqUy1ZmyXDlYquHhWOmWfIgmGkku+dUdOt6GfkMxL/aHD
mnsitdzY+Lm/WB2J6oOcVYHvyLb/F3kXHFOZUA0Gcw6xabnB7NId70iTdCmtWmU2pQNVzpg6zwpW
MY2mRaHdWon8c+CghMoU9pg3Cbi7kEm1Nd9AmeXoofgh+DSFDziX068SyUyU/zo/3f3M5hnx40/9
IjyQ2bhHDnDxxAsCIeRIk8/s3RUf8jV9j6fiJlisn8lK+nbPk2jrhJ8Ig8bBS/wfDMx/Xj1qN2gV
YL2s8zHvSFPC/2u8cPKesFm3d9S/SEdNQKqA5zdq04yZqt9lbrFfa+B7/mbae47lnkM5RbTcaKuH
QyfWfuAVdXJlu80PyvltuZZztFqMqivR+6/i91B7+mdHwV7BTWmLY9cDeCloczXl1ko6Z8jLUacY
hOmewhk0dphWIW4okwkWUbGy8YkBu5Fppk1KO7F8Crvfd8X53DhZm/mN1jOvlax//E4pbVO6DvVC
H2W880VYgqfX0qJqJsNlQgqjIiKF2kRu/VaeNZzAJ0fkN3UZTXLB0u9cvvddSVOulB+eRridr5Sa
nzYwwAa/CYpnK5nmW3f/TRKdIaafMWaovDQQUTSbiEJijni8xOhRT8UzJzWe5VIb7DBpJMs6cSO/
rMSPnXdd0f1BW5HLW1rjrfedfIk4rLN2E5AdjEkP+ll2gaCkc3HdE/AV2Ng0dUdxZ71gpPp3zGwJ
ZcB0KdVE9TW3+XbMw7U40Jw48SH06SRenVAou0MqBI+hiKRDO0LiptIJVAc4V8o4Tddpc8tVAIGU
loC4eKefNIYwVJ/7zJSRpIUsCfBFA7KnZup5qO26XtVMGTAKLPqmVWjoazeqDrr2TtgH5K7v4IlY
DjIKVrw3hRmrXRKBlUR6wdSAT17RifZUrHIB3uzxCdhAD1ZfA2bFmT81g6a9puO0lqyEKJ44WoHS
83W1ztV4FG6Owcs7ha7PgYRq32OWRW9KASp0UYHqautjCgenDXiK2KbN1J3c/l9sEGNoGdcZ065l
1Yt/ZHTxa3Mlvqbr6fxppqmiIb5jbpMCrNjFi5qtTAWNMSc9g/0hCrpGAyn2kKTgkFu5E78NzqiQ
xrhx+XZzzDLInFgA3Sr+DRMIPny+RISSXVo+7/wCwRWPU5EGjWAdn9VNrTlNFH/KLPUUxE1dIqWD
7ubq9A3EM6iizsWGydQb0KGsQZhE6xpN7+rTv+GxBxvjWHlJH2QU7PokNzaGZ0WHm3aU8ItmqYYc
gB79m2F63hKVjaWjrCkGYwd1S+7DUTjJsJk/mUOwY/3TVKhtY8HdQyNMZ/uCm3P4/nPvpRrdKbP6
1qatb6n0J2Hhkxkwjv5+OI7j/Nh22hEyObjluIsWHiA1TxYqp0t4khJDbDKKLVGLp7PGyhEVyzu5
Ua83N+dSnLmPQ1bomU7mXUYf1IevUy7Ufa15/nbuxAOwi3pOx1Hn1XqxoKyl0pa2TafL6RRXuKsJ
cvXmQNf10nkCGh/9hdhnpR/Du4PFJ//nRMAUsSiAZ6WErhEuQyE0+nxmmvnw5XcEZRqeuoClnhwZ
nXIdNcPJj+McXDvnooY2MqYUUDFy9DRdCs6q+sCjz+jqUPgFKpMOkcBw0alEMptrvRSbPHoJaFDh
my+hIQ9JzXQTx059ef6nwSFJ77vN+EvWO1UtECAtzaBJyb1RkbWAVGtGyxg1YJaPpHmJV4xm1XUc
3n5/9UUafuKO6vN7b5+mgNEM80FKmINuoQpc1lXI+gS4StiYyQ5k9JSl2fUOUP28sSfsQDsjSq27
x0nUGtGou+1WbJ93SXgieb+luN4kxl55lyl6pcdqHxaZcu4rv8vz/H6Ku0l0ba/779p2jgQgk0OK
C0hSEDSm8y7xpZrs5z2LfFjNLO3Y76Ico752YHEz94nde9/lESnz7e1BT7UH1L3uDzXjf+AemvFf
FKImhMjzytS+OHvYfxKat1Xl2+Aj0vCFLmDkyAZZ1/Roy2iGDTExb+S8HXmtjA7xCEtTA4mqjHPo
bxpdb9VZ2hdSmd4ym5Jk3+VqJenmfRrqLCWZgYLKrOycE7Df8b3vU87pZP4vJiX50eDrMZgGyKQ6
74zAuKuatukRkoiStRVJ3wXUgwv2DviONl5lgya9MabWMKU/L6Cl2l1nbMdZh1gp6y4xtqRvsncX
p6fLX1gLCTfm8bi9oMxQizm7fS/0sPyap4+qxqdLOV9wJTDx+DLLqQcHUtiC4BE5H5StimIS7KNy
w3G0x82gQrhYXzPRC+RP3IMWYjLZba3RutZ5m00riCEaEVjQUTnKwgbdqFXC/BGLrw8f8Xbqr+GE
RgZqcIX6KUh+0DFU4qLosrPzxSrUpoJkn81XT1AaBesxjU1uEXh8ytCS1OMfrPQCuvLnnMUUxwGS
vBaoK9cjfcePbxXZ8MKdEbpbzcyrJdsUoGeVS5mT4DkXwxWfE8xDRqRhiU5Jb44V5TkqccLkFxMR
/BfAVRq7g9ULUrkRGLw5blQ0ukBR17JG0Zp4JKo/IgxSoGAoN+JdpdrqwF9DWrG/uTEBMO43wnd0
ML/IjrfiDfqr+6QbE7FxUVjVM20BAK6A9EaA3R85C1kSfo8VYtRE8ys4HIsqo2jdNxyVfFr3EOsr
vkwkkGdH75113uw2AqHcARkQSOgvLmx/HWcvn0LxksW9WXfV3e5wXyglEpjpgZnO7vyUPwTK2QLp
BDKzuOGVkBGmN+Kgmt0Sh8+eb7SjQ45vjTjXXI2P72x55kVmzt9ouJDo7pdf9NgsuD1MyO1NcN7x
3S2PdX9gG4TFYjldNPeStb4hPRlfVdPWEkcdMW3R3wrRAsg15KX56HujCtDidURuhN4gG6cCXmea
hllbmK6fQHJRev+H6LPUg7drnAXSMutuAch07M84h77H73rLeAzx2M9JIDIneDG0NGaC7XcPgrf4
fj7a4fUOCOU6PcSp9+0pEHa58GAgjhQIwSsdB9qWlx6wOuyAb9GrMM1svmoM/XnAppY1LRaIRU22
oebNM4oDxUwEwzyeyWdNukpKqrTSTwpB6XHTPUa7CkuNMukmyDYShM8DyC+PDarUJD59e4QIo2Rw
70ZJq5xtAQC1PadG+3FUzxECClbyBs+OeHuf5ZIjI83tK+vD3f8xqNq4S0MBEMaxTLDwWNkusj1Y
T1wtod7I9wB3ZtWkP94vKmvC7yjegykQz+BO6Vr9eUc7e4tUKsv0rXS2vjSOqEmFzTBkHXD5Efye
FyghXmHwL/QCEiK+GU3YlaEessS98BhVzYQ9KcL2PshwOyopHXE7x/a/t+hIWvkvWjdu/+o5RZwq
KyuIL4rK/mFoj1PC2ifJJ1LrF5pcai/yKNbrIAUoZGiFZRXsX6uWrjitddCIAh6PKwLkHQmq6uVL
Xl0Ydk5XWkxEURbN9u+vkkOSTJcjzkjCmycZl/oIwUlMBflU5YV/f8kwPHT3yfB6sLhvkZJGg7N9
rLgGRj3vzEuBhmjfvQahvZ3InD8ekAfDFxSQqoc5pLM1enQu8kbvizHkTtd65D3xKm0BdgRCVw7q
mrcx+iu0N2YvMvxu2IOt0U3wreSFYG3XpROlc2H5tcIfUtDEZ+C4lSIDkjDu4OFw3LGt8ZuzxMTg
1i/5+9Oqcz2y2NHLCqrxUP8HTVwtYRqtL0yNfF5pKx1Fc8I2uNsb6ECHRy4ADKmeydyYDc9e2vpJ
WnKCYh/BG4uRreVL9Ug8Q3GOZE2jwMgLnZ5Lu8hy4jaKyMReyCmEVBbiBqrHsktWNiTQu4ZQGMCc
t3iWm4WoJDgl8ePSUXLcHWkzdMFyUI6eZ+YTH3dD0N2/H5z2ja7mg/ut7Jp28/MEVc9EJeykN48B
Lc/t+ERwE6OkAOOPaCf3XGKEvrnoW4tr7Xjq4WCVQ9bqtO4ulS0y9qkl4OQYlEm6o55Nf0BQJ8/9
s1YqEiZHLqnWyqoNNSE76VPLKjiFL+SyKMPKoc655djdDqDVrdyT9r5FegnlnTBo4985qXZ3cdRc
V3VczxP0oxRBOa8SnnV/J645yFQnHudJvTn0hUT0D30PZIF14lmxyZrBfi65C3y0vnnizvBiDd4e
wXFiynzZwIvDBYstsIllLegSBVgGny8t/W16q7gMFW7TFkNpsGgdt8w8tDFE7QjLsFARHpmn4Hu9
eHA8AzEW9NqwLSRzM8aG0THryUa45Rtef7klafL3+R7Z6pEreXvWGBONA8Fe+qG2DvrlJMxpf0ET
ZT/8mdHNs284jOqUjSBjbihrcTSFiaWSbGYUsh4cEQ+UGMf17+jcnDh3Q3QATaKxyM6Z3rYQ+1/x
lCL5H4euFN7WNGgkPThunwntgZe+04+fy8jPQU2mHIBVig9uKB4VIs5n6GcKY1WEkch5ENXjJEsS
rpwhKDmRujcaxkaRB3DVOf/NYplFGApvpeBgQKunXQtsIohlwQiRDG4CAb0UO9CUBUddlEOkMF97
6SKQYRa1+Q3KAFCt2+9cWIsbFSH+dGxInrgMO/gIVnkRgcznwD5EACtAodHptFNiTzlcHetDm16c
0vSUJMjaqSsvhPkXTpefP/3Gkpvv7BfrGylTRCO0j/ciUrggLZZ/xiIvL2LI0Eb513qLYFUkH9hA
chh9V9pK7as1uFTc0PU8h+EFTvrFqzMFqYhzQ4oHyinVJ29sE42JHFFA1MjmFSmyNXyS7/Fqr0tv
ARD753GbeP4OGGgh1mGu2pfDXiOt5yr7cexDY6k7muJsnaTKn8cIb98dTtNGCz8geSLcZ52LRqbc
W6IOB/0STlI0jFtTzA8gKCmQlX8aYfP620l/MQThtqOsywzxcsr3zSNSr5gQ5tdXLKC/vtE3g3zR
qymWu4mEpq+k/s3fpY3KDTV+yezm7ahIVxrUjXNOI87f2qtzkzkv3YAC9pIfoxtdi7JXAbCbAVOP
UOSref1FpOdec9Og+eA+A1PKBmLdymEDvb6aqkF4PVytPjX5TyIX0HtN0gER0t6r0xY0L+DfAEM3
FgZa2tU3btxHpkrBP3Igg2B57Rof7ww4m14ngs4uMdoPFV4Al4agmY29NorneYG1/3XyV25EhpFR
/xFws/ECPiXNZkX8ZRgFwktT4MOZXCsnAbug5DbKOoxmi4wIp2Cd8uJsqr+b1TgKYm/FuZDD5wcM
NxwqHsD0YMX2Lg4HjShe4OcA0BjOKlS1huNXjQzAnZAFn9m4YT786LiNGMv6BrH3DJhZoBInzzIu
LrWZ53vGy/flzWJuGzBX50EOtpg+TC9TUF6v+NyIdfpi2mxyVGVMyDrRaJ8123Ta/k47HYFBpQN/
A9GwKIZht/FzfBCj3ycSV1ROPyF1P7YHbo3Y6BJJVf4QdvJAVMjHskfXBIutxi/rBwR3qBy/wHux
NRAU23E0T+G4xwokeYHCQNppUwgVUYxe/QOvf24rpwgrEWLRz3oavOfPWM1dG/kjC3Of+bskAUgj
/0sj65KKS+R01sNzLYub6x13qD+bdX85fkolu/2VImT2bBAJO7Kp52zkxrnQ1YwLZTeyQtHYwcfa
scBb9n7p8mjSspoByqb5VnsFxY4mT6J3sqEEW7WaBKROChRGkENRKX7ZX03QlJ9YDEthZkW4Yoie
boSqVUxVA+ZpHq94CPDuwMPy+EDlU/w6UTtNZtZiEB0kUoICL44AYlLk8/qPMOi9FSnSrI6i3uRs
OdqXbRs6zFQ/6BiAQQbhgEBBRmKtrpBkgi8GrG1JmicddsYTNN7rMEB2oJm+tXqQ8UAbTTy0UhFl
8Z+oY8GyYggznstRHoc8B/wVYsHG4QmZwDKZ8ze4pIXHo1ZnXftKCfQmogyr040wKQ6Ol/uF1THe
Zbs4+dARIhNJbvBkCiHRHV8DPf8bU3MCPpBlpMUQCqqwm1CcpfFltmXjqb/CDHKPLhaODcnGUqMf
S5UyQgW2DVV2pLwO67Cv0xlT+VMgQvK5tPVwWVatcJTBJ0nFKDzCPL67+OyE4gXM1jo0cIBkXGGD
QM+CVAZwKEaXdHfcJ8CTbJXQizbfNEa90Ow7GN60a8Qf91gU4qI1U3TB702AMspi1Th0X4F4iZZ+
xfqsGFxeT78EanhTuJMPEbzwDjm9c9QsNjlW/1wd86+59gqjBhxNDPYzzozyzotARQfpxi7EpiO8
lK+lSCvWI4gPvgW5Q/LEg+ifxp547qk3lWI7ib8wZ+09uxtAphPcc7tWWrjhGNWTfLK3uG6ROqia
NCLLqzsorauc4aC3hMsIfv+kg/OoqOkmqElFITlPPxH3YvN6tIF5uLjcFeCmZ67nlAGASqmS5TgV
M5h7hu19rWriKNVZKdyLJlCmUcj8mkGwdU4FzIMpHkAvuRhwftsCMolLMJNk0c4gPh2SIpc+ITw8
69oxwZHH1WFf69bC7sgmAVkarfa1X7A4wjDsyv+7JoxYV7LnNsJs2sc1Lh++r7ek9Wea6al/NCQi
/XKNEumajQyQdMSC/ZtgrSWE7e2v4nsJhVuMlbaDT8sArWsy441EalgyA1g34ByHKWVtStaF6CmA
QbR+xg0AK3l5emDB6MqjHb7oXfJCCRTMVLtuB6Y3LVL3Dki54KyhklyZNpjQSufq2s9dmbSkfFtT
EKLEtiZTrYyANjnk5KrJh9koCizhx2m4/F2YpG4RgTZuMrM1KkzLhDvHUTqse3/3tjonmxju+t+g
4uSkyMJbiCFyypqy775CajxanRNrQ6dr+BaB4ZH36V2/OewUPaMgFafZsCgC2MSZJc9JutrYLNYn
Oq5XywDNYUNRQ5q5Ba9RYQ75n+QeRdOWXdvzD6KDmiFaR+GcFB+4R6ui5kUIh+PUlP48yqlTPGej
Qjf1HH+OhUZaGOejlmk76pHQkmslkmPsPP/fZLjhTgIQgs9TggCWvn19BpYfuZWxMhGGg+Nwo0XU
DM5AdWzl6tyNPTP5eXOsGdDNgzanHki0r+ll+lhdXcVMFX3hPEfrW1Gp9jHplzlgw2LS+SE2kTci
V2hn12SUICTiAuCdmo6fpDka7ugzP2gSsrjG7JJ9a9q8ltBqdK/8PmZuuXMV5C5UAf5K43tMr+yE
Q8ExAWOF4UD/5Owi1dXc5S7KHQ/7MTrEpItcXksbiGAYLpnURaTFZQXXmLB4UPEr3lP55c1hm/XC
lLs/Sfs7YW/LOk1BqrDCVm/Ryy5xpSI2Q1eGmMSiJV/CRuW8/Y7NyZvqL6XM/adS42Vl62lHwrpi
Y+x1QMAaFQ+B2FdKeCAdjW6yWG/AnPuc4gKISXcdsbHsPZ6G1MEcGseQ0MaTfySe+cTzY8tcDTC9
sc89MuL6UZZFGbiWldDCkoZ/LUKTrp0n/WsmQv4GXa26Ws3NPHbamxjYaJ6ZOlgTO4w5e7S6+SyN
xA0u7yOsJT1kiISLEVqzC9ZG8wax+R/vyWYHLXCJzA006QfdbRK5EXIWor3xaAR5EYGIqW8gAqhI
N/q+4eF/Kv8GoXBR/wPdE7+0LB/0l9NpG7LCDANvkTnkLw2Bds46tCS5Oe5A4ddyyvGqn1nTG78z
/8ll0u0FidSt5n240sj+9qJSvVsNixeyDZOv6gq/oS81T6IhI9PikLcb5IBODnWD3/rbUynmX9NP
M/ITWhUc3nzH6TEV3r8dXqYBMJxWoKQ+JutQtIZdEt/o6CsHJKWbBEpJJOplbVkP68y4lIXYi7X9
5OwWN2/jf56GLnRfEZsdudLVhpw7lJ36yGD48R12sY3kO3v5Lh3WWx2qy1auhZpo3uNqxinsWC3B
dFqUjFFxFestEBjiPeMlNNzgm7LUsJL0y8LzQAvzZRaC2mJfnVgG5j3TLNTJdcmgVScrskP9I9uT
p5cf7GZFZf+AjoMUhnCB55Q4WSKELBMk7PvGJR5HruoT1ZLws8z8wl7tfXLCg6Twn93Yc0gtGPRj
aKe/BFeDlYXK5Vgaixi2cJJNLRq/O0mKoh2Yp2/I3632++pALRk5yUIdY/VBcX84LSh2FeSIeKdz
0riix5qLbIoeu05NzH5hVGlWWBji6JK8sXmG4poRyarK590QX8q/AZcAoEGF2o2w1iN/mHzrfbWG
U8U+JSXl6dlufuu2wGOb3PCvSFHtG3jo5dAar+v1dgT3oJ04/jkO+u/hEMt26KWmgOzNHwb+K3kO
mIFFDPbIOeD6AK9VvWONJuGCCe6yvGWQErW0GAzHPZiL92TQ9WodUZWwE67e28dXSjddojOOYzvO
HNkOPc4EkOmQvM2M6cLWPMPL8b1B1eSPfsecIj2LNPnL1/mvVRABnIhBUmL3r94if77+hh5i7SMQ
CeSalTWpSKIQlZu9Fn8zOWkdfXMzeo9+DNlYqU8gMWmmQmPwdxT9xsceT5fsC1z7cSrYv4dZCuK2
QGBgNugRQdMNHFVSXQwCxeSPQhsFp+qGVL+LDAcDTNI/8UmAmtId5gQe+effFWC2OftK4hBhK4d5
T8XjOH7owNWFS5oyGBna+r9RK3cN1suwyw9vsaQC6RBGANmC/4D/izQUhPVBRrBa/O1gPclNkvEK
mZ2Dyz0/EOdyCv7yN97FuC+V1jbxKL/TI0meqhpCR5x0DTUxvt0CMeZAU6CitOYErxRrOir16rNg
ElI9td5I5i2byuZm+bL0EZJwIH6K+4+8ZxbPIbg8TV/DXhcvlG8hWAf6oV8XXDH10427NAyKlB/Z
HiWbJzZeCos+WIZDGhboy7HllTU7Szdkuh7qJDO4bi5t6fZpSdP1SmLHx5z5LXdAUozTVu3F2SQC
QtPf/T7JJtySLmFes3KW2ewK/9P2EbMdUlIjBHFa9kis+SchKdZe6zRxgKgw8iDgTivM4BQFtvtf
TEvI4fkHnD5/nWIvAcQ7o7gl1WJiJ3PmiUMh7kDS/IfpuAdnuSo4l8JtVdEgKCvFo+QfKR3n9pS5
qBvLu0zJLZ7Cn2LP3STlRDXYx73eJisr/U8cQUM0O2/9ruVGq3D9CkUKXp6moGQLdOSXJW/xNDIc
DUIlYOhJWkyv+kOC6Ke4WT33OvdYpu4ytL+v15d13F/hvup17EqJzhEN89vkwIF5Jzqz7eWEJww+
hO0y0SWwolawpafvnUUCuHxwSVeFBcqy4jvY4ehSKb4DKvnawQ/fsZp6n4VRTIjz1TeSp9ipR4Mw
0nI81QOVPEb312+PXhHa0X1/aLXwHyqP0XzsG+u++cobweToMdfdpneBj7nkGMs7sP7ZlR5KHwQ0
FEzSyST+cHmBu5iFN2kQWdEuTB/Li8cTaXkHL8l3dS/uLF9/zyIVE/2JK2h0OZ8Q72QAfLT1hKFl
KgnjbsdRGFbP2li2Hkq5YAyJGAZtZy9UJ/We8i9y5zeEmMT2VWk7+E/Mggz1H/5h4I5P4o/3ezfv
nHiJ7KnUog3Lr6e+GKB3VVEF6ZEVtHQw4fYYNzKUQcAKla6Bzh7tzuJkDc33JFMTEJu1SYISbKSR
Ib00MVOeydIXtK+DyitT2gLMmIOuPbXmZWXlvzJScIYOLWMKIhzzS36oNSjHUWGngkgBrieqcPkH
hqdiHAOIVL9kaecWVXYl3Gk8B4vu0Rteg7Day7PXit5fLX9sd1hlfFqw+CMYk7uKY58qD3HlpHkn
dcuCxfoq+jZug82JjrE9alHJySGLkdRXChlGSfmgUMuTmfWh6TzQ74MXZRHYuSDJyMPhzLH0MqLp
3JhYpIBWcYkj7uyNy8jDRQU1LJBnAUd6g14TxkPh80SNarmVNLYmczRdSk40uVWOSlRGb39HB7ZB
kPeSshMRXLaAOp9/SgOIjy2PDmCY/8d/iuMOcI2CFCq995VbjmIV+0H+eMZNjmy7Rt4LrCL812JQ
t4E6H1aEeGigTpEHN0ZvkP5e6+G+muD8BTtiB7m8Ymwh+8703NQQSJ1zrnLfIrsgcEO/1Iccw1sC
bKHk1ekRlZE56IUtiJxu7t8jZKpV3qm8eQ6+eF+zt4X1YQIXbqQYxVDaG17yDsO5KShCivRATfzm
260y/IzcOnm2oq5jPdmFayyvKprSh4+RCKIFGz03fc6m9ZZI2414WAAut8F8tNHxqIsr5C0oVl/A
s8XyuTBnmJePCQesL4KZ3H59X44yF9FJlMSllV9LijdeFojTwBm3WdSK6BmvmS7kqOpY/EvmTuH5
jTuJS1SXRPGWTc9vdkFEVf0oSq4h6o/dUR+5xwZEILiwG5GB6VYkiUKzRT62KcpX+YbCVZVm5hyd
VWwH1Sd8pHqljskykZm8PwB58t750BO3qgDQB+MkeTT43+XficHCqAtvHMFQ29XTG8pL853NZWsc
NsR7YoyOk+gwYi91qUg5ldP0rBthHNf7bV1EIXU7V7pUMW9Kt7l9nsrjxoIU7wfLeMmOb/BwDQ3O
7CWlnFm/X6zz7D+H1WOSRAwmpw4zcWajtIbT62Xcc/yHRULyO379Tey50ai9q8fYo1NDOKWt40Yd
3XDjxDxta30vhZ+vlOrBMkSodQbiXA/s65fY8PASaF0vRjiz+6R+XqeZtmd5UwLs2tUD/0012O6j
SWvMWZvvtuWbAG2Qe+bNxuFrfOgNhNC+QENxKiZQ+g/XukkDNAWuAuv3qPLUaTuE35S1PgoxImMj
2E3IrShyvJu8sSDthbpcgHBJuCIEogIaO/psBOIDnh6+cRUh7zHr5zBfpN2W3nerUg24cCzDNTbA
Ci6ZSmgYBTafxUPuyxWgoQRJ+od+TcHptUuRiKmFYpI4y0ygknR1L2Q+aaYUYRM1fsbG5aDShg44
4GgvfPY64Evbmr2FZArVcxgC4aigOIu7tTC9LbPzuB3M4nxLUsHALCIbQxFp/ilFVJjKq+EeCbif
2mNQYj78phBvmN0JEV/OAwgGHZ03appApXi2/sWUjqKDcCoUyXRIowbzvuGx5bd551EeRt0Zq6/t
CYRa8rIGio0edEaZnZlJTWIbgSrraf4M6AoVoEdWLwavWXa3jstF4xt1P2a4YimeFEDK3nqu1wH/
2rLYchX9uKzaNE1h4/tYFKuvznrtGiJrxvjI3d2RRF4rmQXo2Fd36FPnHqU1vmtOQPL48HLcoA4Y
9HiaDoHtbbO+2+lk0mRyvWBZ/nXwbTU3hv5yFyZyQQSdFUv95lTrOHSK8xxYO3IbeCmQlZrSTbG8
A9vppMwpMv/hExUd66SvspHjNe45gocIRi112uArLvvjn6Pe15/W3jVh+9EpSwdRjfQmsNzyYiZj
D+0jFircTpt39GgshOwz9y+nvRHRtqKgbsvSSmx1e12za9L1+MDjw6IHrjFaBVdxksh1g1EVG530
BslZLOp+iS/gL1hEuW+d70I+OMcrTesmv3g3ePswapWSDuaJtABHZW1h4VOEZDisx6I1qFT3fg5a
dvOeYMvhOpIg+0HtUegqGiPz1UBKIR4y4STKc3hsDYrTBX7iaVCtw7fV4+MT5JnAO/+thojw/hBo
6Fj1Z0Ya2ybxVmVf0AWpFolAbO8mC/4Txe6pBRfXA1yKK6vQJavakp//aaB73QpFs3d5xgeV3hhP
USabD0NbBwhIzALzf/zbLw81og4iVcCj2RyZStyuDpiIyyUksCTu6D8DnkBYtb+w4iokFQAlwEiS
NT35dVqTshOF//gAzPA8av+Fje7eTocMXIJucbqXTx67FIb9Hcyu0EWjefA+MqnEmbkvzAbcBEKh
3llY8PA5higQQumaD66cjN3RDdTPQef2X+dIk74NlhMsbQLt/9oxCOll7fV4uRyYjU5NDDOWDO5G
MLfuHKSvsXmTa5wATF+k3pRIP4RMbqpPOKitbnRPOApkXm1hemYI93Z/YIfkkvLbMyRCZtClZIix
uqLpGDvqOfI58Nl851vjFatVq9YiV/nXebDsepb38xf716r4m4LUPvSL213oZMltIZtgjk88YUBM
fQeTbIWoOLbtTFUqBXelktt4s3IlvGXP5dBFrij/6EFEVoblph2Rm+aWs+2fyJPCnNTwI3G65TVB
DqtxdXG73qqdrL8NYCClaJSjiOeqa/Hz5g0yiOIEDwmNjEg+3IV+cizLXxWK9wRqMzkMFR6wEHp8
Sc82VJOEIo+7axp3mU7F078Rrx94KaNw6VsRzZ1ZRKB9gj3X7DAnHuq8zNzl5mytByAulem7B82f
J44A2ZEIACQQviHjF8swXaUH4sNMsfctJ3uQ1xZFQx1qcNdAfKXywtGqXExjTM1OKuEbkguXoGZ4
gns75Zo3x69RaW/DlxG8VTauVQZmxKnJ6He+axoSxCOD/LMaVz6R+JaGbr9egCgk2gEV4BVuGEVv
YEEqV+HjY1u2Q0eQp1NUhrbE4vHItHaD7xtgto+6knxWHRdUSTfpazqsM9PusDsrUQt72M39247O
eBwto7TljrijKAZE4j3WlrW5hu5zUGuK/Z+ky+Ovrc3aAU2lAjY1AEu2x9PCM0YKIESttiVbFiy2
lYl2UFAF1QXZMnPc0i5dv8ZEF3UjUNf7b9ZqhbsuR+bDXDrY/aFl91Csw9BjMKiicXu/UdP5/rJF
tJ85KRnO9hORi3V7vP50sx7B1UkGltPXUUv5VQh9LPtEZ+43EuomWgf0xMqlLBkcpENU5iswdDZ5
VeDcXETVC0A8essPJu0bYsLNhRyNxonMlZy+YNdoFaYnxYXigcc8xwNr+LH68SvBaypFNK+j02oM
b9S34RnpFuj9okWwRqpO6pWlsnQe4fadnkiuV3mOP8O7iGkh6LZiznSr8AN0TY46HV9Yc1oWl4km
Oc017hbbtDbAtmaodRBOP+exfVbGgV2hznQmC8o386eZN2rOG71fIvf2XtCdW04hBIz1wm0dehse
rP5Ld/+YehDV3uk08MagQ24J9uIVj23OhJYI+CXB/hc29HcdsPBdu6QAZlgTNKUAuXQJOumwiIxr
hjdD/NpLUrGN/fv6c4ic41rLFgrhjiqFu18enhfHQHffCyNfmftFVdPOZc0JXtWujRYBjKKS8Xpd
QjA//CprMaGYj/baGJ96NcWS1E9SfYOmWCNVSHQK0xQ5nDE4ffUlg2j/zSyROfQkxxF1ol/kguAQ
yXGTMQDmUG2qJg/De4V+iml35fnNYwXZaV3Xv62QIzmUA2qPRe7kkVqEf14X2gZL9F7LwM3XijuX
562x6bwLdoLfJdlO4nAhcRiPmiOQiuxvBK/O9O6wC47FHK8rAOdoCUiYx/DlH0uuT831TbZab18n
eqe/ppypOKIUhbYSn5pbH6lX6ni2qr5IKqMtWFrg3wi0rMqICPataJCp6jdKH3fFEQcm0IerKI5l
YhPzlBmns7tbsy01AqpQt9yxrXjdPy7BeaxlAt6TwLY2bVnO9Kyir6iv28zFnhoPM1jPIhTXpvfM
zVRPVLv69eptNaL3Yme7naQIuCERyOaZ6e2d3+nfnuDkqu7Y+fVWCloU1JFmaHvqFWQ5rj16Zcrk
8uhAKPeiC+P6MGUfk5EaO93KEPFPKcsL76SLqqHyESdGHukSElnwredx6zHlxp1OOskobJmPuDcx
IyiVUvoGHOFOO+7lD5fn6+druulqFe2WTG+nNlYEw87kQHOMBOAy7w1uL5wyconwSGgHBLRvWhD2
QvPSazGT8MEaotFUEL3i1w78Y525HkZpWEv+RIBWivj2UimQsa8ixOPdTCGpw+qsQOhPWK28D3ge
ywJOaBqmnMriVGrHEPwGbbhClBYqJ977EZy88r+MAH74ZRy1rLzY8uy43q2iArlyJ0keKxs8kAjL
bP6W0hIdusdGA832w+KNtNUo2xOnFCDdCNeoSjenhDZTy9zQLvHSotAH0L4Ffnr8F7f2jmKKb3jn
wnNZJO9ksM9GmfvpDZqFAYGKpBgGRY6nm1W9U+giP6Kxpppn9SG5fXxYiUNAOrKUlGy+SrYEtbJh
TiHGify/G4Em3Zgcd0nMDc5Z86nPpyvOY1T8wp982cGq9l4xNBa+UI1mExMoIg7TDBsbhRzh6J10
nNsd7JUi899hOVf05R/5VCw4i5bTIo3fqd4HnNwcfDqbLvQaAbI4/Gdj4IXpUPwUDpaF62f/Njt8
2+jbIBsyqetUWgG6lWfyYU1EkASWeLhTV21DMfvPBrQb56koUYFCP829L241O7EGZ7SK2Ax/PRYz
Sgd+42UQ/JDrCPFMgAmJSR8b+WTb5sIDcADRDqtLZqnZBSJ9AvTH1Vyh0BTg2KKzy4FtUouTo+5A
bb14+XMyaztRYQwt0c8XABWhfV6LBDLnXtgRCwf7IqG4AagklRlCvOlv3t2a6CsqOWty+hGuwcd7
QyuToXvmYo/GUeR9BszD+qBqG0NUamVjMg3cyiow8jNR+zAgnyRsKZYocQy4YBrGzr9fZBclq6MO
McVLfa6bTGMSIYa7wZ6SnQJ7czBVpZQ+DYzas+DlVd+vYJVjQlIishDyTJtIITUEqdEvsNYdVqco
bhzIbaLHmmf5B6cFi9+b2IOE3IoDjhU/f1V0wvX0iysb9GJjp13m4JwyGu9M455KAdeaj3EwfyPV
usKkw3ypm1YuhyqKA3HL6y1Y2EQqqJV3IJGHvsHLzwKfRTcaaOkTddet9feIdJWzW/BsIiPH99ct
3eaXYautgCbD5R5NYwXCxINnZyCQPv4YcMJPXmJoFH0uUdWKJxSAU0Ml8NsIl5Se6WfOm9InyWAJ
rmmQkyvhU9RHBSCmD6a7yYykfdBxn4fnKOfzVglvEfVPuyFToeELLXQoTjZ7h8EZ78fziy4eJ63X
pNVTbl5DSIZQOWN4cvDyVTV3KftbmFyKdosqu6zOWQPpEhenbG9iXW1fjnCD+LKV4NMoOdaQ4Ght
U2juhrzkuwDnscs4UB2hym28HhOn7za9xtJ99hFW+FzwAFH5JSlQ1NcEXMiOamgi52ATi5j1A2Ko
rPndHu9HOkoztyNXNU+JLBlox1d2DVpAJkHnKQvZKzxTwMbzZQMumIhJ9qtNzTlPNIn86XC8Hscy
54vmGqhXMVlex863VMBp2v34rHSQwRQXJ41wCGc4Rao/IPxmk4mqd0jzs3kiqAaKcUC3HUSho182
xpWKMCK5JBFGThjJ0beh3hE1p3S8p67RbTChxR81yTyPqhZsQyeAaqRuTOXhRdSpgZC+lTZxynyu
vP0aM3P+vgeGeJxPLq0p3V6kZh13EzglLpewA0q7riyqMoBSUHEkBwwK0KV/OrnZv5yM6TLn0f33
Li/olcBPyiRYoBYEYVO6WKWGvRFBuV7bpzNqr7c9XnoI7LFQZI6mbHlDsu97h4SqYWKjYCqjpANB
EjbgWOs4aX9i5CFRM0AwV1j9CGVVc6JTBD6k2ooPCnBhhpkZDdpABIPqKFgX3XSGCXjOVa6Guegj
hBuyG9mnzLmbcGGkVtdDNaflFtCPBbv0g+vWe1N0Z7BXi41DZJHIxPS8/Eaj5rPRO/PzYgJnOuMo
OaxzZMcjoP7LjYWev/6JsNvzzPfOJg6Kju8+Jm8HUGlz5HYNx2qN7ZedZkLth00b3ENsBywFaxRW
rujHDKl5zqo8QXj6S/V68Aupy9YjLIby6xmTLU8gmgeu2aQz6AvFinBb+AwE4HtaSQeZIIDBdtRq
hQymj9ulG2un3FbZ6j47OBz98UCXLU07m6HgKpOhHZRheF7atiunZaq+AKe2NoWReV2WF9S9rl49
1VNjZ0RWQFXdyQD/2mGOFwBq0Kkt6sqkxdNhsL0VUafS3dshIYphKLNH7wzzy39fZaJuVmh4Qz6i
r3uGIlnHKUoKCtgoCZCdJ5gZoRNoeMEbqcaMqN/T6Rrh+uA3d5zIb2I13s0Qr2p7oBMUyG2JXSK3
sx5jcSI3GAq/ZofwiS6qZOZkzQwPK0Vw1T3jro8rn4JV6URoKAo1Vd187EzXbyFjeL+ImIuQserS
XkKycGb014TaZkDNPPHPJCjXN3vesehz+7M83db4fg2cgZI6NlfSGoUX6xWxZ5ZYBcnbQUYZsmfl
wxMcQBf6q0f/CiVjUpPXP4SOHKevJcoA8eylocq0QD8rkxsguZ9LX01tBLpSKC1w4YMZWnLeoS/E
RogDs2MFD7RgikKcoIBZQqkjYCga6zUez5pN9V3nOBrk9+qycsTddCUwH1FV5CclmxpHvdHTMGtE
0yag5uy44YLaekxyjCLuceB7oYD/kJL5l2ZvwSu5xGaAaQTCjZWGztX7FTY70NMyuIhyw+Q9N4NS
G386MAi5d3y+IcEti0XT6hK/dSr1MXuYDXD0iVtcK4+6HZUICnxobTHORt5P2G1f0sgUBaK6lZjZ
n88kZze56xl7JiCiPQ23pk61+3krolQeFX7gT4BFLaDj8/j2ZoZflwxxz0ogM+upV7lXwSxkQxEr
MUVZpNa2tufZqIKXamp3aZJbI3WhqBVPoVeZ0HFvwdU37MtTYfyp0np11uGC0zZu9HoLib2tATCy
g0toopkeyT8hziCTDEZhZ18Pgu3lG1vtsPNgF+SHHd6uYSL7nXS8aa91gcLnSg2zQn1hRHiXjmAJ
rq3Y4H6SGYtRT0fzhLZTmzerrUD60MxnrpNglBY6MkuKHbUVrKUjd+bXZr6yH49JyGh5eswTuzR/
3gHjdvOWdyRgHPKP7rMpNXIeImip9H1zIQ/ee62ZrARxTFX76Ig94DzJStdOCYSXj9jGVIl13Iag
UL3ILGanwZBwPYburbKSNuXASBNEurMR/sxQcrtAjRdPGIEYhspMhX1exV4bmdv828eCbBcZyF1H
vs+XsURwdtVpfChnMLAHV/+3uUdRjja4WJ/o1iP1gV268yONUuPm9w4qahHU7A78uNtWfn78Hm4V
Ql/fiDPMQmTvo5KCyDhYnUv9Q+fCfv8I8r7IVDu5Ntp7u1mBLhFEa4VttCf5U4XhCs3AoS8qjxaT
nHaQmpvkS5KE+MyerPcRW+nZY4p1XJIF9pt7nvVF4H5mzH1QObg1ohU7BVFPzUR7QHZzrN5Juh88
z2nxYK4X2M9qBCZ/tfklIfHaDtgUlKGz0jMdeC82hecMHXJvh95iNHTTSOZqncNMK2XRCILfYUmd
DPuq2M9UPvE+kAz7yClG8oUv/kMRTfWLMcD5u/8FHB79T9CRB4uMRCCi0krHFvRnLWF8tLmAvwG0
OMHCVSBnz7t4FJBad1LtsqoikGxq1C9gE4QSyX0fv+9XIu7X88UizbZAAM5GzVc0D0CWnJXadfU8
KXqliGKhUNOzrWHrpJK7a8h2AAuw+DJ0nCbVTX58vfkDIBlrJWoxWvlV05e9GXt9fNvQ6cOc4P1Q
c7zaWu8iwjlgJpxUz+AsO1MU46pvbhUY/IwO8aqWOY8Jz7xkqUB7vCf0RljVVKo6qMv0dqFtZBZf
sl48lp/Pii6d+PsXVCdbSkgI6hqL4j3BkdbTackeyFUCu4udpJctLTyFUswjFH0N7i+h+go3nb0s
6IlJT3a66daYgE/bSV8ivreAGtQ8mzmjh4WfIjYeavJrX7dgvTaiDnfulsip9ggycwE/9z3dzbPd
Z5uYu7WglSgqfUdw5r4ydg+MtgvLSrNFut7vWiD+jLZfqkOn/vPAz9vDd0MnMgUvZEx/jFqZENkK
NfxrksoiJIsYh9NkrZGlnVw9ysK08djVJTdVeDYtL6e337IGnt0TrkboSr+wMYPziCg/zaEVxl9h
BId6QIejxtguuPb4hkTMrpBEgdWTJAH68oc2PtiIBSDGvWx4mqHO9xDvVfCd63YUb9qX66hW8A2f
K9wwm99Supu8ZWFWI+3BXCc8peI+JcKZLiKV59JS/n+PDaQNgp/pJ69JNUbP6rr2UcizWdtFP+oO
NjEyiHBfYqjS2LLatvTygCxytDxV/jl0+EIrgJDzz6lPbeUF7sQsd6B/TOicOtA2o7DKOWMy0U5u
RxvkpOW7FJ4shPVwza/Yd84Dfs35vaHUQaIFiTXi8viEgmcGWhwCHoR3VNLdtyozu6fIrQIqRDyc
2a20QkNqzhvTu9UfEQy0t8ekmrY6rwD9DQEbpG5d/YM20i6T+0G9VwNJuBC7X4Yrp0FCDjNaSPXr
ULRuD78rn8YsIsz++Gp7N6zP/+32cXZNsuE/SJ/NKrwA4+yP2OvEtvRsMH6RyP8X7TbnRnrZz+MA
0f/lQDbcLagfNDWpAJafV4nKh7JRYDz6YTgOCQfilcbk62u5hAZqOuExYpl6WgEmXO9yi0w4S7YZ
K9pNa+PhNLaUZ5wKfAlm3GC5nkf2PxOTJS33l/1t6ZV8ExpXK1c/HT2eS3AdrzKtqgVmiDMVUYWf
cUSvHjXLpU+lVZwJteImsfnL1rpUKb7ku0dI9GC90G93BNbjm0fuxTJtzASoK1oJ6Q6E985LjtcR
I64qaRaqYDjyRrkTkkaFhWl8UqTdsj6a4YT0SF01whIpQ3YsrTpifUF+ylZPGuu6834HZCVFWFm4
ZB7/Ofr+OoCsGwkU6TJVpodanANkw2khyQLmG03g5kvqkz1hZInonB96Lhh9+3Rb6DdrKzhxSTet
BmjdvRkFobiQfqefSIeY3OM2ID7MTzY5+afL/fIHBRPVtnKPVmKMaPzrkJJcEC9hu4hDgNDQXscC
Qwen4/64yge1vB775zKZh0RFvBEhFvRNcqzMg/jLVH0QY9Gg9qJT0D/nRe7qgHNMi7vP7dwXdxwc
4OUvkb9uZD/kv80DxUjDvRR3AbRWxkJyOkGBhW8RehYwbHjq3fJ5sOl2exeHWL7o1b3J/qFINkq+
e91JszBVNTGzBdwMeOE7BxYx2Lf3ub81/k+ilR+Ayx5+51BMXqpCFZ8yR60mIFFpoo9Hk6axY0y2
7sDknyBsYtvYw//38z5b2E/A9Gawe75eKYR86y/RtnKtRyyMqGjxMWU3AJ1CRZPhOncChU0WBsVm
jmeb5qVfNL4gg6jskzWKr448or3i/cbyU+xlohAiNFtKEUYhWunTXDGTh8k7MeTdTi5ka0wS0Q9C
8frA186wuU/FbkbwKCEr+9/HvQS54dM0IVhi6EoafLbbi4wJCeSWDUfePLUaAw7PRN2XG7usNrKs
kkztfXVfnfi8bP5vn/56N5vsxG/fdktVSoDbr8Of6tOwvlibb5UTYbogmwTZ3zdPKw9ypqIEqnnr
U+O1V8OL5D8Lrpmd7N9w44LVyk1/NUw6GTun1rGLD18yHHSWjkcN4nhI2JTsKBBxNLwUYSVOS1pd
8mmP8hvVA/8rP7XjybeLbbhWJc9eVwvMu2pXLN1ARPzUQeYB2uGlJxjY8Tob8joRYulyNmUJ8feP
H9gES2DzUWsky4zrA2NO2xNInki0QiqXxvkAc+lmIsRVgNUrwiwyp/2A4xSgupMwzmYz/E1HlSbt
U4upbnOvH8mW8XnnGwlcHh60DCzL/hPhIG6jBQCnFvLaG4iLcX7JM64qLYchiwuFfIsG/eK969Zv
884FYwYBWuKULs1G5S12miu/0VZNvzvh4oLp5DYFoMHWKQ2+G2UJNpGiFsoPgY7pNuV06TRRkFoG
8kgPxLj5cbQBKToZHIt6w7Mfox7xlUvN4BWXUoWmbK+g2wdx6BNt9hFLawFli9XpUM/edBoioiny
abrDkfnQUes5PttuKzL/JDX++eQsd1VoFTN0oHFqDz/dh3/46wKWpF9FMceKLxRzIj8D4RsiuZA2
weJHxJMVMTFbUt06JTGO7bdCDJ9s57CHrQROe74vstJgnvmEEuX+6YKeHAa+yEghszM1rJMqPAfy
HucTEBVaWDs5oggaovJdlDfdtVgXCA1nZAocqs7r4qCYRbBEsRpOogYXIsPtlQUzEnblisuqrdxy
K3E7jL3D2bF+P8JU1uTrd859/ocOPolgqVZJcIW4kCMnTA/UPaFUTXV2fU0Y6fsOv4wnLaNzxhuH
v7LNtiGofEx5GBB+eJXMa7NHJKXRDBhRWfY3/Obw99B64u+GuKLsysGEiF0FGdH6xxpN/T0QfLVR
n32abrO4vBxKj/NrGoiqOjPUFrRTeQqVJwm63vB5d2Hb+Cmf8KrUhoWQBcGOlF9nsmUeZQh089cD
ghk4py0jt7rJBk4LDH6p66oDSYhIaypws8Y/oPyT87PPWTtmregkid4IlwjP5cqZb1xxGLPfszAt
bxGdfjKh9UfdEAHLBHnXV+0hk9LkZlbXKAiLiIAeYv8toggKeZshIUQSyust4QzmacDIGwGTSIFE
c/nsjJV/FM1HrNuRHeV8pcRVXpBTPT5IFbyZviDMybewMWE9D/rsst84cIs60v2RRgBQJRllY76B
+jxWxssiy9yedbjpdbZdMIlINAJzjVJQN2gs5c1vHNl/lpe/bY1X6z/HlMNPvliIqSR8smm7+UZj
RYhro31/KeJhco2qO13LXm/7NrisfZPrXAs6khqE/69NsyST9QIoRsZvGqUO4CW42aZ+Xi5nAxRZ
8yfUtD1x+fnv2XaS3cy1m9na/TFQKEVvSke57cFawh399aeZJ9cSCxcm3ldHNXM7YZQbukWbOTnp
s0xsaqdaoChGiBk96dZ3+EZEHLGw+t1ATg36GrRzOXzGG+aFw9cGBrfs+Rcxi897wpoRf56yxlEI
HLiqiN0R54qU7wG5JZmBhmtM58RoCkLaPLzrZN+OEPcR7Mafs45Cc7lQV+fre6nU1vbAb3wPRERU
3Huvcsa6tamTKDlquSuMA2RqgczEqr+9dYXS+ahC54bQnodmF1ln6rHU/SE3/YgGz8CgnTQKmVaz
LYsfS2OeQB0ZAnrdb9cdtuTXyzvIHsgGL0GIDyfp2hA7OgjB4AZeojn8+uT7KkTSbU3XY1/AIZMU
f/FC88rYo2+eLC5VdYcOERc1BLU5DqYXVxc6+K/1f5DlENxzaBOfpSCYQxMZm4fOulflJIZaw3La
JXDghtJRm74dI9qPpfeI0Esgysc2TiNyaHAiJcV9B/nLxkGPRmD7bz2uD8gunEdGIf75Axxf9HUX
HWwxAeCa0UWh2S95MfLAePwVaYNYUVNFdP1I1JOYAY9bt5tqtv9fOXws3bx2K39fAukgszTPbM4Z
DEJ19KAG4O3u8m+yK8snV1TJiMDVEkiBS2zyI2lAxy1R9yt4ZRpVk3pW29z7TlITZCKEPZSSc2mm
BDXwl9KucUwTzrjyKWBQEzYk7sniJZtwyWZcNfVIppViccRfw+2lk19GhsQzgO8q0fk1K1yqySpY
9QREOP02AodOSa3p7VPt3VO9b4HQzmh11rFSX+5oakaPZtJh6FVNzMo5KJrl6DlnH9w1wIGoVVGi
08RcnTBR+Z+bBohLPC7rEB0igFLEErGd0/KAJkU+S7xXZuDEDyvP39zoeknzTFlArOwTIjPz+eho
JpRwNOuh8hNEB2XSJZqJIoFi30EcBt4z4K2nxgydqnbsqZEqmE3f+RTdKwg96g84Zt+/tZkuuTDR
B4wzVUOalfE26l8YHsJbMA2vBVAsRVD3g+NKQSPUJJixfkj/hVFIZEjQAJ/g4NMEH0t8v3W2E0ry
jwk2MS/RgmUCG2za9YLSBCEmnnAjtLd9QC5lGqIClVXSWzgkTnEtFRYd562Cotcn5NCg4WfvyM+z
mr1wGavx/zz/C+24OpfFeNpbK0j+kO7saKyHATewjnYAmDZXyLcHvD0LQpfCSDw673Pgu2oxTlfc
jL89o1hY/58vyZCe0M0wKDzTB8NcorcpihjcIqvMP7LMSW2TjejF3ovqR1nWwzY0yFlFuXk4sLaV
jpS185OWGjvFJzedioeBjLbEWlViFTyaYCtEs/gwgOp2b2Vgwf0nDbzXWD+V9OZyAkmgOvpOoIqV
4rAMgWJxmfesws5TxpTQvXqR8QEoA5k1plPrrJzNhwV/llpMWHaJBepdarsymbGxN/WyvQv9PZ6n
I6LhEsMf12kaSH4Yw5JdPK8am5qwwJ2TgJ3uHKvT5WFi+v79nNvQdWqtHuarGTU7IpAiIz/3Gh0r
E9/OLiKajS/I1WCFQwsLdSWvOZ3s9WdPEBhVjlQ9H/IZFKnuhKed4a2L4xcsQZBX27fXtPAjIMS/
MH90B2JYezJDpvoQJ2eEWhkFLJtON8DX/SYUeqzpSjSeZdw8bJvADwjHbOEoCsQq1ownOP8t0+tX
0d4bJdBc0ajK2r/6LE9dXNaVGgUsN/t43dxAo7JxuBz5GwYcC37j2lvZsvo2DoC6mX461b/1ZnFj
CT7gfP+QGrD27rRb1Qjv3Pstl88ORdTCXoqJHOhbPav/2BrZAdKNRQkiVaR/XkiNs/aLOVis+Vv/
nMglY702vN99nWP2wRWwu8wtSqE5WWi9dmfMnDDO3/Cn+b32CQUSYAEkNAhLiKgZl+cH8/WuxK+c
tgDS8cL3wza9Og33LsMqiXwvd1TRP7FIvQvqTcJTiKRlz/GEsPBaoC4au7WwXPtKbM4hqRtL8AWx
IxxZCQzyldky3Piy4Vb4PcL4DzbHhQQg2ey1YhdnKiZqDyu8oIB4FHRZ5w9rbWbdqSZ83d93j3Q1
lYgYEhnTqaJWP2WYegP4TGXIaXwD7wMRdwhPdFLWFpbMlEj1dNGQoNaf1c7JvyD7Fe1jQpkEz20E
FerhIHW0oKlw2UhQ4CehTjBVEooZO+Wms6mY0GxPqhMBoli/iJni45cmqcnpvZI3sWgD513m0I1b
qsdhRx/RsylN9uui5kJxjZUPWkElfospZ6/0SjUTxm6MWu3F28tpxseped91Ne/zTNN/SMN28OcC
yZ+aO8jhBiGX/3OpPPoDRDuENdSzZgVceduIUxZQ2MP/cj40Ux74XMBRW9zCjLdKhT6wVpg8l4FZ
daLxSm5wvOjmUPR3km+eRC6gRQNig2NerPT/LFu5tG79A5+NXaVGKqZccx+b6NapoFOnvyyTxp3Q
D3MZK8SGogOInhG6OBkgqOnL/PReu5k+1WzYZN4eXEd5MifuD/2AjELCBM6R5Eu4CoWTQr8dMgn2
yjwBg8ry5vqTI/XE5uWRmn91MjAgZOWjlorCl6F32X/IgH0DX7T/UhGJoUB+63MVX/TnCX6C8+6E
L/7UFH7vO14ydZVUkpOzA4BN/IPCUBcWC1YZjQUcz9A7x29L8n/XnZg2V991B9/A2YTB3+q9i5n3
/8QU/DQnO8EzIMP+dOBnmglJwt+fp76GD5ee0EWMYQisw+XIlF9oQdiK9j4yMwu0/WBQ+VVvJm2n
4aRAmom1+K3nBDNRFog4c3BykO+biV3j9Hu9LNobee+Ai/cW9VEkcQGX+J9O9fqynuYvMj2kZ3P9
c82lw40aGUgztJN5BcC0gfKMf1uFCv70ih7K4BCCWuVTWgc7KKkMd7bAZkuzD6uadZcR9cqiDsGh
CUEYHw2lhqky49vQtZKtvU2oX0XL/RulW2aBasHHQ6BzR/kJ6f2MkR17QVAwnelCcETaIQ8BhAUJ
TJQf6rX7Hr2fq8QmFdZfpyNCu7KpIdqlR9cxeunquppYbyV6siaf+0G/L4MvelWnNV37DTUtbT0B
tDmW09Cb5fOOFMyNQC16Xd+bF4I/DsyOYc0I6KLgDAMjLQkRxM+Wl0RzscxE9fLjc/lzen0R5Y8g
LZPg0/01bSQYcgwGJWL+s8WywUcreP/IxmgfXg/8HXTJtP7RpUDM2M3zWwf7P610bTpxlzlHSsj3
IeTXxl4595uX0wDE6X56Mu0lOXByWk1bS0ti+qYnDcdYtXPql8HMneePs3uKIPzp7y1LxlcY6yXH
J5hLBTa7pBiiSdDTipdkzuAxS2D6990UQtRCaXyhiISr7qxpptk1PL3AS8CQ2AA7oetTMlo18q6q
A5gMFquNw5dGMwZptwEssEYoM36b3X0ycVF90q+yBpPYhqCbTYuYFO0/FoHbE4s4RTPnY8/oNETh
jfXOTF1dnB4XsXWs4kyOX3zo9EJSFgoDPdXYuYaJHLC06vlUEhK1BcO3e1PrQMeNG/weUXyQE/yv
Un9Xg/n4Zfal4RYJmxYayNWlE+Nh1HTeBAath93NFLkEzlfLmyPaKW9sgS0K1YM8PQl82EpGdA1w
86Q7B+q2zz8JDeClIkeSYi8+C4JHPrmK/VM/00Ve07MYnHActubaPDQzmzpb2/OzSHdWGn6AI+Mo
JjL40kf+N7QynWymoc53aOYrVwIDj17XHvC1YCp0WvXgQw2khEtlPefAhllIqxV+yXCCJ6U3r4l8
SS1WwRMquymCCWoffxCNg+fvUjvK43nMiGe8FqoufxAzYW7Iz1bRhbIiP1/bCRBRCvU+JJo0P4xX
IAk0m72Y7joLrs0b/mB74Wk21nd80+LH8otX5Jjjspn/4XxyvKMBMo3nk7JNwrgYPHnd8YALvJ92
I6LS4XE6Zsjv2B1BfqbKvVNA/WtEFIo+5ytL0z/8nuB+xJEMBXRwUqTyuL8y8MdGbm9u7sjyfHUs
kQC8OgWMxrgYPY/qTsxFF+O2VWDAlV975Yj6TNJuj3Tq/7fp+Q+GjsIzj2WwUp9CuRgs2D0oORnp
WMzVo7Z/i50S0gHil6jUa2vkmvZ8Mh11bHDJf7OjXLMFRhQ1l6HHosQLnug5eGJZFdAwORpmBSnp
81ff30/A7QJt6U15bFkaQ+tyMOr7jttSqHMyr+zeUUIV9tlW34MteJQbknRbJRbut5E2Q7wOqTOz
QnLMu/GfKOcH+S936zzc+veJCbFtgNFigy85Cc1mYbilo89XJcfac8YBfL3kb1w46TiFrCpqopqu
t8i87D15a7gkZmMLXDGf8wCfl5ufBWQ5YS20JeSdfgFSkP+Lo0NjZzBFnFk5xZIJtCo5koTcBk1E
2OPQSVk91FfQp/QwyyyeYctYdjpKc3jhoH0XJw9dTbfTItlq4EWfW5szRVZ/zjH5FQulH5UWx+4M
unI+sRcM1+aiqUYgFSI2UJA+bSpORo3Fk2ntqrCQc4koN2ddXmpTAE9QGaO80X6hH/He5+XkQKvo
YaGbgYukw9+6rvO8vV1q86OwylhV/5OQQRom14O06sb/i/dlcI9tBxFxly2G70+xfpJcH6LOZSc7
gghpPlofNL7RpCOaL4+zgzoZketuCYcRcUCsquvP1HT0QY7xUtfoWtZvJl/VLFXe0wlaJAUjsVjo
4eVhETSxHNK64CaFZhRZU374QYa+KM5O1K1OgoC3ovqMAfK9It9sbsYtg3IM289UsWbQ+O/0YZhF
wFJGeIBezPphzTPrzHP5KKuro2vY0d1+aF6LqImxhkphZ8tiE44cE7oYAk1SCpaCwRrY9n8IMLse
j9L9YHt7yf53hj37w2Wn4fH7SDjWnDvBnj2zhA4hAaNCq/Ao7I6bTU4dbvA6V3m5CtbMDSsNpC8Q
zeto5UqhifAhD3XYPVeFSedrH/AgFN+GyQBaOBc/kY0089CLCtgsQKgTVexpobFdpesN67cz8VD1
xMSM1bS2QY3fh5ll2nHgWgdSCR+yyIMxXdI3ahFY41/WMWHZNQ2lw5LRRR//R5MsfPSTR8VZzgnX
pClM1z0ecV07HoCxKlOhDwcH3aOk2wF7RKDZc+3azLNeyDeH9c8RH3dBECfsRpVy8vO+UF+18KFJ
MRJiCOePNLKY/x6PP3+FMipHwT6U7aibYAOfaGZ87LwlPtX77Qhbz/iIvu8LY3cLkFvG8v4CoUQS
Rat09eczUbJVRY4JTlXN+iCkb/rWHmuhWSfcwXypxMSfChi1X5Opw4VsCJUly9hfHIFdd9vnrPIJ
JeAZHtfgbyzX5Dwea/jU7nl+icV14/10A9+2kqEZm2oIZVKLd3RG0U52H+a0M9DUciCObT3Fnzz0
zu69U+D5mi6DzhnS/HngbMQRJ1prQmx4pmPQOXWUJ/EI9y5Qq7vIZBGdZyFJFHYgZOlPHIieaCaQ
iBkzQ1QnuR/fT4XZyw56xd4Rh2Y87UBHlf5BC9L9jFQj+1sT4AZ9ryBaRFpTOr6NO5M/u+GGROEc
UiNdeOBilhdo1jeANLpJdJn7pAkPwHOP5aLeEfMU8kyitxGyVjZZz9h1/qi0otpV6mrwlEOoCc9E
2YhgiD8A2oVGMQAYQdLLT01eDn5xTxO/zlfAaGC+hhg2ioD5uxuhy8lY+inQkgIcXLiLmmF0WSEd
Pn0pTtw2W8Wu37vYreMhT/mKeOh/rFO3q0d7dP1Bm8cXspU8NTkUvF7VU32Gf7iUb2UREtDEoXrd
GakU56OsBhLptlm840QQg6VnMjpxWzkTLbCTGsrZDz2vraczMYYHNdN9H6pdBREjEIG1/tNR02Sh
nlqzJs6PlAzHw2e3nMUE3QARCSBtY0at1K+VQv4JM6LmRm0pXPwKSvvpa3l8P7ETTB5kUBb0KfaE
4Wyp3cg6QKQ64OFa+R8Vi3FQc/PrWwOUfCJu0YsPxpNLHm+a5I+/JWQBWciZLJikaN4/MGkGnEsD
tvU2VRdrzzGm06sWSMtqJpyBu44q2UzfYC35jqpVDB5a+6kMSsDcfI040HBtUoyjJX+M4sP7N+Yi
1OuvYUx61WHvezd6WKAgae5O16eQDYVVvtzKp37cww74WcJ5Q7Xm7JaQfpnuuc9RI3VEIBdiLuMi
ly8OkZ0vMnTre+WkFtmvjjGnUdn8w/pcWkblMxG8G8Sbmuv6FPvypebdfUbRItHeC1/IIyTZwyNK
O8xTv/Av9p07ahOyEgqGddvjpZHopK4Oq5Y4ITpXP9pIZkSV90xv1Cypcs/qimvGBbc1qmWml8W0
6xbdo+fGao1UwwVNjHt4lVruGMPSqt4aYnCDl31zWZr5x0I7ox/rtENPRT0jSyBBV3HgjzcoUOeN
OJq88rRTwyQBTMkHqAuiQkFTDukXchIKl3ATB8pBgmpBe5cCps/gVzQAt18OAPTsCwSqtf0PPNtZ
yD3KpdbzcFjmLakRtkConvIHhNNwPo2mnphmt9ungCDVcvOYhtgGT/SO5SWbENUgx7Er+UIg0rVj
OcAW7d9eNiM+A2ZY2U2WGKZp7fty82dxoKDk/S0cv0VzDSZWtwzhF4elnBALuyGVewjWCn8Jg0rK
zX7rPt/xloU7j/ubCPuoHJTmRmhcA8EnXIYPQsIFint3KKMXHMgjPJHYBSRttrjHaeBAggau9nuE
hAz3PLWSb3QcKmMXuHFWPHIb0Bfe227mFOVpwgOtDDTd0PkGC73ZwkLsWZmuiVrq+XGnlL4wnRoG
VTscigT4/mZKt4W90Ir23sNazjeuQkdSScd0q6a/Il19iGa2qZ2QHUaCZFhBZSrMP7E3ubDNulFB
PeEHC40FtFuMC1N1B31Sx4szxlXa3RmSqFmvjOB/Zbpz3lvVcYNejtUw5ESjX9DEgHNxi1NzIGA7
C5xeIwS9HAyWnyEWSjI170zQIXWRwm2VSe9ahRctBBj2/4TPcSYJPQylGYSfyKvO2uBW0P89zKXU
iC5kvhIedAA8/vA7Q/HETUpwpGUxH2MPeQY5XS/etXEeL5iv90Uky1PLtHDfVPGA+re9lE66BnAX
prd/Ehsp7KsAyGETrTeCTbEutU+ndGqVCcjA7IdwwJ4nG8nQEUNeSDk31J+0aEgpGgo2qFZkS0gS
KeHyzox9EWxuICnvaDSL8Erk6xAGhyptObs+Icb20CIcqWEbcOtIoIBxYmuOR3SitgFnMNJfb+kd
nVt3vKJpsyzLJeUB0pdKuqV+Gq8QYve5efr7ER/9ipwX87tSB4rNPiJM0djRAWFxebpOtf6ySp/3
2GU49oRCV3F3cssBq04165rqSB+fbijZW9RYqPmCsKyBsxr352IRa/qma40DwwHo16APQ86Ck11F
j1tjV9yMBpVtgYHdzZGiz+FA6hh/s7FfMbM/hI6oIN1GlD7wjrZKJpVUBaj9SVLGAVJM1vJDPTDg
jNaZKtg9RFmRMHX4C4AyUU7Oy+j3DiZiiPPwei8AWbO3F5yJE2YCp0afqkvqAjztgJWVN03hxUxq
TWZLpIZjOuKiSJdfX+CHuz56NMwbU87ne8myCP49UWCe5WetP5402OpodJCt8yDb0sgHN+xygbb/
HsGguD1Rm588xtLJ3mGvst+a7YZkLV3O/8rlwIxd+svN2r5+QQg08oc7AVXEFWh8TXNo2JvsatCJ
e7tkyhVigWg8nmEMwgZJgXnBGbmhCtk02bkUGymrg3RUAQMPcpB5/03nYdyjj7Q87NK9pjGTQF6L
lJafE+99wmINATYDVaNRRMgsFu0Q+dy7HIF1tdMuYldS9UTsGaZ98pBu3FvzC7I8leFQsHHEYPSx
55YDMr0z5pysclloBNVISmey+4mA91uKLv7N8gH5IgV++JfAGudt/EN17OOukxrpOaH/Ih6BIZ2t
eIc4KE/Eex3RO3Frp3+hWLeWzH2+spbGnuI9nMWvKuMUFyvvhg8plLN1J2CWGOvONhRXFDFr4DZ3
YTVJg0hnn1GxJRD4Yddym3sk0sPbfB/aupxhTTZltKDYvYUQImhRRrOrc5SzzPCxsz9aPGaAcKM+
P2Y5PjeuT4DC0Ja/J0oZhZLSI6yLnoGGr2kmPSmrj1iEeoCzJMJXf+7XDkts51pbvnnBs/ZKJeKM
Ni/x8NfsQuKaALjvtUfQ9E5CRx3K3r9DNe3AqGc2uemzYnM9GuyIqer1DJHskQGjigdlJ5H/WYCI
hiK8J+5qE4RsGdRFD29VbGekU8SWoRqJMuwljYZR0zuWSxXd4gAV9nT88BDtnBbPZ/HivDPZfQr5
58qeGYr0GMt1jooV2uN/a8I7UROmwbFOjW62q6hdNyuGVAmJ3ArTfsO8PYiFC2hjaPvZBgXqmiYW
Hjs6P/IBO2h6LIPf4KWWW6L9ooJKSA4pWBuAXjvIrQG+YWhia7JyA1u4lg9eSpL/s+nzHeBIWMJZ
wJShwmiELquNe+7gOwRmRjKG4rtyndVxNqWOImDs/Rcqb8c9ZaCHx64i08g0T+iVcWZu//DNYYha
Df3E/5dV9hUQda4xAtn9+pDWYkGpbJesG9muExBgZyg8lLeob18dsJ99x0adB5re1cWkRlgceb8J
vAbLwOpzkO8TY1VnJBpyk07D47cbrEZZYnM10pzPp+4/1AbMuwMJTKtuhI/ZAo++9IVmtvmiAnMv
p6XXl/VjUG6hnVqu3aE1YPjav9nmVK6Vw/ZnN2AOxZJOptyLNuz7GLDwnUEIpES6qJzTFaYpB0ah
Tc0vPYdwT4eo0swKGPgohf/I4ImtsOl7OX7cnMLVGK65aAXOnsdTk/+H0/hFypd1HfmxFGcr4hv+
kmRUbIziwEaEAghcR+FH4QZF3/sYv7l6tE7LXUqJ2MRFqtP3+oIUQV0EA/kp6kJ1+cuFXhHoqiWf
mOLxt7azwnAcEI7cG9wvnR66q2J6GmBOabdvhypzixK5+7W5q63jngY0T3rjA+nkFJfUN1aCGbMN
+skAUFyeJ9rSnJa3WJFVkakt6apV9AA1tyT41+ExctXcsopNMwmf/psDZyiFFJcW8Fa8QUAiVncz
/xLhve7IlGDMkSMhurBN0BTjkej/4kEs0U4FhUb4m76oNHEhYwzyABIvaDrvC4n/KAUId1Gg34r9
GV+YQ3T7UMSzwmUPyKkNrcrVaO9pWF2A8ErdYA9GpXD7HCequD0EYs38Q0LaKiIA4ylH1i0fEJuH
7Hjgtz3bbG26Kz7RxyNzu9Uqmk5moiQjumXll6xUYS1y7usTUiyEvY7b7e95U6A/LC9Z1CORduyD
UEdWFJ+6vtCU+Z8CU927isAbXeGbJT05QsfgCy6rYAUHAjIswnhE603Yy8kfR9O04Fdb2yZ9315P
LHiQf5UGvKZy/5hze78mqnMK0fYTgpOhY2XpVkdWbFUEtn5e+xVgp+nZnHaK2wYVbCQDDUxo5LVq
Z3k+pzAnjk4xChehgjlYu6Aa5kgJjttJkPmndyA1NEHykz3tyBt2gQMlH6w54JXkHMkxYlj2cbrZ
vJ66h2mIhp1mg8RmjqbJRn1v7OEhCwa09mlFngRAAnHIELcSBLZccKt9zLfmqFO/9+P2ok9pLLk9
izovqGrwV270hRa/YUy0AEHfYkQ1Mwvla5Q0cEk7HaYYv6lrC38e7JDySigCBj7sGLCBt6A4A83h
eZM2O1+ZrX1LAomML1UZUsln2QEIcxQljK4D11E75UjnAz9W/qe9/Z+MV7WJeA4E528T2mtMwl4H
YTdHV3Jvct3E9tK/BRGBA7+oqSxgIwipZT3/K3FcSDZI3+LSAH2BMIkz8JIV/z1BnJzyLqyPUFba
dX9ScolEtRkivsTYOgE1c6q0BiGPnitrgfo2HYqmrw+7DVKZBWF4WOkic/FtjwCC7R4hpJHFBX5U
IoNttzBXw0nTeVyEaWz37srek8uies7UtduqLcUlT9RwZ2MYTZpqk5PznKjxxHdNx7QwkN4r7K1x
kD3qFl7LvllwY2WEiHWmddM8ggwCqYNpudJc7d94evIB29pdhTzl94QEUkYZRNiOYwpH5tY1a5RT
4/ytsgYiHzAylVRmBGBCDR8bf/f36hFTovdhbs5t3/01X+l1tHdbFTUfwTNsUeMzZU0YfzuYfDc3
ytN0b6mlxCtm45CYmAvtTzWQ1SVHpMtA8jvKQos/s9E4MxUhdifdq2VjJcJTdu28dcwToTIeih5V
oTF5IyZIlXnBLM/u74iI4z+9KBdYELM5TUBdHFFp+K7NOzi8bzw4088gK6lY8OlD28i+V+kqIDmD
bGRjZCx8GVBQR1T/g+8SG/Krp7fM+Xdc0NeA2QL6SzRzaiMIx12xEKiQ8d+mRsoM0V03qOaSXGSo
MAYuDtPNj1asfrECVzMG6ZV606dbUT69pFyC9+WZzTYeNACPGnt9RfFprutDPAlNuCmiDjS/He5N
yUmydqIlGuZ8J8Pd11GkQqIlJc5xQYVqrFaK3MQDfaBrKNDYPKLhGP/88GvLe1nVLO9VP+9p9iGf
Z76f5pun+p0q4prUAqh2YfVtAXvRqriSl4LbxA+ccl1f/fO2sqDIHOHMtJpHMvTCI9qQ5IU9REF7
Z8Gc2U8pjm2sYuNACccmf8Eg7DRHUS2qBGklnc47DEw6bryWhxG9VSKHhtunG0wnFkehDSWe3Ybd
Pr3KcerRax3hpXKstYU8Jtwf0kwfD4c+sTX47jL1jiAZdp/tefzCTJ6wWEzpJr9tf6CzMV24bLKn
SnaRmefsmsN67Srie2z1BOwRms9VM9eoIICx7AHZJMABUZ4kavnbpD0n7qNeCripJa7yqVkG2fGC
DmDsffsv+1DsUvX+A+UPVmP0HxdNtlTAyL1DQYqao/YUfb4nBa/wvZS6pDHWaqZfVKka+zvp55I/
ryh0en3Ylx+DXCk/OitT4sxXAo75WyCfFFP5HsT7FTItxGyUU1dA6r4kW6HMDt0MdHtqW4pL9IF/
VwyFzkBHlCVvGeRrcPIaokU7l3W9NuyIsJbuTy2BGJAavYptqJhdswHYcauUBzEpZXtl1P7OEL2Z
iWE1JJIPQY9MMcP+2I1Hox7RFURRwzVFZC86hNM9qY8N8HtoWACKiomNYl6gSRI6BuNoy5kxZAFe
K3wctVF5suePG5LV5WfhkAsVt7dYocRnG0/ndp6yA1r79x37f2fDtXuWOFm3FmN2RnmE/G4B7t5z
SZIVcQivAHQFf73mIn3VzmtJKWXbq7zqfx2H/Z7HdKzN1qL2lrDburOzqzXWtP1krEqJlgbfvaXv
htNxMe2n1SpsVCY/S5KC/OndCg4xLfbIndMvKa+1zJgkFpq8yjF0z2pL84ykVnQ16dntQxtKm9nS
xLfKBqs+XwPJkIKfO3mncQIASR0HOvVpNOSFbLxX3KOUXLW5HjAB8kK5C2942KPzC9NKpoNxURl7
lVySuHO2UyTb25EYVoT0jwWd2V25oMstHI0wujX+jf2j5aTKUqkOG+uncFLGRDJ8Oll6fr/wlKdi
Hz0LUcxhJY/0rrq8tKh7BJu3kDLr7/61Gu2hLNqkDz52FZjnB5OBySXbb2ih72ffOpOQzUXAO8IM
DYQKjIplrvsR4lfJxa3gWKsdv+rGB4ggFUKc3EXQLcR2Dl27w44QMvFfd1DVOJYOYvozJwPbCwQU
qkaO/psN4+mYvYG8oVgq/Nwi0z5i5dim8N2r1PifmKaHV+cvkSm73AHrm/EJ3rConW3wRuEKY16J
J+eCKcxAzk9EJSv6n3gGyYbWXOpOSHRN4s8FF2blIgJTlWD5JfSKdmjlVSKebxfUKAuC53qRZTsB
P8MiKiDt59DKgfjvEMILHpl9lOfMMYQAtgP64xeco9XN0vMX8zjPnw1jcUFEoLxH+6Fk/VTq7tSg
HF+DvtH1s5TNfhBOwx9ifVi+gbjEcxku1uNNhPKf/iYFLuDL58jZufBzK/uiMDCaHAaRtVtSBcv7
oz4HWuy6me/7yJCv/2h4J1ogAkcHbJoGDq4L9W+FF8PF/zQOccrUZgzcW5V+wyrYGJQp5UazYWsn
GAaKHhGtkwd0OT+5xEghJH5rb3JP3xrARdFRFOeAhNotgX4H1xbPB/OlRK4AMrudOEFfoxLB1MiG
DFCx47NB+Kd7UgyFszbS0p4oHH01jafrhzkn3ENPFgCz3jAOLOMY//ecAq5OInVcig1ZpwUxaveL
Q8XanIxJA/i9bv1VTMzeESL+m4gADCS2HLVqp6CflGXP/d95qZN4sMx5reNkMcwY0hu4F8hBrBg8
BwRnJR0NceJOa1P71rk+ue+OXjMBeSHseXCWsOXRuR0gylITIkkDvQG665RSo1QoRstubgQgwoXI
SQIv1XIjPNCh0zW6Q8vrRTGaIDvdZ8QpBzuVAcjgz6tIAbEPv+ifh9uxPFRyTBAVuLFWLwWbgbah
hQLkqzwpbVRFsiXkS8fm2cdGi/rNAR/M/dj3rWB0F54n/apBZaAwJb5eSA8OVboF3wHxLQT2sh2u
Zws1nGoEyWcsscnlskrHF315c5OHO5Z3Bz5u9XDM44YR7E0thHa9k0V9215tVDzz3yk2+jjudNcX
RejZrGBuv+GmZJlcLjUnWbo2s2SYr7UIzG1eFWOzEVucww6HuqIXxN4+a4dpssL99d9gi1BVXDJ7
ODe6XWizoJEXKCsRZseqv47BICuuVcVbDSncCl7jvfeSQdnMXzlL9Zk3jBgn9rKAUZbsKBo4Vf7T
vAzD3c0m1lmQP+utf+vsmdE7lWmSGfOI7mxlX+LtnE6eXSS0LcRxCkjrX73IZn3xoAeqnpLLU/f0
spWkTf/3NaKSDrk3DoJXq9MOD0TyAGC2JmObbSpPIh1+sTCZlw9V2ietEvDSnJxw8EiCKTDHF68Z
6XxrSrvdri0N+45CekSF7Zoc8VMbRNTvRX+pDAh/DOvBfRtj5BBJIMOAal4qGd+yBsO8Z0HTXUEh
1WOdR0pzx9CteCGaovKJdr+sqXabM2y56awwa+3isdhMWSbhno/zKU30mnmdvQ3YEXbgRqa2oQos
HXJsnGvF97cLsP6zpUztAO9KnT76o38pK6so6juoWHtuiHcXujrdtHaacYFv2JRWYi67L3zeZaUi
FBEnOXbvk+XVS4j/JSxFyrE1O5h7n26RrgkZbIngREp36fXJDVn/ptrwYjTczai7oZdYla8XSydA
IfD/DA6uVHDOxc2DyRnzG4xdWQPlJcHBrmCzqCnsgtUr0jbHAIazxrcfzoUc3YUWNHA+58H0TVVR
4cHNX70iL47R2p0c+bNZUzK4GNtWd379h+tqSV7xDJvLin6OsMrzD7EcRgMUFY4MRXMdHUW4/yj+
HdeS0VXIUtIce+3IlKbKXA/18eEDp49NIjC5BhQnV8GNszSxFJV6C5cTYEVOuPcWnY8ekbMdoGfM
BbWHIKjxi/lOfFUFrfl3gtLUtDuqYa0r2ZkMIuIzJpiXufDmbbVE6H2tLJQUcxyjtKGaSzjn4EOr
PbqN0N5NIAvIiXggLeSI25YaEtVoZmO4Cpw0VjqbQaH3UGuLquf5A27J7YRBi28V5/ZnO5mInvW7
28gHoM4t0zb3cDyGhOJyXhSjUKAMLnkewHxn09NvFyYgZA/hmFHm0LrG96qCmJO0MtqbWws0bgLi
BdagM6eWEz7qAjG3C3JTgecUe0Njo7Nidlsb1Qv7pNgua+5qRi8QoFnqWDxy4f/1lgDZDTWNMBOs
96SHH4zPiLhnAcULN/txeMenk8EIOiuCwXdK62mDcij/qtxx7UUngdEK5fc0aHPIU2XhVA0ow4m+
CjMGzi/MBbxNhePn9wF6RFNe9xS1TNP+ZD09YBGCNBfxtUnKbmmS5joz0jjLC5p5dMYmFQPaifjN
utnsSq6QCQCQPgI2sPSX+xOeq0A4iUfa13dJXrVZGuQ8PKq52LI8uEOfDZHZ5PqBlwJpa5//gNKr
j3pDKIEa/OD5unNXZ3Xwc7ffoedgapXPV0htIZrTlMwgHQKdCjI1eeEBIkmbhoyW8gpDsH44iAv+
LSTs49iobbuuCBsqWsCvDWoyKbw1OuAGPsao29KPL+3ls8rJWjRDzVvQnWUH0y4zmKyiJoNrH+JU
0im4twyVn5NaGyMXfQEKmCYCvNslhbvWYuJnHGzugdI34Lxasg2QjUqONVYgxNPTl9PIjQaDwp3x
O1qWIu7OWyrrSeRyhf01/gH2+oLSAOw+UUO7zMj0tXPv2Y71PG7zbRWB+V1MWeg8RdJySYCZRzBH
bJTCd1kN0wSngPIMXnJMbnVJWAhJxtWHd0dnvX5mxmY6epIy2rpsXW01IPyibWT6YzsXLgEBz7NS
u5oceDTuk3CCeZVWSswDQG4tsFSQKq0e6PzhmmfIrDJsYlc1xR+oxzRt9A9y9Pis13A3uIpLfCdA
U04sArsliAbT6hZNuB90114Aczj0VMnwpqKio6qX4ItIJ2/oSxXuMNX4u1j/uRQwNLDRcY1hOQXr
D34WDNctsggVJNSSIYUrXSzN8eKcLoibB+KmoJxTNzeVr1Fk1SVaSmdax/FYUApaIn9g2lPgaWYw
WCr3O4hp3r+F/jQSVw6KdVbzsa4lD/UKrpUwAbXX8IMnaJ/BnWhQuuPy6WTmsWFqXZwLb3CwkR4Q
sn0t+NEQFHhOPhXLmTYFVnO/vWxRs81nlbIQbFXlGkUYWo1TArQYeD8a0o4p+3Pl5nW/g3TCFyLs
aTnO1ak2loKOv6/w7aR5PJKgsrc62W5svd9uIfBjdLpZRAH1DY+m/H8lE1bTOkIJ9iOZ7R+kqu0e
5vAkpDI95bZlXvTYamsvF9vHHYrTnF3mGqrU/UGW2P67tq5NTj9G0kg2YTI/gq64bOjmuD7QHZ6F
2HveL52NLi5+tJUWflViEAXf/QbWNqfbKdlL3uKxgxTVY4GZjFYfyGiYLbbF0AEg5B+LUHX3sovz
iOW7fsc1y2aWiiGhFe78qtydhhWDp+nW3SKjcvz0Lvl4SbdJqBaK2qyRa0ZgSKdcnDIpEMrRzjPX
DFew4awEX3EIbZnBYFlJJwBqFi3PTnpsnj8bOGB5K/WC1E7j/wTnkVjOOriBatD2K603wiGZZ3ua
WpsfMMGxUYwvW6y442z1ulFtMzhCQ0qZHkEoFKTFymnXvar7ghXuRTWHcar2LuWGg9RBtUp0Vsn6
FrjIgHePmwfAcPWTcbwjZ54e64O04lypQGbRODO4V9hFPIJV9KHFJq3g3bgoc/EThmwgKZtGAdCS
DmEoFfiPc8DtJD1qH3Z3qgyw6FSe4a8OaezjvNjN4n6ZXjoaFWBPJqu6y/PT1uK0zA1rMgkpxeq0
ABpFtMJiNql9kniIU1rF/Roa4lRn825LhVm4amfcC4ys8KttyU8TLcZ2qLnBFIY0VhrAwurzECfO
MOdjBV0pVbesyWtMEeqoONGGfW2yUh2l8lNx+R5tGchywZ0sXpU6LG/v2lJzKxaasPUhJECi4ECo
xv4I2tnqMVzrgJpHjrDIdXk4PRYZmoMQioqqkd7l5ijcwBcffcoj/ZVqhm4ddrVQZvL2iGUMDHdj
l2idB2xo6GehrnmYdi1uugbUEVNw1qqKoCMAarq/sk+20UmAPSDcToEIWU4LOUu9gX+W6AtHAPOS
RRfFRI391h4aZQ8Ti+QT8LuTYcPWVQj2bI6ggP2KpmfQUyeji2kOx1691tqvwKmTzjLjSnrn1a+V
iCZ3ewocla4R0AesbVovjvCAFG4AbZUVGuilY5tk+KSzGlpjXDMLJSHbfy0MgtdAr9hrLj6lRQdU
O+g7z9XzYCIfFXdVJmGItMIhfWHi0Cxazxf/FWXQ9CqbZJYSwNggWFFN1+CtHmr/Z2YXYbHtEMY8
W8UMMll2Vjj++DOZS3yhLUyXrdN4rBeT+iXZrtAXFqYntWMwnqAYoDArx8sF4ii9N9XNmsWaZkfs
Mh61zfQg/zcr/EdTt/kM8fygyjNQw0Xth03StlZNsX4pvLvIjL86CbviMGTNUGG25VOu6Um9iGHV
oMsbODUae8cVZvIZles4g7EZ86mEV7P8bTz4gpZFekr1abLnQMq4see0MzqELfCSB64QpsOyItCy
FmHU7osVhxWAji/dar3N0WG5d0ZYH00gVgbYtGgqGUsu6jyzDS2+LdO7oLhh+DUsnwLBwyoOxtN1
6cBmYu59Iu+J3K1TbiX+SV/9MVCz1eEeWsGbpiskImW4ryOdIkWTPXANQFgPR76dTiy07CeLO4zX
GaSgrjgXOqA19+TB5+ADwb6RS61xtDKwKbDBA+ZYpdDnNAc0QuHpDm+XRBeq/AofiXdG01nxXnln
5qBbiXfctk/r/IGW4H1kkTIXBKCVYI+vE45cHfPiTsCHHXFT1/3ffJFOsD4unQj5m0SFok1WLQwv
zBrx6SX33F4Zz9fbdkgtOJSZda7k5oXy2zCGOl6pFRwVdkrXNp/zDEPfLkdLkwx5SkzNzQqBtApc
pCdSB4nR11HFJQWl8qE6dpS6Tj+cqBFg9DydLx/eWzMgN6kupmSl6uw8W73Ov8Sq0X6jC3TDL394
ML17yGueQa1ytHlVDX+0wAKJRvZC17Dc5jl1znCuaO6xgPENYGnT6oAiXheYbbdqoz0DYGttbbOD
tS80Dw8D/udRpSsq3mbGWQRl7yNTsgjzW+JRNl0F4RgpzndCUbvDmyNCHE+/39V16pJWbJMl9HHg
i8CMmphwGVUc5ELxLgsL8Bml1jnBj/3Pw8SzcdHSn4OsY125qtBQp8UPV6DWFPVfJF6QUFJs8ih7
QdOy/bWCu1DXTDLN8ab4CPLxqs9OMLiyQ7uAJGYxTB0hvdcQ1ox6E/ppbo+ZQdY5ATbKq4nQdEj1
wLXIs4nOSlqFN6Jwpfw/mEtuLPev+8ED2RGX9AQZFQzCNVHBBl3gvYW9dD1gzJH/TwwwclDiEU/p
Xgc9HK2r3ut6QA++K8xGH8CsIx1SQn6VQ7AIDTyHHDy/DKcPKb9lavdcdvh4HvRH6EkIISa/mBII
kP/qnSyP3vkyTRgcJUf9nvOBo9YOMjOtcBw03zb0kEl7w6iq2KuChxXF1odXPTnmc46/tISJw/50
04r2XiSp+xiN254l0aSv1ddEomQ2SKQszbwAow3LkXgI9Hdn0t/8J0UK79N7kqUCj3989SEyHVE4
GahiiHnnDPy1JG8Vpc9CG2vU+1jnouPwlVA1r3uflsHCW9epEHgDAWFlt92A6XeRMKd931HIPhf+
YD3aG77sT4r1F+fg5axJGm/Dp9OTGamQSmfnsvgcoLgQcu1yyOlHCFbzhNRWwN/AiH8ZDTfKzVcE
yuuJYh/PxwgjObj91t3uMQBrsOJSbLNWn8C+1Vw0WMcUdWuvgdWGfvSebENFn5v4TuGlCF/h34Dc
oaVLALFufMqWUPStuftSghy6kNCbfYUx07oLMi8hMMO9jK8tgNDpYpWA7RNKmHi28ZANd5U7qChc
mfP76IbQSs/FxBq6H+UwcbnQtwqPdbVDD/CYxYL4EANu6hvpiBxII2BYzykU9dYHzyWIDR5Urt4a
UTjv86tVIV+L9faX22sXvRYvba19fefMyjL4cC6nN4KIJ5guHDPxz8Em8TB5bv0jxbPRAadTBHKk
Arqw6/YET6QGgBzh+m916x7Q60NWb7e+zgsWqiCTsqnspen/LV+RMX6oMV9V3+MK1qyE3CDq2QJD
a7LHUra/pewXaIQBwr89SCaJAWvWyDBwk/761xokW2xbSkO4u1GEB0NrOmQu/K6mqot1//QPaXYh
0Rly91w1RnHQOowG7TSe4qLJuK/HUiShQSkNM9RinUX+OiLOjzQti84n66UrbgYSVD01LDruJuu/
um+fUGrAGsv4VqXAThFOMAowgCkd5S/9D9wCFFk902Ff0KvqSdQb4TVjU4xnmVN0NvxhmwP9nNvE
Al4hKXo7nUiOyjrZWm3UkB9JJ2xOFlW26rT2Z2e0yx1KLiXeOx/bIS2Y+8St0oNrVqw1067Ay3WN
RnAOIbifNpZ+tsPx/4Wg36C2MtudrAk22vHJEM8kcknykHc7lhyvN2jUuDX4QtuMtybRx83wSWZc
vpYzJBJrALTKlVaWVddV4u5E7+uyZg9oQt03CuplC8UV13WSAXfYIsNx8X/FJg9bZlLw4a05PtAj
f8hF4ji6WlaeQHkAggYLT5KJaPzC+QrbhhcrfWR0Cckg2ZvC2d6mD4l9nr3BkTHHMhdvE0xSwgeO
/35siM/B+0gQrCtcWWJsckN7zsKfn7KAnjDtKY26SLH2paNT9wN6SmQhq0Pq2W8IJ+DwOBodDJlg
DPdzN4af4oNz787Tut/jXFan/sbPgoW/KgqLwRsVOjcPcUIIdgEnsRh/jlPTZV52+Ninr6puYzb3
J1Ps21PWvoXmaVYSFGgrQzpscYwXN9GHtoZTs7XmB+1LkrMkKmNZoXD5UXYH6RYeflhMb8UQMQ52
l4kT2c0X0kxx1e/Lw0I1+eqZMhawX3T2+6Px2kd/QebOeSsjy2e8YgltMOaHXsLAdEEOf7WTUmkN
DCldaCPJ+VD8myry5sR39YilLp96FXLVPjOrJ1gKxxqDc1eBiH5XKOW15We600QalyS6TxoHsboE
iNjhn1Wh8OtiCoyqVujPLPZqkNCFeNDRua8xJyDjqMDAzYPBz2bsu/xSzSzA6StjolJS7hJNX/Z5
MxZk1q2EMTXOUX9CHSqMQnnHR06ydPJMmDk03sQ3ByKkUiUoUddVDMR5N38fXE7nmKWkR0B9s2AP
uUymEIbZ7sELbazarGr7FWhuDIsQ3x5uooPWkD7+j1FsHDblt/ClVPLKcW7VXvTJa6Qcd0xgt3W6
I/b7tVWvUY/gaU9UyuxAuc5HeMYn6MsYjNu2Yf53plDH5SLIZ8IEgZMDCmcpU4+h8Pdvok2JHkQm
vRnBKBD/TL/Qx4qJpJtJDU2+NscIkaIoIpMU9ocfXzKkUsdY+ST/3Ulry0tdITWgRurzNPyZoWIj
dQftfIBAjkvN2sOMKR6iBkmL0kOQOQghO8gV3QaakVXPcOX6AcaG6iAWffRybCyZ1ifOKzFIXyzY
rb2ij7ie9gswLucmFgvnXcn06H2DnGfuC960Gcp2wILxYGaD3c7PLCGjyqT7l6sD3eCM+yJspsCP
wP5z8pgrh/waFtp+C6ZnVKAwE1oAzJ9ilmiYTW6Gc4FrejCwKl8KFtOBcejnbmBR//H0nDDp2DvD
6QDyfziLLXkzNKFpYA9imFGXG6Pc1DqacfRF0lCgyo4O0AzUGh/55tZATD4u4l7uVXAILJEfwh1F
qphzMKlFbrEJXq1fu3LMBNhZiZEvRH/jAWiVctVhE6uCDu84TTS6VH6xZGwJB7lXbUMaSjcvP8Lu
h4KcNdSJtJl/dPSW8GgGJzu1WLrA977l0dJvpNcC9HFMmX1SQzNrvJ25u3DhJfwNkJR1uU1Avgmb
lnkRzYvMF6ap4pypaKfGTFoHRydjaijI4ZQhlMYMokoGZ4vsL4K3Qmuf8rjJak87nmwnOLr32EIQ
sBNtFOn8zmeRAsTcxUdO6eC3phwP/EqeZw7ZPfnhqlBB7unqvJdZVfCSrwqUq2lCqbHumaXBupP+
mPvv/wmKx1jLg0hx1u62NYj49LI7BHJbPGVcHo/1xxFctjAeQY4TS5cVMRmTsUMga23a/896flkn
tchJMsusSpWiqsW0rQVGOCP1tMZEvgtxY2DD3i0/Ohn2Ll5yTQSB1hVDNQPY5q4Y1f3j6mPJuyV7
H6jkFtSkoAI3P13/wHDY/6Yxsp3Ze68OyX80nvV7oWvQ49NT8TLApLzPXcTAka7hilshy2K7/1lC
UR9YtTuEpUN/ezqqBC/7hnIbacTTL/DuD8Vx9m/Xvo52kXi1gX6bD2iPKDk0CGyVz8cTQDv8PPl6
sFLMY6Gg3z9Lx/C8bVrIjlXBW6kUiIQkngWdwfU2K5tDffDIQXi0YadBIJfdi3lqnTjMdgokNobh
OuveK/P4uGoNv5FTfkVf8vlkmkRNiLy9xJbPNaSgy5JxzzOvEfMLM59I+jW0r2W7sdjfss6kcRrz
cIDj5618RwzI5X7s2w7dXbdccDKYNF3BYFp5BlQ/ukGRx1kZ2aC2PO06d8aSnwSffbx0TdeVHlRh
2gc9OwA6QFulAkUPhGHQyaKRd+9SnMCwaUVW6pFPWMjObqdHB7mcY0+dk4zP5MLsj0ocAHMkUZSI
eGcRdq+oCjKzM9puq/LKJEpThvSu60KhJ7KtcGV89FoWe614D0mOx58/r7jjo8I5q/rF6eCoXbgH
MlyoizmKydzE0C4KM+qH3bb39YYUhulIkVlclTupbsnNMkX59ld6uGAF3qmA4s4M3HDsQZ5VrWrY
PDSvu+M9oLvD//egGMHhbEBGbyBhfAGVuwTPFsQTM+x7bsO/pK9ePyRlmJNew4tNUQzCmftgwlVx
pbAdPA5x0Zgax3q+MrhH4ztRtTBMA0G5NeYCmQIIra1Hlud3pyL9rQXR+rCQZFEyzkKBupgtYRXB
0D31WIQsEfpXuCCb7clNXnc49aZ1TLBm4V8YmbHY55Qg+FNFn9mZrk/WCN0rZydKMXFBM2yeoJ7J
VNn8I5IPTXC0twsbF465ZUW25+eQqMxkecGqXyqqrHxGUc7ONIzNTyphStSwjfA56hQshp5YyvP0
6vPmwjOS7bGV2pllW7PEquqZopcFNjHIpKQFUprCNTQhq8PzORX1pVgFliAPD/H1+0RO0Xx8aGFN
q0fL27zXpKSXwYW5qnyEZZ+AKEcovve04WtP0VxO/xZAB6A91+m/gQXcClgaR4jrAWfWoksOeG6E
oAdV014DRj0mvZPJeXrf8CKz+2cukX+kx3eHDSmfByEWI5PpKN/i76wa0mYBpvkvZPaZtySLZ8CW
i3BZ+oFpdq6U93NCdW3ydQNz/YPCFFlylAGlJ7VnWXR9rjQeks6RGHu+6RaNfRV/C1jiq8TmIobg
JoFYCOUmjQim5aeitLpw4K00CMcmxqtOH50f4nnTPuhaBm0mTEWdHZXVrdPjcGgGAd/SZT8sZ47V
O8wVHrOF+LGjvwOmR+xnSx6VpYGyH65Utrfl1KFYKTJEPkySbdard+8iT2dVdZ23PncOtt9JBTqf
C9QzBUe/qgnkMKmNSmOvRLeCSkKmu3NhiSQketH/H6FxHh/UewLkcH8wXLh6xT80YEGwN21h2smX
nwZpUapSsZY+EoggtDagCg9veFGfm5VwLARtDEjKEhDELNdOp2/pvUDcOocHCNbONRGLe60EXL9Q
/I01A6p1BvoYDIZMgPw1g2KPQ7uJugnrlGNdJDn9iz9CqaRCFlKqhoLgtLZjWL8+71vhUCayJSV4
Og0vWblIrm+mJrlwf3qTen65xNEaKCf1przYIYR5BDizjPmSbDEtbrzKp/I5gCWpF0wDcpJc+8m4
is2zUGLWV2ilCJWVOoBcNKirIhuByeYAiUOHg3H8wLliJBibi8GNc/wvvzXrbvroby+kEeFIO0k2
hxYfsxhZDX0lSu+b1xdum6lLMZXoLkuedJmdXqfFZc2d1aJCUGabra2mzHNR6m/I1cXiaZjg816r
zM9/DpJiyc6k8Ws9la//fcJzRICbRKoJlxAFW8s4wsURARMJlTcQWqhmeQeyBw/FIWrQ+I4bwiec
Vnb3GY+6/LnJBqQ8nsTjLtVnUYNzGtttfuJdjzh+6ONDizeOROOD54WpvM3/yN3+BF1+2e7bJ+VY
Mv5KGXOkCuFatdk0logaXPBe4WFi5vwkvVPMMmxWl+DddmYGc1twcdGcdajb7zriopRGuRvzsJpe
1y52b/z8twHziq332CnjDJJHepdtkAz+/2PDDy1lsYQFgatcf6Wjf0NpuP65MPuAwXi/BlXIAhKA
DlCKXL478BpPnGH9iiP1kF8lU7er1aIOKEKnzIaqavDY6ALXGPed8GWD127O32cmfT5TpQak8KnE
zjO3YLAqsrlxpvF8xVtIhcnITKIPw+JDCrTom2gxwQCAyWbDOF9+Fel/sAKQ36NyowjRWB4rAXxC
WA+Ru9ZnHs96kKOO/GvenxeQaRoyUvtpof+6wewQYWPSjdR2+EO1oS/RDPFdTgewX6BkJ3J7TXcz
QXbkzEvw1OmK7On1eayLvWGZO8iq7VvQX/tgq2hNAj5MRDze64vZMbyP+JI1e50qAdKI37zJgTLC
nCWuarrMo3i4BpH4gALVLw5kdNaI6fkwzcRBg0w6qJStkpM/C7zdy0sHzVXOKAu1/BwtL+y+EPYk
RqY6tQ+gRT+6Ob4ouPmLwveeSFCZCPKnIGx/ZCCs31T9qorK7A8lA1AngooudCFad07QofOSgZul
0kNUcI6eCbM/wqgCyaK9ARH/nKET4KeMQ6M1T93qLDzBIxN9YqAaGsdIsAEud+p4o49hFFYpgCgV
OgYHzaLWKG9ZUvumDWNc5YN442vopIvy1lJWBECi+XJuPIRaTn4HfMS5gn6XH8EZbT1jO02QhkDH
g2+a/JgaRI91eQEWWl02GqTa9AujD1HqrCziLFqpDG0/YNiaNtzWL0XIC09/6uRaXeWIi6ZYRmJw
vTQHeAMFz0c8N1ObpQnUwqjgaJs8GldYAPhhc9Rqp8Twr7tpv6Tm3xV0s81T9PWyXFnJ6LqROIaN
8vxABc+c69e3Z3gF/8Y/wt5kWB6rhS3BjMZpln1FijNoiADfkuXEAY+MR8vU6gboLg3GL7FzLlFN
jJOcHyVE5axUPm5dGTkWzRGfTou4z4X6VYOVmqeTtjpW8NGMcn3+ydemGmBy7U7Tl/QOPOm/wQ6y
LSL2ntIJzCtKYvu8UKAh926XAqraufgaJCcWG+aFegqxysqMa6BOEfKQnt3x+uKpIFUuUvsv+YgF
rU9YELoE0d3Qyecu7X/nrFP8prLA/HzkpdTLWTfv94fm0aMGAGvwJtvCymdQU8k0SB5muG5oFmx2
gIhlbstWVAuUCCb6drZrMRMWjMAjl3FR8FcdfEN3+RRnbyGzrLj5TgvBUr2jWB4d0VYpoGkR/x3l
JkJlZbgXEZ31umah7fUEDbXyZ0TnVxy0+R+mqRPuC7RhI/vAV2pFfC0f3ZUzT4A4EQyEFEVd1CPS
969SKRPXupEiawhBbKvaf0gNiUhupEso7iNANlY8pTwZ51mtRLeOxFeIS/rl3bqi8AIvmbvYXvGQ
WwhZ8GNwWuwZCVLYlYsLdVtJXCSJvlPfAgH/VOwOAQH6Z6MhqEPYIRVwuAtP/Apy/HkvFBXufK+e
a+PBOUVRNBOalD0pl/gpqCXRh9qcv6larP1zeQF3S8s4w8qz9la8U0+OePImq/KLDaXgVLtdDXNc
luO+yBVQEOgUDax29Q+0MOJp2AKPTKxcd03JkJwPKKwD6mn1Qih5INlYcSIl/vykEiQk6LXmxHcF
qE6MpYYwFESyGas+C05xYO7nZ8Sba88paHWLvAkVFQCm5QhXLDU+ORP2vUfJ5lFyB3jY6ILcXP7a
IVBs7Xrh8oRgpYZvAYg82SdvDrpNuwOlUYMQ+hQKg6glubD3TYb3z7vvsjsmveo6DScp7FDqXxOZ
gKLKuakY2i3MUyKeN1i1NDh5l0ano/1/Y3L+LZOoWaicd8SM2B/druSTTjVkwxyQSPa/QPsbnqc5
V4DXw4lBD+G7lhPdviCHu8Lc4o4wnOlAoAhOTus37IYm8tIBJVypKpevjDzmhm4F1ok2p2ownU9y
WwPg/eK9MqZjuDws1EgOSlKQxHcLoSQ/8sumv9Rz6NOcBbi4dPfVJ30eUNp4Rt3swfVJnJQngyDh
7Nhk7RmIOcf5bJne7QFKO5vmlJn2rgz6IM4ix1uytjYzKzfKQ1JZnHSz6S5GfKNpf3N92vfmhkeT
qCbgrQIPXj47Rq7fUkVdbz5c7wdQTCX7jMGjZhArFAj+5CFy52dpz/4/tS1j9rlvLJHbikYZ4p+r
CDYNj8qZbiheq+g+/uUT1eUaqDJ+/SUaMiIPEPV5rhHAXX5m8HZIscEzmPA+gi0i2bYwWiaZMOTv
5V4hOUrxi/Yd3i99eLzgzRpTVTnBCA+NNZlmWpqqBUR3gpTgv4Z3TdfVGVRu8HmOkaZhFOo1e0cJ
ALxF7Kv/iy8ARY3LNlWC/I82mIz+xlWAGzaOEdkJYkRAEGb+C1lUunxeoNp6o8TXXOWTjYrmKXyO
8P6FsyIveJQlzgkKY0Jst+kKgRqZBAqX6Afw36zRFYJloZq9RY4AmRMNm/5zS0VFipCi8j3NV/PV
789rxfuts4DX3bmpB/Fo+HQZgDkN0KKsJaYisfGWSLAb/FDNqGxCgNJrgMq74mijiX9TlBPi5UWo
EyrTF2MPlwc9NTgCMwMRgzBmzi7qlPDGzxC1QJmNvw9iFSFHJdTY1Ne2eeZkNJd2Y7AcL8Oc9uwE
vyYCLxryPs1Ky6E4xyuE6Z1x8jwEgu/eRB+aY93eNoJlSP5bVjF8ezAFtrYxh3FCkUeyDXrJNoMM
GWrH2oIf+I1oRJVNLOjQ705LWdNIaew4hXrdYcZOOfBMdW1D1caSnu9c73G9yovrZmViYoRxLu4f
9nX6NkpeFxWA7hlNcBFn2vd9Vqcx3unYQT9291bIp0ZerovR2I2u3ZkutGj7FnLBs0O0rgHWsWrP
B6sU3xh6753qFW2TxXrwhDJCA6a7DNUw8I2st4dUTldATx6KpYd3QEyTK6nFpNY0GOtP39xwY1LZ
BGak1H/ouZj1jyyz5mtiWXZSmrGfU+/4NDWrkq3Qjirt9XONdGgw3w87hCZHu1B+oluEq+bQrTcY
sQe4c4nCarRlIuCeA4JdafXtH8tXc7g4/9JhTuHanoO1hm3W0wPlITZnFMgf5GxqUrYG96ZNgjzn
KsJHD+P23YXBK6WHlKvw0wvCRwmPfi5bNqDW5bnSdI3RJRD1Xgg6LT/Chq74qZOBmb7PRaM4jmXW
7Pm1LplCSkgyKzlqFPYlJQqVjZX1oVHP/Evclj9TOEp2t3lKuAKMiX1xSOczc6Vdum7Ctl2tChqN
geBL2dhuV98O4nCw7BuU+cv1u1LVilW+mapWV19M43Qyuyyvth0V9mkglFBCUQ+6gmJYQ8pVYwPj
e1K6U/XZHSp7VXuBMrsSiAUeYDri4xkKOdPil8i2UxAM6BUPkQij3safCGKMEAMGHGPO1amF/7ZH
vWqdxP5oZJrpxPt4E4/EATq5yus4ujOIS0G1yz4qsWcaUIrpaoJB/J+8/gVMwfkR6U2nSssC2h7E
ET7w75E9YqpryHi8A0aaorUG67urKB15OsE5Tp+yty02xkSmgyXm4ecQpBCeIEiE3DI9/ul1WPbI
KITGnY/MGbxVydFTbSvMEfuubC6ufvOVDNWs37PRmnwNoW3woSe6PIXTnyud1vcfpJ//AOt7IBOd
87PKt/noKvb07FoKutwSuR12Dpe9NHKqpS/ptN7fgGSBC+0MYrLVaM8FIlfWFzXucoiQUCd4Nd1g
vPVKBu4R30hmGkHMwdOAZ6sZcMmxUTE6FsOIMwCMdZgzYAuwRra4v9R7D3QJ1kzIaHv9U/463gFa
oShA+KXNQa+19vjWw5grizZhnFZNePKSgPF90yIqYGiQCu/3UkNxQlod0gYVKCk1BbJPDGiGQOXY
mdMxHc8tdlDr3dzjPi8IaZC2ivduRw1w2dlmCV90MEYOMGRywg0p9EMG9VNMKf6KvF1z3Nr1txiX
iz+rmuhO39W6mX+8D0kAngm9McEUXZJnoroL59B7Zv/YeuFBgTaW0j7XE3xDDXb1o6IlTKbNuL6x
r40w0tAcgmXiCeB35tQ674hrxgfUFNH52oFBzvgi/jBBgFboWYgg/AuqqwL4X/z3DPkcQR+OCADm
wbFaNDxzB+jwpVEJ62dgsfk5jHpSaMrvn8mcAl+I4Ahsq/D7ria1TAkLaxInACGXruH23i3v8xPW
LVwRjfVIhx+koH6MILWHF0B+o9RFuXNu+ks096Ljyv+YKEVdWxsLL6r7+1LhJXNvLh0ibRRhmWxC
0h0r+XYuO4llgWG8kelXa9it9GSWGUfnimBAEL9GYcgwBQmiIVPN5gEuuatBqeobow4M7L8HRCgz
TTfmyV9K8p7iVxef0VkkBIhHFRN38kqkgoDYahTsQDe/BEhqbm8nvjfiFRi4+Ltliv6foz6vzva+
//XfyAKN1Cd1K3zHCkxejZf/I7SJhUfwgPNJA9cZn5T+QbZrG7yg//d4gG2IzNSv7SJAVuFEq3RM
Xh/f0STLzPvI2O/EkP2Ve+JWwCVftvIe46BffTj15GFiz/WRxUmkcdEiNvNTlUv5yrhYI7Tl0Vrk
P9F34Nhg2z7jYqfnXWn4w63IBoYhXXaLi7sAxvrvWESWGmwYQOLspfvsIjrPofgVpnZ3O+9y0ul9
SKDAg0gz/JcrmYA/cMHFB6hM1uZDTbinj1uwsCu7nNeXppjXsuLC28dli0LGgZvWyi2WJZGSImHm
B5ZmC2l/n0eby/MHgcC/E6+SZbAdlpb3g+8Ab0xh2edCkzriK1c6IXs5cOEivgSPQ29ny939RqQ9
9VLGHrKE3BOw/UgLqrqu4UWYxliYRpfcNFhUo8WQPL1qXcDbQlibCmkt6OgRIVULA7W32bAiyqzR
U5ckM0Ct8QACGn2rhORrTzlOiZgCEvXL7lKkZaceJD5UdcJ/cHxRsjJ/XFs6i2H4+ywv6yguKVJ4
8HM4GMiVuNKYYb2ib49/QHPEw+lkqo1RK5t6tGKAiPDa33snVUEd39xxRtUsUStXHcDFaMBW2H8B
6xcmZMYoyzwZ9nYV3i03QJ2APQwp9mhWGr3kN/xfNps3bjMJVO228+pXHjJyts3mhZahxMU3gIeV
E5q9yd/VKbZA36M329UtVz4CfGtY3NwEEpNbq7Sh0MjOc9/jbRSPuOdix7lxvvXac62IQZWsENpw
JDIlvuhu5GQCCV8q4x3kry3RJSQFi938vAT8YpQW0HwoNL/1h5l+lUavH1e4x1m1oOPfkISKKLdc
Jh5YbgUe9GkX38+e91fpj6s4GK/sV/k1dubG/0NW+w5jQ8UdB5dRJSsV/AvCLOk3vUSbX+F3Lb54
wukbf3bP5jXNKlLkEp/rq0xrphIPT3TrFq7+8c/tESHDjrWL8AVpkzr1TEu/N0B0k4Xg/UIWROTM
xN2GxWMTXlW8tMSXji3CNefDxhZpdfpo6rfzSggKqMRarslN07b3gxaQ8ujwbLBiAJ5QTsCmi7Zp
gwOYaP3zPXvMkmcEay0v7BeR7SYP5I1vUkQJcFE2kLnrFaPsvJ9O+LhHZDjWvY7bBpGYSawGsefm
+JglArMTAcO/mIJ4ZuZyGU3WXYfAr2h3OgWzWkhnTsmhLPk6u+6YMi1UIlzPJyE1/jC50wHDZwBq
6/tgjjvhVDH46r97qH1+AERbBX58Jtyu3Z+QYdHyP1V8LJBgCHbzB2OmXM1LtxBXAXl0wxf/9MdX
+SQ+1eTSjceePIMBqU63daGMuiD4voQwy//hh1A4hzVyB0wJnTJMgjYnFZv0g/VUzmWiMCR+Fvtq
0eRXa28EQAVM3JrZsemdmUucyNohLBpyk7rACoc6blSQi4fHZjjqgGghT6AbVFeNCqKvQy75AyPj
ITNGlqvFbCUzpqBCrH1eLoq9CDFM5nifxcGjLZXmUcG86T6tYTsggAboPg6hLL1c3J9lwNRdXoTM
QKlOcsz+p1YV7TLnMHuoYf0YnJLjfEEmdkR8Xk2QowvOhCDMfVwAMNklQwq1qp4SpqGUN3hq7jkj
JNb0kV+MHS7xLUZhpTUv6rwU34LxQZHsHhuV8oUL21+he0rX/jmB7PCsR+KAkTyrYHsC0w7iBBM2
6iJUBF1MPLqCEdT3ByjgzCxrJVB/nitYMul/MYmyzo76tLKgUEQM94pmtg6zgRv14aoWWV0FpQXg
KHZop8DbmlHT8V5b27nzWXpP91SaAv3hHpYadwD3OFh/2XaOmQMqWLR0a1wPNUssY3k2t5wlqqm5
JKDveRd6PnniT+tIpgMZnSthmNxou9iByG3qWW1rggfnLD/OuJ4y1PeVycbJ0AxsI59If7/em1KU
clCfOpfaawCKJ9SevwcMEIDvLuN0tL9mqTLfhDB43hhpvIZqzVIp3D3hERsaFvvFA9DmcGpJc0Xp
PYlmi/EFa1oTV+DkF+o8OPcUg1pxzC17tiG1rvoxTVgxE4nt+XmPPBdkuSIpFaPMBSDA75ZKbyve
6QskTj3piOyeIOmSwGCBlehTGwgp3b9l80ZSnFRV2pXaDH6d0F7Hw+H5KKRrtXLKDg340i15NopO
zEk6K3U+NsrfM5yzIIH39/idnSoE9VGmMoM9rebefQHwOAE/OSmGK+MGc3e+t4Vd/WoY3AVQo9FZ
HFiLLR6mxZRNjbIjVLNBXsF/N+KDw76+fu5oBB5am+wFR3tWhti6hmCrm+vWzEeHyuvACtW7+H3R
7jW7eoYnzZNtlf1Ob9MPCRBaAAhjFuxO2gTldSR7K4AxsfgTISelc4K7LlCb8iKw9KwTF+PsliwE
xzEe73wmTkiYn8qMj3v7+VogpymX80Dz/ZgDznOm468NNm+p9S0KSuZ+Qfb5MY5oA8s+7clzCmOs
1/ewyqMKCP1ED8vGKyKeBmIt98AIeXC3f7/Z52V2jF1GmqkcXVMxr2AMIHDuO5KexNgd2pDn7/S+
B46H2wA+qOCvvOI+rOvUsdhqlidZ3VEFKyeu1L2fWOGr6s5kXN9XEUsD5tJ3pT0HhELEujoIwI62
PlsmkAbNf6cymt9fakvLm2cFUMBFSOwpvM1qkASKXtrGocCXf48L7YmT4il2O4A5svHRv7fTJ0au
STrJdNJ00WLegSlvhKOg86J0yQy+NV/+pGtH/ZzragbWLZX+UYWihFcSkFjbnuQgWGXzt/6RcqET
zjmNns/ZjkNs5AAcaHOIfPkLXfErUqKBpTsnC2OFGdTkhGBOFmzJELuBV4UDlnwgBib+txVPIAFp
x6fEhQu33Lys9KlGGiLOgx99AKV1/517nhgXzeLb7UJ6+HMW/XPcv4OD6r+XbDioWjUGEz/YfIw0
+FY4wGkRCTfSUvW/W27kiQAHgLdKFjBFV31hqVG4aoUmKCW3ecyeuvEuROS7Nu14HY/esgp/AZEz
NAjlQzy+o+/y73505UGx5kQ+Nqo8az7gPe4TvsW0jZZjcNdamXxLqRt+32Cqu7ibx2B1dJ9Xy/Ls
o/8NU2HdNZgZIeeeIEY0wEVQ5mIfga7FgSoNO2hRIlo6ak9HwLth7fyXg/6vA9kAVlmtzveknKQD
HpyQgLS+Me/jMaxz150Cb00gdiibh/SuRStx89LBCq6N4swLnqQSG0BdDycwiRsZSk/+hq9JunQ6
iOgdIlB7b7+9L2QY/oC6QjMUODN4i85JnDCEeyHTFEFmPQJf/+Rul2iIQ+42z+RzoqXIbK3j53pJ
FHD4D3S1lF9q+4S3SG1UwESidY6aJPP1JVLbxLq8qs8bNCP6vcKM50sz3GrLh2zgDzbX64oIwkEg
oq6exg2neM7SNtEi2oCQcs4vPQ9B0ioX49Dm19bC0UcoFCl6Mv2gWTcsz2x3xsEk6SNOV0EYMOjU
GIV3a/wmiXG3gC3idISt8moI3oI2ZanV+ijXXfydLnDA4COhlkFjicYWdOpYZxqzh4VyZO65gKms
AnuZLGBWl+dgM4/eJ0r6tG7PgTM3gpL8A60uIDgdiRMipaU9AbVffjAyHEGjs7OWyYMXo/QtjdMG
BvC2o2kbaEtA9WjFwpFk74PqJXc3Oef4N97ngnCU8+cjJhiPq9p2V9AbWykXh5v0BSuwmfSA0/ZF
WvCuq42T1XcMVCxUYOc1aw/XANBCtzkPzogBsBtX2B75AKkRwsZmh3WsLw5huG4WhwHabumDfkXy
vrMvfVhULYE6GnDBYPGzlLCxGzrToI+0zgK71xP9Bdqx/rfYYJcYKyzGCh5JZLD1yLoSMimvc3fs
dwVKIEYP3NlYX2S1f4qj/XMxk5S4CMRtZd4Kly4jl6a1fNHaheB45f/lCpSP6Z0XbXBgEXqVsDr1
chmX2Jvx6J/a11naIU1d0fUptW1c+QnZubloXNo38/yEaV40FXM1plPpKbAcQIt2cIpICOVYeLPf
bzvE8R9M5coDBwGuGmzIi74dT8eURmEXH7l+vyrO0K/PIsSxNIE1VRKgQDUzxzEpAwLeT/DnRgpS
J4/6ZWshnaoB2pD0yyPhQ5t87XaNlRxq2WyqD8Xk/R7x3D2OLpOU6c8zmQtnnbEC5PUVOpQKA8qy
JzX2W9xOt7EV61c8tMm7g74xQ5/lX9vt8ybdhAMZkH2EsOTXSZzDH7fiLc0/teeCF+KDwUALEmF/
vB2MJEYNvEk/VtK/3oDkRf7t9WsULI/If+WBa06Mg4l/IcXIxbq58rNqXOLLMzLNH6vuznbspurh
9KGJh4VVCUFLj9/HMao8fUUzAWJ//38MI92euC4Szst8FrL2V3uo8s+e8IRMeVG7qL3PVIAhW91o
f6txqTbwrZHEO83QP5bjfjaIyBVJSuYyNf4UyGSHVEuhWk48Njc3ISipfxlGjIeEJzsJujLIjX8f
EFG4KCbuUQtzPyJC8C2mrdvd+OpLhSZXKo/LUgp4RQ/81zoGTjSwr9cBAZ4UZWa3oI0/EDsb5iaR
KHVBpA+q/cYNb1WL9skLSikPqdGDlaUrpEXmbo8o7X046Ynv1FSaGXKPVkM5AjJJtfXSn0TpSbia
CNSF4PrnC3ab6jTkqN1E8ygDVYNJA8J6Wbl4haGE1WL0+1mzy4YD1sp4dAnH1Rslf8rWJOYtW259
mWMxVmR0QJi4mmSyW5U26E9REElAg3LHbaXRWUXfOllt+LQklszYI4YhgM35A+ZAUM3fKqL2MZhA
9k1x0Ajg1ltgsKRkFFOFt93E/CFRF/iiGhojUVJ5ZEBJIGbAsJ2UZx7eRcn7KGNmwN4wOMa2SGqk
np5mgGpPjSpaD8t374SXLikdhxjNmtyrjQkFr52YhpUHfaI4WyXHsXUtzxf5AWQUwVzEvKiaLcYg
m9udlAh8wm7bmmKIcZuojkyVdb4UAA+WjB3YqqC7w612S4/RUDv4LteCn+2RIJz8d3fAxbw80FU6
pfMQyO33TyMOjc8TdZxOXRf6rsijjtjqBdnSpXYdCPwP15U1CYBQceQ6u5i20QwVZ/8jWKyYMTUb
ttwCD6Eqn1zgHkrqP3dt3T5/gMba/rnTEPYHMqdV9u9k3oNCkED7gNXX/Vm8ap/41i/52f0njKjP
pzptDg2tkkQKMk93qgs6jEdeFgLRdvzL9ffzxkKlJOAa8eGwKbkZ/ghc1+uNetp2ljbKMjrbUYvf
JCmsV1LlBfCyKlloMeJj9G07hSzmXZFLQpH9+l1TA9QTKFwyApp1c1nDtn1MJhp4r6kvFtYxeyQg
RcHWBEWdZjkUZV13GZQWilkSzO2gAk9RwRaU+LxCY4VXx/UGbRW7VsytnwKweW7hblvIdmcMnP14
iSsLty08uP1Erc6/9uTWvzUr40tMOHOWYGoKJUpPw7OTbPoTESUq5kZd4I1Fy6DUQ3t3cyB1gMYh
Q0M0g/Gv06JoMCJZ3pE2K7cpPNNLENjLabwBonz4J0GCPJtAVUkJcR9Wnt1hlv73jyqm7oyiWetm
8HZKOrxWLJoyHa6VbGxY4o0WnYqod5TEtBevqy8bQqsI97ZFGfXXLhPU1AIn6efWX6MyKGfabjo8
f99Wl1sHEFlJ08oLhEQCzEbvmGeP4f0/xvAma6obMele94bfNWt47XxO0hRtLCvi9A48yTecBXl5
qNHNPm6slOYOkxVLh4HMt6e06r+5ZZGVe9Lyqmmxl7eP5gkFoDGthD96QqFMD3gAuB36fs8s0Gsm
LCAfG+U/wyJqaNail/qqR2sJTZGZGF30HYU47FRCbhtgZnrWG4zAaIDe8OhHAUIpsvnnMR/MpQuc
mOgQaEfKyfNlcAvMY3sojhp7Hi2wsQl1kRQNYLTTQezc4WeiusC37zQc85zjwjoDb/Yd7JTOMOhO
TOxI9yLeStvDWj+DAgp5ja4Hk9E1/rYRaC7Per5SnMTYgRPx5GBHv744V2/ramWJV5z23Qpogxn9
9QyuvUwXs6BYPthuwOTqo9ZFCePQXY/2WE/1nCJF4ii+QkAx6ut2UHaODRDcbHKUmUhYMKJaCC5J
3ortUqOKjLgxmnJfMPtymUBWfCqcRO/tjOUzfOPiAZBfejv9d4hygcyRsJcxg8U5giX3ZGJzE9JH
omLa8ScxUvoMKyPnFtOMpY2rWihsG3DrIQxmkXmh1ypenrEayKngu15VovTUvrIgIa+MtA3sLPgn
GgXwvDZzAKZoaDInvvBCzgoc18/jVL6RHcVqCkCVTDhN5c3j/scumiKaueDxv+401/M/Vm0lVjUb
C8LF24MjGrBiYxOioPsZdb/SPRbsik5LsIljO1ZwRILrhTqTGHPZ48lPJaerIEl0tzcGHKjLQaXT
rGzKBVfqTpHwrmT9k3GvWrWLHpPRY/0dDKBBiBDIWi4tw/J1vfl09Ej3u1nvAuAFOcz/otKlWzmV
sox/k9xRZdrskoMPpoXO/3GivYRDEic91ip7lOiiNm4FKE3CAyVPTIzmKV4gvbQMQdoobU7f5zdb
VrW0gK8A16hZ78/iQWo0slu7rRN7M7XjDQ5o8Hr7a2vsP3Milhaq/IZCHiCEERpDFiLarz836V/I
oIva2Ux6fG5RJk5DwGI84GCCaJHuKwkqJrSNROyaoGDyjnjxP4pv8zg4Cb+JE44GRA0dcZRvAN2x
FCd8tXJO/2mC1Sdg6qQlp9MgDiIequSKxd46nu/dDJsVsh0lH1KYlsyeu1gROkJrRDTs2ezXHVVC
et03QQiGFseqUirSp3FmDSKt7jMcCOEF3VGVnDKadBQSEOvERJmL3wCj7UhcMtM64Tfi3CDqrxU/
w7HnJA3UeVpzWnjMHUapuziOqQBErElf5jo6IcUjtDUTK4ytE73OKgpyl6sblyYsDGfkkdhBiMbI
FYFcQphnmkqM4c50Yyvu0pI2PEKgn0LSqYYfuwa1aoSOnmd9Kxmw3EtVZkOPERa6veNfoWXbaYPe
Zvxeo56YqSQSUitzjNbVmGU5lBBCmu3iStQI/sisE+UD/OQi9sMGcuo1CtWeTnVh0Q6ET4j1R4xl
UlODOLyME15F8fEpruOpgM/f1IPw/PmOz+UZrlcufHwJvBYbSbtp+KlRykzYzuO7wHIG0s+Y3DE4
A2MhHejuD1FAfrTWxbE2YnD0K5lWJ7KdbuU55tZblOo0PpYeMITVSPYNfe0Yg0q0qLJmLdfAji/g
MF3xxeTbPdyKQeuR3/aIocIBotz46XcC9ehYj0gKYrCVZ9VjpUG8d05fQqNj4eLS+yf+sCurPRER
9fFyIEoJxZ0qLIZrxCIw/cAlHmHceUI6YHpoap3YjX1uCHLrrXu8+NFzRWhTi3TJB73JRTsmkyjk
T++3ZKFgS//ZAcwxlmIj4fSiJagnLwMUBHRAGUnVjEt77irSWkimJfREB5gKez9Df+2yBcEzWdML
XgjfUU0RAfQzggYbi7hWjy+t8UdoCkI+9bJ1givpWFXAfIQBjYZvh5G87JI1oehchG2nmOgMB2RW
NDt8OT5GOGXE7YFefK3iLAr0+UcgxnyI5+c5FEAvLTu/INZ0d33Afcv4laayioxp4+2zPn0HWNBq
SPDfiOht1F6aQUdR6unCyJewzOrg5rAc8kXnjqjVBCE94+MmXFQW6N1I1YjQnnL9IRiNXcnD1EDr
A2dE7k6m2RGp85ORmdywPrMUkHgQ9tSxIzQ3Rb9UY8ZUF+fyXDlEjdsf+BJ7ttq6anL3gnrIA6j1
r+TJE5ei2awIDJF3E3J7eWwZ3kxS2UnNDW+MDhC6npW82H6j/Ji0jfeK+FwVwg90T7AngTJM9EWg
TV4PSSRgLGrHoBGZXkTU/bfdBTirQa6MyhTnqxTFPAAvlGHdgu4uH94Kv60rov3ZHI8R/IihOl+0
CRKhPV68F3Ur45VojSJ3W7IetC6xiM9z1aEKAgL1M5Zr6qWm3ZttoPbhExI0aiSz3X02VDlWGlKG
CjvgO26ZTVnU3zkobXkXOif0KD2AeXU3izwrGwF3e5kefiwh0dPG/l5vk5rQ9K3FzusG3rzfzyuJ
fJN4KreOEaAWNcDryviLwCq6Grv0ow6ip3/DmTxy7TbG9vfjwkeHF5SfkXOvCUGGcxzs2Eld+Mzi
G+0pK1yosx6e2Pfpv06zU576fKK6QW6o+97EATn6HGoVuTVjip8G/vIm0yRuNo5pZNl1J9e/cMkL
p96dgLymorHX3uPScz0LNsAuVlDOvElPc3DJxn7p7T3AqkmsXW0/n51aakWkWJb8ohfU5aeYvBvb
T9X3AoC/77yADn+50d1IEyie78NYyikZUPNt190E9W0Fgpgdi/VGNNiUx0CK/nhCWlvctOJHjaOP
sEgmGpn8/NIAhQHCdVGP6X15z9NC9E4HVTclPyiIvPahvguzM15JiAfFZ/qjZ4Hpz9cwW8LnOlUH
BPusvEaT3jvbVjBT6STuLTDUa6vpxefOOvVGhBSpvvLq/DmD4NjM2ydTHn1u3wM6xlW8usK5YV6u
rS08RdnAil6nbN0+xiX8H6bfBkmAH5aRXREJSdOhw3dxanzrFhsUPCNsPJvjRKCGRNzfy3lKMwfx
mRJvmrvTnzP/Ra4eY2uWmzE7qwtZeQAnqa66hg1gNl1+nCJ2R5n3eUCM8S8qFkJwqe495LPDiNFx
ReP/3nSbLosdjOuplK3x/p8KN0C/Pli5L9kPTCSVOoDX7zq4YE+GoeP+rW11T4UomaoLzz/1OWN7
s8Qdg6VxyVCGruSM1GE358QZOFx9Z10iS7aHtItwqF2XM4sHtfLljXZtPRLq1eMcpVkxfus7oX39
olccj7sVpRU2/o3oH/EJdKMjgHcjGgRZQvQ3dap2Qm58ajChjwZPE80+5nU8gf1FIt4DDYDpwBcU
oYthOoJqUd7R5EX5PC+RK9GXFPjclNIk3RmooP5aqyhkcpVYFWpwMqxq3ZYl9YTqb5AsTMag/2dB
l2vKFRi7/Y0wCjU3o/ConHITmtB7XZLyzKD64UHPOPzSctziImDqiXyRooK3o1J4x2Q5RJqnH6Y1
+P7l+Up0g4boDSgk45wr2+31QE1JJ0w3F2A86Uy4gXCHleII/KoAyOAmf+Nvt7yZAjA/AWZI8Iwd
ydBofIn1RcsaW7jyQsiuuCRxMoi3Sqqt7PlSLFyvQOx/9CpCxPc8fWj9DbPzlgu/RD+KSj4zFmWi
yM62svuGjYa9ub4pHSJF4gpPjMNl4zx97/MBeEYFxzQPLCr15DUUz0hE5hZ1XR9v3PlF6OlcuSHw
DYOYr4PVRg3wjTJT8tNm2kLnwJfTgG4xVy4vyyVVRWMEjwzCiQQ1BI27KCheXeC/x178y+ytyxDv
eNW0v4Ro5TmwBpcThfMIOxV67pOOP5WyK1c9ZSUynbMEjiSM7u/AGH+StBIDiy/EJXnDb86AMNA+
PPGTLwnfIJd0IkEUuRpJ6UDfCLqaBdPI4wS0W14FXtJKEQhW3HclbXJlvvZn1Ovz0LW1NRInk0xE
AwLnmIO6w/8ZgndYvrSnWFN5XadNfwi2rK3doyPOFP9Gg84DrObYdRAmFt5mDp1zu9epJj3YN5ZQ
B8957/UqquOUApIxW5awAhWbDxFI8ZvQPoz8kXRK3U/iVHy6zYCY49hVUUS4GjGdBM1qDpIMrlUa
sO5dWyJ6SDAqJtM2w6+NWmWu/FGjUHNnMm9Z2VRyhIrZjzojwWxBPqHgHL/G9GledvYaCjDaxzFs
HCpQwQdZoGGcMm0ljMT0ohUEFjQQ3d7hOBSonIKRu+EUR+vHO4eym7JC923YL5pIxy6Xz83yDQdy
oB97y1U23i1Lsz4EHxs9MssTHiql80CbJIqBj55RHoLd071HBjeHeHPlM6v1cKN7xgXosrpws4d9
9IkT9ik9vkkR61njzKqZihfyxSBw2k2Vm1/Dejc8HXtncf//xf+5mQBmIKw7t1QXtipVtBXIwQK6
PpUqf+NTwVRhxaORW5kevuFgXlLvNPx5uEWSqj9eCCLWb8YCbB/d37B4De2MKA03lCNs/vfTmaKf
FKeaMF6ktj4XMJANUE0N6JeZ2WylHuQ3Ah07Tttu44wDNL2/A8mtO4SDkuXFfZ+r+/ym2f16J0op
Jwepg68TmcIqFRGUa6hHUdhXlQ6eXrz2Mc3G5E8MKSv+WkieVcUKF4OK3Ut2MiWxnA9X0shaGfnq
e/4OKtjBXS0Wu4xjXQrjYOw63VjhRnVtXV7b1SzAjlzBrWuIEH9f8SB3uRbCImi8IPDCKZcshmeP
2QFtjlAQiJwcI1Wge2vuq7cNeJ3XX7qxfOpXptNhe1bFMlXitiz/9f8p/BhaqJ66fyoSKLDL0zFl
jXH2Hx9xKeBz/FRd3y7YtLjQNxYlI18wS1sDe9Aq8ydVBxxd309WMUC5rppC6uQjNeOwaPuGIzq2
NQURtSFlQZ86B6Pt2JzuJcWOA2jaQ4Zf4EQh/M6Wft50V831SCOF/wfHt4IKg6WHZtZKV7yGAEGA
0wMmu+OUZ+J67S7idoXs9E3jrUA+/9+70CEQLIj+60gwW6VVbsSTUqYXE7c2Uh13oIgdetnmwqR6
rylXvyzhmE8XWtbrN3kU/zVggcHU8bvdgvLi0Bu57aYFWMLvJ4ebzRfdGzvr/k9XGhUdbmyb7G1f
cMU7xW7afA0nOwZZmLZ380yNhwhWim1jdZ21unBUP7SwjAwqPiHgSnNMuaW29rCeu20ZNesfQsbX
Jv4pvbWqXsjNNw26YGvsY0DDtt0qTdHzjX++DVInAtNVbgBmBI5OcjKPnbYAq952FPGyBxh2Q1Xe
8mpE/O8Fmzeu51aaJy6jDqEIQnOjSOZX976JZs54y6OkGYqUoz//CGq4TOBTtOW33H81tOFZl8aL
AyFA7OnU9P6CNhJtW5gf8PSERD86vye3hcTIDRD0C1RU3WcYGOqd1AmSnnmZyh/fIc2YVoC+G5YR
JcI6+IvsMFEYEIuzZInLXQwACGVKh0dQ8+H9et8QC6hc11dg5Rd1JNXnif0eMLTGcI80b9YUqy8X
zmRlNgJu7du9l45h/Q1uc2a94569UMyP08dLpXB0ZLameO9XR2D0R4TzScGJuyKwE+Ea/pFc6XMS
HZn0hoo7y9Ymdx9vL+TNCP4qSS+EpQVDfNhVkz8CFmaFdsSVGNsNhL0D9CUdnxazi7T2A5excSsU
GNrDdULytuPXmZ+VAOTY1nqG5PrJIfcKtxFuFczIRzkq93IGimffGXBFmyuaHeXYJwtMC/FIktfm
Ta3S6cY6wyCdxlex/adPQW71hiRwhj9rdiKURGS/GulHJCnihCJyzlTalKCNsLs1oh+oGxfYNp3K
TQkZoKVp4W5zfcMeMMTqXoaaCmaI3JOzE7644jwhsJr56JnUIGKqMYsWTdh2c6xoKbenZGBEEJRb
cvMR/jKknO9ox6jMWKc/DJbBVIB2YpKLa8ubkqgrqgzAHO7PaU9mlIh+6hSVbh7Bg70/ernmElf7
AWD0HEhBAyarhtAI14qp7ZsliGN+3LmElRmv2MEhJSoDpmVJ0LMw1AFcR0U3bRSfLgeDofy8L5xW
GBiFn6mB5yDctJjmn2v/NSxszjnO/KF16Bwt112zuIKVExSHX8hMTB8qMK/HBnwlpjYqIutZW8w/
aaemB2dwhOUBfDrDrg1xhqoD9DGjHyUYoyGo+wqDG1iwqbpbsnkvrQJW6Vlc4RlWrFO/IBbmteHh
zIUci2wPh1ybBovSAgD130Vj9M1SC/k27sdToW+khXlLPOidvy/yqUApnvOnxvki+6OWuEnrMMaa
CNs1HLtM4j9M9kg3mXU6uGRrQJPTjw306lgklaWyECJJ+hNbHoO9DlYvfs/Sph/n/zz5eg2eOfLG
i0sBo2SCsrMjKrm2w4rWq5jE/YxWjgr3enBAlmUXlKUe3J3eaiwCFYN780u3RVLzyYcxojhb4HX7
sqiE+GE/NVlYSjSY66UgDJYTcWpfuL5vBe/1e99Sd2fD9JHT+Fg+ZzNPC8sQFlGDe+WCeG1+JnN9
3RpIC+yA/c9pske+Dikez8GNmCV27iYiMFL8uh6Mtcegs6d2HYELq9IKo/sPUrsA/DlQ44ozWYe4
kklE2TTKd8s1a+SVdMKR99odcturHtdZDFZjrxayHKJ8jzhkA+XO0Nt3jF8WJ23HEewNyXy/mM4C
cHQOL7VO6xNVJZXFMZrQ3UoaoTKg4Fg7yzekllVfphfQNWhSXCxN9VPzq3P9bvxIVaL5X6Wxr/yV
zyIrtNYcidpg6sPwhBc+pmDtyx/eJaefOfkTDs8LnQ/z3pR+pwcK0xaj49h388T3U4WfpQKlOY8H
A1mZY87djnjIx8QA4C/MpVdQuXm82KJa2CHdIwKJ9KSJK/8US38GvFbhumcy/LptIVydEzhv33cw
nDS/SeOuk/SG8GcLQo83TGybkXK3IxtiTEdkWSBTVLbq6h8ybcC4DPDeBTVYSZFooXDl/BSrq7QZ
U+u4V+ZOXTWLl7xvB5dOpeaAMHuQw41e5X4m6kiFjaP0dTCLts0tVzn2ae4aLPj0iGPEG5eRE82j
L9BY++EP6bQ+3OH7AcSPm6ZXl21GDj+1zEQuefFqyU2fnI02GxOLXYD+PvBBPTLmECwYMIRFuI68
Mtwkch0+JHVnkNaEOW2qw6pYTgs2D80hHL17IoSrcKwR/QlvytN015469Xd+MCnTGc+zQgm3rtID
3I84TpVssFfvI/bC4PWAd8hKtinB06xZmeebtvRMVofk979mexxndUrZ2o7oaiNqnjeOPN5tH3Yi
5sgSOOU1JATl7FzJ6drFJT5SU/bYPUW3I1R9TbP6fT/DzDze5+RozPL8pOh1iX6E4lAqlqg1Zizu
nQZx7DJQ9I6DuD/l97qonqgh+/upGskCpk7/86wVx9Vr9SDna7DXJkqMo9sl4yT31FizUxjsv7Vo
huhOumDPdpnkC2+nrFT+ZPg+P/b76OUFglpHD4Su57iiLZod+nmZ/W9wg6zNoLhY1nnlrbwnA6bP
SZyZQfxi0S8Q7y7SlVDm9AWTbEchu6A2b+ojcK9SzcvB8R9u6+KcleOqntsoxE/yRjlPc5kXClp+
dl2fMo+3ErSuoY6ZHA9B9fkuj0q21NFONI4CBOA8ufQc/KChrZ7W2k1gZ6CJ3MfF8nrM2qWCc0sU
8mTo4vJPVV8tlZhtpk/SK1L43T9M6E1Um2na3rEteo4EeGunmZzEQPLX7i6xdLsMf2TKxbOhkf7K
kFNslyCfCiRcit+fEKP+zAyZjOi9Qdf7E4iznxFXe4pumKeT9bAiX71XSeXD+mRrfXrna6H13/iE
rrB/EsnDZomxY43LcYbCPKkf7fkEzv80V+jj+NryBouNgebhOEfTIEGnCq2vkfUO5KP4AyrAzHA+
x81beafQ9O/l9JImGUTBTNwJHEL15KjcepSzHtXotOIZzk5cVc+EpCiAvMWz5q1NqJeZPxLyyDCl
v5c2wSTG/UTrs1tMUKJl944lgp9vPFODT+ZtmPgEzagk5Im4ws8D78/M3feMjtHO6bS4VPblCPMh
VZSa/jl/QWD+r5myON+sSDKjSkUhZGCk5heRv+Xf7zHM9+UGUsUJ1p2KjxJoJXZPFYqxXkucQvFA
W9y3pWok0Vr57lj8hm/B+6yiMKmt5LOEUWk6fFRupnjlvdRPkrg35+O5y+EqQZBh8GIyj7u/gllF
8aef0GnsINqgWsBQTElJxqaFhKVnDV2pCgY7hkrjVNYUcJbIB6DyK05w54Xik/zt2EvCeA0aZAY1
BI6ZJBAAf2g+XZy8jwySXfE9sgwu6ozJBrdK4mjx3My1SLt0ggEACnlPOG86dii5czX9buAAcFUb
L8AkaSKuhdI88n3LINd5mRmky+w5ynPTtOBqE6UnsJX0lMSPn+dUGZHd/KI9qFjnXpWc/EdzWDlD
XFUNKfA2PyHU9vW3wepZk1ShcXbt/ibDexMFrTEmWHZJOgXEPgB+ufIUXjHszuVO8oOK7bBaSyTC
tfmI5zU9VqkG36vD0F6UytOmAUm9VPcbuZINxns4Q/XRPYbf8fwfnU7VQSqF3U6KZQAt/helXsGb
7MYqRyADWoe4uNmRksWq8fAGqyVw7aXnOfxTXDoTyNbSFt4vOSi+l1m2HvdI1iiNp1cJy3G0jAfs
Xu9Epnyg1BOk/0PEUTqKHP4SWGyUiodbXfSElrzFv5DQuwuO+DHpBQHi56lRCOrVxFJ7q1/kDqVC
Ibikmp3+2DHNSodu6yTDSYAjxq2BwBe7bNNm3Nw34g719i2h5l+gU9zw/F4Gd2QMZmcLYtVJtyqo
HgMwzgVUhcckowGwmR1NqyQl72LO5WXIzWWl9IV0HBrZbqx461QBJyOQhrMcDeKI4AsCkqM6xOgx
Q1eRBSlRS7XDbjTTeImjIjWxseNe+6lne3Z7Nr31F8ee48o4LxMf5lb+aw84JFjoRy5N+mG3FVzU
/jiaWdL65qypxnLTuxorG8/vbavtQwKD/rU1F+TYlJP0q4p6b8E5iV8hqxYcNfD2/+43NY9AGuYk
6ccKAySX8jwg1liVBaXBx7noUVbOk0LU/1q4Zwd5GhsHSAGe2qKm//q9GOOuAOYBPcGbqAMF1+PW
jcg2rsA0rPmuAvJpKEUTSeUjmP9jUt+X1qPY7r9dDAMRYpRe9N1qhFPsUGhOFTLXwkP9h5IC1EqQ
1ZKZ2lzf7htYOM1ML24xPirD+cQDPpFFmSa/fz6YtXU1orD35LoPx9tZbOF0ZcpRmdky24h9DvAB
rJa6q9Zni9ROdsIXLM7eKCuiLvu8mag0Y1x5SSZpjk2LJaiC1FgOSt1YjJjM5zf48hXS/jAFVaae
e+tJtl5JaBqu1q293PZ1NREagvPXPegpafJyyCi0QZ8YdLR0WShWkCtzVNE2FEpHUorPRGqx4Eom
LkWTpCc8xl6dM9fYwPQmffZiz5GN7zSMa8W1K8FcjcWDX/PuBTn5SxLX48oNdvd2law0dPhx2I22
TmTtsJerr6E2itvFhhgsEnL7VIGqHdi4uTl0GTJhWm0/bOMVROhKC9erCzKnJkwNTSXd0y7jkEpS
lvN+6i2eQL0FnaOP9VtkvZpmDK579DDmsHCBkiZz+Z8vfRIv7YJZFVtb9xhg8uCujz2Cfnxcw7Gf
BDiJoie9wF7yV89xqobxWj7m6ySZqcDzqdYWpGLMIyTCpHFn2DYYMeLq6O2zo+RMyJVV7dWfMK5h
A18pFBYYMdCiEEyHPYY7E4A4JM8wGqMJwW7hVl6eNFvS/Mprh7XlO4bnH8l4SAGzvEH8fWB8uZCS
Z7YIucRpKfcXGcIBY2kgxeYPVI9gNv6QSqhegxTQTPnRwkcPgytxoq1KFDtN4Sjlw/qa5EJ9qGCO
oo7h7Fnq1lG+tsgRE0DteEGgrlRzUXB3feCjbqGb0IF0KZ75VXazkW95zOVEkGHTnVvX/LITI4P2
FU8E5i3DM53/c3QKsRvrLVqxPdrCpdfrdz9t9ay0fAT8Buw40p6ZBpBrjpfwL23R4U3+GvAUYSA6
9dI92fWuu+oMFy1rCJ+FT+kTsE8JYf3KSHNMAbMubsqb9ant61zyUAiEiaOTLMA7znIHbilumRp3
Aovf9CJnmEaG/2nLEAggEt5KHTXfZkKcRZ0e8PWiAm7MS79mP+idyTv6M0Gp2+z/lFFXkw0BGZYt
UvNjDzrYN8NNXnPHvI2WfVTiwN31aiNsIiYdMytKupI8844L6m2Mh6ozD/cUk6dKVHLgkMEEHgAX
qxcx6RT/Mj76Cgl/pkzzEH7w1J3vDQGbNsx/fJ+95rrT0J8h1v+++mC79dKjMuTdzE4Z5QjgMcyC
jUaweNnXDkYaKhZ9l46xp2fFZniJeM/oLVvCzam/4JVg5UrpPyl0D6/bN5n+A0HVHy6f+EqFITIC
W90Tav2122R51wOc3ceJ4oHV/0ytSgoX7D6IWuJtWLJyt6gxXNb+9ftkhH6rUOQkV2cAUVcZ/O+I
5bvi5vIEaDemxPAUuSifs70b3qbDVGsuytgKPgwF/6u2Nh1a+fpWf2cZc79EkScVjTR8FXUDofe4
quAMv3i1K7ibBIGX1l3rmCqVNHupVPt3zzsduO3iqL3/nSCWtur3tyiTDt4X//6XIq5onMtzlbKk
X4tnja5qw1dg6fqW9QPSBx3Wt1nAagkRcgEELmUQUHVKrBsutbVXRU073hLSCOuoghS1/SH3B7q8
eI1wkecMpqmif4Ig0u2G9U8JSF5mpQgQKVU3YQV7eJbNRkg3CBEJGO6CUe+4V9IAjo4HaHa8PFVi
jJBA8zk6tE18Dwki3g0PS2r2TfaWVjznPqbXsD5Fn0n9h7PmDqJh6NcS1NoU7McvzApxYXEjCDDp
KEw+cExP+37aYWWhdk8p5QiRCm7YsgUlHMYSBwbBlOCUag2Jlw9DLfhq3Fb6Vz0nA6NQmnWP89fR
HhZ5d6G4vk8HF+TmKbdwEf6JbgjgnZqiUku3bkrET3yAVHLt8HKC9XR0WXjUOF97NYZlEG8uUCAj
DRepo0y8YQtL8EiGOK15/Aj5Y0jwcDq4mYUpz7y65Sl2NHAs2FgA7ST7lwUANl257KG0apdq7xxX
Ga+R2rVo65YA9R4lWIAPDOBdll7pANXrHWShjUVXSu1O7Pq+dIDa0jUgN9ugYl6CHo68D7kJz+Ss
1Qaq7ljCBRsqCvIvcVrRr4gUIZCgWKnGlNFkhvwAKU0krmk71be9HRDHg7WjbIIs4F7ago+3zmfE
5EucfDaH/wYvNTHz4+1lIdVcmauoK7K6ZMx/KpsDmVlRmIKPgnXzKm3QQRyT+SqyKv1NfNMP9xAV
cbopBOK8W4V714wNmvTSoGif0vmMMGJzq/6V499EgfWTcO6d/vH5lLN9Qsk0WHt07S/WQpKvJV8C
eBGrRC8Ge06ImsRf9wf7NDMaBCz1CMw81RDiOxnXdClaNqOJnuomWmya0Smwoh4EqtGKTu8SgYnV
dSlP4FMuFnIHo18/0dsE4vonyTm1GolbOrkRzcQwEpAFzoCM3mgwQfjU9N80oHLXGL9fPGo5yBz9
kyBqJnN9re+qe1DmeYMf1ohlvTFqKVnm4ce13bq7Mt7+pbia/CZ4u7eldytSuyAQtym5SeBUaCGS
f9dLTKsZW7PeBOg8jRNqAht0IMCK/mMyBu64wLWXeY1Yy62/QsyG28C4/U2jlxv2TGkvOlIkvBmm
Ct2lFPNgZAnXNUu9kkZNCcI+CxdVau31U7lJvPZUrlWVer1awYMp+KAdOOGVffnqgrw2bntRJx5E
bd1HOLkMs/Ib5PC9l9zjHjyOd9m7tR5hB9MxrdiB0olWR54JSzsUoUK5rtymp7svRn9Wd8ODpHgT
+/0wM0YQlfoeDC8+SZV0EcgWKPMnH1NcRS3dVL1M4vMm+79U5QIIjuLnCXQb39CccxiZ/ZyNsfeU
QxscWieZe8UBCiEctD5dvtBSSGzQg84+GM7mAlo20GIXmWkCPD07XYg5Zn8qvL4EdaZkT5l1ERpW
l5MPfbKqfzjeho3APYe4VsaKwZfKDU4m1M26Y7aq3y/YZOASbCWG6Oriov67s3AOPROTLZDvblnb
pNkpDLiA7YJa1cmH+LjnQ87dtkPi05XEp8uicTrfqU1JXOTlpzAQLsN+TuPttLeyYzk6yPRJcAJC
Qb3YKFT5wijEe5tuV6RBr1O/b21GnsXTnWZKoQUX0SPR3RiUEk6fa9L9g0SkusMmrHSaUFCeRSdK
56yq18Byud+QBsV2PtgeZljuX5oHKAlMraA2TPbSfE82paud4O2sgqYrYxhLVD/RSHLsEyzbxawZ
b2Iar1SRhM8wIOSvfi4F/Vp5CWBbE07VQW0J3iNDYopMjLjcSbwGcMT0cNb1Pzd33HR0zAY4NiGh
9vlsWXgUz8ssGI1k9A6dWq5sF9oKGJ3nyn4v7uD/aupPK1evik5YrMzwP9fpcT5H1Kd+mIkOky+a
+7uMmPUSBwIOpvUJ49SbFnSF+UIpM/3BxAyMpmDc/IBTHgzRbMpfzbS5/tBjfkoCTbquGuQO8Lqe
xG4KBI4cbbC0hvbDIeQr1EK7+pnmRkiPM6OZwwc8r7f3fTVeAYyFAbDJUL+I0U9Kw//YVsalplxn
qijOUE+AKrIHIWrHwHPC+cqaqKnNLiF81Al7ZmQkDsKT1j9QOGV6K/nkFyi3EPKEPL5J63tX9+NW
63/ws82wt2pDBrSxqXkrEylrYPwoOafvtstNewC20Vuy94mLtjszYD6tc1AjsE9EF0d4pLIzyPxv
5SqNkNFjTEhHabwjTzjpZnv/3eVsFIH0/euFyQlH+FEgyXY+rvzGuDVoGNluKn+zedIfWPEAMW/q
wkxtc2C4hLw9SgpjwOZvORjzfOAityY7DgTeRXsExbox6Lb6PKGK3dAc1Kw76B/BEFTmZ0k/wInF
zgil7W/f1vaXot9Mh5OGYh1STtCj9kOiUm7kvsKJ8sZHhwm0TOF3plbb6C4dvhy8T3F5wr6QbVeP
1frpWrpd/83E0R5Ti0EL5PZayh/2H4ugh6bi6DOK/LsIh2MNho9zJ5iixZ27wGzWbX7wpAWbRXc+
08XRr0liMcBpwCN1jLijOAHnx2Uk7+SdrZ9qkGrZCYTfrfjJq+jBEArBM0o5ZN89MYnZlgv1O5oU
L+i6WMnBJ0CVgRMmTOZSb9TGcH2MyKri4VYsH4HKGZqUHJKlBXAYRuIIec+U+t6PGX297TlG0Oht
Au5SQvFaRwBEGa92XO7mW13wWbpjXteLBpX8nrajxGyk3+lqkN+SPPLQGn5qyWHZcb3T7LzOSl1y
2hrJM/c8Y2vqtu55x0z+UcCkH7tSp1z7XJxhKfrrjN9sqaI7kRl+jBZg4nFl1DFcV7bBDIl8NHu0
99Hzt3f8MecWib5mV7J0mdzsTE/8LHFdKm+88lcu03WFK/wAco7SB9l/PfiRY2Jt/kXZUt9A1bpS
jqaxeZk2SMrnQ89k5kfrWqJg8p4OG3HaC+IUl0anaF5aeWVShsqYsfLac3KwoFErUnnK28ZeNqOK
VlNyPdQXPvEzzFx04QYmFJCoVCZBFRWguOhUjsOy1OiHXD0TrCnOob0cWNw0aCoZjtxhkr4oUMqM
2ViQDpvArYnW4b9ahMnAST/aP9IUrsF+iOBy0ewxXmZkCb3JQOndgWB9qr2RKaJwgD5mypgKteBh
60G6aAPmBpUf32ykuK2sq80kRwREvZe6x5/EVfr01ChgXXm0dCH2RPQUylwh+/W8Aq3v8ZQNzkm5
2pue4CPU6YE82rs61RT1Hh78fBK+Co2AK/wF4eBAzDHlMAvqDfLeR8gLU4yo9SowogqjXpJ0HTEQ
qZkMPmvoOgbvKwQLoWNOM175I40PLNFN9lxXHurbiIJLjnwiKsRlLKeBDN5EaONfp/BYd13/axnU
AWQbndf3Lf+KZFh0PNZSGX5o9LXKhjtZu51xhSSxyHeFgIwwy9x/BgMT5JG7P4odt76SE4+sosfe
5cTOq5/vdlmZljJSxfMZlagVwnyXcELEVeifzuc3aQU6Og8fh7lHc1y43i+e5df2dQ3yO5HWX34Q
I4OTT/31tCaLSk/LAi/WUI34/uhqXFzNIpLOnYhaz+mlBDgOcSLzR2/LBbOFa1LuMrggd7tNf78Y
S1l6bU1ii83iJYlcgdGIZnN0nILyXjQ3gUYKUrQfSzpopULQqLy0q49f8veLPGe3hUsWO9s+pbFQ
eTycJA/7Qh/Lnkh3SxAOsjdwhu/moFlqi49q3aT9gYEvBOxB9/PMusa7+4mPjB4VbO6742KzPSBe
moTO4dn19uNQc1yQmC3jx/Ns0gMWNcnAYEnLyVwkQyc31BRt1f0lBn9sSHwSlOkc0S1x114Lq18i
gxfP0V9bCI9Q3qLhlfrEC8M1rkH/2jIhMS8YVVohY6fEaeHEEFOQwnbnp6y+K9LpgOu9hpuSdPJY
2OcajtLSaGgIXSjQ+zPOxGL0Cb9MVltLIfUn/hJdUnGDDMzIwuQd+lwghsvq/mryCPUAEdZeUu2C
ObVneSyJCXDUkVGGtg+B7F4cq3vobvFBe4s7u+O1Gr8g3De0kaaGEysduEyKcy1ERIwj0Wg5fEIF
MsH8Osf8SnNs54KXF4h8pSMIzgx1+DDXl2miMnTl3qa88F2Bk9dGyUbB9YOSFg8LAWycBF+Vki2Q
HXZrheBquQSUnOSNOTjSgGIp0TFaui8bVg+f/ms3tWOApnfv7NVfoYi4FZr2TExNcccnaNzaeNvE
d10ObaAwA6YPfBvyOl1JkdcNOKMH6KOoqXPmBRxQlnfT1s/avwiG5VRNf3hT2DndQlTgQ6DO0y7b
fq6Ce6krC7jA/XMc1O7OG3Mhd29m+v30AJIk5lA1XWDNvuYFvAnLNgc4j9fJ8Qq2dY5zFOG+C0dv
+fMjFwgw0Chi2nK13T33ks8yCBdwzG1tTYn/PMasbT2Qbkd3kZvBzZULz58IGU9BID3Sm6SBFHbh
2exyqVwnleFgl4fOTD29BjU5G1RQsqnLeaxJzYWVYp2BYYrO4olONPrXOMechB/a9idZed18Vu+y
bNhE2WhK+BGGwjv7xk8IUQDAR2XysHc/ABxeyu/darcA5Gu+C+cNAWzxPGI3CwQTTCoWlhPDkG+G
qWwOFVuhJtAUxmta3Af3E9CD+qA9ZVSIfsEvTL2BJ1t3CpbaGTApdnIUxUhSu4imsMpK+vFebUcf
SVRQLyz0/9eJYRxeb0YUN2AtrKiKGYGKTPyS9b93DQ0xHnRL8PTuPPaxDHndp310/AemS0OQ7pXe
stMO7JaSIxsqarkFMnry09RMy82B521qJCUmGVUIvUaLL0LcyrbKw7xmtm6PnK6vo6vToUQ7Mboa
zcG9aiddfjlPw7xrAO1Gt8p34a+M74NA3Ha0bS4Itjr/D+L5qcloROuzM54+Hb+hWFTMG5HxBAA/
uyQMMgFmgZ9QmliU9sRzmnIX/1RjVZ2dd901dKimmXdW5djGlC4pMrn5nMf/4VXequj9rBZObH+H
KJqh2qommzWXH6+uqw3fJfR2S9LxYOWh2gUCRCTcGv7mKc+Z/jhdmEMkXkN3mnAxt274q3UebHuZ
qOgQhzLVSguJhmWIqP5fTDYRnwSUUBBaa2YjAl/N006bI9g4brAXkmMavwDtM021MZQuo/T7tW8x
32DKhhUIMdXtsOviAKgO1Gl2fAPlBzkrXhszrClhJNGW484XH/XvOCtHlCgXv5wsnD3KQ+NgSLbF
e3TavFFhGhHqiXKOVL+RyxMVbutJz5R5jSKfmJ4B0mB9X0Uyc0yqPTZcc1oAMs00bDNox69m6QOp
P27jkiNz7tQF8z7p//GQJzqIE+4SV9hv1/LnRC8uMCOzHDjqnCMZWWvIGJsFpNwyBvlOhyXKT99s
HW3v46Dcdnc31D+tGImySYUBe6sXkUNmC/KCvCSD/Dl4JSHMo6y2120C75ZPCD7vovP5WaQjfP9j
h1Jdw8fX7U14ei7h9F0chY9G6Tz1yZmwaH96QEPyR4XuI+cPLOokJ97rjhWkcPDr7l5SJAggzaHo
nxpZ6vIqPSTx/cLOJRXgyP48jqekkwJ42sD4IsSBZ02J+uo1I6UA5ZDSKMOOyGS3COxSApLZQkR9
BxDuXM4MMA2OQNye1xYgomzDwCfyBc4Ds5UE622TL1d1pLvr899Dtg7BRF2bGV9QBpD6mAOtd++S
n092ao5p/77IR7pOR0Y4I2AfBUvqhyy8dIkxOvTdasFx8R2Twj2V/D3BlsCbzFBpsO+1ybkuUgSm
GT78vRNcisF53ArCauGdEWkawDmtTmj6msZyiDBsZyTE+V5PbcddG2rFCZSfVOh1D2kAxLoA8yll
Dwf3UcfEvdc9E1JcfH6T+MPyGZ6G4atG1Jp07eLijoyYerOO63i0nVYhxLsjqX/dpYGJyLArk7xX
d96Vthxx4b+GGyJZbl14EMcsnb7/TneBEu+gaktrwTD6dekcprYobfPPYnILe52SbBji+6BfsHpZ
aUec05IIeZfsFlmSQNzOWxNVgrES/e7KB3xB0M9LzdZAurQv9S9surXPz+DP0x4HK/4qAjywIjq7
k6lBU74MdVhIBYBYJAKulCg+ArsTA2aBn2uRKuxH518vUmAXVQOjULg1iapCAkiIHiEgFjTrMu/y
zLnmr7IYVb7hR8/Wp4p4i0/t9vKs9jSrSof/uSMZGIhshKigk8HSogdJXYe8KJq1PpOCylqX36gO
QZKAWOsiClNemmSXImn95SqhknHiJUN2KzrnvhLH6ADlH1Dm5V6qRrQynMKbpxz3+k180RS6ue+H
Tv182eY11ERxEZxeNxfZFtEupNNqdtR5hoJkRR6kO+q2CYjFKrf7DlffcD6oc01QbWZjn3B8yqLu
txuINQZwWF4bb10xAndZZoVo9UDQIZt7rhc5MGqAjxnmnXeKwktnHCNtEk0vk9g58wEAQTP2okPX
mt1zby5TS68seGgr9b6b37/xQGJ1ixm+P2wnotMRdgzp1mfbFu45Q8s/xqUxcIf/m9TIFxvzEUKt
T4mkHY9ZM68FmGEkFa4Kp+ZRJfD+koBn2RUYxsbnu0yh2u9b5KwzCmP4R86qwmR3T4AXTHm1xRNL
xf1JfFvXXy5GfhXOoAqmKxhTlT4nU3DUQylyLs1uXBgZ7qPu/NfOMO773rDP0CV7wuJiUOyK6/hf
gxwnVRLnBZIvHIXqpjGQVekK6/b8v8zucxt0JilqxMHgfronUv/l2ujz4TCTsLp7AvJqeZTAsCf+
6SgQay2yGsyIGCP8w4u/Gwa5NrtzonE1ikO/zpgDQXlNqnXdPygIM+i5id9R76Eqc2Vw8tVbf63V
q6itSvH5ixO6sCRHYGHhkjDhaT9FFnyx+TD63dh9GomwkSFbrhBoOvFqUveG1bugBusoQwChsDae
pZaghuR77m3uR4hJLhLa1mH4rqYhSaqkE1/AF7+8ZSfDS1hlekTFH6dUIwAqGgs5eI7nwtroPFQr
Fz3BaZLeDGVawG43Fxr6WPwI9P2TW84EecSkz6m2R26gQe5HBdhaQAdjn0vy4p66ADdDbGsbxZGw
t3fNG9euTRM57sLQJw4nwysPcqov+r20zVhrveNuRBX+S6/M5HqB5Y3/A65EWvE3V2pv0TUhLuEM
BJ6Vz0jDNNgdmk11kKiWh1wVqrRJFvM2EK+MtF9qfxochW9BBKlxUBxqD2x1tabOUam5bmyN6F02
iocKy9bIGnv48kgmrxEbELod6jKIwoWvx/wpGClGBTqrh74BkWKblQFO+VD94EYbTOB5Hx6GqXsz
gWVR/SshgUzQo329XcZWof0J9ri61FAyJcMxInB+tU2pmAWHUd+YORc4RsvxT5zZMOjXy/kwAab9
5aBXkFVgn6Le36Gdf+hGwcaVy23p/RcPjFW3TI9XIbXoUUWsCv8CQ7hQFwRrC6yJtl2uVqAYA2pK
JO7eZNpAp9qufGqfHJGHgxVavy30T6EAaR7PvlbOpRY99avkdmBGUBqva9qbTseyhf+q9gA1/ein
1J0XqzqSAIRLlq98c8igS3HSf01g8Bl7lpFS4tbz5dDw/tHPT0fYEnVhLX8hhXwKM6NY94Qodvbj
nec+9i3IPiD7T/CsSkAunr0Ng+L2uw7jl5655uOzA80O+XKesaTBe6IfJLTN09L+XwAxglBKpunn
k7Ax/BIoDsqNCyupvC2pIb2lBlv9IRy2XSm/vlYMBFUR3ptARnAojS/fdO4YLt/ULIufpDQkacI6
uLH17vaqrmHa58gXlK6Po0LLaVCR7JCaoviAuNncPdYYFeZCm0ddl4fVV26bVK7DCTxU1rk7lp3u
lOr9q0gzJbXubhy+v1i4H0CgSgJS/LTMbs/quWQ983/dMrPAxVKMrXW+9oLUj3ozV87mpNhAhvB+
Iqusrp9wAgfJXg+/Z56UTSBRw2A220EJVOwjIrhj1EzCK7G8HOwXrZ7ovnyWhmgJnyL9JnZZbGnt
c63J2enf2z1QAPAu+07klfZO4CjF1lZ3bHKQcXVqpSdMwgXvgNlrdYI7wM9cgsEYDvT38JYjNR+K
nKthsbW422ziTC8Hj+YubluMtT5x8oom2rh4+IWlWQCrwQupdB6SLqz6e6RwM9p6VDmtR1AlL5q6
3n0oXxgp7aMwm5fKEbc1K5gLOqn0eC6bAyFjoGunQAIaLJdEtjNFBZAllvpFHhA50NSrRpDkneAy
GdV9v5onPvkeLBPsbFA/uiyFfRS6Iv5UmUap++9iSvcLD6bi4oGtjzex037oJpyflpFlwbrFDyNB
TU06RXi5sRiwc6Vyp9Nh0H/a/le72eupHoMr8bCrOAQFSARCxvLOhygmWOgfYWhvUJ+lPvRjHi70
0Zk42POe+lWx4kdn4fZrFv6f5e7tDJEuY3xzQeUTAFs+NHI2EqfM7SH7S91BoGPyzCWkHx61IcjH
ghgxnMOvjln9RhZgB4JUBzLsO5xKFim688ZGmxaCSdNWS1We/iRNgS+I5bQKQ/5OPXciAkGgt91s
l8PLgkU15Z0UEPVskbm9EUbKDavmzdzwIHXptfBi/BepXJPpJYWvnX/kaykW8VD9NBtDXzJJK0fS
K/zbySo7pScs3ybLTJGs9EsvDmmpGgQjh8PxUqZM24yRPqqzCmqVI88g/YL5rJsriNPUTVQv246z
aukBoW9FsFJan+fiZ97guTThuLhKrs6X3W1pSWbrhkEMloM2mSDnZPecKQFalhUauHIO/ANOot2D
rFR+lB5YIGDrARvxC6vFL3dek2KdhXRV4EHpcGxTtAUN6gBRndndnowF3m/5xpnS/YFjeMyKpXvJ
arubOSEsHVU6rxjrlVlmNvxjSSMcsTqaO5UYbOwNVjws+wLPgdLH7d85fbuMk5ZPJ7RaufPP/biF
Kt/KTjQEtzxNw4UpkpVM4bzmDv3pAK3skjrqBJgThYcoto0jxA9xaCSRCjQ0o3wxIQDA44v1JgCf
zHAHnc4o7DZETIwzVaadcYQSrNUOcOS7gmKqWihIVEqaKyXtZYSFMwPZRfryeVL2vsYONms8NoqN
FZE56GNRL/GA4fiK0TW4bly2uSfygSuMmwFmT5664QiIaiw0/eMxHAuTeqyhT36Ku5nGbAcJk5Pb
ZmvkKTZYzlPrr99pmUwLAnBMP9sarpdYpTMBa0nQrMh0FxXV9AiIxAdoJM5CvpHpM6KSry2Xzwls
uK8epbqma6RGjaNGdo91YWUJMylNSY0L0jFxfwOyb825WaSFBn3m7Scj4sYoQr4UZgKOCfUg4tv+
91ganqbljUnC75gsm2xMnb4ctuDyYX61th43sWu1Fc9y3Ev40l2mK6zq9V8jot87Vxx1tgMnOdlV
GC9iWmLf4auGes9Km2NffNkd6MM1mRM+oXr0ywJFwlVyz+cP2RlVohPs7ZtZVQsV4foh4DG1hErH
oRRjmxupqMZ/bujBfKO8sU0HZ8GMXaGPLJDB8L5x1XBAmO8zt6QKQlta/gSx0jVyDQGApiHUXPi5
YxUFbf4bjKpQmnpA0bhfsneu3MfCldTR5HDyF/K8odOlRnwTHwFUvwQmvAIdtwA8dBgpVCo2uivM
7CvvAPUa8ZqPISZUSgAyA5HRrcYcMn+K8d+GbqUrcgCsegFe6lSh60Mnpldk8dL+PWGBU11zMny/
gTxlOWBXAZNk/HR+rVtnVVt8OCaFSQ7H23hDQNlYnS6O2ahkQKzARFpjnYk0jqdXP3O3+kyYkFsm
zfKN5QNdmJt1ixnv/fygorXl3Eyp0qNADHPNsHfWb5gLgeVZr/TOflI+Bz/UKYgP4yxd5E4FKiT9
qggduizWTl7jrGbQVKom9W1V/eVDzcH1EZ4dkySkOOyGxiKNxQ+XZrWeamXcyM66mPOvw8LPmx+T
XbGVkRphutkJzPqDVVhLannTDMCqAz+ihUx4pwpL8vqCBS05AqeuSedcHJeVCqXmrw80VOZ/ED8q
YKenE6OJSYmm/m9HAGXJuwvw7bzEPsQObYtoFoiVgISFOw3aARj6mXSJsKZrYK7joZenMXQXC8EN
Z6SS1yVbwStqXe2JArJyGsce5twzSZQKgoNlvvgSbzyPyLFjXurdkQLjDrJthv1jJtFO32+rQ/ok
vpjbo9Y3lcRC1Ok2UwKNpCX279QKBcimHWwySKtF/ndQcFFqDq65BT57SddXCMOJdOBtqXPzcNLQ
J+sodgChu2Uvc/Xt7uwvuN9XNE/Ffo9/fI3AjbehUmDVIS5qoQci3s04wggNopDiw5cGDbmFj3dc
Q3AVHiL0yidLlFXM7rGdKv2BfEZmfmWlxosbPKkbVVMAH/rLfTRZl8gIi9Vvg28LfXAbGz+lnAcz
fNPc+6Zmv4qUAQXdS0lw/hHBIC/KSqN1MKLsOuVnCc+tAdH7S7+VqA+lcjzTj+bqZI58WhU+GAol
EXPcIIjrf8fl9JyuX6o7VSuPVJj4ChXiNh9xaBVH7gs8ytrLy+9e/sI9ozdQF1R5tNQr5XlW1Y+1
mN9TVHgwxzxv0A0SSQuE+NPl2ZQTqwF5E/G1Ad/Ibk9y+d+BU3En0y5nj3zLDo4jqjizraIMm1cW
bmfWo4TF3Ak9SE6lLMCyEHyFkBdqPp+M+7giH4ytNrExW7bpoh1HgtOlR4ecklEvz3OW3EDiE94y
MdD+hMRQAgKdlYRFR71G6//WmLaOzt/EiE27uodRIFAnvkY7hD9DZCnHFXLeI2/NONAKMaMxGMPt
7/imAogA3l7ac2muDJ0zYRtO5+WpPwFoPV1vGTmD+gWcAvrSIq6CFxMo9+VBYaiD1sjNi8doXHgH
tLLV4E4faCNsiaxn//YFuOWFUEV7hdCKu939hxCXWvBx9V3YR8OByYPeP4bom+Et7gCzPR6oxX8O
2W5ZHqckVxBe9K5g9EvqPCkNxu23mZylLBd7uRc7V7qBPFElH8BfHzP4Wn+M7p+/6JpmHqg12sra
qKmYJc2TQaENnPJzjiZDCIqv+TCrCNQImMx+nDwy9a3Hy2elvveDnp7ZkrFZdK3OXqHbK4YQVZjn
dqLQCEB42SSqR7hqRanyT87b1VKuDArKWwSf4PuTfb63M+bjalYjpJ/7/Vkc8LNdCYYS/1PaTI6v
weLc45h5FipUpXyuy0NEMWXVlueD2znG3lc7yybsmTFiTTYdWMg3ExR5HyCs8rxxv9hA+5PIl2jz
Is3sMmam38GQ/XsA5ru4OBywmdAgkNxcyKXuOYcWcyKrkjcOcMuog6INTcK6hzW2FrVF5jCzyILj
LCvtlqETezeW+3ZwKqYLbPE3xA8og72StVBPpi8JSfzvSa/AHSP+YKIkg1IVKnrBhCWsIWdRK7mn
RGbXrBDQKKJQ+UrOgZJTCuJYiVZRfGn75N7/xmtl1JHAqbrQyYja+s7c2sJ9MMMlbKILHBnu0FdX
Gd8PmuRpXRcZxVcnfwmmvK/xwLVpvDDQeD9E6vfL6ND19GEiqJoEnYYBRuQ0LN25EJ77EVVaR6Zg
G+n6i4wD1Rhtj24aiQ4VLqByo7HM3ZccnQdXGItfhDIbx7BcFy6NgsgxhRZARbimqIiXaDr+vQOl
UolCQFfMejXf8cFbjTMGd/sj6RAsXZ9c4pmD+UMhsar1ylJ4g776Jk9OuPaQV5IJQL3kBckPViBW
tpM00b6GAn3ywrP5iRlynUzcjP9x6VjhMqi02QSFbXpzkms9uWSHrhPfkosDz5V7EVSBsS0NvTKj
SbQX+uOLsQjLjMOMDSEePW1Bj8suJ38jR9ttmGfT6BVd51FJancp2iG7xIYeLydYxsEwQcRxvj8g
8q5EvSrsy+ibwvgQCaae6LNhY9Gsfso5tyawquo7pnsZXVI62wGbQExhfbjBo9YcPWn4Cx9X7a0L
ARAg17Ie1HgsFY6QYciVo8TAlaTngXInPIt0aCh2sYr/rUY/Ah/tGOvJNExT2YQS8CVkVirIBvFW
W+ik7/4HWQDYABini6sq5q1cUmUrfb3sckeyecz4bP7xtqv2pXoTScyc/Onp+vDA6flqsWVRHI6L
jm1qo45Jpgd0ub1p0LCo7wM2/DwFsww+8ON0F5c6K3ODkyTo3y29oEEtoJmhhxXpZB+FRvqKDIhK
+9UE3hjRjlOD9AlFDSniW6P5dcL9a2OxG1GWAC09SgWB4IOy/2zrBwdSD3ChOChYdHe/5K6hpktm
keql3Gh9sQLaHh4rwb8c6tf/Goz/bd5Fb6SsYn3rJsLptRB6gJLrcx9lEYV2i6HIy90V8c/f5rWL
ZUnN3oK8qO2+PG4AgWuibLWI0dX1zutt+geqCRsShOUNOXKfXoYFCJny0wuQc+iGcUG5FaUIQugz
m5mZ6EoTMenzlquq8eHevKcBLxZpO00h5ZAm22nqRNAZgbVX/KGWlRZwXFsEF8pC9jURVixGIw1V
5GwxXVkUNOUHtJp61wA2m+pMarSc0fBoGUctHyEOh3cUNKgYv//B3FEUkvfGj431voGzwxOV6Ewr
xFfk9fwo71OLk/Gxh9N2FTM3epRzRYPNk6WtQeHyijLGvtaMxU7spCo7lA00B/AkPxkw9WSmgasc
AXEdWOOjsXa1pXHdJiBJvvvsk08NXVLEd7JcPyEBzOvpk6i2/m+mHezAZLAKtKj6OGcMZaQAK3uH
D5BVXv1xLkq9277lVgq89o0WTenKHHTvOq0doBscdPttB41rWNh6ctArdPnivbU61p5RIKfhTKwI
D1ZaNFuMqZm+WypQKr32a3Xwzv8+LOmG8krGqgExc/3QlersjAr7ShR081TcP3aP7rM/eWcY1ljb
d8uPhFVyrxeH1toHt6Vxl33MzfP648oBDaKcKUwGC87A6TUAkox720iBtNLvcEzQTePalyocnFMO
HVwBuYvc1d6+LWFgOvhlPI8Zfa4+odh6Kw3znBQ77LAT0D7V/tMdQOLPvwhiGC7XpSCnJtq+yYjc
D+GQlbNOiLioIuyMeW5Amf4FouqDdnIVQSLI/IDszE2oFoUIbFIKoslOiMPo7S3HiToqkW9wsIU7
v16yZKU3BKlZ0WmEpooOXZg5+Swf7sRtILwLO3zdpPUktCF3AfZgGA50x8Izc71A+xi3XXl2Nbcx
GghgMglN8fExzX7X+xVHvhVnHikvZkFx5RvXPvTdFRlxfSBNScX5yR9igX0UZtRQ41/xCE44ZUjL
cCtFJ+ceDqWacV6isQThgatQBatW9yRQWh6kAJbZnBcAKPXlifE/FmZAa9ZtwQ/sw7wqZMzejvuj
fGIFhaUQlAKw0h6Jc/Yc+TWuUM7JDZ/oJ6Ktb/xn17rXkBbGV3Umdn+01oIqeKHcjQvYCIfqMASW
oVSONGMgI8Xnth0CHJph7r/qIs28UFyL+qWnDWtjBfAIMG6mxJbe4PEjCJlZTfdTRo+9A7p4bPQY
OT8DzRDF8a50ImP9108D5emSmLMpE/s/LE7+q+WBG/JD+OUv/nE4UMyeAPqEBlCBiI5FTh9Q1J9g
Esci6sP2S1s0CJRZCKOBdepxmvhyQyJzb7z0csMA6ZeOeZoud3Gt6HdRD5aBJKOMhYTk4b/gSCek
U67Iky1+y8ivQVkX6IeJLTIi6OvvE/0aPp0WBLm9ZgSBI44Nq5GtV5xgnrocdMje8lZZsoVnND3q
KjLnhhrVes96Xc63psWIU+fcE24X8dlNM6F0iX2yo7QogEFjjNJxMdFLozGY9vuHyomBkjH9joLF
nykKjvvFwRePrQ3kXIjREc+IbZZ+8o7YRehJ7EcwUa4Icg02MUAG6dwnkQhnSeoQc3d1PI9yVy39
OUNUSie3BhIKUVjOyz3TqpMOcDJLvKEkh/udTmysM20NILZvJuWJzZ/e80NvrvwgFaIRl3Tn1wmE
bYqm6X62ufGAt6oSzVyuymOTCSsmZ2a1pWhFQgTNCoJwpBgxojKWtqgeNhJmws0GlzjUbPmGHmDL
YqoSOShslvpPyHeaWy+6Iuq6+pjR7ztayPK4RQLiQ15v195JxzY+nLWFF+OPNnwrSocCVlbiRyoo
fKG7qoUKPANQSapJvas7gug0GoQ+49qW2+ch4XViTN2MjisTTQWBpRLP2DLa3pTHDhPwmhoHoDrE
HltgxDuF8tMhEuHQGZgVICmljfM+aqUD9xOErwJPYSqhd82YJSGWZfntiWYgX7tvdRoMGtKH94Ry
OCFPthO8OGAKY4BW1U5/bFZh2wAEzDJkG+WQBMb8MImxPNqErDfCqBQEPdI0kzRYLbgrCrBtVfi7
Aw64P69lDMh8CbWaWGGDQwI50dmDwg4QrMZSgVduflm/1vVMq1uDOvmTqi2yyF82Ex9yaHx5mGM1
1wss5DVJTtNUb3hpO2SVxacfKrrpc3ghbGPWLlXpFulh2Z8YsbyCKYme3CKBC2f0U9CfS6fWT7GU
kGLCBjHsrBXbrPVAFUgqF086fnJAAQodxycKuLSMurhQH7zR4SzBM/lBPwXYAYG7wpmssmcHZa0Q
oqremf6m1JnW7ua8NKPX7/AD3Mi9dridLUG4YdZGzNHSx3jIRTEFZ52XrSXoE9jHuEG7p9fufp6V
8fi6xsRh1ViFnfdpKu1vEu+x/gsmkOMIE5+TvDK17nhOI0Elsojee24ab/BoSXH/bSURQhgaT2+D
zqJoIuViBi1qbxYtmSNR6nR06n4Oc1Z/psugkI054J7LYBdnBp+SmcA/648lnkxKl8F0ASqpUGja
5JMdejtqMOpzTL8+hs5hjbH0SB0/NE0q0JIpPdkeSffPDnRNYQzkZJlp47cXz7jZ6hSEnsEFp4Dv
5Qs3wF7LSUdct9UYw0YDRSeAs1SD95Qf8hfgO+nQ8kIVis3gzWORUd4SyhVDIJfRU+7gYRvti7il
UUB1kRheFMj1b3L/BGvJxZbc4wkkIXTpFRArgx8RnFdsA/6S6lGQFemd/vq6OU03WGOed0zxtN94
EgcgEihyDTkGUQnu5JjC0nrUvqzTUrSjCvOF9+mHCveu6r+Ma+pfJT+I1vQIsTsG/1AsVnixro5g
EZw4MDe2aIW0VoEBf2L+lEXnUK6GTkOI0NpoySiY7+qIxmwHirTdvyBpiTDX+KrRC7ajPxfsatiY
S9He8ax3OItonw3YIBIVt57xgOOvq9CG1UHorlA+6nC0bxDR5SXq1s3Ji87PaokP13YL8F3Hq/Ho
qxlTTi4kxdd8VfCvcbj1lhdU7zeuOasp11wjCAFbE1g7yHRbaQYPTnFlO778In1alWGZg0aqNEl7
UGhPSl6iSzMehKQxGJPUTV8vzdUxnFuK5Uhec/iH3lkW8fymylt89pdVlw1fB4jUMQ8us2BqtIpB
Z5Ne/bXS6pWlzfhhpI+YBZ7s1W/DkVUnIQIoe53HXOmwLXnqB17PzXtMQSB4lhgM4PsJ/7qwtAO6
yEyundlJzS6pAHXiBeKbRw9C8aXo+RVL9WdIP0N+njQr8q3IdJ3e6EUEHysNTuS1N9Qpi5Vq9KJE
EKxUrUiWMpFXs6nHmMur3rW7A17L3iN9tCqNM5Uq1YfdBHg4d6TE2d9cSiZeaP1hd5+s42sdCkPN
2uzz1nr/Ykm+V2SYshf8vf3LiFzNH4hrnZG6JUBKbXln0NHJe/TT0Z2Bn+bNzvpHQtIO2hK7mYBx
qHJH1K9+iDXkcHEK/aSahtb5Zx8FqHSg5Zqgoo629g9b1P3ZNhgXkTbowyJ8VkaEg05N+9+C92DF
wzKcms9K0VLCXH/114DFurLi4ClGXynjtLcMahevp//+U2HNcGrjbJB3CKuFkpbgOeTBmSttQJN4
JXBs5CSvp36cmakDmGnmuXtc/Lw5rQJVJBueXcn0nE+opM1a50uGNQqT9nKCG5FASytqI750wYFi
BEngPMzmH98dkkrxbY2lgZhsrdoQwNeDsfuHltx4yesPsBbd56bv3PHYCFfqxrD5RSA6fJBzyrO1
0OR8Bdh6oE6ylDiRwWTVlkZ2Qi5MtnGf9VTnQhP3EKnMN3zioQ4mha/gyLQQbhdJQIw54x4FSKyF
OIuqsQBkyPq5qgxmKU0qqAAH6kj/6vdkwbhVWLWMwPKzmzWzDNvSdAI/Xnn+xGkYFHuQTj2nPcYN
9wNK9ED48tbRZIo4iDRgo94VPlNNjKTPecIpMqbi26AE4+mK1Es6k+tySbQQK59dxiaaTsqVjBFY
Ms7YgY0zDDhJIhozs8Y+f35AJ0uL4UELcH0D2EGAMnzwmDjDe06OBA2ZG4g1ZbOxf6i52b+7MfoQ
B/Db5F5bxqs5ijHKWwyaW6wpA4bAf46C8HGwXl34Jj4zBYxoSpNSjSd54PZAA2wOFms2SJJJum6C
9vdON8clS2R1mH14yY3xzwnOl+EMndbSH/ukOIF7hvo/gHn8Jj2EiU39yglroc3NFF304b1LZHTf
M4IoRSIfEHhsTW/7LqGFqCDN3g+5SFGj1JupjnESkdGLkxTW0353lNc8fFofjmggBWswkfem1oLc
DQP4YA15vQxWOT29sq1CZRRp0sZBwB7Qg8HTUjYfxNwVcW4tLuLSsAhilGP1xDI7Zz0ai1lnCy11
1tIx0p1gky/4VnLsjeOIRDwsukq9HowPPLpPE0wHx3DgyNglv14mk9+F4dSD4+Lp3iyj+B4me4RF
oNB3onnXHhwKu1JFC1n6u0bNS0aKNy0vX9e5H2QBdZZ8LqMgVTsjBh8ao9jcNZr1yWEJnbluVJeX
Aqs3KQT5n6oa4Q2VFP7hAOR1vpv0haCFC/TUJNK6wgGqqGjx0OzxIVksNEt72HG0kaw4z8XWXjEt
Jy7CyrfzqpQqozJmw3iFDS1/PuBo7vS4ZF1HYNnqGhOiFrNxJHjL2Favgt+DcgaIC53MxuEjbRjh
lLmENgJ2b0iTG7o5LuahLJwZMys2uAwlEUIY8bsUgsusLdoNszzgw6jfLzoVyym1Xy3QAwJvAdBk
K1Z8fZal85QiRC8gfyZGBqtxYhKcxIUp2kYQu8SSf9LpAHZBtsMwR+wcwsrr9jUIOiqLyanL+wqg
etDkb2TENlWnAOc+rLQlBtCZR33wOXaaR/DBwQxRCaXIhkp166RIavV8inQ+WsxRL+W6otzUnH8C
g471yQgA9zpB93WkQp09M7zSzvo/SYPA3HzEjx/zWp3CQpRhPcVojZkyS0zZeEvWoD0WC18RJl6/
fTLi235BnPSTxFsTLcwd2B8xZvpbsVyTWPAWhvZE67hvytp03q58XjFWIVR/Yi81PV3QeiTZjRXg
/76+if10Ei7/auCxD2uLgCVVmNHaEeZi8VD0FjMJSC2wIE9RD+A6Bc/xq7x1YNb3lnUl49sWPgCq
f62x23BAvNUNhkiELKRTk+hZOeJ57Hz+AgpbxEwwmJmxsoyMIWTmzUqd2bcZdKRehEeitWD/e6wA
hXeBB+1CifHuc87YmjGpHVMyMbhMRNi62Yw2fVujiO8rJE3CXZU+1YV7oAkMLVqfgCX3L1RP00I7
VluWmnZlAX6zg1j5LvHKS3oF8GNuysuL97DPm64YBoJ53szvJgz2hTbqhLi6W/+5IkIX3nR01Mov
0Cgg0QXkJdaOBMDeF+aZKcCEFmrkkINeLyHwE7Rv0yftXrbWSN54tdwnLbpHXWolDOo7rNmBIFA7
qAJcBq+/F7hsa3tYupJENyt70pHPoFvABReS60wWrHbH1nGI4ppumuPVudMYvPOG5IEAyWIGf/EV
J24L+cr5zCy5VUs2Qhz11iLGBMOOsniE3ZPcpx8eXIb0G6XUJh6kpYdptvQqssf4AnqlNssb0/n+
qN2k8BilGfH6V1qmjw+V0UaZY+vL4UuoA6nSRDijNdLrEgFhoW2Me23W3QOsZU+l5uiPQJ3twPMg
7/9MqI+OBeI4CP26gm1M5Hqvrtb6gmvf0HsS+GI1/K3j5e1xEHVs6HG6F8RrwjDZgUXR1Rlc2Epg
qTOzDukR/Mfi0Rzd5D+26PVNxeg9uvA+Zo76oXpiEFeAnvoDac/mZoOYlPw34yGU4VuBecEfK3AA
LjvPDor/72yj2oELrUhVtFzj1JYLaqkzBQKJv8yGdLIYi8WUeyMRDJMSjFqZokg6qzkTvitTKYh9
VZeoLLGkOPcFsWLLOom10wbNowVfRi2tYazjb8kniHamTf7IeRO/qX/RdvTrpBy+qJlA/3wcrWp7
iXKzGnd7HPBYxHqssGVULdyMiobAosFqEgtWkEYDhKOMwjiLmZMvmdChqpwxiy7Rf41FbdFRfMVr
BEpeIMJgMOv6Fq9sdH57q1caUjnJdkWcABGC6bzm5ZC6/9QiG2LLSvCxrGKv2RW+jdQUdJEpyFNj
BYrtj+IydZfpeObHLig+WyiFIwZUU09kAWXrfLR0k7PpJZWM3UbxR0WjwaSJmqfBY3o+VBH0zhgN
t2zmVthBhz3tW+tdx2xcqOAa5wDDq5vSPIg5SQTk+qKAWeLy9kZ2h6JAjXGxgwiJ6pVsy1t4t8cI
je/SWoGCJ0h0hhrrmzXC8P+R89JuQzE/StDKakgLQpfkUx95fcSF7cMvCDhtPH3PIJcnwWRWbOS0
VIGG2u3SPqNzTnCViYwXiypTfp/2HlqlJINYkq9+rL1O/Pa0WvR72hTYYsyYIeg06VDwfU9xsSjR
ceBFve6PolVsaFRs4zCtgJ5gVjZ+x5SK78LaIljWEUIcg7+d1RYgf5bd8gIpyj+l126Zvv1wcHt2
7E86Yy7OmggLqcD0MXJntkzFKQhSP39zZGUlu/XgW+I8iYTzzvMSIXIXGv12D8RK9Vvi7n8FhwvN
P9Ps17j1VMTl2qa/gKy9q60cOQkYyJ5qbix6ur8EgV6UtKGtGkVeINFDjAn1JPYLwu7k0txol1ol
9bIYHs44GQs0IOkO6HO3wa25gn96+wb+Nf7o5ZQ7IMAqxCf7n2JhhZ1DuaCidGGUMmDSWt//BnBw
H38prnMROMdzth40z0i76qxbRbzj+FBblj9KPwp9p5q/W+6YY9Atm6zgN7f1iDhyHU3WbYEjnam3
1Npzi+T0YI9f9WTEaVuhzSI/w1l53EkLmCQ5n6qXtYpRA87oj47GwvqYhRihn8+RJiO5XiYZuna+
3dkE9TtY6QFtv9CeK07x13Ug9BYzE9HMKElbzpPoezVX6Frsya5QTXMTn4fu77ITNWfuG7lhJH27
Xy73GscB0h9b2tzPvKOclH0qA8z3SKZIYPeyyoWhqj3uzn4/Z/fuD1wuAjkDkyU0RZP+GCHnRRco
HlrSzgAQ3qkf+qSrvh26dJ9v561qgYGsW4qs75Y6IEJEJh4wJV5e7/zJ1DWZ6NiW+fNz4yNYy/j6
NzTZTxrObUL4xiQCzkh5TsjKp2QewrQVdZ161PqEwyYU4wJ0LHqJXTzDEeBGdlEiZOvmKDM4XYLK
6RpAMTMJVfoVq4J5n0Yxnl9awoOC/kfCCBrVG9DUNBlVwffPG3qTmL4HVemJL9hDDCBk6B37Vhxv
WC5TuMduEaRzRWya/NPAUKbdpcE+QE0qfSYuoO+AtYy48gJgE+i6dokliRNuZReE599FcNhr/2C6
EYTrQRYuUAqh3UosmCJ73E2kuUNEUa9p6OTV2GMPAaDnbJuxKQeru30C0CqTOh6JQUgWtLyr99Ty
8c0dPjsNf5yCuVbvb0MfX68SHi4lQkCmLgT+Plqtcy38WWXd8UMgP0zvkujplsJbQMXsXBjR2rlo
9FxZydGuoto2mIsNTo8TcSR7siva6/FqPcmLyu2tgGUHNNvtnrs7S4DveqoOiHgfWWA/NiRNeY4N
APdzAiVNps5YIUPzQkW/fIK1yExWSH+7G5Z9v0cg3Nix7rmI5siBMoVW0VND/PO6pasX1fHkSeNi
dAONqmBRCg6iDnjBK2+79NtYdhIpiCWarrKFzkE3ROO9peNqnmTY+Z8mILNoFDBGY8fYmyUiw99W
VyVX9cP93YRM2aOZa1kje0KRL/gsYv0z0W8lAzoboW+9nhaUf6etkBBjrNykz1sji6sIAbCQ7Y9T
tmTE0rWR4laFjaquen+JU6FcbstmWSFhT3UMgDRwK/tmVJDGzDG0EPrHS0ioWn056cmPVOkJx5x1
AJKSW+fe63HP/NNE/L+vhIoFX5Ysd9atPqhDL0bfgdq5WCwMsByAUvBOaS2fpkV+HLwgLfMh2N3w
SGDW3WGppybpQ7KDAdaZRwEAGCUlkGLPTNC5aVH6cu40OJK8dEAaQRsbDfUSgSW25haveAvK39T0
KPVon3lJ6ttBnZQN1Qb/249FPlIi31IVaNqs1eBT5hX6YzpVJuKwA3+uf6afeq1HMqQ5EwS9LSuC
TbhS8ZKMdCkHb8RJneVMFGR06yz5grXpRaLBj/yWdSGL9GV6x9diGouxbZi+/u6VS8+l5KGYUQ+z
xLj4G+Gej28OItLANFBGYiNv67FfN2nK3R3uQFHdPwQjzCNNsadmywVWxrXMVO8nN8NtSMx1ccP1
Ey1mPROWIxMiy/IvbBwvtfkrc0XzDm5kSpUKs6afT9Zrg59ofkiC1f9SU72gKQtHp8N+l3zYBE3P
So47NQf6R8MhiZzH9Tga+NZmjF5j+9resZwPMEyzIvobHYDxRZHK/oeWMjasmncWrbcEcWf3tmvq
+c743XPGO1cyR1KroQuhqG7dUsPeY1g0zIpeRiUZCF88/F6xT0fyPl4Nu4osiPSoCrAVM8ynA9Jg
flj8VDT6uzHlaP1gwEbQjiCHvyZDEfPUKr+d6D2csJg94yuFCKRzMUTHtqlPN+g2ZFtBWoYlAFug
6OupbUoHDDOlHh7U26BA5ugFCoDqG2m30T2K8CgCEt6V3zP7BaSUI8wPvziby0tui3hphWp3m/AU
pr7R7OueWTmGKMqoKSfNhOM15AkwD6PDfFURD1ah11Hb3p6n9D4wrrFGXLM+1BfI9a5+CVsgMmYt
8UnDHCD/oy/8XKRRoSiWc4+I+BtH7MuauYye9DVSER4mgYZ4DBFHiHwAftpqanTM7oaX93cGnMar
BFWv/xdSUorj14pwoOW2iattwnbPXMIwvMbJIiuU+zErcqbD2MWuuiMWbDS72/DgSRTZCblYgUr1
tccw+PqmdiisNKeNVHX2REHaSzYCL74l3+vcMqchkmXdV8Ca87Amzi9Z3KSLFHmr1+64BNtJBgdr
N8hFkGkcFmvDPVCK/l1SADAK6S1SxRlUTvkMXaLE3YrrkcW3mNPfZx4HMdEV+dd+n0h/BC4oaRUl
KSctBAw0gE6p/8gefacfEIKpR0oSXLROqbWsUVim/Vm6pyccl3wwA/V3nX7hmEHPmo6xNtDnBzR5
2RUyBTaPP8Ao8SPfNHTjWXd+n4AwiOmuHf+qOO7yKzWoBXLJtayXs35fOQupI8f0CfodfCw9VeiT
3/CSqxuvrFq4Sc75U0WLxNz2v51Jt3tbxg5ZjI4fYXRxm3G4Yo+L2KIUSdhgg8iQ/8TEEdYXqsCz
lmSSD054k8bmfgGwSrRb1swXUKxFO+/5VgC3rOyfO3WFxe8rWWZnRH0OPPmg7UBEOGAZSp8VwzlP
ItTctrUJa+m4+WZ6YmhchqQQxH7Cb9xSh5dCDpgVHEVn0su4tKOK8qdVyC8ju8t0XkpmzE1N+l8f
GaA2mw7Qgycad8ZPInxsXdoTFju/vF+bsn1Y9XqcZ+QzcmqmcgPDt1ZAhXtJx7qAMEtf89GOAHNN
oXlfInIuaw+NwpFzJjE4OPvdqXFl+ei1nOgqSKxX9dxTcx21ujaOxKeDWq/8armFudGN6xy8g1xo
iYH0NUxCg6wBie5xvo6LPI7aeB1EA0kDa4fnFb9Rw2BVqj3cztEaFlAC3ZlP93jIPR2Y4gGTFaog
svmWXXEqamthDS11evLpNEJDYh2quHjvwcSBxzJ1DKmc43/oTOH23S6p5KHCe0ZIpSfaq+Yh9gQ0
LBQ4RwVo6Gj3LpGju8gwiMnLXN8dbzoEWAYLx147QmzmeGnn4KxLNNmLFHJiSpGD9soFSS5TAuoQ
TEccvhWG7VlLj3BPoHUihiFLJDy//zT+zoFNIYok36R9YjbZGQrZINYXB3+SB6sEr9mbQoFIkT3Q
9PBvLT28/plNpdeRzysJ3ippKy9BvVXSHBrp/bM6c4jv/jDUbCEVlCgy/EuD+cnH4RTwciisE87N
EwEFM3ZefE73RJU3pd52ijEZ8eoKRrL7h/n4yRyKJCahvirOyWmiwn6HyCC5bnTi0XrpqpjliMFB
NHE1eAn2rlpev7wKRjW2P+j0gPBDyHBQEpfn+e9bK6I1upya5GTKh9rBUlFWpP865coYfynGhd7f
xU16yjuN43997IfhEjBsj6ZTjgx4tSOjTJf/AajeM7MwxO2DuOjiK+a+p4Z4rI300uZ8DO2lgzWO
DdcmNGQNn/uAAgdZt9/Ps1R30ZYRM82LzQxq7cpVcBNAs3v71Aj4asaaBg4iIIdXNW8vcrMrIzDC
h3GShQV0ke46Vr5qoYx0cNPs0Vf7sXpc/EBNF18R0I+Y50rB3pTFK0NnXE+v2iqM+P8JFWUVBZni
6i3qOIFK+mW67b6BIgdprt2+9I1LrDCQ6JpL+N79C1Vz9rzn5c9IfNaS6AXHBLFZrlO2oOVmR2E7
7VN+bgTKjNXz1841emT9rh+AklMI3wQXiy5QKI8ZS8+R2/DUFxPK35GrD6aqWjd+h8DbxwBqzjgn
wxBdJ25ii1LdcT4lYQfquLFTULPJRPrO+u5K44Y9Iiu9D5HNnuZiHI939rC8n3/DPDuq7qNhGuIo
lXDzKOZ6hyEb5KEbwOeKsVZLbSig60p29N5W4nTR5St/AOp6zPmUG3DMhcfSUnBBZe+RNuJsylZV
6R9aooSCIa14h0FM3IOwdMCdT9kKDsxtsdwC76RwEaDyZi/w3yj9ZvkHz+e3yLuHwgWwNfH/7/0W
cLNt8I1JhVuZXKctAwPbaHEqUu4mlbMel4/G9U8LySdrwIQFFknyssBKXqI1LWXsk1PEPi+V68ot
ZKFgHS0u/6+3bKWNMxAaVIieEiYVpDIAhcYDpQ/KfzHAu+IpCQiDqxGPDoGgAQXiGzw8LC9VageW
qy9zZ5kxGl4ECZvaG/Kec5hi/ny98RgM4Rths1EOBec4NEiiaFnegO5GomqHvA77DqcySn5gQ5+J
5137BXac1xWPtitaNobi0P7PtZUC6YZ0edc44M9PsceauX21LwxMODiBgkrDgy7mS0DxjRTHBTND
676n42ZEwsEEK1zJvDUK5b58Kmq0AHh1lStb5Lr5YTYcW+CAXs1/x7zYxFOd7xAoDwlje4thbZTv
EakjOVSrOBBnR2EmJVI7BZxzoGjPp0CoEh9lo3yBODvPJvJKDxxtg5E2iyFZo6pBwyIohLRcumuM
nRLQOlIYSETbpJ5C05GVO0q6UMWZm2NpUnXquBqWia3hy2yK8aREuk2mBvY4eDh3IjeW4pagM5pI
t+FweaXV4yYXZ8l+z6NOBukX37jPVE/xtkIzmcs9800cXoVhn1rpg7/XtZMfffswfhqhHIp0a1Fp
5BHUYQGfdQrYQ9NOKcxYJOFthBmyyz3DPg2bN2x8UujWBVMqXSCX6LMHViPbQe/F73HNRR8vxX/E
cm6Zs8deFrMl9n4mIbcPz58+LtxLFlKEpH9TFyBCV0JkwRb4mZk00JLaxzNjotQMNqakvSZ9f7qz
RJr/ip2bQOSPoGYaaTi70zZhnQAuUhVF/mHDI+sUGx9aRerwuuh8CEIJuxZn1GAQ+NZMzqrBNvyz
tLb4b832I91i9zjXQ0/YBVJG+qrWooGxLrZ3danz5hKjvywrnAReBgTAe5x9pftWUvY/H54P763/
zg+6fL4aixkgxS6ELqFxk/XHKXWDMLieQGby6Qq4v2GQLbybXFmiNayOi1j4ZV8qoMcLgP0tvjg6
S8cIJujLzC2MQmCxk3nB7GMDRJsjNFheMYkDaJmA/oifGMqkzL5jmJcPcbqd3Hnb+3xNNLUBAe7y
Jh5D1QShnjOfL3tLAmRQov1NYqCwzhaTJ37r29O7N8d5aMggcMyuQKsvcpXoEuvcB3YGxfQ9EbM4
PJM/wUTlnyrEcbdyOhpm+nmWNFoyeVBqZdtB8X/qkoP+/Wi8bGzjsoijFOMr37s1P3B9cHZcr1RY
1K5mLCWgKMWxADV7RH6CrrEV/Gb4DEuAe33VJL/5K0wz1F3vsUaaKogJWJTduoH48jDcsn/L41AK
yqk/rQbgrsPW023U/GRC3SZMITA6rgJCdO78EEqrDkPGTMGaNqXEGfYazcH4Wo/xN3XAyePJRLkh
+/aVwc/IPGsOUfLfnmnSAZabSDzwspeQBGnVpYqyEzffZ/JDF6X+f/vFHPMGdj2qnW5/jyzhAo/b
Kh6oKla5xkfe/EVowc++zyphkyvSHD8SDFPPtU4BR69oNSNujSiwdj3iQtq75+HJXoIvZt/htBx/
bglNGf1Ys3Pw4dULdjpZHU910sWoCkXywRJGx98EGghDsOeHagr0fJ8jbw3/bMGmxNyZQ8zN51Es
TSI8nrK2NNmcZpQ3bUs40+TwdTfDFXjKph/DOrMyFIZtKP/bRgSVTh0DV0y6icYcsK4/tN3w1jew
sbYl1eUa0BJt89fiJpH/WywXCvq2FwRtkxaOfTpOZGaD2Rwp8EIJs6F+4d5xQfSuyt7YpWhi7QK8
PL3usCgPtbNIsEJuJtFpnkyNCt3ykBauUmgyT0VUpBzkuLR0HgijFN94qmipQ4uLUdY3ZM/yP284
1qe+GDoLdL+qfdbTf6xJylg396pQKY9ijfc+/V8QmEn088aiWvKZjNfPjXN04FcUwYN6oevq8mgv
Z4FledjuOGXJpwC8ftGbOQzyqwF5dV3Vz6IUMml0XNQmjlm+qwtv3OnkwnjuMB6oHR+677IQATQ5
c/egZRVqb/Qev34ajMl+19HJSFJfEhyOqwsw1SkM57JMg3BgjFDK0pLen4OnGmMFzVpWgRhYuv4a
nxGiWBY9yacmy2rur4iq2HySyz6bzpgd1MVPmxpCGWye+wpoCMg9ROzN/sqlqm7fEt+LzgC4/E4H
YGTzerw77In/aBDF84HDN2yGQgrjyiPcNaC9z0eXzLWEG7eh+jQUrRw14P02f6xq5Wdm9wlA0z43
BnaxjmRt9uCN2x6d82dkCYx7CeyAllts6FdiM+zhwHMUTEL+HGKRTVlmjW9uTgdi7/F68rsRNufy
hjk2qvemHwiW9/Ot9NSE+U4ux9uDZmcMjeEQ85PiHh2YIBV/fasEaegdHhcfhj4LR0v/MqALdwwX
tOcmp4C+jG69331+is9yCqpvGMb2Om6LbjrvxQKgXGlx++g3ZHEAQG/Hhi26rCXIZf4anSrWydzK
R0jx6sgELGesyz2oaiK/ISnmfFtiWqW8MK1r9GRWFYzAvtHtQYUccHhC/dWOE6/MyghhSfYf4BKN
V/NoIaIOHL12cdoWt4NBS05g+gop/IJdFaztCf2gxIbQuMe/UB/J4pdNJGk891GAQSqjfueK61RX
vJpLuGK06jYKXbvTLuvD72pzOkPjZT+wRvQ0FYCI90K1GzdpxMKd+bmvvXkoLkQBzq8h8PjtPvV5
nVGpB70gRgU4zgMT2kZB3XiyGZhCWN+h6KqfdUZZDD/LAOLx4ycYite44sDyvGr+oofa3zso8/Dt
T/X+K8M9ZImf+KIzJYJQwUjvXZ90O3l+5rdnN0wQZwc87n6gUGUcCKbOXepxeWi4Rvm8653tr+Dp
VHDQK/P9moeSovIGpvvOdBlMhtCdqGqh5f1/Aa0G4RWLg0ECqCqBv+pcECd81KzDo73OHsOw95wX
0FPRk/d0SShAsWJ0vvpKBzSgPiOpoZgDUqnlM3sj65DnE6DvbsEA+E6owrn9b2+QU1vbwVocYa8K
/PgECHIQs4tEC6XWMNDqnbSIQZPPMGpObwP7S42EOhlmEzP2on0I7Yt+VGaShS/n1yxMNbb1yqod
2CxZJn2P8CuwnoeDI+hkbY6UXVwfBD1O7kQHtCmORAt79SGEasFQ3YOSZ0OfztpNgkh/Vka7bSSd
1EpjgZB8xdhA/l+ELtndocAtsX/R0P91J1UL4ZtUcLNnRLWcFbjfju/eYhescPjPAWsZE2EgpS9U
wqKzyGVWi0XehjLX4ZTjyS7TVvMXgFYmGViEYiGIs3OoZn1zcJKE6q4CZtCuV6NI/G9SpiQoMN3A
OOiwPHJHJwiAXjLhD06OGPvpySVpBavs5/5P5CVnCoDQrRNBk7aruPy/Ay26Zx1ekzaFQ5g6Jylb
iGyekq0/ec4X4NKMy3qRLiCQ1bB0oZZtbDYMKjDE/VOmOYfCrw9lqh2DtFbjI1kaaIWTAlSBWlYg
8XeNfqZznBwebqdRVWN7B1yRFCEv75PqaEQN1/OwG5sCh+YcxzZOFcZeTBS3hn4XCTQ/gA5/jq8V
mmRmeNSjnV613El7BJfoWTQ3EEQ/VhhTPNIT6Uh9s3RdhOIyR/H/3qqEWXDJhY+JZ9JaXVDhwCLo
rC71U7OMq+9l40wg1C/6ukWB2kt/YMx99JsOm4c2Pp5yZsau+snNLByATbL7dEgMb2dl5qV+kzrI
g2puDIviuapewXaqUnLOCS9SySAuYGqFsKpxDw+lbcatCSyWHu8YcL0CcL/Q1LmAJTJDzfjl508l
GtFxyq72Rakv5J0sFpGfCDiiBf8mII6HZe1fKFML0GwPbQzf8J4Q0fsNHUT/odxt2ojGEAniSEiZ
R4zdOyu750vDurmBGf9kdP8vlaN2Q4FHDByxBtvNbIbcWLRHZIxcoY+4mxAPyqFakGfn6TijBvDK
wgkWpYoKuaxutxD1pkmR3ZoE8hJXnjqxsJgZKPzfe2qZHQRGVTRwmtmKj/nwYqWTiSSQI8awJTtU
NPwPiGxY6Jun5TtA2EJ1vojdki7WOHzDgaglLL0qMyiJUAPaUliO0KUUX8eC1XXj/mdeuzijpMOx
JoLn6GXuWjDg5f6ZKi7wEcXaRh/DYtwB9fLhkDQFsR7bUKErTAN4eR26V3fl6cQnIk6kj+pi1cYH
82umPxGEhCMwtZ0sgdy/0L5bq3e1VHpID7p4asESSqvZmc4AMJsn15xs1+QICQfcwMwGMTpZypGN
/ZLC/e9rgJkOBfGfbPgUCyJQ6OUZFCtErktkLzvmegPoN9xSLBTVwcAzrV7v8oFX1iDJ3bEWzlwQ
wZNsftjr37JOicCUKvYzSHKg0mCpLHpCDiZkIX67sJxDEaKbwr8IIpBT4A9RLm3xCkuXOc7SgNtD
AWS6rI96aAuc3zkUY+8c1LVX8DCkggngaKYjm5jpGzIaM4HdG+rrb4u8gYufNDMRVuxtfVF3s/wF
GJuET8vmyy9K4MkZtXIY74g8xlM1Y9QFpP9Sy8BsPaD4UOx/B+lM4RoRTXppBbinYtzR6krPjPCX
bFPsLHTU1F0zc1LRb12/vY8hyAMSAZHYVDJXt87E5Lv/ZIzyVioToUhfYer7hgjJ0WJRfuUuj0pY
O+a/sGIBK2uAg2eROUrkjQ4T8cdQIcOPKMXtLtTzdiyDXoADRs/6gEK+4cxD/oWecJMMC71rfLQf
F54P3un36A9npckaJKlD3d3ABcRD54CAMyMdIrKJ8F7hY3i3DhQYdoUWGDt+Y8S46xDzCSbaVG8B
7v7aIXVyeoM0CuNaGbgRI7f5p1PURJwVG+LFerXs7m7NXRyTMTDbWugqkpDppuZA4J5sf87D+G0f
xMLJTd4wSRcnGDpmfcRUzPfIDHLlAELmVhHQGSuN7sDgqBB5JFRwrqtmIvcOyDIbxQRmsOJ54M12
0kV/zteNbxDE4y5fU9BCHaZI3EHIrTEsdP5Q1cj2sTihT7AfBdgSPZh2oFyzHOBpQDz+Ndv1aMD4
qqq2x9x6bgS1eyQzbGCGOxrYk6oCNYmm+gmlOveBLQk6eigSXU6EJuC6IA/gtnQtsKbatjRQCopW
Shjn/mhFS6kNYus1UTcW9hF96ZEMN2k2FuedLEdNBYYF+6m5LRy+B3/+8bF/EWvG4g6CXov9zur9
9jW/j1fWP5LQaisK10CfbASNcf4zX1hfMQNujoblCQX+qWKiigd1e7BJeQ1fj1f41LMbLoUyyTpM
iwanyCXBe7GA6NLp5JpQriQ2JVgLHpMGZcvdwAye2ngXb+DQ0ENUTVn+kza7yv7/qnCkl03NeyNo
tDgE+dA6IasAGn6T911IJmoetB3R5G5IXUrO3OjoBSAPBhnqf6WCZxUGkuZmmO1wqnSAj0DxTLDz
2GhITQvMH2HrEx/BiEdIThReXtctTkKFOAK79w/szlxilTlp07sgUsBWZ3Oc+VUVKvCPMS9rtlHp
urURNE2Gb7TIw9xGqK82qpTFlvNcXJr1w2xSNAYY+DhjvpqzINvtP2+IwRX3U647iO28C01WxoVo
ABfi+XC+yQ6HHVy3ydrjXXqIv78E2IXqUO5hkox+jA3SkeAYnL8K0n6dpQWcogTJIkyU+tftxhjn
qtX3p079EmQcF2wF/Qh6IbGwLbiumOXURd4W9Rs/SqkZi+ZdjmUKln81vjz9sXnM5DJnO28LCSco
mICy7/jo+qy87U6kbWbvCWCfKk0+Uw9I/zGtncJe6aSBxCq3UBIdipztvUgNiNUsteMz8NHjRpBn
vNJlZlPRZxCSL4fNbrVK9BwZIvrDLZwlv5l4rF2OBGXMhOUmx6bEk3Vax7wmiOJ4055YS50riCu5
V4mCz/h2LZSo0uLViqDRAF022WR3dJ9VBETbtqZWxmF4KI9oxejdFNHqurCLZox9B/m+ap/ku9pG
V3cvMUPBQ+eUGPWzDhAdmfbB4QQErumPLKBVXgOKEHuR3m0KffjPSAYYcc1kqxzha7QQUe8VVtTA
hH/vv2I+VL0/VCsYT6qEd/4hKWR4Vl68xYiQWKl4Sw9BFpHRfMAujbbgthnL6Le3YINbtEH0I8Fo
nl573tH7I8S8BRkxfM+Si8n8Nvk6FAWqriBaQMXo38/3BZow5qp6n23FbFIq9UNbkkl8Dq2WJHfR
FP48YF//Lm/dqMFE25Wi2bO19zVBtMQCOvP+h7JnPxYJk1NcXiDr/NI5MDI88WMYO142jfqpT3vp
phxMB5HC3RM9GE/GzAG/boZLqF6OFq5f7X9XQYf/fSWvRfBXL3LWFXfzESrhw1UKUdniWTj9ckq+
kRheUJkSDoNmzKTrGmLtrSmD4bRD+SowKKma4f3K3qIMXiV2qk8IsWHTc/XFeS5AosydEYh1Vztm
SlIpjc/rI2qlHrDUv0n0v6TNaS+UEXNmwjyXw21qBiMBjh9+O59J25ZxflcmDmQhKC7YKpuvUYjb
nqa+EGCEnw7jmv6gLrOxGLxvpcV0ZMAPwMDQ1116ZMTPmaAmmIp26sDVz73lFs4Qd00y4RcmjhsQ
7g8Y9Zs75sGbPlackWWeDFFCMbpa7B1A1v7T5F8tG6JsgLUJ5wuX/dDxx4B/oNI18WaQthFgYBtg
3FKNNiZ/G4qYNd0O1uBTun/9qobECMMXg7oE/9ov2KbgJvACgj3bvvGbu3CuMriqxZFZhMBBWSlJ
QIAKYyAhVDjTLmwZVFnDTG3HGgywKlvjFzUZr4aV/CeUqvj2VhLkmnU4cjvdxfEB4JlkzTMurkkl
zZgG1+TrjB+udUz6KF9QoqsfNlQ0UwT3oVeNo3lbxz5bQBHA5pRz3sox+m0x0X/J7A+nS9vqjsd9
ICFGCx+IukaTgPpW9eUbjFzF8m0P3GOpYEy4xVgZFT8eqDllzoyIvCYAFsBGjK29fig3OWDpP2IC
qpV2yFYXNdJjj9X7GrlBLJB210kbOf2oC+t1qTWIhl2j3SvWjHNxSN/5BlP+cGw/hBow59Whxerj
LVdFzwwbpDJrpPQNPUvRoQH/74Ced9FDHajjbeVQU9X6rqJIZv2+nF9yZcgxRFGT8OMfN08jmDEQ
iFoCs6USBd4Li4vfibbi2ek8M2VOKd9AnQeuBoFl/TAiwwsRFfYQtddLT+TFXOUqoLENyRqhHbss
4aUt+LfdWStJOSxzYylyiihfBr1x5YOw4pkuhYNYAmjJJRNM2TCPkGbRLhKvqy/5yX8AUwDX6er3
5SGH4fC78dVZp4tCBhAd1hgzkROJJF9YbLRfzNxEOqYJrrYnsYCCHTABW/l/B1v5v1aAInIIBCtf
t807dzoAVzo0h6UL/Vy6WimrH1H2VGfv0iaEKz2g0y63Nxe74Dc5GBwWie3zrnsV/JvCqLeIe2V/
QfnIdOzr/jzDHiJTlKY0JIffmY135Rq8qnadWe6UOMBILVmTu10XkqHfPtm9dgyekSFDAtYOa0gt
1JI9ybZIfjORTuEPFj1c0Aa4uBuya2eFa/Z34YjyOleOcx+pfnpRBr3VAWsMNSpeCuZdKi1/wHzv
m/zvczk0fJBCHAEv1FrzopBZQvPlSEWOpnaKa9RooSWb66fDafxnwcTDWz9xeB77DsBotYd6cn7y
/q4xtG8g+n0ydIa1c9h7w3qC0i25MiCqMC7CZCwJRy7DUxez9v17vzp+cgSRTS71ci1KlZFwXVSK
ZNERifdGTEHp8kjDtR9MZ26LWUEyE5i9NNbQ+c2+kiTY7hQ6gSeP47Eb/smJ/qlhw3AtxBruyLTO
vQ1qL6MBEGEthYNm0XfbG1tvvKygteQaOJiIDeJ0VjxEV6PkQ5Zrlt+ZmU3fcNRXocXy4cPdTW70
9GMkAb0h+RoPBS0FM3oDpByjhIKVqEWuOgDtsfVrcRGzrU0YAyM0jZh3gTQY/QIb6nIE39jqrD+z
5unpIevsaCrp7ujnNVdKSxrdd179ZLRYLF8fQz1sUnQhTZXFdNu5PMVLwekwuCr/TNi+cHX6x6Fy
pfblzV4TeNBnyOcs2kAZXLVJ7nEFZiDx1P0AfwDd+Tsah9ZCYh3tq6bEwZcqzaD2TDp1aoLC821s
aAzXl8MLVu78sUo3UwjA0lGU8UKX2oA4PYSKI5rBOleSaFpLeFpq1FMXHoy1s12zcKBK89MPB/PI
TDcA3n7xcPMV9vz5MnE222CvR/G960rit5p9GdfsDET6R+O0L4vD0i5C2fA3GyMr5AgdhkaEC+dU
BG2NJobamcPzJzu9IXmp6hbqmk+jgD1oTG7z5+81V28nET+tHwSq+v5GxZXHiBGLNaJorI7V1uMr
nztmyKLGSZfxzWgYXsn5I2kpmgaktzSpprxN07MmhxwnIZSX1CKy0M69HVm3NNNtIoGYmeFh132+
tGjT0HVrx1EnR0EJsrudfr9XZbwugkaSqE9cuU3/VshEAH9fS+zTgvqmDmcpaJ0A7+e/P+nPvBUu
qB1FA0+cIGuTdfFS4LxnR24EQ8tHIh+KQizG3RR8DWcAo+DxrPbKDMsK4TURNUICr1M2psBFzQq0
4bwH6NZA1k34ALp0YR323qL5A75WEOr0f4aVNQ2t/p+J/EJhHxQB84P8hWX0UW5G+G2DWbOKRA2u
VM17rbVNsp+ryCQ3iejMgsTIL4S8zszO/kxV+S+eb0FN0f1RnuMRfXQ6I1SF2EAGCfAjkl3v3kEH
sFXAqpxZ/zP+ia9hWWcEpx4Rhxck6sX4JfNHALqtqt5p2DewnTS/lQVEIW8K7bF355Q2ML3gn+BV
5nleUy7yZThWBoS0R8RCio44dBhiMw0HpuKhm+568g6FJXuKqid6k9LVHDeq+9dFDseOzUmv4EPk
WR9ZLQ8eKC4XtLmNqjpBDn0cnfDJVp+9WvKbdVv7DphZIQK87fHvnJapVv3q9JSxs3JAJCq1xEhE
a4nU0TZqP87AUp6jrbO+uvhLxivXKtMA6uO9xoy7sGI2GaU73BBtV0OjnN7acd3+7ihBR1qxekDM
D9nxcFx63uZC2SMjqXsFxZrQ3pTiA7nvhsyEOK96+207niwXpmOcRaNoWTtZTeRd56SpANpmpio4
kWkX/IKDO5H9bKhInP1Txdo7T8MWXV0FBtaE/gIfXVtcqUIs3cL3iIxmv6rTqIBFBc0WedKia73b
scqPLLmDbWQz/Yk4L1uAZ8QDTWWTktXP0ygzjkwsVIZewY0ceg7aSPuPDUcr3RyXNV5EQ6YQrmDd
Y6oxDR2vJvKLJUqfXZ6dNtX4ko5fQYVJXkjTrp2qGfj3iy/xYWGimJ6w/5lSHc7DgKj8zL/43zRi
CPbNet2ObKHi3SwckHIe28DnxioZeyxjf9dQjo8fTYGWYkeL4i/bC0r8IwW8ln6fzJKI6XVNDuUH
E7FYGf36G0q7DCYtPA0lZXcOf8qSWYThsoRna061xKrl+zVJzPmy9Mc+yi96gEgX5AbHb+6dmN/s
/p5usbit5EiJ4fPixPlOB/db/zqrO5/Xfl2Pdnx5HKZ2g0848bqbcVNFSQ4OkfncBsY8XwT6nYQ0
+RE+ijaduiBQUADtNjwHCWdKKgShUr4CZbk9+w4X+eXqYUprkfpEsM9zX/JDbDS0H5uBTqSIt/tA
icfPvYLt/xd2H6ZmN/Kw/XeNM0i1sbVQNuDo/tSiBkOFwpsCCZ4p66ORmnNhK6mExtrVakadkvw0
IQ85rggZ+lC11E9MBYSRFoYk4tMrLzxMruDbAlmFKDYSoeOQhtIo98qTpXtDIxQNCI4YQKSrG8g8
kqfyYyjVIAyjQLaf4f30vvJisccGCJ6nawo3MIce4OmqegQPdZ1QlDJScDp/bF3sHL/j20CoSZLS
WtQEpFUTWXyv9Sv+xjw9d25kxzwVc6f28gR+DwijfkHYhVVpmi78g0cM/kZcyR+91JfoQ1ZPZqFV
pMYYj9QH0Fs7mlrCMdwUqFbzfsBhtL6ltAqZDyvypCn7BaxorPKmJ24hxvtxoU2PIQqkz4E1v5Ju
dApa46JCkTg2FeLUg4xMsksCUywnKVPi+Vqq6/TTVYKvG3hpgiQ3SkbCdCsw7y2YKAKmAkD2vJfI
qvknJipiBZ0ov1JeiHlQZMeIKsgjL7GTkYl7MvDrA+XOWRV8U29IG3j7eJZgC1uLzWhk9Ib2JzDI
6wl8ug6sOUu7qa5lljbS+FQOBj9WjOLp4Arxm0fWZ+FaUnjxONrBLuAAVJwO+Gkve7SrGw7hgAzZ
zTuiFbcypKQqT2KVokFdupjP7pEIvQ1QbLpwXey2tG5zALpFfSTN8h53qQQQNwBIS3KEjDlM/2k1
+hn2rfEAn03BFGsQ7iUulXs7e3jaZAeklsgb9nDWHeZk4nIriG82RutJwMZ6eFkXm61lL91YsaoW
7bOtPW2ITu5iCiH4V87dYzJ77TdLG2h/k1pz6MSXMgy5VPNnfYps1VGZRYMwoXkCUPBYz+P15iJM
OcndFP5YxhBc2OXuo0vmpDBZeCcmMYDts9v7fX5yE/+1xYas+vWp7dBClvFPatNRG537+xV1MoDK
vOgvi0cfAyjZWKNJUujK++rOz09CZiYRD4oeR6Ay98GE50GbgtveSIpWjGRUJLTszqyQcdAd79/T
DaZFCWITg7XCYz2waptOQWqxC6kk3EY4/sWEL08xt5JlF5QIDmkRsG+KHl/zYDi2YkifS8nE+yeK
IkTHaBZwffqVLFJyU0BQI8rMhUq5EZkcYjNXtRfyzj9pwEgPB7FhTVDDWeHBqQxrgGK028Hfm90Q
HdWljBfsES9ja5eNeProUCRvDG5ErR/4V5EQAqnDuJ67e9nlNXq8uvTBAOESnpvrQc4pCPJ5rXEU
gG9zOEZYwpu0zbs+4E8R1iX2zaXApqC5PqQ0Kr4PISPX2nUZilOAczKOOkyWWRD/byB1dTrV9vNZ
D1pqshODag8BNuCPz/oHM5ewUqXMZ4vho2xr04U40YzXktaEWRTP9ZkcMBopPUgH/tDJl28XUO/4
sVSx1bReg1yzBeMjcWjK0swP9zzFPC9a5FLn6McWWaACYla7xcvWLw9fy7TWDq9NC4OU+FZXNOn5
PxAhl4FKdTehjUxqeeyqJkzH3qxyFPE/2Q1l2HIZRx4Vjeiaa+6OUpKsduQRhyit6Ze9uVWvbpOq
GBy3G5iytWWKX/083JeQXnCX4fNqw84mtMBIrLtSpoMlxoUK2+Oo5wJVwinY6RhVM5fdw9hi61dq
dFE/o2XpoD8a+uL5SO3c1dlhUoramGvoR9eTpzMQwQFJ6gcFymVU+5CVdpl505EWMfIOPfPochN9
CuxzngXMWOQuBlxXSxpes2Pq3VBYTJfXF4qroEPcM3xrlQtrwF+PFTpr7AbLKjsMW6bs+jJrgW/H
DVRUbuf/1e6ni85HAdNaPKbrEcTTBU3XDLMU0HIhba5Jzd4bG+3h69EO8pCBp0e5b9r2oSBfaMZY
7WNkTOqUxh5xkjNUqzdL0XYtSfq/RlIDt5SW9o8K8CLCy2mtKWqPlHPGn0RcDkZvCvdxUqJGTpUQ
955tOY2S/MrQe0l6clkQaTAEXD6JWvxW3c2aGMdlk5z3Cp25jKiYHwT05IvYL8bNvJhvikavVULE
cnz2hPG7NrF056MLiDWClNXT0593jwYKZziHALQ9+RCAQ73vUSY1G+Vg5X9iXhAU2laK62wD5CpS
AdHJyRvAXQdDzy35l9yArF5Ekax6LicaN0NsqEJSJ1OiOL8iqaTViedL0ZbaxJCffF6jae+f/3Dd
sWmQWbpOKM/Y+yKcX1YyCNzL/Da6GPiKuvA2rtXwHUMpOEU8VOrWifyz11G7B6zNm0LIl+kaQqjU
zKzSLZL6eGVpJWHgRWXHo+wPxOBGwr/eMJIru6xV2M+uHqw7GMUwjoz8zlkmJt+SDnuWOvzBuUZm
1GSWN0xfzqusCqQN5/Wig536qqSqtH6NiMH/FmLBAweI2n0zAbzyYadS7IOqvuHzFAQoTY90dzob
q9RMhxTRvCUBiu8IuwmOJi0HVQPWjnYgaq/OwyDBIpsrmaNNgYGeOHMSVxFVeh6uLlF7Uwgu4Acq
n6M6Osbwp8cWc/JZpsSgmrFH48zsj1v1dm96cAeClr2fWsjuEQjB8tv47BKYkJR0Xd0SQuNroUTq
bjP80NGKGFlzcSIb4H5rQR3ZIrf+mqcwxQOvUOVfGBPh/TsHfU9TltriRDX8fpfPNKswrrALuMNe
4UzJf2GnOgylc+UsBZifdD7nAZKnw7IfwLbqm7KS2veZbU4VNEB5SaMnA7/j+X1mG+IizAKjXXcr
6ulaaVDdYwVAt2TrVhUPZ5zfrw+MFU3oJw0r8iEtEJlsqGCCdhbhz1D7DOJ0FmCc3i0iEJvQyqNV
WVI0Wgrk58YjWOp3wzbAr13FOUeeKa906OxB6u4d87sAvrrZ/NJqJSq41dfF66FD6AnI++dGCk1J
UPu6pdEwDk1xBcl5nAcO9diKHx1lSwapWOq8uB+ER8EiEwI/QjkxZ5Uj5zdIcEnwqOTiSIzqXPj3
c8ykeuJ4RaUXFqB62IKUhXoQpvwn3HB2NJME84+QaLdCgUCR98VypAteL1a813CJiW1s8PdAIPUZ
wajbxpBreonpr2ZLWhRdA3Qs8dA7cZSr3YVXES9ypNfJ7J10aifBeeDTnZamFZxUslEUlg9kQcGE
wBwWDre6WJVC3RFd7Yrxw+yttrhPZzOkZuH15G4iXVwI2KA4DaYh6n9I16CgiC9GdKhewHWedV8S
6s9a8s5G/jVdOwh5RYKJ0e3nu1WlmHIcNqQZjh3/Yy14Rrit0jhW3cYYtNCkpX3nu73ofdH41Rui
/7ef1FmhQZv8b9Huec0qBLp9GTbPbTqdzfObaQNVzmp0eOtibw+GoFBXJe1wCUHdH6sNEtL4HfGS
5QKQOtx8wulLXtFrXk+kEv/nMhijteVAXfG7P8NOyCppjEjHHySQfCc1qjNyATehwUPihilS1+HQ
tL9SMokecWKGKlvATy7+y5om/AwmZ8eS4giWa6qIMANr/0bd1bJNuXh5JRJAhVBKGW8ME5sjt9+D
M+b3TmuZDc5Fo4CQYdj9KsvXDmof2Vc0NazLUsKUdSAvfytmAGZ6V/7qdghRNVBcsepTxgOsAIqw
OutxDsV7cGyK/9tZoogMW0n8LXgtYrsoxxMhttf1MWFv9u1X6z+MwuOiqObmhm/NY4rMxVyETokf
QVdkL24vKr1nkZEzxazPe06xEPEZiwaK7pDMRfgdgRB8aPug6Vud/E1Ja2N8RaSWEMrFVzCXsnhd
Tb956OvB0oyWFjI8EaTS9ZZZqb5UOtSmtLgjkDffe5gD/5geTZzMTdRv517hYovQwC96bUKexWPX
YuucMmQEoyhsxXukZhZjNW/g+I/sOL835JVvzlSNZBMpqjCFYXIb3PqDFVdnAY0NGdy071ThG1OV
lJiT9jjM7tjcXtcY0SKMgfen9L1g+iLvxcrc83RZnU2oa8/M0wev3B1Z87iiok1Sgre7OjtuMTjU
eGfm1pnwyTvknBmBD2W1MLJ/33c7hjfrXv1eBsq2jZrRXe6cXk097gl0uvRxhHfQgSMD87Y3HVQK
/k5Pgw2EJRrBAqNPPRZ8tAARx6RIfFL8QC7VDbQtEiIn5yL9EYN7/5oaNZvXS18B6Chj9WTH8UoZ
MdTRYZBw/epae/vnF9rFTQ1lW7XCXki4Y8+TVVNuzk1vyb2GbYkW8sUnbEZ/HFpgqVyk/uEQoju5
c9kilQij9MxHEeOLlNFhr9JeE1g5oIF4AKlUiAzCxhRaI1VDgFoKtw6Ffa1g0Hq6gosSYLVDXvXG
b1kQa/rlUqmIFUMJ1gPkalBsinzqTkUbksfc090L70FxfnMb3OUaa8tK5hwDkT/Xm6rTW+Hh/Wpz
HH3vxFrIKPapKRadHVuRpTm8Np0sU3AOwHYoxHGRA6XQ/cNwMu/QeFGlHBM0dIFka7bpLRTckXye
dF9RSjxfMvqHsU5Guzmkyv6mh+ojsugN8lUiTZjFKoeMoTyXr3L3Ggq/CqxzCVRSp3UhfohF311U
rqWiaDgmvrJAEZqJVWsFsSA5ylyRzL0qcsszHzVXar+BwAmDrdGQH8tCbl/+/48eHGXJ1nEkqnql
rlLZRikSUkTGJvrapzJrLF1Jx4MADORtN/eemRQ/ING0vuUepl4bUyyxT6pU1kTNYVFXw7SQsIO9
8Vb6GgX41wQipGaVJ0Dhxro9IJoRAUwPh5cK7Jcy1JFvK0Y4AB5h2rJl9uvCc5pnBPyKGUVRGKM4
WR5a4GtLwiJDlW+jYv0jtarlWEX3CRhxviTA7hpeUKiQiTIXDiF3VXCbFFIah5gnxtdU5tYHq9Fi
HkFb0qXrtrOZqfb+z+3QN8ZpU8bhqC6msgI/gaTUCq6sPRx+JmwkDs1KYSWbdMD6rLea46taduwE
bikb0cVkzsPUDn6W1DOp/y0UtKNWDAEhlbKN6oP6U5/LbBvaWNoxV/pkA6GMrcNZBhgbhcuo8qGW
EEcJdDgEC6SE72EitVFYHN6Y5Z2LVnaejAarau3nXMcDkH5XZzl9sAzpEUquWrvuxj/xIPF3ckRB
Nhu0DhLG2RepmaaTDR8ck2KdVcWs/pqOI8zJUqKdxgezuPdf3Vlux5MlDPGfVgoxdaVaQxlairzt
VZ8D3ykUnm5kZ+PfT3GvAfgN1whbvjZgOJJGq+Vvo8H4Yn5UCSS5r2vL+Uwcy+fYmOj5n15PCWAP
e5D46RwOI08I7grj2nOuewotasE1/1ycqce0OjxEAERLhIgQ48jtdZFznooryMn2HbLZXzIhkW49
4MW3u+27Kq0H5nCz7iaIgX2brOso8B75Q6svqjAp45Vady0qx2OZqiKoMoWvQBYD/dbdiReiq77L
EedSd5zTE40nL69a+8ICfFiltPQLmGo+ID8WPwxOJXLYXiGvP3pyqvL7FvGJmOAuqi52O2wCLD8K
ls27yocB5zS6u/bWIGhmaV2i5ZsW2JLw9Bze0LPppBd6SUwY5cS+/AeKITFSdlvzuYqViKNHrFrb
sgZAc1+ecw+P1hE+D48BaGoJ0Ws5I2avMnihnXLcWW3mEdFodBsXP/QvWcMPNh00H+Am74JPnZpN
aXxMwT7uXW6KfhVqMt/d4QZ05AGyuJPtIEKOX5ybKl/v2xZszdyTrtDhV+j4kbgdfoqkUrsf07QU
UZ0r4+6AA98Gkb01nwrrSxwafj9n/CIiXOAUnUXryHo87KLJ6m7PmTbrgV+d3vyHHalZY3IWRAz9
e0rpA+vpQdtmD4TZBYuEG3c7Ys6Xn9OSQ9be9j4YCeWZvKHg1KlSBmQzn5qCwCPaMY21y7GBXNpy
fBKAEZueeaEi4MztZ84Hf5+GTIDuj6fJhc0/3Fi5Nk12556UDbOfjBYp5/l2SAUxCBJ7V+XrrgIK
Mwvp4oxC0prWlGE1PREL2D95emZBi0NsoZJGnQn5mAvYDvJE/rXPh0abfKPY5eUjkrwTGBfkglrj
abg9zBujvhpE9/jKKILF3Hs7XO+K04G9bzXHBpG/5tiXrt4oa7R+81KG1s0M2wgPf0MJgfvUWkUS
OWPydi8zXPR52pW73r7QXZCogSKYZ1S9SuHv1/gWUqZ4sa13Ji9R4M2JBHiZ+TEfpvHYOIS+/rw+
lam1I3KwzIaMwcX/YdBkwrmOJy6mrm6QOfzd89hL8hbIQaJ+qd2qrrWCgWF+A56zfVDn+qPUOd4n
5Gkai26ngGrszgXePz9H3vWj3O0fOC4sKvhGI3xEkyrQldL2H2gI0n8uGQGQFyYwiWSRV1H6xHNz
qepsbD/BpF7nRrMPFFcRnyKQoqbUCJhSBAeJ2himaAsOkUrbkv6qZrB+Sdd8uLAs5Ug3vrlM+p7x
eTHrxtK1E0TuEQRXAJb5rLvNPGZOxWhJpzqzQGwgK2cHviMiOGcsMNRuf3dORO4TxqQzSeza2P6g
SAmuX9yz6i5BXQ/aDQd5E8Xhhrb7JUcp8w7B2hRuImK8d7ZghdyVfVCYGwry7oNqiblXRGlViTIL
sOjHMFoLgFWY+IA/FPviLx4tTiBLWQFaTVLVLQpFPrLJbBmc//f4u6ZgcAURWiYGY5z7icVo/6eE
yyuw8SoEqvuMp4/d+tfX7WDx40anoIDYP1OBvtz/u7N0QjC0gnKhQCNAbRcAj0u8p3r6dzWPAMUV
R64BUP7VVAJ6mPLuMcSajfv+KvT510Qn6lRp9o7l6Vaxa0rsXNnRCzVngcE6QoFS8UN5EfFCoUw3
NkmYD/RKYKje9Wcdf4MyO4BKbhTgfY4a/g5y9pE4K2b1YyJY/HxhmHrHdpBtamPidOvxSTim3PTV
yzqfasLfO8GFMSi/pPs6JxzBYYyDvb4KAiDYzvBp3vfo8V9K5Mp+MQb6PLZXr3FiDt1HMVoUbPh0
uaBCoAMksQB3tehzE4KWiIFhPeBpoe0McbEmUZrCHiP+IRhmLdwF/Yv5m5XGHyDHmqmZMq5lMivR
rgA041vUWNbEXiopdwB6OH+xBxRW28Q0lnf8J/I4NPRz7sZp/bWSC1rPMUk8SAw5n2x2j4fGhrkv
MbsxGxewKwF+lopAO/ka94ov2e65CpWrxKt+0KG21qbg2vORiZPHRKWwpoZ4k6dlVj2NevV3rUHw
FuPYu5JcUVay0JgM0kjCKDQRWtmBd8SaZ//q9R3HPkqhAmUDMfR5suVjSrr+B1BKJrkf0Qg2QNZZ
GL3mMo40DQpVpce/DU4DVa2qIsu+QVJCvK45XqpvwasLHwED9nATcllJY3aLBaSwxcIu7dqco8Ng
A3OdCJQRn3qWiXV7IUd25x5yNHP3yZzy4k+qpPQHl2RcMqcyx4jqtj3Vj47DzYqwk3hNUelS8esP
m6su9IePmxI4zOlNa0vrxZOisuXi7ewynJ/kJ5F5+uvrfY8Q9bx+fywRD1Z5S1FLIEsCSElC3eHb
phxVeQI524+RPIscC2kwjYwjjz1aQOqrhG+yKrKp1XALwtSNHpKcDjOauZs6TwAyhfRF1lcEJTFT
J5KDcXwTCxU4PuWOvWn9mua7AcfI7VqEb6EK/8Js6RO4Nq+HaAQMMKpWp+3FgW1cYif6qLNnM/Yd
105vE3nHcm2kSIzchcFY62MDoLAI/OaV6auza3fvo7dBwT/hGu2IfGKMY58WkGJ1Cw58usrDyNmw
Ze9szdYIJryh6WU001FvKZCP/Y2XrWqFmBRUd8yoQDAfV2Max7O9XvKit48ZwLH/VwmEzf/Vpi8F
wIY/1P/DPOrwJ8ZEGGJRfq3HkLAqMQ7Kdb0JTVRJsmYLcPuPtAZxveKVfN4tmtavzZMn8cq/pqYW
rx+I9Kg9ygWRFO2hxPAHRZSyujx2qW6+L0ODhKsLRDMeZDOrQP9uusPtWfdcFqzHwxKjr5P4rD2W
gqIg3yRAtqdFxdTtTOC6mBVbDOOQ93AxwB0MXNvQdUlOTE2pxOZJ07G1a22rfMSNOONsyfV55zRo
JRaRNa20yaYLG/Gc3iyYb+5hA/ysdraRc+Qwwz/tMgX2fKgnBMn6ZMnAt9iGRP8KJRiqyo7cEl2h
rsqwE0kXTdHcUrQXrPIqxXesFJpTZ2fzD2h4VV7nS34k9RTrCstr8sWhHVzmM4w1CD7R1Lf/q0b3
QByArh8/FbR2FARnHFwZ8J8eh7wtnam+HmNWi4AjugccKxFWdhDCFcMkCV5QBwrP0ffpl9iifh5q
RUO73zptsj0qZVOiixKW2574CpGmJnreJqAtbnWF2PKkrzI82i6rH3t7EQbWpVKsQxuElOl8Ci+u
tvpd8cArvTq3TALbuKZ4dKSo+cmbvaefvpQrkgu3gcXjUF0+vOaTVSBYpVk7+0e9yvz8nsSNllsx
8B0/xrGrrC5hzRirO8LDy3dCeb1+lSRAfHXU6avDxWjjrcQ3eDKcoz0myEVW8ALKHP/lIr6CEDht
W3vo3A34wK47qgwtgT8t2QDx+9vb12no8ni94Yj7RMo93k/GKm7V3aadoqW03hUOzk5IOm4SbUr2
6gdqjDHdq8zrMkUZXImZTiJkUIdD9gD5wsrDxCMlfSBrHF42mBaxuXz5Pdw7aBv7vaEm7GP5d5+x
jbJCgccP9IKe1MuxKkSafiawFjcdqRV/KcBIaNeeJMWLwvjL5PleZOZJjWsgCJqEIMBmOQZbKVx2
2l1drg91nL3VGNxQKqUEDgkHm8ME/JxMUibBIk0twGjJznbN+SVUZn9Bl0XE9ME1Xisxg0xMCQ41
I2dYyDOf73z2vw21UCCFBh3RxpkSxdX9RnjAOhQO5fLgiY5blcYqgtOmVd7DIq7WR8UyMNsrw287
w0+70Rb2EyCFh589k07w1Py6R2KeXI91BMJRN+25GPEjDmKlPfUq9dxDCeapyfQNwOuYoU9AWgFj
rNyq/mJ98UFCUPmkLTrBFM+r7+xNcIu4w/ErIBL1C+4gtLzSgwQheUz/4GIZGBeT8tra8awhC2y+
RiWIydf5TtCn048J89AKg4T11nPDh7G92H70yVZC5fS5QcHpK7klfUjziqX9NYthmdvTye09zNnw
VAFkr8Du4cyUlv2XODrHiAQ1+3BN+Wqg8Yw27SgBMjRO7pI9VVToBxDThjndgijE8zRzmwWRnRnX
gOb4UzkdsGndebuHlFkKgagvVdG/+o9wNL/Z/4U8aOx3A0tKjoHlaskU0YiRMG5w9/jcJ015ygJb
uoM5k18ThfhB9ji4hAJn9bBCdTvL1TZLfPbhwM6l772nH11m5wlXVqnaLPYvqDy+ynv+YQ5xtppv
LOjrQPpte6YK1vYkV7iwfg8z+FLruPWhMu+F2dD4uvbSN52O8uqL0HYZvoFKB41+Nii4j/b7WeNP
DE/HntfRR1yeJ/rjmBSW5Fx6stw9Qmc/RD2LeGUUEA/TKxLaYwVQzqTZYQ4EQ7hP+SluwbveJv0e
OaGRg6Yvm8d7Oc0vY5O2/uGm40IbfSMhwFXEIn7eb2BcdZScifZ2cBzz+Nn9pu2NoD2fOXJfXm7m
nmTF5dcXdBQMEdR+oK5uzfU9J8F9eKdHGIkc19FAAugbq1AvOPWBByaMWKFgRNrgMmIJ4LReliQ5
h72LGodWpOBOYfGA1tIoJCjyrG/cYPDNjAYua8PCbLjTPgqNotubl1yfpVrOtQ+O1kPqA9ytwuSl
OxfsnwP96flTn+K9y4NSIYTA0yUQhX4eqpchWgbkrNC4m1fsh+fdG3FsHpQzvYdz1YgvGx1q/kdR
/QlcIAd3zKC5rT++OTkWZZvjPnV6EhzE/UghtoBUUxLnush6e6H8aixdAfbZtjAXRaFbTUtirAT8
HlVZm2T+LNxzGpj2esK+JCySlA48JCo7ZEP3A4xLUJpCFK1+LRSDfEAWADxumKPNiFJ553HrTr3f
MWwzmtacoCrbaH6WWt1ySqazO+uPkqs866HGG3scdRf6Liw2TuzqhyRdnGqnQyJBUan76FLNpUPA
0B7f5BYUixV6a/rwnHVpzbeoFxgNl7o9dP/JmAf06BEJKRI3Nci+NkrUZ5mV/GHxsJyQdMGHLaIH
yk6ggVcX1tsW51fvnHeVlEXBU8/YJyUJT0LHh/ZPs+EJpCaT23tCabY0S9RfUprwroV+6wU+GYId
FU++6mMV1EeiMH14ENZPswicTq1q9E+pFu8KTGQKOiej6XSWugd1pXB8orNqAt8XiFBUT3j5Z4u/
bKWHbrafRAODWQ8DvCUn6C4Sr9/Wua47HpuH5ot9HFaxqRpbxJ4+opEQ34wsdG5gLdf/023DNS5E
CcQOGv7kDnfrzLUI1qXyaeM5QH+gnqD75sfN4jy7L0iuySPldzEtdduzQ4OljjgxBtZpwvkdwP5e
xeujTp+chX6fzQ7bTfW7pvBO9Ak6+CcIE+B+HB2oeDfs6Wfer7gdKdDKVTYr/ob0eh38+kDBfPmU
lId0fXs03MWdooHN1Uul6inRndxJqpxZvu60sw+Yab+EeYYIQK9fQyKmPP6rIyB9+zzqE2cHnfDs
tv+pKgr4lNxrIqTMArwKhx3yo4VK2RiVCvYpNLIYNaPBtH7tgaheNqeRpRqWPqoMYetb+oZnfpPN
8gdIj5vEFOPFgChg8ZEY/04wT+DWUxftNdADlG8yaIEDt1qCxX/I9iIbvn8mYi3eIJuD3IOinVrx
LgNCZpwOf2BjCw2YphUlxN0KF1C6nh7frodnlQJxzOSo3V1QT5do1r4SYu0a4+fRzR767r4XPMxz
EVBk6xKC1XG9ypl4CRussxtvFaVftXbjmJP+a1IaJvfJf/PDDOTJwbKuVjkXxQQzbqWWu30UZBjs
pK/aFe6z9yQVWt0DW1ck7nynB4JPcGbmDJ2vBTG/eEa0lJ2msnh/87tcmHA/oPt7Jo4KHJQ/vFHU
IZCvFs6x9iAYAF81SopUpj1ItBO5jVf7EX8vtoMKPVkO0sheTYOeG3BS5vMeYVGO/YA5CFTZehfX
LEK5K8mTNkytoFYDXberg+TirtsL8yk5PafAfKvR5Rcq4hvyD41AZjzhHwun955cwHHrg2Kx0BKG
WB5bhGF8f2e6kSO+pj7hjpS7y/gjlyWNGVpj2hhDlpdkvBpJSkJGhPoArbZwh1TSojXdCgWlWWQ4
PCIg0Z7F1h/yXoWpmeg5q2iTokbLjsgAwplYc1PVRIIFyu5EK9p9zSA/0+QmaRCdrQvk8HKy/Puz
NOJPRqPT+CO5KuyhVnWFneNfn1pF4lJrvM9/1+C93vq/fJoqMB8yJYIAPRdQTMGKqWya0q8GlgJ5
e2j/l/NAjlNlVlAKqI6FyDrKfYdXXsDMisOj83reS7t2iA1Qs/Vat/X4veXKrDkcE24b1A4sCkuM
acJsY2ABx3wyu/FSuc2qgc/z6WpZ8TIBZ+FWsPaPrzabUnRbYp5ucncFrTkZRf/jFOZW+4n3OHIn
Yzbnuf6PEva3J1ZHvrgZoSkVxpCooyZgsnDp6jjElrLYB7ObiZhHlfFvKI7AYcopTfzxSjEYC7EZ
uflhkHNwgSgCzvvbYqWZuUakaFTvu5yWuYl3mcyHeLwL/ojCyqEl24RZByzeX4HI+ySxOLX45ohr
BQLWeP3hCEmGu76TVQTxd6CD4AzSrjIF47svN3z0wiSbYWlNBnRXFV+jvBDrxmzpzyhNaGf3PBk1
QZLaL+07IAXQiWT3INaZ5CFM7yJ+rjNyklDK9G5l1Tnm7aBZaHcFj8ocW3iRG4o+8tIXw/09Ecdk
E1MhBKrikB/h2DlrbUJsMewvZ62/O++cPCfSHjVSP634MBq34POHV4pun7WnkmU9cxa6vDFE367N
AkOr9Hccg8WFtmj7PRBS22Uu3Sy03IDKtsVMsBndB9ZLjNQ51RjKaBQyu52a5Ovu9fq3ekmEfT6l
tooAuBggEt0TVz2GHUQLEIXPC0GG5/yq9aZR1FDxSAewRe52SWSQg4EFxvgHooENIBtxJaMHQxSa
QQqKn4gXkR3fW54TH6/w3Zq980HcCPk8fLRjawFj2M3SbS1l9b/l8rd2/LG/Qk2ySHf97DZBeZGS
7FDttcjN7t82d+y35GxWRML8BxjEM1OPEcV0MbBtTQT56mmw2ZJ03i5gggKe+13c/ogBaiZDW14D
l2hU4bg9drvw3dmZd2uNU9U8ScaQJf+XShl+WSrT+/Iq5At4jGSmusyONxyweiV4T40mlcK5S4R3
6L5RM6/eyvOo1W9Clb16j+ogoM+j/454TPD1rVViX7fvB3cYV1jH65kzkdOvM2M95JEOqzaapVhj
dqYWKrNknd8vOjZnA0Bik4VTCYPEYwdJIMzycPjyP+0dAuYRY9ni1Aq+kLrAVWtvF8ynXDWSGajv
7iULs98QWmVct5n/YUO357FDHfHjDl0cVcVd77KLJYMRtF2HkyZrByVqpfP04kU6fQVnuKqWokX+
h4w4O4WFTYLudvOF8K66zBz54Zj4o6MIG/u7RAs3oI0FEmJOI/wJus4R/LbjM1Dgk9EbpnrDnAwr
kpEcoAJ1MR2YzSuJLOhRQyoT05XhLZhdzHrfekG7SY9Sk8j81rEcj70qGGNRtYM3XjxzSyHlEMNr
EAt11l7cMqiP/n22LiD5ubrjx378qaxRXdN2KNOXskF/Rd+pftguJwhUQ8kqZ3Fu4TAxTMdOnSm2
EXR3+4wcdILRbMAff1NVDXTAU/feDSuYas6ahNqG+JJqPucu08n9xIXiYGjKKpDTUbWJDJejNOEQ
5Dp03BB2ACd5KxOE90AoiAOPQ6Cdbl6w0X1eSpdrHfMc7t+wRVecXKypWFvS+nyb696+zyj6VYl6
m8kgbk3QIH7UyghcMn6kV5yZIMwf9cb7m+C/1uRcraXUaoG37JrZ+6q+Ul0PjtCWJH01V+cRf3vp
gyQS2I3hv2FT1xOGjvjzRI5wlBczroIKQwVznypAT8qATCgkp9NZTfO5AM70VdLODz+tODhIoPKX
Tl9qmFaV6CKihYg2gyDcmnRilmhYhcF//CG7DoagaHKvhoIs8tQEokJe0QgtUCX0XkgZp+IYCF7e
91J/RA5C3UaHLRedlvwcxOgeb/xha/F2UPEacPiSIQHmicknlLDcnVbNAOIqKRbMMpLcPy9Za6M7
8dRv+m3PjMxMFm/N1dpLROEgWdYQpgKQPSMy5Dkmpx7YCg9F5kUd0/+yZdxGmVFFO5PrAq0eVQ5q
zvwG/xUhaL2FSouM7UbZYLl6/EsmK3GEL4xEuQ4I9xI4QS/6jzWdiTeJ4jKd2uFCr6Q+YPT+d8nA
lO54N7h07pGoMLb0g7+0EbYu17AK0+LiUTQOXDfDcr8VXxLXjIvstYnryRIPqx+fFsrHmS5G5YeR
Mxe33mftnQ3z3c3Zl73qQjmZ41EIuS+PosDAfERujpyc9Dfk7wV8bqfij03oM5LCnjNKLaUt0LJN
4ePKZrwXTJFozFtdhY/wBNckDVm2m7HT3/uq5RBHDWfzD5RCP5Y4r8RrMB838f+IQX6M64NZDAdU
lhUw1DNqBp5pzJZveRMI8fkZEggaXWCEi8bD/iYPAzJ3ybhRg+fT0lAtS4bU1LyGLKMXZhtfpIfA
8n0vHANLdAN65EsYtdEQVGerCZjITvaI+sN6izaQm4a1v7eqqkVlA6tUlZwACK/46OO8/SKgRt2X
GfrgxZD+DzJijGrgJdlS4lYq5EW6YJppTfGAfL5Rdm2wOy5h5rBRcrBu1kriXkMAcgsM/kC5T9NM
m5upNQjIn6WFpE55WNWfEnhyYfXKePkGWn5ayGNgk19xCkLBZlVK2324WhQ/9snPZZg6MK0JrR2D
GXIi2g+BugaKpx8ofNFh6q3t+02MiDN8LkH9HnrpbZ/8zygNs7rdEW+c8swjJdez90JFcnm/7JNZ
7tqtQ5zvAdduAITj0E8YfFjzqHRR2C5OmLHztBjSDW+5mNiQbIr9xjVud7QTIo/lSors0znJWlex
QkdT0LQFkKFok17vMIMVlzFYoS5VjZB1eeAbTuZR4nvKMNzJu8pIaYJr+SzGCs5c1MsNlNWKVfNJ
CbH5nR1viWxj23Zi02ivqnrTUJL3OlO/MVd6MvhgMNLHEnw88hlEaocTzBQiBr7V7TLccjj7Z0mR
0m/OSjfWg7wcQcGUzkm44FLFSrRIxT1Y1wgttfA5Pb6ze4k6k7IVjzVyvXuHG0hbeC4LrZedG5Jk
oRw3rP4Mmqk6fI6j35vC6ip0Q1i2jonQ4ujmW+sE0EbmO8AB5oIuLSz6P11g1rDnnRWh11Zq660p
jJufAs1tvZ01EEPiMfyDOXsA/mJTK+e8VxU6ZAAjwo3Xh/reH9rWKwUmMH4Firs4I0Ceqovugfeu
V6vMlCaapysRHo428MM3wxf2gaGq4tWsM64vmqRD6HSfmtywCijcD7wavz/kad6R8DmmopknkTbA
47FYnvRbkPSy6xIRO2JForga6miOg/H1ymW+NTd4dl+SJSueQr9q5fO/BvlTPDrPk7HRGE8Q3/6O
6NCYUtxFZu7XRpiSE1Lj3aplcPBwe7DibycIFUZywIPWjk68j31mh0bdWpfKVLQP8uihytTbCgmO
sAs4Im6b8+oErr91x/9yYTRtFX/x2wk38pljg80+Qvao8nRTVKhZw/R5UD8dLscjHf3UOzGnuysw
9InJONDHWGPF96ehrKRpw9F9pXpymQ3YwLPd3x3JjVWKySdzwLL5PXY5EkrjjuSk/VvOt0wWOBM9
1IIC6+PTGokyMgRGQCK5GUHM7iUxOqSPExI+cl4ZPZsAd6toE7Xl60LZd40E5ZR20GPMMTyaSysG
RJHMgjf4z9ipWtZA8ENN9e+ZdMjobnO+iGdnJgClYi9JDMlHAFhLYGUwg0H+8EDs+b8ES0yxsu6z
KBc+NDMyf8jMr8e1/XTGPb2QXrM8it+/6EPVnvHvxxFGzSQjHE65ZrRPuYxGwhwZwbsb+GoqMUo0
+QXODBN7eNspEb4uggxNk0mw27xqT/ZvNEdGZ5KWcwEez3E//LV5IY+tADUXtZSJtB7753jwfo1K
4S0pybo3MnAqad5pg4bp1e16wJOXtZLAea7m2SDVdpjehA2S/NA+hI6jQoEd8pyeWqOIRLVpHhel
ksWtJGxo3t2M3gAGxBBiq2ezo69jHTIEVYpDftxlRznYnixmjlNOrtE/06/0RRTZVth3JsuBc4qa
OuQ0RV9G3EaecFUc96rwHR8hfhocJQYg/KQiXKKFHSkBpJ8oG6CSSmTnHrvAxep6C6vy9uo8yWZG
IEnKCJ6OSyJsxwGEBYWAcoG/QgdeNnpcQl48YDPaG+jPppcpatynsheyc/GlgY7ztVO/Qj5uPuKO
eAv3GQITBq4oXw2bXfv+h0/mzQmjy7AEmTTimzxCDg6GSASIk4lb4iFJAo++UQULQDM89N/qfP2h
XmF2SELv9pCjrt3hsU8Y2nJVUgOiCcvOof6CU5draBNhlQj02MJpwY0nAC+8L5AFQbcFx2ejhKjK
pDHG8tgOUAMCSOfoeZHRDCyMh5Z50hg9sil3B6CYHUjN1KPEc6rk57fJH11LgANPsnPqCXemZism
t3TynpQvAi2KpV/r8sHb80PJXvr+EHev2TwQHKCKkXTZh6569KfULrPT+9AvYOeeIwy/Of1dY0EC
RgZAo1cPG5ch1ggt7pHtF7imbUd/eKPFZn3eeRfY2btGafPHlwOmRdByU/w9+FW2rfCFAWFaOCxa
PiULoXN0W4ZPbupx5toLsdPFqpVRWH/4XqPFNpselvoIjmW+2Kc8N6iHKgaz/Xuvea1K0AYBdeqO
/FLX6HL/jUnRmsb8cEUyLXht5MAsPHACIruskCEPhF4CK/uOFgDOQenhx/tqd9de63mJFi7kVZUj
zqzbjaCtX0abNeT66sw6x6I9MWW9hwQwWm3Ak+qfp8svU4fksUv5WnjS5lCxAkfwDlIqVjoDiHOk
7Q6Jd0LwSsLsBdx/tdOwUtzFsWv/JAJCCAMGXtV0PxhS+Y0L4GC5FFKiFuS9xF6XPL6LoamvkLKE
YmUzQ8ow82vbqVZnJrN/2bXpbcgGPsN29tTgWgBi9HeMw4axA/+X27OTWZqHO3yaw3EZiJG3xj/G
9wmnjXr/nx1D8mfmtzBj9JIz+pJYWTPb8ZcfM1eKHsKD+YsSaHJKiwImZ0KbbOZUeuS6gCz+l6zw
sULsjKx08slUMlh0evMtQCEezeDQLLOSFvGQQ5J3e8PRKEywBnxaMypiskl6DlJsyeUeq3TZpd6L
lLVW8ZPrjnfih9NpklgiPC2HnL6erpLZTVH4TSgYd+QXMuR3dq+bQMS/mnOH1AYW37f2qm+wt+TN
GqIh89twpm/sdMcxp3rNo4AkrME/qUhIElJVvcMskmmBaR9aK+sT3VSsI/UCv8HqrkTKG12vbvX+
YzHLPTPAOoxIWhMioNsdjVaRTUFnm7E3lc58c4WDp3irUxJEqoxcz9VwmcqImwrbnNWASgomBnH0
J/gkxB10ner3hWrEYp4L8pMvksp1iN3rhz4P7ZDx3RVr4vqfnDRvAGv3Kxje6c1N89X2kAS6LmFc
gX57nBjJVoQoqriU/T969pce8VwaYavcy4ncZsO+f+foP2qV9SxmTzphQmoq0/Zkh+UTNqxH78sK
AlhgtzegvaOezhYj6AAEFD7clKHjtoCXKNC8kkvsnbL/n9SsV5TdfcmHgQmQpvxERNhA13iC2/eG
6kNN6dCQ9tS6P3bVpPP8f/c0vOMppp4RuI5HmCuHi210sOW0z3pB9NJ/DDY/TaJ9VeVd2+g/aACl
a6GvrQtSXXo/2yBihNbLyO2yDNLvDPFOXbgoONds7WsVWdncS+fiaT2PTcAgakyrOmWDRE00x/kd
JlAR/35Q6u7r/SLQfmnWwNpASHD9zQBmEnZ1CmD1XjhCD9aBZeWdH0c6Yv2tgLB4FYXZN03BebZf
PTH1XfFWjW6CLHxhrHhirD8bzF4LzE1VYfdiUMSiBAlohfue9qtqXKI6FOrB+QgXYxr7Rpuvkg4Z
H+Z7XHwlh8SseKpQ+OKOgtRXkfs/5RvcYj94AlV6BzHfOFRx+gAleNbamNF40JnWS0YaqhP/Wdl6
hjTGALCRjtUQ3LfDGl1qHTxcAfGRpFUMORz54B5kbwBWv+xXMKr/bz0LojhA0JXFhq7HZTwVs2Y9
60UxFRANcHRPwijgRDc9H0auV+QnVXSHhSrDDeEBKDzjTvU/b6M7BlMQFEAaAl2Ym9niki/E6CUk
mR+MoQE5g9OKHFOnAJaz1nti5Su6OkqFpORrmUV/V+ubaVehcAacdOG+smhz9JtEs7AFdUy9RdoV
hcPygUCbwzUXR5M8EWuGKPxki2ZeiIFv/CtMhTP9jorQi9vZ+rL5oEIKcES2bQgoKQ4Ibl3V7Jtm
XLhX4sw5iGgU++nP7krYAi3KXSu0vSVAQVKnhGZq0uVU6nC3afaB3aysr0aWwQgMT9sW4nbpLhtl
bj3puPRhljOS5F98aqg0ArgrG9+G1etuYP4J0c06aImjelVuD5+VPcCdxo5jWCENg0kJLEGooR3H
PvTA9lVnjIxDYEtEZUrGQjkC3b30FBrP+T0DO5A+mO24pKCLWDnOZuFY0GdtrVTVs/Hx3i8ByU9b
JFbGrZwOH552AJvVebcVkaxhk5eaOW6/hK8fvvK3cX8APk+Hi4/cM4uVTBW47shKTUkWXJmqJwsP
AXoaXI+ry1+kz8xCoWXum5VfTNaWYI2S78qKHuiMMmKf7xqkhi3Zi3dcVI5HUA2Ydu8hBjdHcb57
ldNwr0ummyR/5PZp0up7D0oAKdrgew6sKUiExP69QwqkLmKJa9kYDGtZP/XxG2czJIkgdOcxnx4X
/ZyW7Ly3sg96gb6BK8iTIU7CDVD0oFU8MjV36dN761rCHhARVcUHfZ647kc/TxL/oGOdTmhBZFBe
hTb3RllMebhmFd09VzD1J7hidlTBVp4THOrd4NbEMmFFCgWCHyYG8e9Z15w6LGFEMvp+ggPhkgiS
LpXc4Y6BK1yTUPPrswJqbGN/SoA7buFmNeypHUkIwocrEaQuDL60Sz4Rr9+RaM64BxZOkJReVa+r
pNLhiTjknfTK1WioRT3YELWKJY6obRPmYtJbEPBCp2fnyoUsdPToIfChZT+EIbNXFLZpKb44XRGD
9h9TcUrXw5O3GjeUOOFyItubL4glIex9ta8YoS1zMYuprEMuWIqn93Qe42o3X0dZ/lV4Y1hi2/Wl
ABP6tWSv+AWUE1hSDzrqw0YrXvmFqdZoc7RAMFjzXNGP2E2W8OwV0CJgwnslAsMiwaHeSE28sGTk
y1pxucChm40LSffUrb4QNM9VwHEjD9Wl07+V6r4NstighI0d+WgeaFYSoeEIM82d+ZB1AGRpdpFt
LnmYPg6CLwdUplFrHMK6Hyhyt/QZlMb7BPUozD0lVWc/0r/8Vu6UaqffvccEGVnBMtANTLzSSrHD
vmhX7ciUnLuPGEpFlrYWbaaVBoI3UZ1IYHx5uMe4MzOOgx9oRy0ZqE+DZs81NIRp3fHoDoJvymFu
ABOhhedz6HLAjXBTy5XhNnXNugKw6I1HSckQUenMWxKiyNW59hvihM/aWNGakqOxyD87keXfssXy
VC6ytiLBrM48+SAr8e8lawiqpBDqekJX+0aa2aMsdYvJF9FB152jBxtOihuSOBCIsXTkfnSba6YF
Z4p0UnZ2MIMzgt7y/Hqi7fHTE+JEGtEf+G6ReoE9opq3gm5y1SN58t0HjDraHmkzibgKsi1P+04M
/MOAAr+pk+NKv3c105+xoMtnd1PfqLhY2CmBBx0W6BaiXbpU6x1T3g3r1NmWXTmVLqGNimGvJOzk
o04sY3cVBf437bRg+B8b9zH7rs8geic7INo9EYN1lqrYMGMjhjStRI1brIt3PjAauvhdv/Obozj5
k7+YJdZ4LaE7B8srDo6eXrx9I7AfbGDAu6GJvWB1WoXvBICxX4Lkq2v/GpEVexs5c4OMsXueSPOb
SXnsx5CbrP24DaCvMyfwgHEtrnzQCMGqLjJU1l42lE5Wn8RBnlusuGFqVy8bM+DqURBqSAweCqbD
kdGVi3d6KEJ+LFrAGKGMOzq+9Tp9rXASJsSTpsra3EtNRm2fl2rYXCwRpXe97iTzlGteRGpA6Vil
YtVAMbwassonLJR2bg/oDdy9h7GfWFPvzPdqqyoANWq3AxZE4B9t3X5zRF97pceXQiIsIdN3/RXJ
1bd7ixCIClNVJw5E3wLnrDmrX8jEfrmyL09u+TIjfUvBfR/mjqsChtEXwcTIC6iMeN4nkj0xovKr
+ZEKmZuMSeKry2ZRL3ANRSXbLnQOPOvRHHb9p6T/Hf7w7wB63+lbacYSYMdLggkD4QrVVpNQ+4nx
E32jx88eGC3plHO/sDIMkrJgngUhd1tgroUmQPCzSaPjQS4PKGeqXNGBiald8SUaMB06yn7iWNGP
gqDN4L7nMmxYPVI6T4wFuTGYSaFk0KvPO+jT73ImbfkViP2GOrH7+pgHLIe8daM6HG+6nLGxgXvD
xwlQZEPBDzyRzqiSlhpXgk1iNbb60zJXcJDw/az4ODcDibcJTTAwkIj1YCs98l4rMXiGc5G2lWeT
/7GOYkzTHagGXCXZ5to3bkJ6blqmepv4AjgypD+lFr+NpddzvOzl0fBWErx3PSeGebEQ9nnsesyK
fBrv/Te8/d0oxgxytnqv7K+ulvq1FTTRWLpEZqQnhzwqguGKv/MVjrOxq5zOZMjUnhMyLNdJC5Ne
VevB8fX36/qJzePpvthRC1Vi+W35/6MIxloXAVsaH6vK9oHylv7HsvGWJCeZdkp2Em13AdO5vqXy
EE/GtLdsE9Ub00En09TZ90del5T+QILFW7zHr2BItVFEdKMKMaco30fpM4nuwzIgkCA+9W/ZLlpk
WGKX5WH7oTzzQj4WopLlhhrsyZZ1MiRYbGrpm/k+BJaw5XkIi9FCsV2OxzCdxuTMtkv0mcFQO8HD
fRcH3Q5YVzP15ZizxcIojKrfeesltKwMIjd62d8q42OflmvuJgkSVYRHOZErQ5eZL4Hc/p1Xgftz
vV+kCQsACuPLtnyrd9j8A/1GX+SxVx3g66wPBRuJSbJsBFncXzp9AJ5ujM76AcsCXMeoaY6xl8Yu
6NYpIg4sHONwDC+rhl2JyWKPqDgufCLgk4YM7RO39AwCQ7dqpNSrtRnhK4hmeuSs3srGnqD+l7Qs
Ifvv+Vc5+zEyYivSXQutpOd/AnRI7kKWf3D/3Mm/JcjkXHeJ6UUUMpSuTC2ohgXUPuEQhJFjVgCN
LBjNiV/rEaLJTk+89rDDgtr1eO017y0Mj74hHqhqhmHBWBzFzwz6qoIx3KpCP4pnfVEB6CRS2o2S
yc56eUOGPTjSNhHNe/ku5/T2OTRpDt86YUi/WVDL8eskJBiKEZtcmg/vYVsikCPCE7kDvr7lzVog
r2SKxvbH/JJTXQETL5LIvUVyvQnBzDr9mMD7rDWTgL8uA/LxL2YJUAx4/U1O7753sX0qw84ElW13
dBu+x3GPKoWrz5VpjBvBza9cuOVDKNikOgdTi/yCaPBkADS3IJxsvPjy2iLGq5jDZKFvDd+iU+WF
ODXCbPCeFBpgHFLmtB4KnKEGxvY8Qn2GWuiX9L/B8patDzG+xibjnSTK9JVAsecr90C18V/UFT/k
JaXhf9Hu8A1KeQcU26bPQ/KWQrVbDWv8AgOgbu9HzzFvtBbMuzJMhyucDsgE9bFYp8gggyMsgG7Q
Lr36khT9KpPRb1sJlUGqkRk9YdK0pJA23AEQgTyeVrJIMyDYTbqqFTwc/Lr3TEXMRIyjjpF+KTwL
73Niz4GjJ4nLDZLplBJ5ZTUw2P8xWCPbCb+iMeAaFFKs94FNYjpeV6RidliU4Qcz2W2mQqz1X+xh
5qwmOfUxjDG3TmgILda+SVolYMMMbvi5Nc18/2lp9nJrlcJhx0pAkrh9TnjLfn1AQe7u7w7lzYJ5
4yNJGNzDjYKCEATsh8Ne8fTzDAqBlIP0FnTh+Gj6pG4W/U7ZwBBFOWaIARfb97EQccmdKCFUSwa1
PF6IhYJiTP/HiRgWBYi8+ds6Z7znxOuLR6iRuP0GzrsjBtfKKlbe4jRsZx4v6YSONZdIChDPRLBL
lENqCZKnJ6KBrEx7HjyA7nOa6J4++hEW3uoSZYjqOn6OcCKHX7UA5+tNBRngqpN1leqZjca6yh60
uFARwGKm6DOWKI7UBKiJnFicK1OFGHgLIuLPvRC1Gt5BsJp21pVJXify2eYvM49vCwXqfYr6L4fV
pJXLHETP31LNncxYiHChs/qxTz2+Gdw/VK6hguW8U3WjCFiNPiS4ZDs6BP9vnxAfSRE4xy7B2naP
umTj8WEPUYP4pP8M1X37h/BK1YdvisL2xTwb53VsRbDxLjfTbmq2h6Ku6bLU/JhHh9+5bE6Q3Jzw
d1dxTmogUm+1BCZaw6b/I4YxShExWsFjiIsGvLqYEi0j6BUJfxVghFqppNF8LFkIFp+3y+cMFO4C
d7oEr2XMgEpsuzzpLnVO+KuubC0FJL9aXPr3pwN8NV+ZcZ25nv6CfXbDZIAAqYv35BYZlOOWB0wt
fyDl50NDRKlpNsALYZ8Iwkhe7qJkEM4one2JZ/7uwZ6FLaC1isEUKofaqN+2fvgWlqnsFOGYoNdI
tamFFSqAclRqmza/59DmTZtzsTKM2K/EOuyga4wQI6TVSUnjO7wT5y3lM3PyytZDxtn12f9jRWek
H8zsnNHRiOt3UgJtxizomeS74MFwiFWhTe++EXDy0Fv2+VnXPk5q4fmhyS4bBbXC8dWB7jO6NTyN
DxZ3bjjaYbDu6x3RXxlthNfDpB0tGk1PQuWMe8BMT3SDQQt7TMH68qvBME4Lp/G5yQtF5WHhwYL9
AWwXrJxLvikzf35juQ1AwFpkRcKRXLTgfHwaYoqp5S67FoANvGlqzRq9MyspbB8PRvyPUTfaYXqC
1gYMV1igAMQu7txxTKuhiQVTCooVKoDSjJx3ETU8Gjh3GyPg6V5zFuCvWNGXr72lxE6PH2ruY9S9
kX6QmEqZ0MG+S0J1JGbjhLQ0jvwKUwJXDGgXXsFTgavqZBtd8ELV1WHOOT1WzfrBcq8GaFpwMPLp
mXjHHccinLnKRl3p/C5mupwDduw6b/Zk1q/HxLCvNdV6aoe0i7VzdujGYybwwhHB/giqnpZUiPXw
vAEILRs9hu7Jco8woHszxbphJReZRgIqTBT/27HS1M0ZV1nQOty9cLp2uGZ32hXUIZZdCtZAlAnS
oC/YFZuean+GCF+yoNCzJP5GENE4omh+9c9JR74fq1E/1ONTGGKr7NooksKi4UlAQH2lpqFiHCB2
0H/z7fy2TGFN+wAnNmpzvRyyn8pqO3kBmurQuxz8BG3fqOkzYPzZq1IoSYUdcCmVVzQOgfqKSvCT
BZcnXt+tEUn51xRAh8Uey6BJ3sHzpPDcS9AhttcTCPIcSoddFeXk4GU+Dmx39tH2wwm7ZOpNPELA
cfILLmULL6EOFVObn0HmW3GE9riv01y1bI0L6IzITZCoF/GADbiJYiuuMGtcmbCppvWjqIn4emVx
kuFIyJ4PkuFx9xZo8+jdQmZ4uaD0P8odRiXAGI2QyKxcpACZWF37pkXETwrIM8xwlSt9QOoMsRbw
3xdIEhzSW9bgep8/HyMow7FtNXbjRC2qqIfLfCNEyP5rjheNJZWm/X84SFqFG7y5TGEvycKWFPq1
ZDgK4HiUWauUd+RyFIZ4+ktbD88YUCtVgVMm7M/9PIkZsadA7H1YNGKc/Mdfe3C17o00Nn/u3u8S
rKEl5h/NEi8fTRfmaKDnLQlgVekJBXT50PUwgVgDYhc3VEOcWFGL1WXKEDnH48mlzEppI688Mj2U
QWQHJMj+YMyLQtlUVrvjCe6Wg87tdTiage/eFc2RpyvHYOTmVvKVT4CsFrnaFQgm+Ul4DyGwBYri
cwDS7guN5HKseoyay18MgTeBZ2NZXxD2MFl1yyaI9od2qj+Iuo20iNUhA8ofOpA28zmT+nDNTzOK
XNhn4Gdq+eyW2vxfCw4+Ck4lGQqv/hovJwaxc3WVu3LURykP2c6qTiSH8tpHzQdGyxkg9h69YQ/U
c4x8jZ84iLoL8L+eIn8UMqe6LCtHZSyar8k656zs/u7QDk6U/xt/s89A6Ttw1oM/6ZprBgphhe2p
xhB71+6xIaERtHHKXNllHTwHU3LfpCXFsHD1y9HGhYRa6pp57fMCIkDhnrKgClxPJWCQVkW1o9+u
e8yk5e1tFkduGF3y10G4436eZd4KMm6oBO6ZPV/BCafDkaokLvOzuTyQORHAHAod/UE7goquvaZ+
AuhFQEV2wBP1HcxNsvG1qPaDUVB0nUO9mXQD5pqcW3GDGuBxDIhuZJwMvy1q+u+FdFJEw/0atxXk
4HQeJLdWJMgE/bT/s+sQ01Jc3cZpm/S8IOS93THN55rGUUktz5a7T6Ii2/qYeksX6eWnNjpb+KVJ
x2JDJKv1QBKirJUzEau6SbklAaXM6ErvDQAh1kBonf/KQXFqrbSwKjkEACvin8b33FhxAfaZY6mo
S2KybYANfdPfjgAXpfxvubFyeXGmtBJvCoyDnKkqjYLBz1iqnYFOhsSmag2ERC8OENEBwU8xoye+
VSythC2d2EMj8TJRXtQVdf05Ng4vfMhOwwvTtqHY3PLsj02zDFqrEzYWFT4rdHixPPDQbpqznrbi
5BUcSx5ZQDs3lCDYK1KgI2Zmp3/OIbVo8/Poz2ELU32hO4W+m1l/8nX6A4P3wV03zE/kbUfgca+q
63fuUVoehodTxQiMu/VwapQkoTXQu2Z1gF2pvsCCZJsrEfPEyYOxXMeKIjyUGc3OZdcd18FY9vhT
uDXglOwVkvkBiJepVEit01rB+bGE4cwHCkhjYKpjatUL087kA9DsO1e/UHHEqxASRAl9704pJBcn
Cz138Rlr+yuEVXUcX6Hhqdm+XAn9LXsP1/eIO0ZjgYodxaGcNDkncao1LxirqJ4Sur7Pc3/CmGuP
eoXg4/D7bUiNb1vx76rhIVkISv/XeAT6Roj7Z6RLp/5Mu+pyCiHnxHjFGOOchr/hSaz7db8dLN0p
gi0Xvww4M0V/mgC+L1I9D8JJiTpVhIsdpJZTK7O9AGEtE7apegwPOT7N8wUJL7Nll1ycvWEKiekM
VNnDzfRhodDMFPTa4alm7hfhBJS2N8iEPjnyrO9hqn209F0dueO+BB0BnTwKROxAtOZ6tNw3sGch
QHXQtlvWZ35pvhja51yF16BwEq7rzDSXA2Y1rXZtYDVyyoMnug781dpFIMqxERSIJt0ItbFw5AI5
eaD45oA247r0rrhZ3nw2UDQ7fFGKSDVCPl93xpWUS9JsAgB2AGX9KvXb9Rx8sWYgrULwqgVViD7M
4scGyV/jL5mKA1h1klJmEF8TTl1HrOGTfe19KxuZvxV2ZF7vLdYjeOsBOfXbJbiaKGGMcs/1C5XN
xFZcZsgrDMWI77gljIe0nJGGNEHZeV8yyenh9tHs7fP3UgKyFqkd6UrmJpcC66czGw635eAEkJOd
eggXGtBv1VvM46Jdz0Q75fkbaQ4DSOif2weWCeFUBSdLCCvNs7RvNN8hI8e0LJOhS6r6ncrrA8ml
GSnJZMmX4xjUvyHNuudXDrLYIxEXUwS65e257Ycbuq+QgauBBOkPstSdMRjRyNem9TpfekPp+oeF
DOkI/whNXs/ixJJq45fjNk/IK0lOLWIw0a6+l/Ojex0SuuUpSgr9krhBiWVU21QfkhjNelbcbXUx
WuZAVZPU2XLF+4crkq7wR1FhdOwGAxlU1tR9ChKLTkY2aOIpfk1g3fks4aUyUV2x6EhmxvX7qNME
9lQMVES7zZGUNuo2ChZXl5VT+uUS93XK0n1AU7fjl0c2RRLcclx3wSgAa5fTY/OVusiHoAlvVGKY
WUlxA2qlmtnDYZu8jyTUIOI9yQuS2LmXEoHFvjKkKd4yXwdWZxRZf27NY2jZLe0Fh3kLIoczQOT6
3h4ZtKLLsAk7fKWSwhRVkpvkt4wycqDxsozPx0i065DyzKnMhNAQ0dpVuU7DBCjJrTLdh6Q8EN+8
NJibMT0DV2inBzIhTIB1FXv3LJe6tepMogsQFnTG5WoN+mNIbuy9NYbMwnPZkJec8ngrZL19KydT
dxCK9kc87Dri+cMIaaDdIuB5MPGPSTzvQtRaYbA1h/RqFRq2TsfQXGbI0/q/4CEK94LS9sMXvFbP
dD68ay2G+OZ8QMlXnxGdCr2Zwq1WBaTD6qMvMtn2jAfQpIcfUtwHcgp2GBOtfd7F+Py3klohSDAH
NzaYxTNQnznrkyo/ZGs8ll1BxHNoBphqttQAvaT4mrw/NhwwnCoydWKx+jzbNgjlo+fFVmcNfECB
fGDIM4DnuIIuuNacK4BWQ7Efp6WWWnsJgC1ht593QSdrRCdABwau66BjQdtAq2JD45xZZcrlsQSb
CC7iTeVu7RJF8M4SrCgRkxD52CR35d1Yz6gNpQX/VIhsvc/EXRDv9yqN3sPdsTianEuV75J/6Tn2
vKzsAPQYN39zlT5UVTgULpPyqcq/wYQdL+YX8UNGwKoU45Ys4ZfJjBwAuPnkyR/M30YZ3xRsT3KE
k7TcMCwW2LUK6oarHTr/dzyYwMFGcyBs5WNwLGM88tsD59Hw6T2K/1oKyuhWnLdGcxP63V6gZFhs
5xXxrNSac0ey0VFjn5rufrWR7ucYtqwSKYDXHJKCEKDDBD4VYqV+oV/zDvNp1G3kkp2O9jZFXOde
ChSH5DJ4+cewu+HX0pJpoxi+K2noURrLJYf53YDP0Et9JdrEZrHMQ7JpBx/94CVaWGjXF5WpR7Yr
VhPZhfjhug8fRuLDnAFv9snXpSdOuoBy/JhkWJDYNETeXouK38vwhJpllrs50XL4GVM28cGrLWmO
54FaD5obr0UgJZ54NNzoOp/4jOOqDJiLxU4r2teaBYd8Ku8PKE4EzW5MvtD3DXr63Qczcgp1zEfi
tyHUd08IjkAkCvBBdmWa0j99GyMIcoZYnNZBBIhaIQLkgp563+ZntGkv00FY9hs03IdGihCxqph9
SQAbeX8u+bYtmawZGVFMrnqOCITaN0p521P5zGuaryBK0djP1b+QGFteGR/dXGFGqmDZYm+Q+Ava
256Pm509a3fxWaNmRCVDt7d8hKXkxGsRETSQ7fO5RuhK8LKgbOvkWTOYsgI5vFQnk3Ybl2kpcWyV
Pt3tgQinuYRSamKZV8Ms3QXgFhInVvVnFCN+MkP95/zbQqi4Y37pa07FsPe4VoSqTsTzNcKWWxYx
J25j8mGs321JWCPifsX8rD0h7ETdiqLzVKJLpKaTUqXndX7SHOmNzTvt1RU6JJ6e9Q6NBfzCAoz5
TtvDiejqhZkWQL6uOITBjoitnUu0xbwneDIjOR5u1kXEEKqqsMgIk/UoSr1wPPdKUA7TnsBtQ8Gj
uNHLrb/eTYcOKvWvFZSO61rW1v43zrk+bOSinPXvQQ4idd2Ghz5PkqiCsLsNMLSsFNvkR45ghlkw
sjF7G+yA52Nz3HJpjwfPUEBOYr3hBiJ/FcKrCOayjRx5PYUqYnJ6l7cu1T6m6UKVJKVCXAIdEO+E
hiwwxrDjZb3DPq28KcsY4pj+0FPx5A0yPU+8onqFdyCIcWScJxHEZc+3dZLs3/Jn+GZTGV6X4Lru
dpNxwpwM7pzqzL+jqopwiaMToBWbIGuYrMY8v7Vt3lj1FpQwSqAGSNuCIgKZqCo30ppNzOGob0KM
Fq9YkeaUtkhBy85hSuXc59UXqL7vrvLRHfAqTFFGX+f6/bBXCSd/oKudEtj9nLFwaVFTqhsaM+3L
yzVjQmz1IKEIPvTUSyN2gWjbRZmqKkkZ/rSy8s0AArhebF577eYRZ2o4Sy3bwr68VTjEtlo+JbGf
APfUnMuT3fYTwSeyzwXBOP49sVgR9YfJCcbFQBQvnLqZbOdwJZzz8iXVXjgcJHToqIhiCT4hqsLk
tdl8HcqYls2r96KBO1U1uc0TOa6SBiAr2Mtrj0mG6noLltPGNYhH+Fui+ORNngFCp862PoVy0SlO
jY27V2NQ8MTvIDFEvF5yr3uq6KzrBMRzQOL6FAUUKZ6j+Sy00EiU8yQ2BHYcl+4s/j/B2ZgxPT8A
txZZP73EAxHunpeyUX/JEFSophk8I/1FPMf+QFabxiRh/VsiQKytOdhuE85wcm4efUjvcrirsF42
93Hoa4kAw0/nOx9GEtfQBWOjKB1Cc3pMVoBylYWwMrU9Ow1S2IU+KZPQ608VpQUyA4ZZQQa0DvrG
Xek5NVLwH8KFSP7ZSR23qIdfLqZmebHCOQA9/pkD1YbWjTVqZWN+MzjEqNtQRw+cR308FJkBRk59
fedM2JoBdZOAIzKl2ynecE/RH5GmGbtYfRAvrVVKuo0fareQSOBZDsU2vlRgjszxc1kbZReZiEeT
PyRy9YxYyZqQBcCm14NAgEAK0BVXyxU6IXr7Pb53ea82tS18k7cU5XwKDuXHWY0vTIqbFG+fxwPu
2EjpMK4hCmkh864mfaHlvUsxeyAdmpJGnlbG1OX7+Izb/U7KP34VBM+XhmQMuT7/aT9L+QpGfplc
d57rz6PrSo8tUZn50rMpb1Qf+bjSrJut3CNrxn+e4esUyWudgUTEySxQsUj56FDbdQvqU5cT9SkY
ln9HMKyO2/aBqJ9dC4/CCsyTE63yBzNb6jfnw2gNfy6v5OvGWA0YsUD8GO2EdT6qOuyZ3FLNAZ4B
AzdOpofvhW211cNaGyBm0Qo4fFgUs9KoZPT3tffPnztqI4mN6/NgPda9/QLDy7W88bG+7AaitKlZ
Cbh7WnMkjBhtnx/kYiJiRSO9jxCDQNzXpnndO3sK09jqWuTK8ACnNL0xWzD2xE+L1vYURQkoRUhP
QQTiJMBxlYAZTHxkU0jnQZHXTH3gSWlr1J9UPvi1IebZOnpxikGaYuUDYrhOobR069FehXP3vJaJ
kY5pEc99OiK7C9wUgBR/dowK7cafesb2yuoPAkrSR0tuzRCz86GLnd/rhQAmcibCLUJJX7zWxgcL
J80SMoJlhtbPu2qvBvorGMJMkcItVdyyim/K5OtnLYvzMigdVSUwp6m1dsTWgSVSL0zSldmRQKPR
zPllBjhHWrXg5gkAbDHDbY1mqgiJtyQ/sAjVXhukB7PDj0oDRX+fOjeoWphNT5zUzgYPMAwQF0Lb
asfPjkkkTVGpT5nGQ1pmT5dhSZOAdeD9fMFq600oXaVyNdgfJ+kSEbtlY9UmQGNVL8BNHECpkWyK
ARM8TjaZ9IqbBcz37Ysr/Cb2JtlUi0NcmX+1cbGd88QQb6WAxTuOVtrg+C1HM7ObcH8lFdPAthnC
DdRgt3q6BdyP2ymDceUSy3GS5pwnFQiCnvK6u5xwDwmxNAQ1Q8zFXzDmlbzSGY0/kDDpfXqDWzDO
gOg4+QnxPEsSa3nBLO5Q6ofI5IOAS0rWS7ai+j1YRAyzbelblltqlcTN2zF3T55myo009JiFXFmV
0cv7f8ddayZZwZzt5J4u7YvtMlbAUnoNW6z2OwEe96wSjh9TcUPorQ/SMfMgtAGwr4jS6hDBcXft
IRtNVSMSDkCIZ6URyk71zMqexPe3utoAw04T+DLAuyUcLXDttc6/8aKDcysOvBcMyT694T3YYnAt
VsOz4cT6FHLsmQVZsuvzeEyHdi6bOYfoMLuupgIulmcanwYb1MAyILGrnl5ztj2Vi56xtMUzhjUE
uHfYFluJFf/7kAML01bLIMsfM7zGABPrdCSl74x3MJ4E6RV11AMaLxK1A8/xWoqBHlbun6tNElX8
ZmdWN88v99Lv7FoXcrqI7YKbitQkj8qtvqeTu8ioF1fT0flSt6GhxaO0+WzdSvPSJz4WxdAwHRkV
edRCp4mndU8QGT2qG7Z+0qmRQKFyzlkmbUzQbF/KQzvz00xW64UAgmXDikwLgrh/yARwBPQKX0Wx
Oc+FowZ2oKjxtJj0UKMND4EAEXSueQHo7cYubnwyZGvYRJXYpEwfxKxtJ7oJpO4xVVzVBhfi+K9U
4yav62aEcodDM8cyNpCZn+Vlf79idhq9NXTw5Pm89bMwrqyUqA2a20Fl0EUz+aWnbAj3EyomnmDF
slmBM9JB31D9jIoGtyYQlkU5KjpLdKVO1bLfTv75YlMkm6RR4iP91jZoeR4eXkgoENNFRT8rifVK
IBTJcC7ZiVRym0+mSvVSB3DsZ95lwY8MKI2WBSWj9CeDnesw8CXiyqxrv2F43AKZ4KlSOuxDJUOF
y73b5gKMIqY7caV3VlgXFxFh7hLteRUz+kbRBQbMfmyHZd5YW4lliysuMItCbLUEjSOCVy3G6VDY
3tlLF2Ez2WhS51Rri5jM3sS1Nav4fwVvfFRydMfux2C3yOELk1T+Cc9uLFu2eev0AqXarDFAFU5W
/x4wdE5LPQJUAqjngUfOc5sJc6iuAmfrL/AzQ0p5/kGb1YXeUBfN3hi/tUl4EcyKCqg3kh4z/z4w
Ots2MbEy87aVfl2WbvXLujhhsDm5PW7hxqs7kChON/scwPY7+k2j6dO2QL1b7kThkNAY+CQVr2rD
wl3s/Vhsq4apbPMI5qp75SnrN+vkmkvNvdoblW2vMmPe4dmHLQZRDzwR0NEHNkSkM45dHxyeXeI9
NnXPmO3e0EyPx+3IFbe943Uhaw9SU5Oh2DLaJsI3GbBUyZRjc4kjkG8jbTPm2shlMkIzIvWF2CDp
5+hdPXv+NEqwSB0Ofu2pTJy+86x4+BZ524JmgNTw+JZVW0/q9UXa8naRVOlqxxqAAt1OSDDu/n51
bPp9J4TDIppcptnh0tiS2jBVTT0bQ1RsKfQmRx0m3+tm9P4iW6z8S+os9SulpT9zF7SWB5Wc1RLK
SAFz8Sn+AzUsdNUlQY8tJ/arWmH427+MztbffbDvLNtbU1SYmRQEityS1+O/CffTZXZCr5aFmc8E
myo+owAbW1kxb2EedcxazQo8ErHmbMomcLXNXQbyG96Q3UpLGi5ZEx2ouLFKef1gB4PW9TuV72VD
QIEKfPc0Z9fntsuW2CqU+sPpCMOQNLG14lg1gJHrT14CSKR2SMRdB3Gpqrcs0pNkJhaxrBBhGmxR
gd86zfmErDe0XcLnAVPm60Li40gkWp6mozRSmAaLB9JirHm5qKPiky3YR5AOzN70ipND+cnaL/IQ
RP2UwQuhDxBrO/1KfCLuPE57rNeJ91bFOoD61j+QNgKXpQLDNk9OmVP/47IeUeuHqLjWZEw77VVb
TqjnLHj1cowBh9W+Ykjs//CCO2BuDiTbAb8ySJ47hj0HA5gYTkvua36lugdwQirA3QcuaPvJYxky
JOF7HM0stDblK2AQcY7NF6Zk+Hhpf71TluGo7N/5ruJhRTLZ9FsOK7+i94yDDxf2LwqRaNEo2C1y
0lQhSHI9P1EH709whmREw3NyWgynpHJ3MKvpcq3iuiEqUlMRfshLjeUm5JNoq4Qf+k8R6eFwurPb
S3r/Cwac53OEu5Jtr32fIX6ydLf8T1VQG50etvg65quPDsrl553lWTkRNz0fS3Mr2gRCyIG5Drod
+5HKkhEv+/nwjXxJ1VsmwLplPb+Id58UVvtJcMzTrLKNPGLbjwPGsYg45Yx5MKlCujHDBuMz7ziM
xTZBq+76vQbJ81t6bqfHOOtkCfuH5MsCbSxIgs6H+/NReFqJfj99HA9bwwf2Nhjfvpdh6TuM7Z7s
oFL6CpYl6tQYWsgVImn+vcJJ/ziX6Ez5dgIzSZC2OeNpJVRPcjml7BpmKCmC/RhpG40ca+KL87vv
zHFlvxwWnfqYUpoPLQ2oroMedWAMBC3lk3+qmh9dVJZ6SipAtB/MlYmi3HRGTAV5RGSRqa2Qb1OY
cML9mwmrtb/Ya0HeEx8RIyktEakNDZ8crlng00o79GP6rQg0TD0OGgbjOitRJt7PObFqmOWh9NJP
Fj8ccr5YKE38h8c6KLRGuEPn3mwfFdYmGU5vCt4/CBIZWW2FnFmTv6eiGAMtGaZVxbXC4RaUcMiu
r4/GRuB5Tmwe77m+F3BWrIT4IG85kVf+JTq0yk7xzkQvv1djIxdta3GqpW6qsONDKiqP5eTHvXtt
vu/9ynUrAoPlhhYlmwgK1zzCrzXKQamJ6R+wkMAh9eEV3IDeUCJx4PEJkHoiHndAOQW1YafXVURN
31a7p6+y1ar+BhFNzMmfi3l5rN8+sepV14MrC72Q8uOJL7uW2Rc4bISgBfVQVZtWf4ft0S8c7857
iiGsKjHVDjlYDH5gQwzHPZGK534YrnuwpW9TT37GkRUD64Bjrdr8pXSJeZpC8SankrM4cZdU7MkX
fRXF5KPGwhThC7j6VSc4RM2JtO/D4mJJtncFdbk+8mkSf0fSpvkMalMAOwil4wiQzfTBWZ1Ei4ea
0Bx1Fe1QYiVSHmaX5PQpOAx6tv+1ev5mZhacECB0BQ64FrH+hQr+UGjOsclChPAfG2nHkBWPsnYk
wCN3ul/8JIW/9bcGiWRsklCAwTB77adgn1wEe+LgHzr+V/oPdvYO6uptytEeWy7xCVJp3MmGnjZz
WiTQutzKcENSSaU/5X5FzrYDkGSjTKGADO+nTcv7m1JSkNxSdXOxNKgb7urkKHoN1b+1P7RMDMbY
Tw2qB6gnJXemB5ehjq+dehJvXiakagnteUlWi2/+T+5wJ7yah15DjENUTjB/24UkHyhjy1nYrFRP
9khZ13rxmX4Z5yuzziUXqhOBoHxhLhE6glgDOFRwxofRxBDqduYYeYewU48wOZWn7oFMwYjUzSg6
nTfqpXzcgNfevZnM5QVX866S+eBk+qjZEdWK6wut80WTxNWPHOmjdCdyRDdWpbDfqIYyWF9YLrBk
V9091TlcTQ9nzb8lTsEodczyc9C8OSTGjU3JnQ/U4wEVwtKqnTCH7CcU1sGx6BrnSeMpr7bxQoUh
pvaNZDCsS10wMNu/wD2fNhdjsojG4VYrPOlb34XSNZiZrAzcAYXSGuiIQZnb7Tk+X0JsSsFFmdBC
d23LLNU9sqxpie4WXYDrgZR7w0jzAkjna6wNTuohkvG5FeqLhRAipyv0QUgDJ0laaR0J8Y8Hn6on
AmBlECid7puVoOubctaCkJUMISuGc31YV2Oy/7TAUDE3W0UDwHe6sRTqoAyCj5Gc1pwSAnlLGCgU
h82myh2iVWNSa3egu2nCB6kHVPtf1KziP4gZhklgR6xKMQ2CDSkUzBYrX1GybI0+ZurlQjoBS48H
O/ys9Qu8ZkEiICZoZlPlWx3C2B5W+qoRXtlGPkbJTtZmlBqahyBssy5FvHDzfShtUKxsm4AETzV3
ccYBjQM0YxyaYAJM19vOQ4RYWZGyZv4ImzJSBwG21sCjjTGnDrpiJP58ew77YLZ3H5BDssVjeuu7
mcvJdS6Hj+i71KXscNC6P2QXK5xYcqc99SQ4C8m+77wm0P2C9iglzi7oFcC+7Go0b39Yi24AFztN
ebuKmK3q3/X8JnFjcRuGXeNJr0PebIgXqvUdpJ1r7JB8Puf+WsFMNkh3RJTT2GdXTYGFh4whP86x
RtCwYWzPLLISN+O2+uJEtz0HIaqjfKTgHwFe55R3AhdswSz5QM6JjlBqq3oHzc6US0bwjXg7T+Fi
5o+sMHUmXcfRZEHEgn52qeSvSw0lf5cXhnSRCvie4O0ldBWn5utAg/X8ltkbXbpHmuMxxgLNRrlV
qNlqZB5EFmjk6rCSI41/DxC7AcM43dCCcdYIt70dixkMyLMxFx11iRZ97eTqStzDJxTqlmt7qrEe
omG7kizOrxfunpr44RpPoV7HI9NOfZbnWQ6CrMQKyQfKtNLUiwTUmA5UFoiaDxQnylEQHRUY+Bdm
u46pgR5ouTpaUUIMXSPuEpySqVwRKQCjt5OZO4MhqcZHAPQzT7WAgXMsIqPxS1S8yie0wv/YDT1w
VVFB/egNIUkQQHWN05hlyrfYk0qsGxOuzWzoSfhDwKoPip6pCOV6Eza+txsSnmpsAIAhJeylgxtY
hlya5K+aClPPOnvR+zsNvka+tzfeNxttTiN7DQBMumpZ+ghcuOgVegs2r2L9sB/H1iUvMbQumsP9
6XQVw+GkppBQ63vw0psAUSu6oiqkoY6VkoxdSSexS0S02u4FvG2LPSO8KURqsV2SharMf88mKg4G
C7Lw5jBnP8+Y+Ux44gjDsiaBl4iMJcgba8HHlMmDCdHOA1aKtqRYV69UDg+wMUeOP2XTwfSRhafW
f/6h/akHMeDLSI4HL2DfKwR5k7rRlKoIc2GKQwxTEtuFqi7uYa+EGv7MZRPEY3pFGXlqnSMC9oyT
1L5BkOa2Im5Na6w29dPZ/9iyJeOOqc7Hj73lt4iHhqciF+96WdbKeiNAVWs4uSD2PGa5Mmq/Y1HH
kZPnyzFx1mk2aYp3bsBSBGUhTcdAIYI5rGfxflyN9XeDd/2P9NR8fjprFY4HpmWT+t8ZKne9g1RJ
jFcCwdDVB6j7oMT1q+gM5mIByPBMMEwUuz5Js5u7IpNhUX4Mi6+rzHYfTkRIkx0NhLhY/U+RN+N/
KqgU1Z6c6Ysn14i+NWsTjfokCXUV5bLdjmhfq51kxQ5OAMlC2LYwTysiu+fohzkPHW41c2P4oT9D
gjx8Vsm5No9mWrpMt2zSmVMWx5wWP7oXUWK92T/1WUfBWTNhgJQmuyCE/Xo7w5J90lOYrqKA8wQl
gAq15m0FSFTwgZXIbeJVE/XzdCf5dsCZllshI0IuWut7LqDDPgZ7oM19Mo+ZGZMvwNj20TCmFufX
cTil3YXoBeF13GOCm1iTLWb96ecyNn7ZlwZKUOJTtSLdIwA7BpsYApptYgJ4rSJ04P1YAvkeZ9i8
UJMMNIecuzri5UxkSNnG/UqpMSB3rH7o8EsWUhIutUzR/S9qWVOwJiw7nRTmSO5Pa8ARevUv2F+V
Ztomrnxn9pXXHnX7u3sU7hixR1WgIaDyoBcxqaoAgLhFLBfTRoWV1XZlLQQN4IfMG1vu4p4lPWgo
DH/WLXrm8NZLjZvR70EmAcoY58L3hc8ySHYPupYzkK6AKZc5ONN7k2bIzDiXXLI4Kksr+oupS7NY
5l5kbwkBoKCXf+kn8QkwEN2xZJ+VMnj2t48vdOHlI6MjXzbU1xN2JlHlBCRZKVH/Zn2gPDm6Beay
1zodmUn6wKynIJ0V75L6IzchIrwm/yXpPwRV91FWG7b2gq/5yr08Ucwt+HCgAEzfebuQl5JHuj4e
CBbM01t5ONVLxZS/9vK1419YFXu7B6YKxPd+JmEPIZO/H3cfOZP4mkTWKu/rmXZ4C4a2183Bvjz4
iygrplrXREAuImI033VqJJIH4dUbaUxKT3di41XMKH0JdL8C0onaKBXv26ljAlwqHVDikrjzuGdc
Pen6Bvm40XvMl+2OhJ7GtFH5Y8Bggft2HxavNoiXktKOXRfLq5f89ityADtICB4e9Iyv9m+A0INU
ZNsfzdglFG6E/UfcRnciJWXMVCUOtX+yX3FJOFRBDW7Dvno9e/6EficfxZ4fy11mIo5J67GS3bjt
7l3DR6CdXLCr5CYpECv+tYRI5iZw8mvIXXFrU3NtdfTouJyllpqKRbhJaBOOTnXG2NUtHcScYPZi
PQn1NfFaWHZlM83psyeHxXSFanbbv8aXeuREGWe3X1urGvHNNF/G8CgZw7WaVOVTNNgKz9y2139h
s8mLnhR2Czw7TN6XUVOuKiR8/BmyIwbIRYVkta1H9K4ZHTSlMtWmCxbJvC9Eaf6k9gh2QfiEZqCd
humobxDLv+CMtgEmFKrPIP+rVeMthMJXtRozGX3FMbX2XMTh9n4Po4yvNFlCAAthiCGvymwK5xOI
UrifSryTdO8RoerH35sMRTTGtdT07N4Afe6Sh5DucDTeoVD7sIi1mu5v1S7ypia2DQzwDReC3fSy
8Uz5JmyaHx4vHm7XPfkO+35akwfHDGR+tm3bkTGUJjVZ791CCVcQWiwP9SjeQZKx/h2KyzvdkIVe
jTHjrhBCqwAPnxuopgX2omNfFP0iADpTN/g5H8JaKKm5Zh7VPJMKtpzANko9ZqKmjRsekfMb4hpv
aExPm1qC3e/Z9amq/HKK98If553KOe19XvCqyC/jvPCIPO7v2toC4beK1uoTd1x13OyR4ItdFCVj
DDkzc64iD+jm+CvJpxHsIJNEabdYNCP0UEN7SqWcny6u1Z2ikRhl6PynbbyIDSy9tlUB0rFwqwdu
Z5SRsnBv9OUD7yfA6qQsXOwtvJgava7+JvIajAqlRJTqt6Odv/XMAwJhuU5/SjoswcK7BJxMN1qk
sWsKV/P8so28cWafjwaV0jnhRWPI8iLhsVhH9lKTQa47AXcshjNCKdqJPXa7j/8AadV/b0KE5UgF
1V5vbgzARA2oUUXKBpHTjHpNUYiBgC6o6H86uiCTvQrEncbo08c6o3mwLS+YWbXIbYQSartxwjMx
CGvn6QdOWni/bhkf6d0UbJZz+7X178INKF7p5K8hQUYp9g2WOV5DxjgbecGrRFodrFQq9NgfkYPx
eMgoJFD7EuE8cbQPL4e5g2is77ENf3lKBqmT9refdpWvwHAYHOgNx2OQA5uhTDHJD4Ql+TsWdHBw
joJdlQijwu1slaVIeH7rr8mzVejf4k5g6SzCizuF1OqImTOoGplc0U+aGk6x4fvt5HHx0GluVtiV
9FxzmKpVGnkanV845BwVlPKWDFmINcMgdbpUl7dSLr4yOKEOuZO3ks9IoveJUOtL3A6LCGH4aZZC
lDhoiFoFJzv9heOV+4tLy/LsKSW/m9CieqcmNFE9rzagOmGpvvWewvZ38bT1xN1Umi4giA1CFPua
pyR/mCOtSzxfOWfdrfCb1fGA00QBBh+0IgvUPrnpGgjGSuL+Kaj75WDfp2xNlLUuzNNnrw5BN7+L
UOOs5CDkzgqBOBMz+zQDIAQ9TK4yJ0d5UnFM/ZgA/8i1rdEdQTylr+rq1iGkuu/+vV9y17hcDQgl
CNE/y/s5z/bt27EPoX6UKxS6zy08TUvxev/aaYl4ZNyhsyP0SwTDr9GZLPUYimSzu9uNQUVlRhlF
uDC/X62pbxiqbxdupqC+MABsROI3/blM7nc50pamA88/Iq9KGGteY6pHH9PuoQO0f+pEn+VyazmR
goEWyb0W5keo8aSQ42xpy4j53GkMTAVgPvGCN2XBbTAt7o/ywoaQWKwlADTQGPywwsOmnqP1OJv3
BHvS3gfXdh5T2dSC7iqRV3E6xC10yua7O3ubMYVgx0K/7Dc1CBbB56E59W/xektfx9k95uLiUUTm
QE6v72m78YgLcs89iDtq2W6+pAG+OMoI1sbunrbeOVMmHOu+SsejQWyDb9izDKn3fxBCYwTemkdq
bkPRjdbaNHHS58Pc2lGXb23Pgezn/kSzPp3Zv6GkbETY3EGIHIftrLPr7GjCtJlxF9o15wP2L9JG
biJ/aKcsIkTUcDvQnAVNs/xxjUsdesi/5G/ana7WxdWfeXTNYAmuVm7CAgM78ccGyfyy5JuT9WPr
lbmv3Gz1zwBjIbdfaU0iLJMVfupLYgvooF22bIZ5o4T+ZQZFiD7kLWoh4PoNPRDufyQuhj3KGnty
Aoi6fkfctMvVHsEcvEwW8jpcFYLXHSYEkjCfr0PYx5g/YUk1bS+nkgdSRUhn5XInhU0wm+2QyWT4
8tzp+Vqi4qAqhU6MllJxoG/xkkI6u0hTWM7C3h4w/L6rVcB1LWlayEw4bCBDXAYmVwoZzneea2A9
taqmhLMk2TX8GzT5aOve0nXsTgPJtc9M95RItfmpB1uCt33Tdv5Sc/qj3L8E1g1yOSWrlvF9cadE
Z9sv0zyWw1LpBVHFfHkD0uWSZDQTnXclKq387L+XRR/Pvd9ikOfQx6Tjdo69KOBbLLBpNfUbkc0t
Vfgp0Ld6BGFxcIJOVy3SUZd9yb1MABJrOIVi6ovr88AaiUe+ZcvCCxp8/Ox2iRtbtMFdiv+sOtqf
eRAsVkzyN6Pyv7eOid/wA5ZLR4M1+pXOrBAKDbZt7Sgx8UlNFHhd2IyLQym3e0I1ZNaZ/fkZ4Oa0
8QSiaB4P+j8yq+bHiZ6vV+dh55y9O8d3r31uFUvNNCXH7FXjI57V8PzyC2MhbDcjdp+yyi5vIK9X
wNLl+uk67fuWkaxI8OgohX26DmrgMsLkBeEf5vrA1Q27RcxDA4KXRSO9kvscIPDrbIoHEf2LKyrc
p1IJGQ8MAlsCZeMncBflY0ahHBaF4etEtG0oBGEiMD0Px28pHeMAgdL/bnhnZAQsX7ERqVBm49tn
+tsgljLtynLwAnsmIuj1dVqD8vhCOIQOeMnXwSM/6DOjlEFhAWVuqM9KgezGbmf8uicSkISfImzZ
/PoGRLvrIN3ZR0QkgnS1RCY+IdHSV0KzBjGYxZ/urPXEedBmBGY+waqc5kj89Ki6yFONKXm+5Dbz
newinl7/fFROJ8DFWIzQvm3XWvDA2nBMX5SXPHSgvf4rSGTof0OppZblWy/Ip33BLDok278fc3NH
H1E9lQKqPfMmluA+Eiem+kAnPbrftIGr1lc+dkIfp1lgfb4iBrbegnjjA/iAARjBYRWQM1QsfB/m
2AZOmk495E7NTwn3GeVHxXaV+SzIEl9w/wqcP6YmodqmF9XhiiI32fFxLU0NbZdMzum8qIG58TUa
GXm4hEOVR+kQG07h0XkCE9H7X+g/lLyWuVXx2QsvbkLBDFFGnvMimoz69kGbIPWzxOWJ2SHeOMam
Uzs7E/0b6chVZd6Wiqm4RxQbLOqEGrZE6AHzqksNtvDbBWrQrHo8Cy9RIoFPsIhzm3iVRycRhbDv
hXmfnY2mzuN5HfFo6M0AXARJKEgy+/EGE35TsMO3i4xgyuNMZPgFFcVz3+pmoA4Kdaqz2St/pCOx
fPimFUGHop9gbbx5XG0U2gW4cdhce8ajuIZvbh/Oeyz/DTCaue9ux9GEpJY9NhYotILk/+1SBGeM
z248IyANiyRD14vc/7QzkLB1+p4qYIFhiga9kZDntRZ/rVnfe4buKKjjRDBMTHOnwr9GmhYZMRKY
7FirbxCgO81FBZvQWDKB1JJljGL7fy5RYk7jLEhqv2b9cHu5GO83ql/o0+2ueKmj7CnRlsJXpEJU
6XCjdX8SJdS9+d6ZYL0asTchVj763phixLXeDAn7ZwbFg4frJmYwIiWyRWNwqXWrVin2LYOx4zC8
Vj0DPr8sfBj5p9p8xDrpT2TEhbKgpMHihtu9lgEwGdPHs0XdLMfn0NWy2BJGujGfZwtqvprEOznR
f6Bt5gEKbe7oYFK/pxC89ofvj1DUq7/yVM2KEgGu7FjJnJCoBF+NZFcOiH7lVglIRQNfDfVDOWDI
bxXyWtJgTH81TlrNYq0IFb05PfErSczr1q2xOfW2vrjWD66NdLnFT1QGVZAkOSKVKI4TpqfKdt08
cQLcVDhx1mqQg64LAqNsxb3Xvk8mK5f/Q+crrj8PoT70JKzOvR+TVU/rjZdZ/ET/I931K3lnB18W
qweMrnHHIQknEOPDOynnxkbDIkPkzNHHSFdBuJRNNwPP3dun3LuI5sDjx1xoTpx4YvcexzL/58pX
03mm54WJPrt/85qTMCael863lh7OYTXjXALmNXdKnAdQuZaOSP1MuiTq2/Z7ufBd24ifUuD0DsTk
qMponVpnmIl6L7ZUMg9LvokwSqpjhL/kSzlwTyZsrHg5fg2nzWCMKSHCjDDT1nUXl90rH7eZn0tg
XgE+RF7I85iFCdwSIgtGcvIMDscOfXh4PzGlCkILjWo2KcPME63u88j3AX/7QIqZrc/e6VJHr/e9
2IlKiYdzYAZqE3bykhUEWgpjvDD12uwyhiiX7gzGjQzHk/HVKSRZvGcGHJnDTQ7UAEsQzg2x+mZm
okHA0w6H69lqakowpYEza1aMXdJazHk3ukwxs8ZCX76O8EDatvfL7hxMl95TMOoLeewi97q1Wnwy
6f0nq/NYW9BP+PR7B0dkPqupRHjh9apO8hg8IUMt5649G7elpMxhGpJEAv00BDHOURRLgkUZY+19
N68fmHR0ffumlIDk8Op/JBtWFWphJe2H7wekn8qtW+7AUAN1rBRSGKt7FXaF4oq6ojmVNclYwZYE
zRF48ZPqH7c+W7vUF/gTpRkSuNNtOucZKiPBpa6BijAFrlFYQxN8ALvDeTm0sqo7AXAgLSV573GA
dzJAMbdX4iWoHCAwuXEpeHeGvcUXFOjC/umItiVIG/wXOat09gF9Cn7bqR7lSvIi00gszY7669pW
XYjzo2Cpxa80Al42tPN5JhNBb2gwPP7PYOcbgXbVebN9a23JKZZpnKWSCb6bXSlN5JPULQiXxHED
a51Y2LmisSOD4HnJCOJ7dTdA7AewY5TuLsP7tB35qihp1Udeao/yYgqpj93cWPC1riv5Whlx/gdc
7DAp3kBnABSd3qtrxM9z8LPnmAn6G7rTPWvHakotVgNQitLLqMY8y3IAfLyROeqD03i4aiIow+1N
1VfqFPWelS4xZe5jKocll+Asuk2GHbX+ZOoya7Z1JJObEcFqV7QBjp9ugI8kto8ogRFlpp2p/O9E
ahimbfnktNHZ50Gpv+pwhR0yovTfoebo7RLbbVsg+PJE1zfzEnEKKMAX5HsRT8QN5c78Z6YWsvQY
7D4aHfzCyzDn7J/wYCL66PEgBbAHX3QXaCtEdwmqdwzYpUNw5sYY+6BX8zVQ8eU5Re4F/j8bG3HE
w8wKJPCB+bE3M90M16rVUH122eu757bIDNtxTVIEUOAVSZ+IdcQEPqEVM3LdoXzh4syL3I2RayRL
PxsGTeuP8K/OxmetA0gII6SSdiI+3YgpAPxrdmRGtAPthETJs3g5oUPeHUemgoW3w+1sUYzPoS9T
E4/c2si73TYATohRTl28Q4R9VU08/x9znI9eFnW0f8xGp48mYuESxq72u7mRlInxfrF9Gfx0aATJ
D66Pxx8p0PIlsaPdyoluIPdyy1M3bs7ZQn9sop0+YX+IJw+lZqOgRCgftBZa0fbgmJTUyFjDAQZ/
5Y0mBdBrYcq1G1BenruwPWqDswQneafy2IHyVJ/f1xnwxEV2TuENKN2Vhc7MFGDCi4K5EIvJ3RgE
opPSNNra2IloGlsC850SYlbF2NfClRJJnkC6wmrQBS2H7w2UdgskjDEef7giMSYmBmeiSvtQcOmA
UYEOwcWOLodl7wbtszAV4nIXOtBLnWF0tpnFEejYGYvxZozosxgXFj+a4eBzmXo89Iwv2jsWas7r
KG9jM7Zp6B5NFB9inF7biL2O+TKUJTpGjXT3maCLKHlaQFuBc6x0n9rl4aycNX8nSkYpLRPf4ga0
p4u5UdleTCsU+mmr63kHLYfK1LSUb/cuIrC58Dll7LrQC7qmLNHeXfqIaMOJG+QdIX/RjLWY4oda
2snJWpqFzwLWRvkaucAxBvEzXfojnienbnsPRxXn+KGb64uJkDEjdNyBHo0Hk2RSubdslhnzDvKy
9tPgam7eVD7ckWcuy60Pg3htToDc1+28xECDOSPGgFx3ENhfty8ulJELoU7zl1Oq8VOH2g/B/lpV
bZAvKHpnE/1kPQxh/t6F8fjfRWDI0689mtm4BfhVfT2/N3tuudFoTlFNfzvU1ysIbqvaHSHzNaab
tM5FE8KmfR3H2K+b1k49zU5vliSZcXUq60ZG13uuOyRuebEW/7PPNqJSLLEq9qENGAoI5oP+6njX
UOc4sdRNHeafADM5a7am9TsghwzrlhQNmtymHt/J3qQenR6VLDR5Jcw0dk+TpoIYVqnFd3qCKC16
dX4pYLeDJIGSJdi178WRdC+QGYAXDJaNp7i5Yq8IIyTKrVMzBtq2oW508rY/ofwjSWVsz18jU267
UnMOlH+PPV+0uZ6yOan0bpFjd+mb8S6bfrzHRjQOdUyBogA9T7I6QLJ3Z/jpJaghHj3vRiS0qHON
qNfVlYSDFHoV/1dl3GQJpiAjcLGQ4kABJxQwAe5YD+Q2LEAcx3NT/nz/k3OJJdv336vwxzbLvKEQ
ECXtwhswW6PE7CXTtbB82hMlqtP8bdzK9br/KDRkPNBrmKHm7G690+6gv2pSvBS3kM6lx0O2/70s
qjlfG9O02uU+HAzQ5sYSpCaXUtJkbGdyrPQHRqsbr8bUSrkaiwevNF4ISmHV/Qjce9I4RNcgPKhF
x60lgZIkk3ELHPgGDyZ9ARnIGAMhoZk92uNevhKjnxnFIZkedQkeo8a71kmgfRqPxRzU8qLR4/o9
scJXcot4sEUPnAgxrLhK5A/hipRryKca0L6xnv5oVpAbvgPbCQVdJPRm92PWvDZX0twcFbTfe2ht
dMAtvQN0rTBhrq68sxxsW+OWx7fmyxuX4xmqkB8nGCE8bE0VYFPJa1uOB5OiYvHIrYvO0UgyEA7b
xn9gIqTFHhRM07x6tRzApJfBXzZR8qOJfPQYnaQ6WAcoLpuIodr9DYkTQgL3PO+vsI/gqPwlImP5
/d18yYv0lcTpEKYw5U90NiMTd7KjXSTK88w30xzbXBX0D2OtMmammrK/IyV8Hs7v0RURA56JmAhr
GLKN4bjp8XXfaO6fZw2s3fmcoL79OaF+V1LJqbsgolcyGFNUhXKo1Yl8g9WPi6b7sNB0On3rtxLK
OwpevOXQj+Nj5RH90E5xu/e7UvMRqkle/OX60gtHXgwBadjvZX3W3kjcW2hg82DUEjYTYJ4PuL99
wIMdMJ2uVO10kzUCBUFbv+o8TbUj5UPFrSY6s+L35eaznOycS3Q+oyt2+nFxWE35cBfbw4/mMVV2
PIb9lQ2Eem3eWcVtQeiKNE+erdBg4cM66BOrkECpfHuAVtayTbEHmyei/RGyug8mNoYA4nW6+saZ
NbuomZrL9fb1CD8/XJ5d2TCJubVS7NAdgI47JyZ1Fe+n15aP9SlgSPF8PuJHOLzPjn0nevr/8maH
KTGhHOHgDH1w5e8ECgkFpKifimLXqnPICae0nmhF1ukxsiBa5APySZA+m5cAt/a+1Yaz2AH7Q5EP
LsJWvO2zIe+pv9Lpt+jBXu40LSUWhyh6HGPIjmQBQ7pcfN9XkftC51tl+HJNUJHai7rhuwQ9fW9b
txxqUbS7aW4kfp+gEVy3ugNxYJi1Tqzt4/0hecE1Bd8us/YhuzYtXu179DpYOI8rV+jWXmjEOLOR
pRYrMe7CADu+RVucvAsnpnMDKeABI7w+DgaN9w8smBmxZ32IpG3Bwp8E1rUyPKJA2XoSPygMSZMB
MjoySd6FZ2eeKnU4ENVnB/Jx/UwYz54jZW9UEi0oqo3eCkco+Jxris1BT2CXxJHuaheRCaPJv1Ka
gG/S8VeFKB1TbVRjjSpQbXKieuiOZvmlmyV9J5v2o/37+29g2YRgttjXpdC0mf3SJRZjd3eCEiLT
pAaIH4uo5077copIEaX0eRtqhJm3spfd7AoZikyD5jOLdtB5/GrihHlzUOWPzmgbVdv4LMAvAsp0
6Nn0b4+SzKa3HEyqsSVz6QyMAACgzEUNxYrMT+Sk4A5jNgBYDGlXhw4n8r7H+ojJhx1m4xFOYl9E
Z8y1WWfOJnCXC4SSv3F6vU8nfCxt6oO8oUkAGPKzK6AR0ePAaH0OncfyMkD0EajGdH81oOx40sZu
R7MyN/Hj1Q1qD/Hh9zewE/kJxwXLqsTlh0tTPrDNUBi7CAE3D8ptSpx+cy6XSUlSXGVoBJmBWd2C
lH8dQJ3xwiX4EuyYPPsXwgB1V28BWx2NiQnrXFHjFKtQqTRc9x54HRgGrODNH0LZrmqQE6VvdL6I
8wi8w7wCLrGFbR5KZRYcXN260l0IAxTOkRwLNiiGkSb4Cf4IS2cyrMv1vBaeOOxVNFMk8eaiwpKV
blLn4vp2xTX2s3ys0bpfhx16gWWfGRSgbDs3Yn/AJE7DUrFVjrmVkneaHsB2v8298F2whxvrMe6M
uTsJG+CExIZd/+byuNCQ57kBAZSmETid8wZIsWV6jGHCwaDZbkMmL8DMDMwwCz6VnWSG7IsbbH67
eMI96QRWXZGjTvZuH8/U/YxU+R1MDLp7AcgiHXkkj3l5a49Y0R4kYfyl9xms84DupjR74c/Fu4OW
4ixJV9Q2e7M+2w+72mnIJDQ43qaf7vqsBKRGGTf0YgwKA/59ct36v4XMkQnDQyJCfqf6Q4CiFzKz
ObfWCMhU3Tu6IcPTi32mRcFTURawFWsndby0v7/MJaNaym9VikJ01YMvIFMppxtseFuKSYWVWwhx
lCOPQhNBvIXVBYYzcv+ybew6pz+VEyNfKGnNDFbpwCmnEnnyD5Gg4KB2SzvZjMXBt5l/hr56TgNW
WvlU5meIz/orm864aYd1IcKvFNHtTVGQVMsSFopOY86sMeK4JHUypBga8+0J65vFF4fJjtFXBgvZ
nh55WdDXnwA2xBEI2ir9qeS8nByHDHnDahfSeK9YfDHGzlaKYg7ws+0igc0/W7wqRtSJmmTFNLqd
Mce0sITLKozLtSk3juQdRKPegmvkCByYbwrnWZneJdkWBx2PCXMtHyt/sjhgX1iQ0OLvOvYvuUBa
d+Xkg1Vu0v/JLgRZ9FUuG32t2FTJyOiHdec760GuVOaT5liN0ZeZabEERHO4dbG30oPv4/027VVS
niGgb15QDQOhrNy7x4IWe7XHCS67SkPJy75W5lyQkf2Qi2BKqkdiecsGLN7zruiq9/d7X7heSVdE
S7xGcCfExtG+b3LiKjeSvHOPNsRgArhZnmBx58pRnxIL7yY9BDFpXucgwMf7qjaLuSsDnVSk8T2s
KTJg6rOUwWfvYBfkUUHYJqMsctIT7D44G99RA7IDPsmtyPHtjCGKd2AxoFD2nQvv/yKovk/qEI/q
HrDyuYq0iY43gUAhW5zWDxiWMpU/0ZFve0fWzIWsK57n4ZjttoII2K/rlCM7u7oocOqR9euX0ERG
R15xOSJeWNUMcNtdACihCk94yHyv3BKpXnGyAjE2Fjhx9uVrW5haYZcDnT5Q+rdfhc5qY/yYTYp4
uqRu7VJUxVjN8SAStjJP14fnKTdY6Hf4NALdiCWzKKrHMKxh1x4GytoijoXz+YR6Upm/YtsynEGw
vtWlGhOSiibbw8g306/zDghVoUFuk/gR86lTtXlP5WBbzK/7AA2UucUDdyLwy0AaUfMZgsYZCek1
KnKbRVUFvmF08OEvzk6gjkqJtBDkV7oVOu6GQPto3Q98SqCyXsL8TI1N3LS9nxtCt4EwN1EHpTJ+
QPP8EykaOV6HAXuOrR3beIjxb14Svi3EY22uX/w2/0nN9M3VP+lvcQymd3Nw7rYGFfWjaWHIx6pV
thbmWQlELTz09/EDKzvSGMd4ZUOHpo/MHDZvbxwkDKU4j9jsX1RACp8Nvkj04WcaZvQEWQG2RccN
5y1E5voTjY6pXW7auG8T62HDEB56KW+fJ0igzz0HNcn71NbOMUC7UJ57fe1pcW41GvC1pdWV18GF
/YWKOa5kiDO2LKDRaJwQSx+euXkp0RLf9zHUTcgYvPKYWx4MmfZSvAilX1Qeu+w0jmc8iNkPO4b1
ZtUjn5/cOjxiyy5cNDCGRR3qSrWh/Q1vwv3/89i2t6ZlDINnUCSgLR0yUSDj9F3b5Hh6QoSIOuOH
jGpfy8doQ3cMQlWW780v5gBVxRX3jVySbDymajyWZLCu3z+t3msQeJNIch6nHc10xYT5Q37TkPNq
Z5cVyeTK5qFkLWpswFS9Beie9vanKcZGBziTnj0z/S5Lb/7BItuC2mDSLQvwAsGZyhqkFQ4j9CPN
1uTh/JJQmvbM513mjTjifZozrBlglZxg3GTcL6LjUfxQN4vmtcuWLLqTQA323yCR9mgT50dGxvm2
kKp20l69ygY1a9jrZZ7H6m5IaOiddzm+mOIHAW4JamMdPUeX3pqvVmJKgM9dpEC6RQnuOvbae+M1
9Pdd0dlRYSmdJ3BBlERSnJjFBom2itVM9VJ9a9eUCL/y3KxLYl3P2OyemjyQuugq44hOPCZ3QYug
SNzWiBPoTCo2UKxEQXDZVp3y40phBPfEp+drJPgaiecfB/+FmlA5sk5YVSCGXLzyNktc5kCw5U+P
1ctvlHLKuINc8OfK3cekr5M7Ww1uf5H+OFh1IxpaCmSODhSfZPYf6VOWB/asjrCVJznXv3XAJl1H
g3JvqTFdCgpDlAvUq4gp8CkMxZld6hN/QAJVWBovRry0xSjvsanX8sEHJJSN/fQGMD5eCC7HAGka
MxHkmNNZF6aMXcdqggYyHRc4BPiPceS0jke9c7+uDWD+aacSYvY8hhypXw5BOhC2e9JAvafviJGa
RjkBr4aA5lHPu5gZQvbKcZ9BVzVkUV72dUhC6sn7xvBSUOQRI1eVfHMtiqyL/TGcqEX6lcK7oOcl
fbvsWz4CiKxuRGDp0iR3B9rNnjU2UEUKlae/PDy/aQefav3NnCBAZlIOZpQIJJej3uhwi/6RYphw
4wsfjTj8XRcH0Vt6Zz8+lbmOBa0/XdQPMZEQQh7hcPXOw0Riub9O4f8ovsvQytrwszEzMpl2kpe2
I0U7nLkTwua7fADp5G2PmxxwVZqUfPxLjXBh7IcXDKgjNpb0oxh/gEHfA+MufONq0SYJuqtSmzLH
aHwyCidruQXP1YJkzYots5t9sQQkWdcR0IOPlTSdH0Jrj+7M4Oss4ixfPfoJXiv3p1QR4495DUT1
viW28y2vZ4mlUIQnZmWmjpKBcVaJ7l1H+O3iWraB3knlN7V6m8nBJ6bza0YKQlL+JXny2kQqJSjr
k6WkE6ccgOzNXuoRlLx4LUu3S+TxPzfSoMSyM3vzkubBudCAcuZ0OlTAQqkqjZvsv5gnpA6HV7PD
usqq8IPZtVgY4p+MtKgBvYs7ad1OPNisiRFk33VnCPog71ikb/rtTvzaj0Q1tLwJ56o5kjbfG7Me
0MgX8NQw4qqCA4SNvnoVNC8qo2zJO9pPAG3BH6V4hQQp3+8t1EvLwcRVDkpkgXI4JF+YFG56Ft9m
uPQcfomluGEKzG3+vn/7Sg7IC4COCygf6xWxgxaPWelU9XaYz7RtAtZvSzr3dwpdvf9zexgQLuXf
JZ5TUCHssQnF+sr2mZApnVLkGgHVo7USXvCDA2oS7tUe2LlUz6mT0dRO4PspIKgXfm6fKdkvgDpo
C3E/gcHPKsgiujK9GZLpA2IiQRf2nCVLnsnAjKAYV/eDsQ2AVojOCtKrMZ92p+dbuXWh3u8h/sGZ
D1M+FpF7z35A3XniRcMPD12/xVErYLR3WCsirZzNuN4I71HCQhNWGiWH0AwcI/UyAxW4kuZAKljB
4sfL0FPZPcLMCYFZRajdKoSBg/edRSIDG0A3ShppvZ2ibzpgpmnrANfUzZ0XPHIJ7vONNn/jx8Mp
9yBXdSM+QzVyexBPZHWKPlcMwK0YQOv1RyRUeP8OO97JsRT9aBC1hFICvpH/zpFLZGxI+CCl0u1I
33MuXCKu/bAjbqU7YUmhpkf+2vvKoFN0HR5zKquE1qPct/X+mHaAxzl9nUwjh0NgBctXCOTshLzj
13N0sw6ksLs7VxX8mRI3cfMejm5tlB9RJLtvI9XdXCMsHX4dZVRUI2aNv+Oe/LFde7e/kAqT4Hug
STfFH9paczb0zk/jRV4kLZRpHO3gL5KTTLFBBB4VOPNvIcVT5xdli7XiM38nHOpLk73WGO7Ziuh+
t+6cXlpdk4RtvgMZpXyY5yIEECMB22oz05ExXpKoFQstkspTkNRFkmAWM750h3yKiRDKp+TStr5W
I9Sr3mLfnJSjSz6dm+EXlXVLcPQrNuH5nyTfnODUIppZO9A0tEC0UviHv1JK4kkxPyuEzZvh7nHc
GNyRXaJID2mXwGZ8r21rlSbuJn5aZ1EVO9iD02l9TtCzXSAXodfwuBMlc0+j0kKMYilz+B5AxrZ4
4iGIPyV1NoOXJ5jlSh28d+oUnNW91SEyFKpGcE6erPajuOM6WQAXsWco9o1xZ6IEXRg9lGaHkdpZ
pT7FFIPYSTgNR22lSTRjlozYUCTL9fseuPo3Fp6mxRy8CC/wP7xrOEchCfwEKpl5inCErrXmQQqo
MHVdh0IzTFVlvEntqXRl7FCi/Xwgpi5pfke8gcF/boR43B3O45V5x8KuTvqydp2AoWEbX6JbWKbg
gstiw1cfTKGAzq84k2Ev3AXEMVrE90/4vH7I7AntnJlNFsD2HI41cfrXReJVl10ssKzL68QhFcGN
E0EhTnE3NzAM4sSBqcyNZianvDQMcMGSUeDW8F+RQY01/ymEFXOgs//n9RTRKCYd/JbLTpU4MRQv
FPGvSRBT84JRx2Lg1Td9fNvPbwxyVbHeAmrH/u9HtIvNrM1wqaj0Xw5WpRvIG+X12GoyJFsajqrN
bu6R5ucDqC4BDGVaaT1huKiAzlUW1185W7K1t/RVaQCCJaL+TaIZJcYfROjrSqqaNmJKUdqjKMex
o0dD4z0ffU3S16eJPPK/F0U87XJitqsCXm6Q4vjMXeF9cHCt3QMBLdiYeuE2mIyf+a7Wqxlhq6Br
hdYtzvQuTl/I6EjQgqxJNluhfilSmkUyV36cSZtwBFUnJeJzCkXfiHgti8nvFbfK8w6yTfvdvZmp
rvUXNYr1/7ksMobWLVugXgBq8rXjzYubENouYyTmhW5ZnQ03S5pI0EUnQ2tln4uoD/mWMk0k7fTO
7qvUrposkKOVWTiW76Nsa5P/jO5ITnl/HNK0x3S9RjqKvYy9saCu8MLTleAJa4QvyumYK27nVEr/
N6BAxFnQBsu9gYi3aaaiP8Zs0jo40XkV+hyb3q4EGtcRrmemg3rrCA6NWEBtA4NKVe6uX0YD1shL
/D7fYgNPTdWdxJ8nLVn4YMaXl/7zyM8YfMakIObSQmDb4zESNcLQL/nf6lEMknPpCjXepy4CGAL1
+VSaBP3s32ZZ8nsUD7MCqbnb4PyEcd6AC9TtmUT52d9ovVEGZL/qikXqz2cPH0Jh5GoTRDer2PvX
vlQovDeY1uGQgrGgFB0leCOICQzB0L7gc175wuQYbhjw4vJNUTQVGAZe6irm7GGVKSmXvMOxsqCH
rHfmPFRsibjEmuMKwbiVNi6H28Yc2GC/9FEm5utuaSPpKqBOzfqIiYvm1RwgWT4L/a5cpnY06Afr
UdvyKPWmHrGwsszh8avgiS8rVAZWzjA6JfGeh3PHmUkSKYtcIUTv+noYH9QURLqSwYNBZjFTM/DK
haBOTjLk6xPRMgqK9Qvm56PWomdlDKM5UjN9qm8CsNU8hWFqNw+mCi4e7+kB3Y65I0Ku1DdAOcKh
uznnegLx2agJ94yuhO+AIqB4ctms4kKes/eAmrtUOhcwtVPiMLdEScfCodKrwV325MZTumPfRKC5
q3wzVquipYhCCP9Akx/640o4oxKLS8CNror62GZOiNnE1UhKxZKd5FzgUQamGkad5/9Xd0Ioaiz0
pa7+PlzXCifHvAVSxQf21Qj0EaAmaOS0r/AwwFnK0OX/zkIr46zC4pyKJKP4wxHFnclYt/WDymlD
mh2kGdrWx5zpXCSwMw5f1QFB81lJZEbhvchzwXTGio31ooNCu0mJ/qnVB6X8Z2hsqi5uP6UMgGtU
sMFx2N3ugM9id+eHmMvMYuuxMKCmJwk11zg3q01usTR3dTxk3l4/NEofE4Zgx7ZNvdQvnuoOufju
IszPMiAO8Igvh75Pm1E/eOKch/Sb/rv2JhRAzrktdR82hrcwzXAiVDMSQJ/ocBAY01JpvGJ+aH0v
Iph5guSHfjV23knFt3FjD8IXAJABt2zCAS/TacklvtIGtrsusp6CYIZ9tHc+r3cx3axvrpHUspAv
eILMNzKocjqi32BkgVTf3+b29ntqT+UfJ76s3Db5tsOIUX5XtFK2K4m9bnxFwVZTJEvmmePWz+Zj
nqMo6f+9kUmoYex2Q24tSfxHjfQPgVINFuebeE0uMVZ3/jb0kdBChWEJ/HDaKiyCEQj/5/Gq59Gw
b14utXvI/Wgcm4QsgeTDua3RJ8NAIm1gMPqrCsNRvd2WFawZrT6qn8TxMV1N3DhoBso5j9uQAaeI
ZW2EY9gVLe60XqkWs/jQ7kvvgl+Gikol2SBz48JWhibxMAuCIHjNhQ1Pw9p0YIrHnWMU/2gfxZ4g
dK5jXcD85i/6ac8bIv5jDJ0FVhrJ0Lm266+xviuZIsuB+TnksKbBYLX8m1ZI+z0TCU+pe2epB+Sj
TCi7JYpDM0Z+3Q8DOgobqrxBmZswhjjAjwsFl7vk3eh9i80okU62pf0HqJXzGwN1WpGSCvNsL3UI
optidLpdQpUBo5uQUL4kwwu6TlxjYLy4UlNYaZvBqOO8MXOlq8OnO+bZaZ0eseaGjNHfkmZ0Bu4J
DqgbRDnNP0CF3X1gL3R+pCDead/cg8ouIOpkXfuRQ3EUpssBMiNApfQceNxT//5UNJ5B0SpoC+AV
br1kFlE0YKuDJ0isTlSo27qXUpaMKsx6xlNQQ7PdXxJXv1YNni//VYgkZgazABfeIhj2/mqW1Vjy
pJ0Vm6iA+kTxPbaWeJyddOjHZsZH3+EQXPbqHLZtyut38b42xq7MqduqvKpD7SEASwB//OoskZ4H
rjnuhczpO2J2hD3sZQXxZXir+rmAvqXG45oQuDGWOvThSsuQqe9hhEFFp/vq/i61RoCIA+JyhOyw
FJAF5ENStX7sE7sufxqWaQfEqTBl9R5zoze5lSdhDRgSH6sFTNp3hDchiqo01SdRd4+3Ho+JTwqZ
dkWjfgaRvEgIKpOZEwYAnYbhlteL6jrG+5Lh2F1DStUKk8BRphZeCnbFUBBuSjjGhrIjdutDqf7w
Zq5dL+LzBUQd5wvgAmfUmbLKu+4dFR7R20n+6JqFguFR8dVedxKrN5PjehtNvCAb3RfNFotXsoK8
jvtoZvT0CSBZnuW9hcOjGUGklo4GBHCZ8vAL3VhZpf2oL1suIf8XPgKBKM+QVgqLuhu1FeLsL/HY
TIn+aCyVjvgl+NCPmMQ1RUKcyUYTUtLW9UuNRPtMXzhQH/OX5toUibSyOmDFOz10TUAFdI+An2HA
PY6sX70w+BdDhUrRRp5QDTXCM67Sl9qUGEaI+MS3pad4Rz3o7vl4Cl4eUTeBg+KjUbBD51Eok6Zb
p1Vbqw57b8zQ4c7lU+QB7iBPVyTxL7VOw+szN6gk1e0Se21AsUahB9gsLzTMqgGMSJy8gZaXCY38
dOWenoEfTZs2HMaS573QFb13BdrPw6R2Ix6Zwh+IAEa67CsANHzA6KkqjuStiEVrlpM6XRSBM/X5
hEAEzAIyFhpPgNO13HvqgO9nbS1uA79ci2wDSjKY72wzivAr6KqClE0fFL2AEiYjzz8aDWIYq2Yf
aXi1IH8ULwcCkSnZ/CaMDY9tDcY8c8SOJh+V/wOJlVKUnNE5SqddDYyiLmWS0o05lATd7JMKcLzL
Lw7k1jD5cJnkG3dGupIq6At8TiikVoCC4ikB5pGO32Z9bmbbJW0EoGhKISybUJ32kKG7WLiLV7mQ
q090c0tp/nSkUfK1dZDT65zA0jMCSUXusteRBqokYzm9pPKUTY9NLfR9yn+Af9bA/+4aQz6Fbn2y
6ScPLaV3m53B7q6sGRNt7akN88BQbdvvvLAH008DNyClnBvnWRfTovsJsFStJVGyuwXCe4mvfmD4
fkDC7qa5z8DK/j9/Q542Rl48ON/vBlUJ6vO+wMrBmvfvq9bnhdB9UAwNcNLrs5OFUa50ldsil6Mo
xyABQwPBrNdNz6CEQkg4Ba7yaRTYJKbgkUlaTF4BicxGMduXwY9aViBmjN5mtSLLUweScJCoBzVR
kd/cYmH/vfCzFM2aE6yMbKj5l2WMLx3q5D+QD7rSgkBnJTnPRuZs88V9EGdnafJdNwVIOge1fUnt
vpI3CCx1+OdJj/+Mci6uXRoQp0C9yk+3ekOvH0q2nzBSCtSPmT3vLmjOQqitbYXU44VqooX7QwSI
iM2fe9ovNtVj8UO8sbPvWfCopSDdeNpKXy15RgIGjkVWrqytsqmwD3bFF0oOENlEQoJbxrzBGTnw
YUrwBG4XFc/CTh1aaMvth8C1HYa7UJn6FuavEjbtfNqp+069ODNF9zxUzlYi4ETvweZuFvwxoD9z
kKz9dl5OkOOJNqRqR/rBnlC6VsSMbIIpAb7pRCtLOsobP25m5MKYU+dyWXxYA4gHgq9Se4eTq4+t
NaTNGr1y1oqZNrXprdiCZ4auDCmPijBNsLNFfE/lvWOm7MBL9qN8OZFNd/fdBXyDDMH3VY5Pc8ZQ
6Eje/BBacdiVVEDARwV16vsPOn0AyNX5C42+LbGU/99W49k+AAdPdhSI1jDTGLYzj0GfqDIJh4kX
ghTizBaF1yQjXIylIti8pPV3IQQ6iLyZ2C/vRppv70GzJRqYdRR//SKW+p726SMTB53d3KHcaKBh
o2OE1JXME8+FkEMjVaXcAvqW+u3WQdMEem2d0ktTTo4UhVn7iaszSQI7Lxm4ozTmKtjTji3IQWui
xrZT7+tu1y6QJzO0RAsHo7sHPTS5zmdkSsXKuF9QbIVTIgYGiqm8o03YCmBDXV6JYIVWRlVq3FFp
SJAc6cubmXKwQpjHLXgGqnYKCOsdKIZLATMecZcDrs5vVSHa3LfsOYPeQ+70bH3QDnNsWIk5rMy2
SfV3gfSmJl8c2xDVxSUvzELsorxv8rWnMLU7uwVNKuaGEkJD0Ht5jjavecVWOkjE5cyo7Pk/zgQE
Z+M7xgIZHHZwx2UifZR3fp3mb1Z/FvjkUc2v9eeKTZbVynM8lbkuajraIP72i0sKCmd2UgfKQRyC
RFD9fhaXrUdmBnveM7oO9/rZWOzUcTO3O581gNYeFLccSBt0/n/QyPsyR0TWKilTTAMu0XQ+dksQ
sWX/3SzAsFuBReQ1Z43VxhdH58mhC+VYPhuNFyJ6Y4AC/0h0kVEkF4woaro5ybm2ri7lwi8ON+m2
ZNcoc0GGonqAvM6GHnCBwgdyGeeVdV28LsCAK9PVmN5ye2JrbDTeBcbtYBO9E/3ALXqdDQVF69vc
U8EDJJFlm5tybCU7AAQNr3c5kVzp8nDsCVfjUEI1xAxrrlIHfeo1SxO5jea+TFSYkgCG0R4ZQVP1
0tVZhemETPikSesZjL8+jUEAIaK+K15la/aDw/4hxuaMkC/Y7uT/vVapamwYPFpMKlpNEDq54r9w
t4ZE54stE4Y+0iOSSGUSkgB+BT5Pq+ZBj8z6gw074e1DpCL3S2u21R3IwZrJF/r8tJxd+MJAoru1
eAMBmHC0WZ803DZTz2v3Qazo0Eu6WnDlrrFDTejbjTR5U1g4Ua/o+hGyxZg0vT8BfxRCcbtMsZMv
4CG+JxoQln+901Nsnu0/itYw0fu7OPXqHDaHN7PIKUUO/vv/woImmAAZUDxxUi4OsQsP57qFVzja
iwQInU+Tt+YEz2G8a/Ss91vzVk1FpUNsZNyrRW9hertz425aeowXPlG+PyeS0RF/I90hAEOdFd0R
5dJ0cLwSINtaInN91ALSX+MTxPogwa+8HPHNaNuLA4qbwRPKCpbcRgQgHHhn9Vh2wsk7yoFYSfp4
dhYMB9DjoORdwF27SrrZwVmdQjh530VLGu/u2rkP9rqQGpas50Dd4skkgws0qaw3v+qtk3il76CO
SXaNyApKLd4pq1Uw/OQbH48AxYx9aDc8IaeW+RtmEF+GbOcFK4vd3AVhX7ykbkCUVvWanPTPWL2l
48n35yJxNFE8GzGf0eUDdGWH9AZKw2ckAn9Ke7kmJ5ccuO46M8NW+LQP8Ntbwm4QN54lRKMCLXnw
Qu5DSJ+1WQfc1KsWr0owXPtH5JT7EAHcmazCePfSj30L5N2hA9QjDscCapL0mzsLT2nd2uMhaM5Z
3yHcrWATn/zaHl/9WZQNjCwcu7AG+MGeCZ9Mk7hBaE/qrHbwoX8fUlyGxMCQQaSO/nYAx3XldrPK
xFiU2u6eUK/6pT3TACveXFd4+v2taEvSzwzYS6qAg6flkWRNemfJjmdMRdAgKmBHT8JIUzFyIvVd
PhlF7cFJJXZyAnf7sz/sSRb86I90+zYwLlvv7vQWlrHLT6obFkEAqe9eO5IkpLV5Qvpf6MG0Lz6A
EH0ZLgsaTInJ+uZ5sTP8hILw9AnstFL7V1CAuz/KHl238+NLVSABOfwr05wN2BIxNd6knRojxlx4
a3d7w6ZZxCpoQvstv+ELC3CYnUbE7kA7fXS5EWisrzSxAbvLNhhifkyltsxx2nb+3QqRrcFRnUPJ
mulN+TJiW2ltN93La8vs8lJZpXK2eNCLqIX7xrJPgWPhlvmm8+F3AeOZFUbxWHSjy1yfqhCnId6I
cBA64KpNgDmPireJeGgpY7J+IDPiAbKw6meMIeq3imVsbcIG5lIbBYC7Sj4xs8CZ6GP54cbhObAl
UwsKpFbl/m/JaKq2ududT7+3RhEzSxvFG/74crVLtkKXTJ/vbvRAyb2g5tNPb9ni7YgrVx0rqdqO
pJY1N/JShSD+bePLQqUkgbBswfxZSvZKOrIgrxDWodihvvuixAUc0FJ8WWYq9JCVwlNDgEVloGlx
g9koECpZ9K7r9v4PQ4LQlEtrKW1ULV9gJiJI3+ILawtHRFgEgmGWzjJ2rv1LVxwubYG1Cc4uAb/R
THPjm6f/ZhzUb8IGEgey5R4a2dW5aIjTkJyzAm1XrNBgasSv8YTyPcc9pXBKgJtkwztr3TbjDZXU
osK/il/DYbn6RWCZrGcylBOsUHgQLv8+aQZCFwSEuZIGDi5w/qHzLlCIWd84W63u5IWHdsz6RAD5
OhzbPWQpkSMnD9vhhyHWQyN+Mw4vBYPvvZuOI6BS449FDKo/ldvNRl2FB5IDMj4JBTFScnfsT91A
3rI4n8riTjEhU6tYJNeQ2q1xvPRPYwfAhY6fovNQCA8wMfGBv8YgaHPbiFmtJSiC3onfgyLOuo4f
Bt65eqDmiRZI+u75TyR3M7n4Wvi1KLPtw1F0UnsjILrJ2La45dKGJG7YzXWGhmLEy+KDeIzLeZWo
3cjZQMqxd7s9brmCJ41MVltf7T1uki7ihIVJuRuWpUCuX2lpRQ/7CZZyHjz8Z6aSwPCjYoLZ73aG
9uGhzfQYMsr6Tftd4XTZYuOo7NALVGhRhawouyjxGGBmO4VXMloOTfABXkrx2HdyJY0Vnuk+sjkY
BJGo+xMKFdM8gHZVbyvDMJI2zyosHZo8J9kelnzN4cQXM+fvSZN7zh0S3MPeRSinw6MXIP1Emic6
TRmllPhTSZG3Erk7au9eFhpQAbCujTo59wdjlOfY9GQMeaLluD08HC0BbwUUFrlZk22sksUYBrVt
IqlFV81O34pjs7/QCoJN77qHG6CbXOzGVX2gvMVSZU4uyVMTHYtpbWcbtHr/5owjJv237PsE04gJ
t81ldzlwia5uBOck44PUzjAUeeXSLPauzNHezKlPdiC6q2nWh5M7ViOXPucqPZdnkdOlZHgC9vx9
X7eoyypiypbq3Gc/m32CVndokTz37PWkROAwh4oyQym5UCnsOzHp/bS7RQ6isAZ9eF9bu1cnwcby
r5Cm7q5GsFUvFHW+1vs/272LfeUuvJ6CB+qFB6ussadr9DJVSTYEVjuq40rqVPsI1/wwlXL5VsXw
MiGiuEnWLk7XUfafzaC/IuIHXTxxav55WDR5dpYpVAAcMVub7oInFbwM2YLQ9GiEwQXA/FyNNyO7
Q+skwJwe7aB1cEBaCfVVMqYhbadorJ3h6Uf9N16noRXky1v/8TBojwosBsupX6mFwlvDD6LjESvr
+eA79MrEnM7V35RpxNuHlrYijZ0fi0mkmmE73zS7UKRYU68qmq0jhEw4ahelo9BgoWlFOdUt9YmG
yxifEKrf7RJ6nV7y21KSQGjnXyIBEnwg+FnlVtAXDJr7d8UWQVLY8S59FeAeYjIELO24sST8gGAT
iY72qRTJh/Q3uzaOyE6duQK0YWdoOERIemTPfUBGH/puQouGp7xsLwPaHSriEgekl7ST8v/2xrZw
eYB4too9pnx1BTG6QU2YY4yTCDeT74fBayMuITW2x39VqgkL9w+YJK8ayuw9x81HyIWKw3Fj9y4z
YUedSsEG6CKzd5evmH8/PRo+rfAdnl43cMwcmX86Nd7rbjS1HVj2RhMH7Hnz5FYLSfoT39hYgVIh
45EQE4EA4hWLjvt/DH/WntTut59LcDGLDV5od7M6UGd2QKuyaw/G6bg/em0hQzezThOslcbH5eZC
fZ047f2N7nQHbZNxDQMo7z+KDi4lZ0L6Q9ruySdcdH0XMwEzhVcD38OJ1VAo5zBE97mwR3VoNCOU
xBXmaVVfIWFdH4fekq8I0MM1X2SNrgEbSCqsJGAu0Ax+0VVguMlboeIeQ1nRgx4aAC+Ds4KRse19
2eICOmxbTap0wn1EsfqY2tOMlrK1d4BKVIueVjoMBRj+52exbQ88RCrMHlC3e4IYknlGHX71ezRB
H/dsyqWP3EjFnXkKJ7DY/UvDWw0LYIDg+L4P0LHmt1cWaUKpMq1ZW0tcjkQfzf59Y4h/PdO+l3QF
gjVW94w7z648xjO3tsV2riCICrtN8BcFv2SKN3wB03nwqNapZLTXN3A4JrczvPxoERUznINfFbgg
tNx5DBmPBJDHp61RdLdl39CeIm6nwHj3rSTR/pr8+3T+PKIK3CGxpV/RNklgHlktDbCbusmwg9+Z
SEtMAzwcVnZ0PLIDjnyMFDJAE91AnvR3tDFhQIqx4Y5e1moH2yzkJADcTJ43J816eRp2AqpF9DL6
noeB/Cp+/uSgL9wDeg76DkGnJLQuPG2Qo9cq3yWTR2SbSrH/X5nxStdI0bBY6cvKsGzALWCMzDX3
RY0UdczHiA+ufxMKWA35+6Ji0uOlX1AhkNupNkpSkAe4zC7pRfHGA+Zf1LCwsC1EAiHmRUqjHObf
B6Eg8Kp3fItChQmQFPRTuzS80f6br0q0lRxgQbXTMxgE/hBA+fsm/NVkcAoU1l7jv8xb/1/pcPty
kxqiPhVxjyBXI4l55hP+TXzF6lyocqYAUjAwbUKkDvhnsE6jUHXsfxOvBsoKTkDlvHmtEhHFqqyU
sZEewgAJwLHvU/0m4S23R1ci2Da41jVOwxLrhKBrUw6BS6XfMudxFo48Af1QWQkkUDE2xVENjpkF
Uh7IBYOng2kYD0+1PO7xqjHIuH0qMuNdqmcSf13SISfZ7lqmRQWabmWMT6kKoriU2i1nezNRvAmN
KuBQV1RpB7yHxETFPAmUyykO/hfYYKvy2y093j3oHJ9V/p/kVA2LfLdY08OvlR80Ry8pTKLLBiw8
ZD/IhUboGf04noPjH1c5KZ/Klm3+IA9XaHwucKg+TzAtZk+WSp/ymeTLKqAOMgAg6e3Jp8Z2jFxF
g4sRQzJvYb+hhdrgqYMDNCOYgZeoiZoVX+/JbvygCyoczYG4APa1L3iAIPN1OsIclxI48B5WKVyl
nbbuL6s9VaNTBe08lHevcBi/qyMAJCVN78Wg3skoP1bzLq2e86XtVs20f3SlMruytZnvaheZ6Vkr
GxqLR7l3sFlfDvhnwfv+YlBpsHYgY70iOgQmvTkypo7ddwP7yMVz/g17SINZPJ8bAtb3Bd1/Lzbp
ByO0wY6ebMOPfLPq+Kj2UN0UWftCnVO8EQv4JXnjRHEC6LAVr0oawH4QlUOqxKHBa35qoiGlmIjf
1/hw6jPCHfI6g9MxnzscXPQnd88r9gW6o5tU3PoGL4XPhr/nIgVCcKv760AqPFB0sWgZRjQv+Rw9
fdIEAdpdcmbXoQ+3+E43zsjFsrGnDm7ITEiqEijVnhVYmL3eMmtBI23IV+Hkoiy6DSu2vqKPnEl/
syOkK0r91pBY+EFnBzTVnVKkZ5XULaJL2xRiOImmPW7WGR5+q9tmXvUgNtTALvoEHvhiXOfpIBzk
Q0MNGCFIb7qH1C2MxTgVeVum5xZmCDcecok327qzqkez1KHR8H0f0i5Du1ogVkjOy/oTz9LLMBrS
iHuooix7isMWdxOa4fJq3Oi8yul1Y3nyBdSgf4uSrYoSye5iDBJIrmTMG2RQ3M/GLtm66Vz6bIbG
SFA0RBZxds3uIWSAkHwSRFdMJWH9WdFpHpo/WyOguxc/E+O1rcDfSF8D7hZ5WwilZoo1ZPvqdBP3
sYV5nlNtN1N7/yicvfPald+6y5jKjBAWj9TAFc9vwP8dU/eYyRXi99Y1x/tRtwiL5mDHSkEKedjc
AwNztAYuoovHIJPlTyvWih2fGHLx3nyXtdTRdwwZWoUn24lYMk+rok/2a9VpMqP9DOXuZAEkxqQT
ixkOBl5Y0k7uSeE9nUjbFn/98YaGe27+H4yguqYHx6FpBRYb1Nr5wUsk/5yVBuVecC6u5Yl/irTg
gYzb5Uhsqpt1N9J3ani0RxQNK/qhBiKKGT/vjbZnwA3VDxuSfc+r754GtZ+rhnE7I5xxlt9hLQEp
1GS4mRkrGHSCvn2OKVLEFugyUq4mWL7wMsxO7+NnTce/SNnmRbXHDsbvZqLHBXPlce+889lbUnyA
kVQA2S2yTJQHO7yKJJPMxZlf/HmI8JUEPzGFQyfM1ja3wwBayrE5Sx9JoAnONq6jjkzc3KcMclNw
u9H47nAhHBozpImGgPXYZbZrZFhyIzFiFJUS+sqI1VJBs3q4Q3fLOG/4/32cUcxi8XXalAdh0f3z
ntxMw8SWPLSMkFirg9xuXLjVHH+a2eHjVofZbohnz4RDemk23F2+SEavw1IthdZXSUGvZ8sL9YsK
8ns5H5KXUfpTlbvLvQtCQmaMNU9HT9XdW+5J3JHoD46PQ5ZCKzBUo3tOZC2S73DhoxpXUnFOkcfl
0h5nFGK1dDICnFojqMr5ZYaGPK6ASpbItrkdeXPqzochilevNVzNhJyk5u0WXiBblliVTBhTtbLP
kadL963RPrcXBMv2g8YsyoLz+6LzYqixNmV/ypO/3ddVFPsnqPFlHdjH/Os30QZvmD/3/dYAQZMa
LmwsEhh/ijdoMy+U8rVU7kDsTmCGm7DXp47O323zchVr2QwFr7LmNFne3VDXBJ3Zp3HC+Jee8IbP
3u1zl4PGlX/SYGnunkBvzFXx2+FJvmvHj8SqOvAw7+mPipEadZLu5V8E3bew+yVRYT8I36OLm7YW
KqPIUqBA8nITRtBnifK4lMByVsrBqG413nqWxPk2MGZlPZGSB5AGCTPWTpbMVQ9VtVKo+kKC019E
RyQ2x69+JIYgMfIdJDBv680rCZKYQGravxpm8/SipNLT1K7Xt8qb9gagaAH9erfK0y4bbnFzC2dC
Z8qynM2Msb0n1xW5U1ipkIq0nkMyxt24YPil1aJJwyE2waBajE40He6W98PfCOTibhZzXHPBP7G3
XSM5EG71w3RLH0nlHd+s89UteNWho09qeQr5kUBRBkBvR1/wjQbpRAz2JiH00PsAi8upD1+FwY3U
1qjsc1c5XZxgmepy5OT0qboVlzAddxVMq06g8+t1yQ67m/O/KVo75ATSTqKVhsR7WMtRFgTkM6LY
UmrepT+t3ZvN8HJZ5ffENzZxsfHNf5EG9Umx5q8vL/Ysf0SX827lOIYJAd/rBYI4253zDBWVbBaw
eqIwhf/kGgp3wiZyY68195DbI8JC2YJWch0a5tNMYVKohHJhi8KwK5Lg2la5TLIhhtlAYslb5tZJ
Hbt8PClClikkvLOGydVCGlGG//obHFJk2L8s4/ZRdjy4jQy3fozlH4k46hbX/ON0UKiSzwRQdL4e
0+dmP57+KcQ3r8Mq2V7YZbb4vdge+OWrxXkY5H+hY/r4qRQhmoofDNbZj+/sWw65NjhjYRAnCW7/
s+GOlYDypsb9CmBcalp95gtOGWiRawE1U2ZxUwkCmz2gNizcnCV/OwF0oHbqtUdoOJPN6J7Ws8Du
4nBJJaA1tSajUixL1jGgp01+VzGaFl048olUoOfzPg69UlRf/SYWTG6VudH8KFKrT+gCSZALCJsP
BAxfHEBPub4/ghzvJuUBPoJs03DNIfRJmaoT3UPaID5pgWoEHlWtsApp7iJHEM1owM9pHCPurC5u
R+xFx+M6mPyOfArgJndYE3XqSufsXFsJD4UNhqJT/XBztVpCwraHPsHMo601yPNEQj8l0CiRshLE
3uH8Wtjge3IQ/lKXfqYPZs59/gY/IiPag/WIT/MFh1T1Ctfz+cSTokQK6tUJ0mg/QE6wB7VsLGj2
EJkKF9bBAEcZ7Om3BCwzlPJBY9rq2jGgCaAaIYfyYmTf7+zMOtrUVojue0RXsfggwCX0J2GS07pd
23ix9PnyUMew53EPDMZGchwbBqc+bAzHHbVAtOSklTXnbCk90s2B/I3ih0zRJ4SE9XZBARgLGdfX
yY1N1H5HqJcnqHyV4smVke8d5kGlUxBMxYiV98lwNUOZyKPCwhvIIKC/oVQlb+VYXOopqinHvfuc
GymynMyY34z8oTAyN4WRAmwadAX7mEtbt1CJEi1aJoALcdRKjM6I5+uGthLEj4NfOdvRNgAageFK
GDlLdBdF1GeWk8h1CR+fj2mX0g7RM1YSdYVDVbov1OiJpUc9WP4ljqkNb+5urNdPT7xgN87Sl5Ui
wpXD8uoRA8xJ9ZuqgOb+KLZscyYl+ibRDb6vweJneLRj6vlTPPfUlc4wq9HxSjQcVtd72hY8GfoM
Q4TdpiWjLauXPS90VAAdHThEEMjUntAlM5ZAmt5s2R12S7Zl9JJOQa5vnbjuGYHe/oanPQsioXoY
2ZKSngRdchfFAy1tRSWgdeu0sCa8TqMMXxF7VQQtnAC8U6XjVcVme1HWpHLDo00Sw/bDzMweKBZQ
jOegjDU0jRZzA/ql+LzmbdbI6tPi4L5THaQyf6oPzMfh89CyFJ7hdv+yhVGfRu/HiL+1Z6weXFaH
wi9n5Hre1SdqDrHHxcW318tpYhr3f0LALZW0uqVX1YN6ScPTCFdebr5opnvUxg6WlOzyIZITnR1S
kjNWJ1+KlNTkldJUHuR2Rv43EAvXF+nlmxSba4wqgGr7Hl0KLtagLs1G1E9rkhrN+pIT68tGlXOK
Wj7PWmngNS1HN1LlI1ZzRlwlmaLkh9++tqHsetN5MBvXAj+1B5GHu+EhUvO553XtZoafB92dLbKx
w+2clOEiuvZp7a9yPQM/8WMf1foPAPUqXWKGdHn2QdqxH5D48ko6AOZQgj1wCqON4F2gjuepccbZ
BjQQ5Dum1Ea+p3ieZi77ZUlBo9ZUCxFhC7AytX25jNehv8Bu11QhGKGvyA2gTswdx6xDoDzizkkP
Uv5eP4q2cSr9xYrW8kCu0L+02iLVVrgwbQYBmdFHKckJcpVqJlJ7zXOG/POQjWvRQ8IC6P8asly9
YF0UKsuJkMWGkx/wqUuD/8UdIGolOtfi717LNUVweg4fXyJmbVIv/fkizebwKi5afqWywbyk8eFV
/Kn+zXB4xjYJzSJitqtE6BktX1AgD9khETmU2uJ3qnN5Wb8fjSn5IRyn9RI29IrUmnahtYjOB30w
2EACPCmRw/g0NtoIeEUbyPhWvaA7qvZF5/m8QzKouI86aA/xVzOlNScHbjSFUnP0K/BIORsTuCgt
lk9NodPWn7xd4MJmyjfix7dhMW2m2uANqfUFH08br1P7ypMe32luNtTDRpZgxcBmig4Vp9bYlrJ0
BSn6KNtD73UHqpH2UtalJtqbwynD3ZDrykLPC+ExSzB/pB01H0dBfYFlExu6eUgLlz57MpzTMBoG
vaXY21h9GiaTGLyAczFDjfOI6n/TtgT23jIH2laIlty3tKCfsDGDNZ0x0VoYS08Xl2PJArOR0+MA
3A3f8qa0NZmXMOmYhO87m+dvGykCD7C7QvGVrVIMqxwTWby923SNgWiPywfnVo5SNZXL+29EvGbC
8etHan6+RE1NCNRf0JQZh0S3bzjlh672a44rtaGwBw9DSqRjBttoYuj3nveEkcR0fsMqGcvzCe7L
40XYJrgdayq84s8Z7d8GgAMUNNGoPAa1R8uYvropfV5LHsahJ7+MV36XoVRCjuJH12jtal5X0ZlP
D3egOjq0PrYmpqWEwmodfxlf+Ez1yX1cMjtQXc0V1z43Wf6CWRyHO/L2aJw1SdDzreYHSeC3NSBB
LwtdJN4x4WFzmlml6hxgwxKevnmnWmB6hbYrCS0AnwVztbccnYe7Cjl7kmRc6yqedU4DpwzrbM83
FGjFvJmWQFDG3g1eqQzew/+ySoCAoHc3MUWS73vyJ9NfsshLVwXyCyN8uG+raM4+MNwM63twEvZ4
o2qnVnK/A4AS7df4ganvD01jVd/D5PZQkUNxLl/GqE3P8vUpx7pvH7UAi8JkjOaPDu5+zZHkZhWD
odLC9qGErz3G44eyiQmHBhUsKQzXNoNtal70zmlNu45NHJuDUN2/n8w2NZzNm8FnUq+0pC7DZuw/
x1liFUTmBWnFpr3VW+I+AB72pJ3tw05ngNdKWNO2X0+tnutH17QHj22XywhRo09M9vs/4j1xggu4
0nJ4EKNEubcuyUzq7eeyiqiYC4jLm5XY0u71BXT+zmipOE/avSiJWitDtDMs6atzKGJHdT2YUnz+
boLu82d9kfFR2e13tRpg7fuwiy4qste+Fawo/ONHv3YpKkUDxAE2D16Ha7v0woLAQEI3lgUuqItp
DK3vJQupjmhGfW8g2hQn7HX5ocU2D+LYn3g+cN8xLjOQER/PY8x9uO+Uv2PcBUlpnsYxZWu3e0+Z
PoRp0sTmMYkRnNOvAkooJxYVtJ1px2iiNu/8fwXF/VkGYiZ895DBNYOms49JKY2EZ5Usgi0LNrfg
ceEWZ1gPimTM+JUT5RkLQ8QJxb/aH4tuyTZ+yz+m7opfMWPXky8DcGE7moa5+B4n+tMkAwySDHJs
U2nfHF/TZJOzHuYAq+sjvCtw/7TPdn4j8AAKsdHPTG2GCYYgaSV1J0L2iSVgW+UFGtYkgDEFYGId
6bvuo3rVG9y5s9qf32PwwG4eTFzNJkYCO1oQWe434a45MXSj/gkobF4OMtxwcJ14weHzOzLCERnO
FjZToS4GBxZeAGK5IovznGPeo8ConarcHb1RRowAEk9oBmfEhEu1b40gP7K4T6YZoHiVISpmtHvf
R/gYArCVeD8cVz4TewExw2HQMTh6kTjn9Fp03HC+qXNF7OKErZ/wgabXk4BzFqOWxE7XgMUIoQlA
oXwLSEbXjlC6uFkPI7ECuRyMPPCR7laR++yxmcrZFJ9sE9OSGOQiTuS4MNkAD2E+tHFXnWp052pV
dtPSHK7NpzKihpxpkBhC2bzz4rqJTF/W1Y531uIevwmUHRotC/aBJHRRIMLfA8kwN7ppB1GBgzAA
HQZ5Pr5D6bVVf44Kk2RBWAAwPobRnAtzl2AA637Z1DKFRVwwhSjqVu9dSl2d3kC0p/5q5cCjq5LS
UYKvyCTgLbxLxMjuhf9iehy6nvEu8ngvFMoFVDdSXQTipQ8XIlLuhW/nubpzz0GTHKD2DUAPcrCT
lh9Asxuxk1h1vaVckDgCn0uoX2q4zeq61d5BVFKYkTYyEQBBswy7cAMiX29hVlNLzGsKepjs70e7
xG1CoE2nvegr+1shvNX4rO+SI9v/nTjfA2KOIMLUfZQu+atje7rKWy1kMnkAotvQfmZsA7GdsPcr
tE667HIOF5NIAusNxibrtm2bgSuJ5fLOyv3xpk9qIvq6EeE18+LicF9j4woyUvKb5H1VEATj8hOJ
EZbjWSQ7M8n4zYWRglyry8z3DUO5GQc+wxh4XXDQ+MVjbo343zvmIdWDjwb7Jgu1K/EviDKWzTBB
hZhJFam/IT8Ee0ChyapwQiNUB+KGt8mUZ/w9/x8L9DRnqBJq5Plr7kn2vwPJswwn7GeXv3njQaWW
nV6gd08sis6TX1sUgXSVRS5+J7KxOCX3T3+CDwYjrUarDggtCmcodDUDhTp+1HOXEZdqu842YCSX
gCRyZNvB3ZbvD6CMtNGhqkrZYgi77WSkQnT3a8zColYMz5xyajftqq4yq3kn7i6NSNKwqDKODOGe
PpuasJyZGvqybsgufXNzgXWPaR3I75NK0T7sLJXyhMIEYbqF6GA3SHl6wfvfkkqoGC19qamcZ1El
OrQGEfvVeGOwxIQqQmBj86nV/S0s/KZ4+WZfQi0PVtQYOOBv3iWIwB2s7FXCCIx0mcRL5qaGD3ib
BjPJrAvSppkSRPEkm+vPRVTyaVdyN/wJvV7VFTnRqJ4iuC/RMBIroKACHGBdRa/Zx+L+waVx/GeY
ExtcVqwDDR3r7GrACMnYdPfLPvR7mKpxomYqzOKOFW3JkWRkwMIuum0Pbg9zUZGYWYMCDQz7+grm
HutInsDQEFkkWNCx3thfnKZ1QggAmhPxPEN4JWyFGlMBxVUTVc05Y4quswpVrJH5KBuFYRr5qmLL
lj/T5fAl7nC+1en2rmARLWQYXnVUl8S9KTIea95Q4zAQFbh1tVEhtpklj8ZUrWQC3jDQKSR2EorF
fK8vSCOkxb/qpi55aIh6gFOOuk0UybDaUPyHiGyZe98/sCG1DGVLxWTo6CO7fPBQ6swA6teOGzyw
jxwCvRKW2MtQVqMPGsxLTbnQd87EuhRf9D3Lp5NYbRt0Z7nIPcaT59GMa1lGAJD0glC8xR/wD6b/
/nKZ2eRV+7CWr3AwJNgRhRVzEpt8MSQhnxkW+JQODNtfLtspFv5q3HRqxS+9yWwv7cfR7w6Yo0m6
TIUe5D3OJSI1hxWVQgHfJz/3Ty/zIZrDGOEScGcywIlzcctURYuQoTv9RyFjcBOv6sanP4oL5pwD
/k/K2oFJgQR1oqbVmyzcS2sWfFnDlqNgTBsSj9lgFBKzGTZPgyXf7TGPkj/s1QwxmFXPFsfcA1B+
w1vGwTxfTTRjA4EYO1ircfbKvzdRYAMy88nqAhaHjDxXW/xE9c1jvd/QhITwHe/4B7gZJI4rVS0S
qFJPZXy4frHjcJGQ/VDjahpVRc21CJ4wN2LfZ0EslrabLW/nyp5qgHIFN7H5+yLe4Ds97B/kJqmB
rx1i+EVX2JLqwY/kp8mUFRiZzo2KAI4CMMnPh7vm0xuvoW+jcRFHdRJITEji1VbUzydC6E9fotR6
fzca1tReEOLL7wzkvLqv4ZIRSDojXpMLLBkWBdd5PLmN+ruFQpEbf9p25kJak7IZnLxckOOpvE3m
J6BkLIOs8coWYAighDQon17achp4my7FUb7T6JMP3TN6pAK9+T+UP95tzwUs+oQJebnkZIYW2waQ
kO/YT3Fhp5Nlh1kvMFoMqbeiArzv3XJQmnRVOod194LJEjf8ZnNr2lsENFzZ7VewYj/hkvKga8ys
HSJs33l2sQGUelikIugwIyrUJUDiwkiWPdgm8VXBh7jyPz2ohTuvrWSumHcDzznrycskE2NY+d2y
zXNhZlS76rICGWo3uYrxNa7hrxDcfIDRPR61Pl1p3gP5OjdAwX7CExQMB++fWYc9Tv2/CFAUf2Y2
STabxiHCKllh+krpVnnvsjIC6tBIz3lM/3ZvO4KBKkbgac+vV92U3Fs88xxxp0dwgKqQtR9YsxoD
VMozdAieBRL8GRbs0T5RqPO0gfkCBbKOgk7N1agTFJf11orotLhL8D0V6F4jMMCgMtSHU2SokyMr
aaUDHuD2vH1yyLKOTwNWNKE2P+DSxQvFV7tKuwrSoBIuiKqtWIxgGzBDdFCo06698zsH/Y1mlxYN
T4aREKx3MDeGEprsqL2fBmez8A5R1ofgUdnLkPSF2kBlQOfDLpgSCMrMJU5CYkP7w4xMdhh6RvK3
v/V0daFHaeFXRDh28Ujerx9MZy/gDpiEaqNTzSVMX6jmRjU0siRFMM5dohgvuprXvTaQCHaegLGb
E1bDcrpesz8k6mosoQdtdYoOk0jFvz8HFBs0lJvd+6i9VmtFht7wZDbOCn6EbcsG7fDYUcz0kwtz
i8liXSU4IDoaHO6IuhykZ4eGUsZnFqOoA+mv8bnUHpcVR1IX4b07duBv5X62ADtiCy43q3RLrIWs
itD5TsVikwR4Xye9GFvlDebBgpzG9ya+cNWV7PBePpbTClhDO4TE5fdERc87O8bnnWzL13JTovgC
AxCpDi9PGqJceJyjwMgFxLGzKXD6Gs0GNuEROA7Y54zEcKvNjK/mh4oBKozhkqp0s6nCFEu2u7CB
KWffxLZaL7hRk6/wuDIAhQYDHoTOMBZ1h+yzw3mC7qfhqsgYFS1jLmBADG5VWkTpa5H6n4soUczH
UTFxP0zo662wSGwW91tEN/v3j1M381+RMQZcyuFXYx+NifxicKuz3Y9oAYlMj8607C0pBgFUAisZ
boZga4ddHogJFCcNELxuYMer+kO3cCJF1uMGl6Mv7YD1E75VGrwo46iQiFQ+welEJ1y6MIUPlO2P
0MpKAr+TbztXmlfkDcc4BnCcNTC32oXcricKRQ0ir9QlUKdn55XVX6kbxuur7zLcvnXWOzxYyFXq
M+q20DuBuZfxPe/A3uq8JD1wX2pq/UEObeI/p8v5BinYcOGZHQxHQFQ6CgqT0AQtCA2TgyeIiyky
XAs2EblSxM8wfk5ek5pXmK5HEKTl7OZK5rXgnfbJR6uKDOAKtOmAWM95nofelBtlnkJ1Y/U7Dz14
0Wh0yAAxjBsM/Mqo2zi7J+c5R6cmbNQGSwLcsFP7YGw7jWfuzMhr64RQNO1e8eiFuZirBY3N5jki
66WrAHGf8zK47pi5XD0DoDpkwEo1Of+MzCn3DLUu5GtgmTn7vziUx66xS117fAdGDQE9cUpGPuw4
BFveozeKIgAVZDsAgLIKJ1OLqG9uRmMRw1dK6gijLPuqykxvZ+UIFxP/YBjOEES+dMNBd9phifHz
iyriyJEEp6B5XYNZ4y3bOqgT2UreOLtcDfX/2UlrT1PK+NWo2LDJ8Ii9JCSYHv69yrrNRT9OqCko
3weKYIoRwGBTIaul1BXIUBAxD+2ljaJZw+HEopjhC4VqTrY6MLmMKKVzDJvh1BQN+k11bm1Pglzw
hpqo9Qp/htKP8vb14EqTIEvkW65mabbFwNc7WXWwr3+2C0J8MQVilz0n+4EfJW0FM+TYyclrNwFA
WNnqQlGeaExcRtX2+Gi4S0cZPqD4YX8tVeP5kt/Mchb8WFEond6CU9afGqMIkCPVd4ki9C15jhBd
gROPlFl98oVfYZnOeJBVT2ZBcHBz+KmFr8JcBy6yBC1NwDgZkXx1kVsSYgQrA0LS25wxyptNK5IR
bLiRLwNQ+OviGOioo2m4+SEukCq5sQPZrUnZ2At+GKKui5Mwgu9YV0sASfjGBjegLq7UYSbBJ0AH
ChrimBR9bFyuw62/bIzTIs1pOgqVxIlbjm8mJ1RY+w9jYYYG+xlvlTqQQSXBR1wqQzxaJGfQbmrp
+uOF5VtL4tbUZeJIuLm0Y62GnaRfE/FwipSEj7QP7NJZQSx2qcqiwfaeYn+IMZ/QXFt9hqxn8Ggd
KLcLehRTz6oY9nIf2rN8bRKzr2ILWG02qEHN3uiTXH/YOblKxBIm6RwJgZnOyTSioGl1g/HP3RKY
qRNieUNsHl7gFEuNznqHN2gYR+/rbBcLRs2t0T0be2brw6KtFy6iT8cZcWEpFw9m1cCscmwL23rL
KOPmPUtlsD5fQ+z95Mp/C2TVenFh8SHGjGtnKg/RH9/7ygh4o5yCv/JqTbd9ay2m/IjE5w6wf2Qd
C2P6EhMcDfLsj1dhXixYPQm9EGh+DLETMXHXJrJ0zNntdBY0sEBl6zQEuH4nNT0WyT4VmMEia70g
khvTvV93YfiWan3w7jQi+6q1fcG9xcRaVhWCWfe23R4Nr054Fpj0FLyH8x4OLNSd2H3/7aO7Smwv
LrYRuDHROA2Vw0aPDGtx+ERkLeUJa2y/OqlBDG9fCYJXKe3iJIiiE5WSAl4ooByRmhn5e6CyG2Cw
d9LNMO8M24Dz9R2imn6KCbN4z36KuwZVGCvSf+KF2PZjkgzs6LIPfuhngPfo/vUjWbpo5t7vyUbT
r/o8Wv7DCXpzy7BwnGPl5/rgXnzl+l6o8alUrkYCOzn7nRKwP4kX3n2ykAqTB+dK1weKPcsQu+5d
ncxo3SKtv0wjZGxHP7nM0X5DJzAMYIftq0DNYcRSYa0e9Wjey9ISRrkjQdC7y/XFAYkDrZjof3Ii
1PKges0rth5s7rca53mrFp+Zj0rYwKrm9RwkdzX6LTEfhBrZAqHPLNg+bVoT/+MH+cyR5CblT41v
NlGa9k/2/XXtZOWemBF08iJnIIne6iWog4tfQv6kKM/C/K3HQbm5+I0O94yHhW9bGLnpU0L5PehI
++0svNjfrhCP7/jSR1dRC+a6fiN3BA6ltdCnCWj+CDwDkMB8e05yv0gvm6GUW2oOaw5WnD5yXTHD
xEv/hMLOjf88bvInZPhfJhySZVEhNdET9Htjx92FAkh4SzVWZma0CmTD+v2Feq3Pj5DthESgRidA
FaakFff3gl2aLojS2SqfdgZddpMqbgyfwcehTlQBh9B8v5HT8iVsBWT9BmBZkmNGTUKy0qXe0YzQ
UFYr6aJfP+0RuzPyzWMywE3pUrQuKQj/ZO15+u4/hR697hLHbrpUgKqRpBwjlFeEh88nU2EOobia
W7QMiaNzP+S0kFqP1KbNsv6axZ1aGPsGmYEQIhvdHC0XJ9FLpCi63A7nM4zW8bTF8bXW1oz1cFRN
pgqzQQrYfRo5Z18BpiBBiskwUbBMR+FIgflFjlnv1fhEtedBk79No+MMr5vqg8QdjsLy+nxmhJXY
MKzZ0wBkEE2D6lvtsp+8bVyUVewGc/q9oiUjnYYvrKFlEHtjzJqOoy6nYKrKANvFI+0082dJhr+M
ayEyYA/UMi/w+O0PaWBrwOfLiePvntQ5DqLimwD6wsRPYPm6LaHvfKDinNXI/MEu7Nf+wbCtcC7o
CdAoudZTp0hQBO22spfj+PkwPGMB0jRkqWCHG2vyqcPUniguEkyxWQlIcGEL4S9Hd254cQiLFP/Y
3Z3qYv4RDgduNdVbGbbD/pRYJFb2HMHqPXhar3Lkk9OK721zZ/txKMc78QHx2NUH2tSg4SuZGX/L
oPRh6kF3gSwVOJjTu+3R9KFahr0tKQg/+379JRdsZml7CbDzYpxJaQvtS4tKelchtX39WoZVYaqP
B/bAjAg/AO0IZd7F/0PxnYEPWxch8hegWeSKrcKaV8F27BjkhDbecQL4j3q/bF18Mr275vY5Cz8M
FRm9QhAIQ/rTc0LB6kOWpNzShXC0ll7adGSZY82VHnQhz3XtUh+/VfIOVr52bUVDiL1RzZamfgF1
6rN+3lGwEKx5LJQskWhbtVxqwwlVkwePgmaTjKeardGtH4SvGVQkSl+AE/2wieOSAPGCqsl+42Oh
eTO0xOt6bPnpVFZYARnZTDXsrLzRemScovkOPKv4NMnlXBHxjP+0jpeK9i87VeC0dViboCk82lCN
1cTbu7LC+QboW0M5d5YUC3CROk0RJFigT8edn8nh0Ds3E87ooqOpNE2ePPk7jCo32LLsMkbnKWbP
kPcKF6BPNaxrInzVlDvlBfHT6cq8dJJD+u2NW+yleLWiFXAxV3dah4GOT2Pkmojg2uu1Lh6LcEpV
m7oLBNnkoWV6neJPS5ujxLvJ/M15UJRy6gTeBiHqwWkZpqIveGkIXUdHpaY5Ih2jPjqZf5O4Glsf
GCV6duAeooH6gWo6lNsLtwuKG8zPFgliXTEptrkM6Ju615d8w8nGeg/7rxoYqV5Q+uVLpZtRnA0G
YWZY+du3cc6kVAUProePrMdYuiLXRxBD9VGPVkqEiFrDcNXSxTmjiuR2JK37AhbiQhIOJlRmzaOM
Wz872p6FZ7izwsL1rrpOm4duVorLrf2D4pCGaymOTvvxYUCccezCfQBomv0VS/rG0k18thIPhxN3
YVUeCAsuOmbrlW1hxAeIkwPzs1lSIMas8Rv4bskrA40ihsV3Dv0KrLd3COb0C6U+vNmPijaPDv+6
Sws9H9mZ4txevKYQaMTUujbU7Q5yvv6/IHY5Zsb0YK1pim6AKzmgwRpxQJwAUTXg8FvFpgEyQKuh
Gqi3Ns7SGhDBpR/8QMNgKkLnGqEHbTF/rIPK3JI8Bn1eMwG6f3yeZdYNT/IPmericUYIjGby6n2C
DgKxTp5wlhAjMTLSFmPrgnON2iDoGgdU9SHEhZY6JvB52upKSjcJbsuwzrILIRs79HROarf0HIen
BaACM39xmpAWatdBdnnYYbpAxhgHLiW8bfsE8+lwHgev4tmmPtrXNQIhQQFBP90zdJf+E6BmVMRB
EY7qEmaXB+j/T9+rCLpvxhHMbyQf7bSSSsIePQaOFnFc8sdywJe65mF4tbaj9/MP+s2B8WPkIo9+
AuWTO6ZpVHtBVQCoS+uhnouc3XTcaTg5QQXq/QBnwRFgGTWx3EBIwts2uuSmN7VD6ldRMox3w+ag
8LFiBnq+d3/A4lu3eZ7NnXUI5HvmaFlMA4JF43EBTX5ODJdjLAY3+y8XGFOiPeeRkgZ65/OKVtZD
SpgCA4ysR2xhG6M87QcqTz/GHkxeQGmTzCevkLRD4kXAzqcO3sLVPW9RfDvFS5VHO4xKdXIHJbbO
zoadzWVzdCBMpgA4agFJdDUU+OZ3cZcM8O/FhQn/3YRVNQlHbIi2IjUDy+FTAvISwraazMGknMsL
4LVBOevPMm/BSZOSfzQQtY+64dGJy7DP+FdS7AY8DEt6Digkg/g/npBK1sJS+TfDBMGXq1r6EiwA
nJG4A19t+yc0uWKpIIShSBpjxiIIstuhGibIQRNmPkOIw8RN299yGQ10ITflPNLMzIlIm+II32a1
JIaSR7rlR2iZN9MKPNIkP38T7p1GXCba5bxvrlgDQFkwZc3e06m2QIhKtcYdDLh9CmEZiU1vHZ5S
ACpgtmuey8dgwzXqlo2wzWxzgmqoZZJhigfBR4HtmO784Lj7qP1CWQKvEpQmjDXZ+cZ45wx2hknt
4uNiu+OeEU8L7zg9nMKI0aJM7V0gz9RqaRWNFxICzYJOiHlXu7Jen7ipZCiFzcBnTHg2mW+fZ/O9
T/21K+URAfdIus6rmoLglNJLx47GXS5rgaXlVWmQMLzP+gPh8Bmo0f8ihZbLr3kX59i4vruEbI80
Ql7ryG/tDH4n8JYAmkaJUOERJXcznFDVU0i2OtTSQWMhqxFmtTtRR2uEwhs5dsOmmhL+J94X7XvQ
8EA2ZqGy0yow+Hd7ak6/ovvX1tZVn7Q+weNejgis7R82ZRgUIIN1Mox0cPGE8N3wh2XBEJduLIif
Ychzp5yV9Aiqxqh/yyWEzroVYPYs++/dtwFGUtWW49Fzt5SH+O0olhWIAWR68Lt4/6YQtoqFWby+
qyM8KIApv99QAM6E4KJpTYOuAUncPeHVO/FfAg3DR8YD9FK5IvSgzq2HqZkjTURpmNYUM++ruNaO
d294ePzReLKFJHTJyy2GjYSip96SMtl+C47/BiFQvCRiL5v/5vlnh5Q7PJcm6ZstDdst28LzEB2F
BLHXzfFHXxl8hxK3hO7tW5cL3xJLa5mUujT4CJaYHLCzk+lsRTq+JoBDcxKJ8V4FgL5/k/JChGAm
3I1EAdyDgG3Sulm92lgVGE6tEIviRjuLUvbRgHDswJ6V7Mjt0lA3NBi1y0EhYvqMk4RZ0kNigNgf
OxfsjeX9Wrsr8Z0JjaoLNkHReMOOn+4k/STZP0ARuzlhnb6wtkdbTi/lPKv0wSqvpvuK0z69HudC
ha5bIyfv0pbFXywOHxE1jooZsZs8pENPiEvPH0DYK6xmR5R4o45epVD9NBpNucQJEfMvrAd+UM8o
m+A0HCSVnTnqb3wjHYEP5frJjk07xRnE+puBsRiDgQ1Ugbc+lIGLSK981ajR+rrB8G6JyczK7kxO
Is+CHwyjv4/EqvT7npbLCFmw7E4VaH1u+JPKUmklPWYSiva9kntaAuQhSu/z7OVVdZsUQkxIataG
4QB+naCxXVFaz7xwrX4UvE9jD6tGukNdAni5o2z9V9NRKqOQUQKCLksplHcbGtmqiUTWcJ5dqM5z
4z9x0eamWrQtukolxK42lz9jGsF5VMTWidgXD6Ij3td3IGIplcvWCzT6JLA7l1wtHUuJf41q6yPX
l7SzN4iS452rHruj+T8goTbhyAixA+8TXyv98pcsJdAi+TaMmFmI4E8N4ujR9jH486otLni9G4Qq
FIu3+b+74ODl4014KPb29DJRtI+XMrSZVhDi4NHirYw+j3cyqvIgtZWNth+E8LmM0sgtPUDDGgXV
OgTUE3NWg1l4Jiavza7GJffbphxwcKvzXnaRomCzsI6MPJKToVIJoyl+6GXkfIOGfcL1Fui2lcpF
Dmv/+lICEiU1lBHlmebIXfoxIRK+0OuGMPRmyaSVZY1K4vS8smKG6y7cePaoHm7p29ZR0kgHiW2U
qywTuVoXG5py5YE2GlUhJlBu4tZsfXJ0hTTgqqsXnOFfB0xqv7IauK2Cy66Q1oO2a7dBy4rJXGhK
4my4DC0RnZx6PF+kh/7DQkI1GMfdpn6p7rlrtTxCxwClQVbCJoQCr+2Hhcpo1O8KjjWrLKMS4LZw
Z6mQmP4ZOEhG+jUSxxY7f6xflz8Uc4HEBTAGkzTA+3/YsqYIfY81p8qoWf8x65qlSgxinVLoPb8y
D6v35ujH+bebLvZFO6C8RTSDkFNFscITl+b2FyyEA4mbvQsJpckp6T6n+uOretaNAdtkt9rrx4o8
WGXM+p77JxeWl8WCnt88jUby2OPm36AUw43gLmud0JuZSKbUShPGUCH8s6LXxwz1tmDgk2CLnjfP
bliCroi+9wMlqs+PkPn9+nE1w7yGgLSG1OkapZCtsfzMAxg3x8dbswf8POvdlPpGOVjyMDjqRk8w
xFTc2X9CFgYaOkuxsNoXQlbzKcfzKn3JPNIo45/3rw2/a70E/USilrsVL2goaRqWFWCDuU3OfLYp
DJYFRAHvBDizymk7l3PzO8k32GjcHQvMKOhXMQMHKYKmeSE4Z6I55pzj+WFVAzx5APbhtp7pPbPn
WqA7rzJK4YZpP2AKwjrbOkkFTEQgL91quE8Sg9x+Cg2E1Hvybn7BCz0Tb+aKHR5ULIvj+NoUqBUf
UMLZLJbyv7VnrpptRujst3UiOmw+WxCCLE3sCfg4JlIinuB6VJ9byGf16r8MfsOgkhPgRAhBz/wv
squFPnl/o0tZF7McIW0c2I/3hq9dYMB+L6yAhyW/368ryxySx1liiZGvsTT1ylcxQum7y1XGm41Z
S5UeyHRfdrhpHs6s+O4jW0g0Gh6oIJffGuIqf0oZhAvAmzVUir98p6LEGvETKQ56tAZIZyz5bvru
KkQL2D+3dtLSQSRg7150+M8m+/L+X/EJZXHGchDxUFjApM+Jvc6xKPlLS7J1SquFguMArESX+elK
CX1a/EuMJPoOIOXEWr0PyPAvePxJz0G468li5VsNUOVcBa5a5ByCLTanxihSV64+vGp13/Te/z8z
jWrQsypiH5c38oODZz7OMWa0TFSbvsmhFMNz6xpe6wGPm2uSZVJRCPXzBpSYyr4bCB+/PV0wROJO
1SxQwGDbDNRolMkRbSfaEGSvL5uHHkHAJSBVPBewZz8RxlzftOZZzUiJSkw7R4SeAcDYXgyPlTxf
dJ8aBn/vQhgXxv/GPawe/7BGVblkR3yAWQ8q6MOFYgAU3++sj809VThSkMdI1Vgc3UYvs9nOUjqc
SoXiiT0lKiYA0F3/BNQYPxAYiMntgdR0EGn0WMUovuQx0TMHlcG05xcVgx8aTN+717enygq1n5nL
DvMNl4IUKo1GVYaovATZ1GMNV1a0/QaK/uSUEOypO+y76fl2dTtcm7cnBd6Ichj6+DY2ZHarilKH
CZuBsxu+YF1qKzxePg7scJI6khx1z9fKfAx0vRE5i7+HDLEDwzz9NXfj/1EbUownoQ14bYO8oRHM
V9QcoeMGhQumb+zW53dUUNxNM38kV7Igkhh4xngtqtwQVfjfMYwgSophQvJCDqo7FuHI7ZPm7QOb
mzxonYHoByp9PHN/L9zDZ80ElJrQwkAMvZpxPoSnpt5HqGkJjFSIMn/JhprqmWfYOhINP2bDnXVX
v5w6XsV4wLCFuKsfkvfykQzQ5kZr5CwN4nTT+IEtYr7OFwTRaWfcIFbacUuB6TH5HzyVLnHDhNnC
OrAj9Ly+m0F2BsfNEnSJ7oV09MRwfSk8K2AD/QrXnTqW1uQUn2srg0UXlmXB0mOIC0F/wjez/4+V
i9ZZExBjdM92xiBNGLU79eJBss2iy9XdDprVbVcWEGTswgh+Q08TemoAGiQmd/pvcJzkJ8Ll8kMs
hlH7ZC7o8Zoprs7FfHU5E2uMHM7st2VqlWO0XTViIesgI1nG8T9T7GYtgqe+5P9NkxUshS92kgu3
R5OaXha5rStDMUdDSQLiHfZAJ1bhjItUApLV/ntm8zX/xBaG6ZlZeQ+22s6MvDrvuPy0BpXK2MHq
NICSL338ZjGnsTnmBA3GcwLIwgQA8D7g0bpC6blOrBz9GG75HWZFPSZrMB0B7Gg7bMZSTPo4maLy
sVOwv49tJUiVZ9nM1PDY1EvcyhZ7SOzM+YZEMr9C/xNrKVgc9IztXnRd9+6L/s/nFn8JtxbqDAQx
ZPNZ4g4sXxlmui3mnI7lnELrwXACiqBF2MZctCSeI3JHSI2p42kjFbsrPxbYE4f33vikSSVY3vmX
hYwg/OXI3Xna8pXe2tY+t6t9RzUIa4G70JsFqRLfUAIwh+ypdsrHVUEZ1SRmrJ7la59HO0cjFjqU
Jm8Gmo6GOZ97mZm80iTkBcAf5naQ77G/gRMBcAfhBtWK7VAXDOf1e29/48s4PMFuQWZRu//NqOd0
6378Uwxhnv9UQB7yF4sfrleDfEHyqY0Czfl2KqYXxd4cgUs6QtacTa3VE0wWlY1fSz1SBq7MQVFW
/zj/a/yVitoiGpHGDcFfeLRnS/A9zvjbibA7/83yvlHURD51gLLsw4+jxBTgEazbN+8vtTgG/Ay0
5xvDEWiEdrkFiHrLLhkkbUSqnVyakULpYAns6QINNDkqldYlpJ/oui/kfI9oW3nPGCE70nnGD/3c
G2NQBR8OevC5UKZDHZHgBw98hGOp6xmy9ITR6IrZGmE4rxvjmUP4jhhB4bpV0TrZnvUcn61pA19f
G0sDV9ZElyUt87NRs7mvqod+ERIMDY5kwlCiYum8BKTMXu76j/gxgkTI4nURYzAM21WedVcrjR+9
86eY5j5LxEOxgLP2KgsDKcVIgPBNzeK1LdnpLm+CmZEKNiMjwUs1OxoI0sX9iXDgvSLtbztXboxd
K0Sp9H7O2ysvG+EYQf/Qhy03L8WNpSo0Sm9BrPldRpewv3kUDVzrnQqpyIZfvduooTBhU5Bt4Bfy
EfhhiatuH4+mKxtaca+hUh3yWEAlYDDHmee2j8pgRCMBrEpFK1tzWUA7hkX16nXiWbIljNfMpu8D
kKPbmxfPJyahiYKyXDrI7WV5+dZFsJ95U4M38COh1VmdE94Uitryzhd7hUMgUf0zL+q6JSmB8MU6
8uRTY2MO/aNNGHPWwshxykJV62nMa2yl99zL4xZwK7lSdyT4m816bkKvitu3r661yXqiCGdWOisY
74EpZnYCf2E3DPX38OI9V7JWUg7VT9nQpFX3sJbg9EHuPE1rrxZ+LQEijtuBIqg8usTQolFTeBDK
gv+bXcCq1674ahCgsd81x/gubunIFF1wCD2ad/E7f2y/z1mwdR0WYEspmWJ299OwRcsEd7sGrIDI
ULWGWXevGqK7OOQHEUBsfNYC2Z/wAMOQZV2PwTyC2GOXF1t/IcgP/W7YTQZ9iFLDTe7Tu3Ul+t8d
ipmAJrQ1MVyR13id6L/cBlSdzL1vMMvn49X/iK+4EX50BxGwZtpdgBRnCqBbNbPIvwL9HjC7MfAS
8rsh4CWldtM/mYyIdkDy2zlTJsOETJCFZL2C2sPW9VxWo2v16CVX8XaKdAvbp5Cy+1xhTbaIPSKm
69a9MZ01+oR5zWj8ByjKIGcH5lpoA6uUP4OfSEAuv91IxWnW3Mh5FmA2PBxOSRH+BMUGKPJCLmzI
uuNvaG1MrXJvI7D2Iz3EqZBXw6no86fmBWTQUHo0Vj2isttZDDjY+18HHUjPtA+sbCffsMp0CJmX
FuIK9V3oENTEiyNMvp7REfJOw6l2Eb562agz34mB72hMNOuYcEe++43j0xdszzhgJ9fGYVqAqDJM
WiEI0zB/oRA/eC7T3Em3/KGVddrAB0iucWRU9igrXWabQBYZoaPMXRlTW2Xbt+BWFUfiIlAuZylR
zra+o9+zuaGlH+NH+VxCdHIwDt3SLitlMjncVjH3na7Oqj/5sn2u3bQUCp2WNrS9De4jfk9xIPSf
P1d/JbiEKkRzpGG2YtLL/GtO/DC79SKG9kVljhz2KErLLduar98bGSPN9NCfQff9NqfpjWMRkO4E
dMttLE9t5o6iBzL73jNbppCGWqgcKgOAO63oT4UOyi/41xXg6EXrUeku5u+07jNuoYAowEG9Li8Z
7yDNpTftgllCn+pjkwz/5B3VREbfdhI6gCZJBXWvSAPAF5VvQFUzmY2gaoIs4gyef5gzQ8kKnGV8
BnZ2kypujnl9FQVlxQVumY+yKa//dF+FLWeCv2K/dgM3AdjG+08F+J0Soitvl4HjpPF5ad77CcCw
1mTEkB8f9anOUlhPJU6jhG4B6FTKgkp6CGLj6eR9TmxfR4AG1GDWuGDwbBT2sAbrGFpBO2IMfqSt
i7RiiS732whRsZ3XAOasFoYDlcPEGoOHRPqLEFXXz67EYpU2nadlfHhsn8ss/8HqfZPsjyqQDFO8
4dsiCDfPfyUDOsASucUOzjpLuwWCFIZhPXHwb0t4dqa6A0aXpNbVnzhweI2FCOFMqZqHBqoNYa3w
Qvnp7leP+04nPNkzKT5d7peEY9Zy+ftpPhLCyl2DkpJab7SeSJUJg4JU5Neh/7OYbna4gNPlm7yk
P8SJYLqz11W5u9HnZkR3RwArgzf6aCKuYxxMMRIMlUSLsiRZa5mEz77rhDfCoBLRg0nK90hpX5JX
1x2unbMeFpMWr4eE/1uOVySRuKsBoGgZmRPUhhzoMtyLh4c0xtLbejYJDEs6dan+8sMAK9966III
EfuKh/hECxruqxClf3DK3jXbL134yly+VXD07EriaPLrh19HJD9N/O4rqX0adIZVuvtR3DbIAyPr
vtL0+YhMVNtGLUOTKn3336Ws/9uMr2BI7n0a9BcVQU9rZhOEldeE0JNJCqjdhZxQoUZyjhwuo8lP
UQPW73dmxN2zCxuhJNX5+heFJ+9bK3jtpZelg7Y3KqJQLWf/GNH+bvihF6CgT664GHOc7O71cr0d
IkD1jVYZvDFA5is8avDFK2VvskvolI5CwLL9Op01+5pkiJBf9hYPJwN4l+sz2OlTjcyfPxfkL4oh
b7l6abfA0unn6WeTTShlU1ZM4qVCMvoFKgJbS6TeqP9YH4TA3BJygEPhdQ8V1k6jnKQZoARO3PMF
ib6azs2v/+qQfwWCOOdWcxL61NDKrWo8PGO1LKdTLAO9l2YBVnMdILTZNCxZDs+X63fgfWnbqiHb
Q/zsK8H4QQQ9mnb7KY8YPHOefxy4P+pE/8Xd/AVT36MFqJcCipNNLrhZWed/yq+pGcfVRa30I8jQ
Ok0jF+gCpScH+9jUHluF4O+LpyXQjkQDGiKr6IwKm7okWYRAKeoSAz6C+eojPJRqldmVYVdTRzzY
VOWDSrXMEFKvN2oq8yVw/TZrayLKg/yxZZkLWXr32i6HmaQhMR/2yyeoKOKJFUQrL7YaWZK4MqJ0
pzdfCU6ETF/b5uqvBQQKk6DcbvRKLvsSpNiyHRLfLEE5nCFV64pDaSs7DPDyjaPtWaNAgpsU4a0u
MM+1cW0nH6hyJhvZavL677Z4VQHIpkhHJyHi4z0PrQkwkalmrcvRa9zav5l4PAxcpquOsLyU9N46
09t5DLkZC1GKr+JLxmM+5d1eqtYFkzlhd6yqF255sLunetC1KzyOJ9/DwV9fI1pMS/p8qbrpMgg/
2bJ3gdk9OXDKlOqLiQPjtNFwk4MvhBaENDfFzrBjsB5JjLzUPyToFT/jbD0peozstdTn2i/absm8
gc6Z5zq6OoZ+jfBROr2cRswzK505C7zqEm/bzFJTCWzaM0qi5vNg/p0sQKFjPA/eLrwiSWSjrPyJ
exfhMQ3k3bpQvLvgz/zvnR0c1LOEWYY38SiAwWdtjcWdO0iMcsXTjzoRPlKeDWlDWDbZzuIUOz5f
k7sA4uPO17uYGD2Z5HwEFVUV7WpXKNgt7QDSyCLpXkicJkb7bK2CIgBNQY/5l+TbtLdlTS3HteqX
3YJJqH9f3MHnAKPHV+lt5P37h7FdaLg/XMHTA130HuyemX7IQDMOzYmcqQ1LEoS5o884/Rcd2Oao
zWWi/69+uy/RIFKTGP7ulnF2ecwvTcQ2W1xvlZU1x0fIrsy70pDXhjjp3a74an9vrca509v0GU2I
KgoVLbJzBr7btefIIxtpcamcOXfCeGrMBGL3/P8oQoMh/Sif0w4iavoAyUC8ZsNrc3bCi9CkfedW
soDLkf+4aB8Kr2uGEs54bMvJ/3oEoNHhr3XQWykIEfL+D0R4QHnHq9FwvcqgdBHszNOjIWaVf2v4
wEMBZczPpOxXB7lgc89kjnzEZdfLUkEnhxvUan9KYSz0m8P6rrdhXDulzwtV/Ej/GRZPNg3bglMV
bTg07rBkz/IH/JmVhoqSGNCRmTbHyPKUQbiwvC1po7cOdbezkO499EBtNq8I3UI/NUz/TtWkpFBZ
FbHaBBHDOlouR/OLx5rLXQ8opRRB3HKV2xqtVYV8IZ/SWE0doFGBCkA5EDESDLYGH07mxeY88K0Q
NXKu0Ivz7DHHQIXaEgCmlH+Q4c6HfEovKRWXXrpaAwtpbhJ/NOn6tt6InUg4l+XXba1l2CFmwNpq
bbi1hLeiiVKgFrAolTPp894m/5Hgk+jSWvh5oh9C11LwgHK1fxJmDEVE4Xr+nVkNMw2EtZKLhawi
CxbUOSt9YyTCB8JT458Rrh1jX4SZANhXeteG+xxXL//FyNQ8SeHTikaK8bJ005rb3q8Z40cRT2AE
WwoiNZmcy6oiOp2rvNZvulhMo6j0QurPLLKuPLmCM3BR4xGScy6FQF/gEv8gdPo2E+YMqI3zMH35
nc/WJPIiJxZQjh+HHtEwwm2pibCCmU8414zRVTUND91OCDY0IkILBNyL7ax+GdDEU8tcMzI7JyhN
my0tWjpJxHi5DD1Met77Ol+cMPZoOewUnPMQY2k4swaXxszmcaVzuXD/32j2I0AxT+KVX8EjZRkt
I5dXvge1e7bCUY5HoCcu4QTgmxYr0GzcjyV3kdNinM5pjiumTAhyTe2LPZXfLMrWVKIfCCOcBsBZ
9XPc/f5IDoC9Upw8GbZ/Ot988Z6FTODzklIMKTEwNRZADEzHmMqEsMBJfnAkvA6549QSYDfGrnhY
3XSJ+rGJc9bv73jxzqs1BTKGxBaEubt7scEZZSaoLtaRD7tLz83JJXSB6bRBDL2Hpi+HnJpjFn+B
feN9/o0i9m5TYO9LcUjj+QXUB36JijPGl0ZXv+Op+3eRWk+Bxe4HWcFm4P5CZELL+zB1rHLYFwj7
odkZZV24ARfiYsRITUe+odmFTan4ZV4MrPQbOF/KH3hcYFXzZF2lpkxDaP3f0uA6JN0m/9FNJGjx
EAOfovxxs4c9gCBzmdC6lKdpSqBgcb2GvLOJrYr44hw13PrRBffB9hfBO2ZrjuuDsuJPlOO9S5pp
WKCntWimr3MoCGWSdQ0tps6BB/xHUu/tH5JWDSn079YGtz8kxZY1vslON35aTgprC36rKWs/Vqs2
udHrYl3bN/EI3dgpQDC1AlFjgaQQ1kyu9HVEqAdz9tar5ww+I89U7BKmAmrhA7kDOVWgdBlftri5
x47am4PqLHbmE1OWBjXsYEmUBISD1fb5EqhFQMOv2E86EUIZ/aQ14veZFvGAmxmGSiqtomkpzXer
zSjddPoeYzfLkW/M1rqgPCz4sJ+bA9+R6JSE/uRO7d7nujUbpW0UhtQ+Ce9i9vgbgECRCfJHsPfn
YqLA5XE2Q7npQrPSb/Jb6HNGzLcUVS5ADp9cTBXFQmyRmt7X7nd6QvgTivsKUzOFIS2MJe47OjZc
u0XKskx3r+rqWbPEPS7RiUk+Njl+1YSVLcNzxItuAUoLbsKGdXKESolY5vQAdnzTT+yw34hDKj0Y
Kjz2k9WOB8UHdDRn69yOanFs8FzhBhMnmk+9Cte+Bpto53pkCjnuAIUMS9xeGwemsQFC+9NEIvbH
/ieCtYoDek5M39A28OcfCCeOsZwu0EgcNPKY35pON3FcWRFbhE/cOD4sV2RJnLCVScIFlzxq/l+9
lw0eUl1B9WqPFAlGwYK8ABDKOj7MWu17SnLgB++n7worsqm3fPYkJncGGAJA9nk06kE2hK46E7t5
2QTSND95Qp8Vyn8yuTVR8frmD4yb7c5csDdm9hFOViC7uY2JGy/PZAT9xfC1exW9MLRqHFis13Yz
HYgivSA2dXl2SVaKWHUnmHcPxmSppQ/2RJWyzngvPGm4HNAMlbHNGWMoDmRTmz1jxu4cHjb/RZte
2SwjsOVCyTK0TNeme+fttIbNkcuxUXp4g7oax7eT9X3+dj9YxEoj8ed2tFMOZqOZcf8saOx+zBUY
CDT4lREiQLfNJfSGruHnsy5FIlO7gwxHYOWmxiaD5pkO6ec7XBUtrQ7ge0q0u7cvCKZ2iyAE4r4c
y3lWcQgl4uHhANv8sF9KR4PJcbIKX0Ialffbf7Xvz+xenqQJnQZZ7rWpn5F50PQXYWB2er5fc8ua
BHM5AWBCJsQDfhmenBytYQBwMZiuPvkU252og7/pDmjfP4CNslgeM23QkrH3Rf+4g7Cq37tgrv9F
HACO3H2vJ+SMXdgXKq3Kvh0l/aP6zNUSMvL3HlMTZ4AIwab1Pl22LnpUgvAbO8RJAi/yh6lS69ZP
Qv9tiLbrp+1A47LiK23PFaaCZG/PpaLcUWRfYabuLkr/4fhiX3qOSrtfeJdETZqfOqX1VqoDpwBQ
haY+Up1+VuYssPgPIybdFhKqaQWFeycs5d5Ombzn1pTkpuQk4I4+OTgGGeP2DcQdStJ5d8xoopXF
rgnpkd9SWynllMeV2m5ivat6erzE3zghIvFUgROzzIlPjhmHLspl69++toc1wGWc3Nq9K5xydipA
zjidYFYqPk/0Sh2UficmW/z+CYktv9xaGwH6gwY2Tkyo+lliLX+66oeiNH20GDcyOHeR3Gk4UEOD
TR1UGKV+LCmW3N68COzjTHjmG8hV87gftASVWpZycYx/xfp73WBmGM7rBP4yOo2VvMI4SUKfd8rX
2eQVDc9q8TGO+Qtn9ABt+RKzH+om7CMwhpWUZa00CcE9zB8cVAAFWoDLxGVgBNh/LoGWzeBMbEbN
KMf2OLVD+G5/bjDwAFZ7H6av6s+BCEab2Fd7Jt8kT9IWugJ/RiWbqmk3a8o7vdkIexat48PaTR8w
KkhtyiOJarSkRQC6XmO3XLbBYkW7d/4vJK5NTCwE5MBrLUIQGdVpFWBZ1huKOEaqJOrY+gn8G+qP
h55VMy+xZIEhDkP1rZeoyKjdvVC68prHhPGsVVADx4IyN2zIEY0v6bc46PRP6VPyc5URb/+uas6X
4065x7yUg2Ukp4U29UW/HdAxNmZfNlKa4xrGiwiKAEiuNI8iTzH/QWxZ1NY3nUzBaaYcKOWPB/A+
DQzdUbTMIsO+NF514AgHswQzkAGl9xhMdMbGZCeQ5WvLF23WJLZ3a3eBMLxEoCMpNc/sfPvSq1Gk
nzIibrvnpcu3t5BlwLKS6NtzCMtuF/sBIcJ/hvwUB+BX6rorKqNFi2438hR0NRt9yoACQbB7ZqpC
lMUsl2etCK947SnD2XOu2tOs1HYiH1qF9+jLeFXgUMi73be5rHR7dubqAb4I+CX0/y0sgFtZFICT
D/2nzVMaM7b9+r875VHMMm79uXPJ1Btar5UmrN4+151grDqUCPKsAJ0GdiHBfthweWE5dNRPOtLq
jLLnrMezKkazdRsdTDF9f8w9BAk/uPoCyEcKpwIsLMq4O1VRHYplTatwVBUc58EepocPp6K1Hgdx
L0JadS+e3EfNRRDkg7QvA5jsdgJTUCL4jdHMX15WUAg8vPvqmrLKw7P3FPJL/Aj4xbMKruMK3syC
dLxNFfKaFSo4bU82oQFTy9ProsmLggelRatZKzlPJLfe9PCKdAmc63UbE3MaKC1EH677caB+1zOG
iO5rs3r+tLqu0lZuHNg7xGAx9Kl5JX7C5dxqw5LnId+TMCDex/1MSclyyaFACjln/rXOWwGde0Os
AqxQz9uuuExlqJpqTKEOh7+A6byiJKxPBYvpNnS9nGr3lcNvcwFwlWFUQu2MS365oUHHGdelHy/v
jeN0zPvu6xYlP8Dos1DWM/m0BTzGf5cBcNlphPLYqY7v2gDfkTo33qKUFf5r3mSbEo2cD4izy8eS
JZp9HGRNgilvIxnSEqkKZaVulJPo1wW9TBPr+XOditnKUpYVQ3fsWKB6rH75iXvMvqJqrjC1s0Ny
uZ8M89kS57xLaIvLSgCDZWSxcGsNd+m8ddRKB7e2ZJnuGs3bv7f+PWPEAPE0rexuzBdUxiTIarpL
3tMucYdowicEZbtoufPBOgqzg22rDadu2bAYUMRMGDojcItx8sktsrKve/dK/ffI+52N9KKykdSu
12AYAVIXflVBgw9rWbzUDbbeRYpH3lGvKYRfTTLE3kOEL7ELsGAZui5qCTX4K251WyIyeCQPiKeD
jSPLVOeVnAoQixgfl51PBbzC4beZaGnkhcmXuGBBnXQV7JluJOMojTH6TqrW/kCgbRM6JB5hKZOs
HtGeMIFGTiETiPY/BAvvJ7Sn2uXw0Cm1SGdEwPk9/brmphxBOQUrVBPxnyuZ/hT0pxVHMt8UHUcx
EPVEBxUG7sT4kWkgkZ/sE0zDHveECEMaC6Y+enGD78LcVe1i8w9YyXCdcU+jRwRVsw0HRAx+y3br
KRWb7e4sDnHx0KNl3HJP1b7ze9Kq+AMl7iRcHpbT2XCYRn2DIiO5WQ9YMzSuW6evRE0ygurxQb5F
US94SU/+D+cEj8WPkc3yeJc+RmK2Ir60emIEgyKgYRTuIBFEIcu+k6GJ52o6/Rg5oIwmF6wE+7kV
F65zfblDSCNyTskAG0lzfRUmLf7uBUGXh4Rl/SuZjIV4TfOP791jdEv/zAnzu2/VPU5y9yYBQZpk
dUUTdUSNaPaRkn9Gp0M/a6K4dAzXLxfQrCCat1hVRLEgvePpcgIyvFrsjS0FeGsFG0VdJoRCJB5J
tiyHVHsCxtwV9tKATnKXm3wBkmAiJ9WZ1DBgjw6UD+izrn8GH8JYE7pfl7IioVtXRwA+USzdHdkQ
H+EdJwKj8KPfAPWuh6ZGdmNX/Vmh1BVuxlb3mDB7OxUdVNVP/4o7LxP7oHl0H+Puy4swLXU1S001
IBTMlqd+5+XBivRjUMtYo7p0k92Yo6LPMLdW9nFj2zjq2epgacDIKvDPjxUC87m8ulgNis05iWTb
BieTrbtZj+lJI1E8+elp3G6ouQnItS+U8D1Zlr/nxCKkaOYqO6zoy1LdyW+sZuLVtcq4IuUkWQzT
60H2j59gOCnlb8sr2Ynu+I9RFTD07xNcvlM72VhTPxq4omKdGdKXGUGcYWLNIlBZSaQyncgeW3dF
uDs6cSNOVaIdLbM3gsx1oXXk4Eqcgv9QMCuk7DsKhtrapnrKYLqUHO2FDpgi2a7/yONFJ/BBGFBy
Rc5CYJn3XfZpJVZP/LRADAmFEfSpr++Ig1Q1Z2XOaJ8P+OWm1iuwmvl53JVC5E62jjqaO4f4qacu
HoWweCBxzFNlP6I+8wHGeTOljx7jFuK2wkua9gVfLRf/mAWEQV8P/H9BY4xwYuY7cme5tsfnTcfN
1MYzJW0g5mQNEmXwJydTfz0BLzIsK3HhM/oc7u3AJOySU+HQiiBy4RYU6l3fn/woYU74Ri2LjcXC
1SuX7vm6kRXRQGnlp2WFqOffYptqHlR6CMesHGzeCA5vwgbNAMuXgwWe3A9Tt1H/t7vb2SWp1U64
pv3MyGzw8XNb8BETYdSbdimVx5nKUPrJ+zOb8HymGgt4bUFjOkGNrKR1SYKo6sd7MwNFnlISUH6+
y48giFcMAarmbgl/Zev+1ypFT671QqNpeFdXipsJx9NAo+7bQcdGsMW4fZQnBzjkVy0EhzVdL4+C
8fZgH1VEYzG5wLGfjNfTdJEQraykv6ytDzhVP7+SCC9LPWUY0rVI5z56jV3Pw/DGzy39LYr6myUb
tjdIjJX3uGR0J68C1OJgTNwnUfs81LOR+P1QNsMVM/qKiVIDbaXdASSVWi6vkyUCtp8ffgcqLMFz
rzaQK44AOh4+ZuG4lXFR5FIXdybo0jGj4ak12MxFJxGbTkmfLOMkPFZkEEZuFMhXtEKD571v2NCQ
0aUm9r1pGY7V9egoclcQUa+qkf1LiI7iPVIxoiksDETKoJphY7Bz6OQ6w4wvylgjk5v2XKUAS+62
zLoR1vy0O7utKw06yTvzo00MTFsEAglPtv0a3G04OpZkm2yLaq+4xAUsB5F7YJeEkhdp9NQdwxAO
fTtsltGe3+N0/inOTRO0shVCQ4UjdQPtN421kmXM4ihj0TVQr9WFYtZTzWrWV11TPooh7U90uDM3
HIEv3zmOiwoXLSTHoVRL5qWu9mZr3Z/FIVypVdB2sTByjHRfQaQLD8cd2xtlFwbGD2UCOs2bg935
3k5+XViFaFVi3P/f+KaCkbhF5XapBRo+c4+j+4DI+KoIYnG+20As8TH+tcmyKn9io69+tu7zlbGq
Z7FYPUlT7FXYWSYHgtyXIHyll/1NfZDI9Y02Zk2zB5lje9nYhm2bQetndzyj6OI/8Pnbz6Mlmv0t
HApOCwF8zQumuXHINhRsD/YN2JeAKBQEMYiMOyIcuUCsOif2doKPCCxgCaV9LSkGO+F8rTa/1ahi
e+gYkbsmsyZdD4JPUNosQBYAw0idKoIjP9zyivZIV9H83TotEvG6EDWnZ+6Awm0+n8NtLfZk/Mgd
PzZ74YFfWiigUc/rvrdwkuJ10bhI3CI+Syrdz4hfBgNYkCNJh6dM4Qde8K7nqzbstn9vOh8QvSLp
TnL+JoyXyf64gSrCKe4GnPMOknCuXIXBBFkVWEcPt8HJTplk0W7db6doLYR3BTebrCYtHYtRI5kH
P39DiJWppXCdgceQLu1mvXUOJtEBedHDsOzAO+CGaMO72Kb4DnhW+w27dRikzrrWSCPN3+02ZPNe
p12+L41gHabZDCvHWgq5HhmJxJtgP/DawWc4sp2yw1NR0R9IRvzih+TZQS982fywj6cIri9r8Aew
0M1A0x4GGbx73c9R0pLeL1OBZWmdUCAh6ILBcxeF8XfzBiuMZxXuq3b99XDQhq768wutYFjB4gXq
RsyePaGS19TNPRv7UqYaBld9tyRC4Jp7HzWd6H665m4eV1L4PX8w3dDDplDQ4dbWg8YLOC3zeh44
u+c16nNLmEbiIUqhuPHIyWbMkCybnYCPPtoFNbO9BdGHqscJUAXAg/KP/hg2tAaAVRH8rqJiZePs
M+jR9rWib40NchKlfE8ZnAyc0S4Ii9GA0MKZD6Wd+7DQlIpfQfPSvNhuS3pIErUfWBGgRhV8JwS4
uXeNcuO4TbeIkJAr2XMaXHr87lXl3O/aGhufaVXPfhVZyFFQp+NkPFc3hiJ6UolD3Q8p4E57oy27
N8vVH923w0xsVWmxhbZwjMR5XAqrj9836OQMzMZMVx8aoL8rRl1iAxQ/B+ebUrMsqYFUtWZScEae
MR3CSGVgG0L2LHJSAHevGXuX9dLZ22vvBBxyLSQaTsSFky7O/3lGiBa19pPxCAojxzufZ764+cGV
mT+8neiWVG/bDvWYT8LZwWo/6/wU2XX/fPDIEJQ65FHSzVzAg933ItCnCNOKH8U8WW9NK++bJtZC
UdUp0bQM4a72HvVxQqjPccaAUOV8uzaa6keLrK7ZnMzwJkJ7V7xykuU8NUnTY0u8Vquw1hcFNhYA
Ahvmprn841BBlM56aJYg0/T0PaR6kj7t9xF4V5yzKl4izC0/RvltoD/nsrJia9n93/Vfh6KCXC5W
VK5Q/odap7uw+Ozftgl9/omBcw91ZNvU1/aIhZUVKFoP8V8jQc2AivaY/7mCE4Kxwg2qHqW/CiMw
nbN8BPtZphJVCM5Ab9v8yk5E+VEXLgc6coFSD1PmUHvIpLPzPzVLl1n3r290E57S8uMbVwrj0LV5
Penwxv+e+TADLfCy+VBaUoSLsab4IA8amtsgzyLPFIrDGxRXlXX9F48dr7RNQvGwwUlZHyrPGAfg
mVjE9YMufpc0nhl4GGxFphnNJAGtFdpWgLtLEZ26OMwNkQ9FD0LOdnMP/KP/IaeSkL7Mg5nXOY4w
VUblHxWng7e+23LzkbqAkLd88IhsVGp4j0WPGReyatQzPYMkcxDQckI2AZM525LtUT9K06ETcDZZ
dyBtnvjRIRc/z2tP66wSytpsiMAtZIcUGX/S3Sp/sTbPezjHxQhyHddklOJJiCgU+lu4AlMiJ9l6
F8nLxfjBTQinFr4ERLC/2zOincOm7S4v+X1+xkb10x270R6weCw95Meuw/d5cGr7DXunr+MRYbjQ
I4Bn+s7TqtLiyG61zocX6L9OodLOs+pIPhexnVN3wEA+8/5ZU1WSqiGY3oH5RRn1PZpOHcDdrUmO
EEmSOmFoSO3vTZYQqNtCyMLUB/0OPfz5JerQfWl1UAh122ZGBtZ3q7bSoiphXgV4nWOSglhFDFKX
p/Ta/g4PJxnjjSFrkrI10xF5o9pdFU+AO3v+xpj6BRazClM+4LD1mF1JiCz4a9svY0YpFpaFKDgl
wUo7uRFhvFwVMZrrBT7beEaSvuAvBkw+mz/g7+aA0TWEInS5zfwwnJVj/imWELdTuZF+coQhBtWZ
UFhPVQ9F4IT07NSp1LgdjR+iLpQMrHUA2HVr9myaBW4R/QMzz8pSjO162bFKD9NU6be2JDXIrYRt
uHUB8ksQfoqna260FJXEpqIX5GsSCA+IUiS9dCBoo924v0+WYVbYnVQNzGG8jK6WBt/rCHuxtmkq
3SXQ1ZwLVvsEkwmobRfJJ+hLsepVEoFn18Z2+U1rUd8SRqcd5unYY3+7Ss5Vi0xnIPmpSgbWOGrN
QUSevRUJvOqRjUAeE/kVBuP/5sdId9I6gaJpODLhae9CBCFSR7qJMyqTMKGVns8kZ9IXUOCHyRhX
SzC8N5shtxQDaeIbIX6Zgz2T0SAKz43186rMcv+MeWDAd9qMEZaed6M9qLJbZGi4t0yknSOdEdfz
muJ0D53BekyDZkpvcPca1X4xYuIV8+/Ih2stTwe/fepc/4rBuVrtmzXCQTMoPok2Tt84AZw9gy+c
zeytA0I2ui+DV/TsgWkNhSuHqwroLe4+wjStlD+ADuxgXRq6O+ydpQGLuUiHIghlGqKa4kLaaiaJ
6okZAaPUXinXWuM3BPbsWF5vzPdU4/rhF8lVXbmoUWHkfSAez5oJnOJN7+W01/tWKn1GazwB3BoE
QTLrA8frR1IJH/4OX99/mF/UmNwVeMM2wQ8/1+oOkjxY+ILwXMdwREeRJXAMVqhAOVk7v2ono6JU
PXdVWrBstXBxnZydVxzSq4M/ZYia5ojNYszo775pU1hZK95gZ2Gs6dJJvSLWmnkr17psO1Hc10gT
z40T9OaUXuubeBYuo9dQzRukOS6QTC4zYz1KBh9zQx9Kt4HH0xvlq1oG6JAO1N/WWcDOyTCMJ+mk
/dTxrme8qup+ZI0S9L3uuvwKymuICQXIVRVZ1kDiKOauHJfwm2iSqU/E0sIINB/UAVyaMTGq+g0o
0jZ3/XiCPVVl6xJABNRyEfOHEB2WhfxEL5YTufQ9fuOMyT569zjtz6SbpBadBLIL5chOt746dAal
RMO+QZXIikz3/cX9xN0H6EDBT8YxSrIRXHcplVNYgqCd+HIFTD4RWCEmz2QWlLwCfDHG2eo+/cMJ
/ZHYVqpAc8SKkK0hdde9kvFs3R9ywXCI4T4aTeHohVFb+tWq8Y+1UWdroy1hbF+XYzfJ4mdc/c1f
PSTJL5Nr+1c4efIcIAcYDjHDT77zkoz7JV1RVQ/cnE7QSYCOnfKMMKKA6gT9Xq0l1XafQZ776omH
ry9tgW3gtLOABNItI1dBhytJn+u4QC19FHXMagSDNH8xoZw4fIEF1cExMkyT2l7Rrb6yv2YzxMhO
PNYxkApFFUcZ28I8GlcjpvEJ7mJjbAVXn+d7f+++5I27S0HTYKkHPdag5YGs+6xmhIxkNxPGIKQ6
JJjaOOujDhHPf70+7iEijpp6HkEMS6MDHV5eI1gPLH17QDDJJXJrHgO3+TzI3PUG7lqR6qCQt2Ct
PeMFIiKTXEEnUjztlWcViC9Dt13pKEfbWPFGVYW+mKlQYRlj2YSSLNp6YtEkqZQnps90kRGFfKHZ
tYnwB7wW5zqC0U1lr0gXsJK07UZ6QtvF5f9lfo9oW30EWfyCl4kfziHiU+ojZPeu5zN0yWiAk8Wr
Dek35lBwXX4rRMQpLutqXaes9+LfZyQJhb7JSPT1NdiRQVvyBvw6wVxPwRccP/Ux+0K0Om6/EZIj
0KmphklxqUbGc3r9noAeCeRuLE+bO4aBcENTQe94g1ROvmmPuSP/Bf0f1/XYokXzdeIg3FbyYguy
cLZPEEPnp3iWLOzypfJURHgzJGgH18bXv4hHuS08ZF1seOPmTNkOx90WR0EO4BNjnOWqLS35k2KQ
zmLouxd/9F+gFNLBs2YUaJ/20fwaYSVLdpnnPfyZ9B786G40unAgNbw7JU8uH44k5ApvdtzbNMm1
5kSbBblbMKtkS+mvvXZhr28qSbcXV9xURwPIzktK24mBiCTxAhbdt+RlBr5cBeY7X8Q3Pe3s+fhJ
AYxmMVw44aKau7vgpPZ3jxxCn1snUtNmx29A4c7QHLHxWUjAUaPy3BQJYYyGqXgb1h4En5GD99YZ
Fa+/o3ZOlQWXWE8gtjNSQCo9toNZFKObf5kQJnRpU2Q0UyscIpzzi51j3dxL6s+Om1ffYen2HE8N
uJMVpw4kuRTl18YB7DyDHrw9tLaumPjPp2EUdfqxnVLtbCVw72ipmf21IiHRd0/2EjepezIm+hd6
tkz3TJQncodsYU367XLMwAtZCHUZEOujCZudovW29erenmJ3YWhLOfwJRHyx/cToIK09PlwiFtzW
LgDBaB5/nobvu7PCH/w8mZ7R+hmFx6+jtyoOQqqIJ6n1mzwlQY2y3BIeV/e0xFuUGBaWT8XlEYS3
0CKejAmzY+yMQ+pH2hZ+6+klHfi3oBo/hSAWbVCtR0bp38FZWYrq+m6KymnznbBN6ZrPMhxbq14i
6sXfgwEK9RH+wLgjCvCdz4LG4lkqgxMLf96AOGYCS29tNIEP2sFY//hL/vTnrkug+5PgI4YkJFGJ
V/yICVpK84bXADHblGJysodH5njN7GgzGfd3Y3kz8ZjE/WqgXfpo7r5yJ37zp7VW0fH84UC81bZK
TPy0xaDR8oMlmi3/PvE2N3GhkRCxSerpuESCD9JyTYjASucCUHpjEFkwi2Hw6FyRKyGgr6HglPM8
dy3FORu3YmxWUHYcE9e2zMnOruxYpj+n8VJ/fUVXvSkEcaIW9hc8stHZ/ZFd6yHiUJBPucX08wPg
M/x8IfAPv3g3xXqE5j2lGEf80rMkHHF32fhY2NoV1ck9hJC/TIzR5nPA4w26PpYQEcUh7F7QmWti
m8MPBGsRBkXtkWf+g6ETPsnuzzPc0p6gy7ZJJ+d6BrYTPvXVsOgE6R3MeLvIXkWmoYekfYG5fNiA
9yqplmZT+J9X7weRgvr/+aXKTmpHXx6LKxzfNgXXlbdwK6BlVIQunYtk3TUo4BsfPw7oqmRYfkMT
tESWmawWuv9MvE7SET2Dj39XTVwZRYFcVm9PdYCGtYU4ZgfBBhCNSLj0xne2J81k5stc+90+9vb6
W0tdNFlNWOMXuMz/PFcsBcfCD1KsooDfZlnujgnBQQAJeNPGpvv2uN30JLd26/H+jiPCXCk3Pdwr
oUhLf+WXVzV1WpD1YerlnsYlms4WIbyv+vss0jxiViFmIGmH7DB3KrK+w43LcxuO5iry1a+lxvDX
myd3csw5/rREsP7RYWVZr4nhtNAzOC6oknloVTCQdRg67KIqbr3g9vhKzl1yEoMpjjeq180kyFD8
vp+VVscgv9KBixEEotE9+FZFWuJjwbAMmsp8pTQdT5yU1UlAhAbL08VkOidQhIwVAjBb+YCDtZtx
mfb9Ps60AupQmrU7todE4uWUaHdtsWSDktBzIB255d9+rlQD9yX1ftZZMQ/SIez0x49SDzoO4BwR
/cvJFPsD3K1ePHh8pbTSH4jtja1sOGmg2LQeao2RdnI5ZJr61sW+G1dcC79hhyPhl7CbVyBUEkmw
F0VCAKmmG6jy7Ek+UrxM1QMmDA6kL5WAYY6z38V6b3VGVVh0VGIy+6mBmv6so4J+SKeOS2n6ZikI
dfODZ0mMB1OG9gkMYvWi5ETeRScva0GuAmppZ5jwRlpyqTk3CPS3y1tp9G00nYz4BMS7en9mx0/q
dyuSB/2xKkBWn3To2pLt77QWhySH5+8cP7dVGgeoW8mL9dGrLdGuOBK/JiJyz8aHAG//q93zTKS6
nSZwRNlOMVk4iFAe/Lu3Y5zoCNti1ejNZQnaQ7BBFyGochxRtrH4bP91ewRfOYI4PibAlbxIQ0PQ
nplgP4pLUwzS4afjbq+OVL9IUw3+dYHBilsUlNokJt6LHxaHoIkxSitkYaNvzHT93CUW4acLtF8D
0Di2koUAX+ESw2OAIAdQ6FRpRy+fhmEF913bEetJHk7y5DbVzaij0o3j28QFHt0h63HT7uh4/kg/
2sz7catRFY4LKfoOfcEiK0t0QZjV4nj+Xp5SlLpQKI+xopl6hBnNkYbNoh7XceQ0m8EZ45entxQK
CntakBr/6y1+kuDS4CawalQXKYy3J/2+WON5dObn1dhML5DJ9+nMij/hhbiu7jPPe5vFrCsF1GJc
ox4hZJTNA4YA+U68CG5H+m9TiKtQk/UzzIXWLwoN66j8R05bdxRI8oaXEKCguQl3tHVAqr1UyVYL
b28PHEn5u8+IFZbu0Agj471DHCxd+GhI9vZajhiqkyQbynFFCuGi3QJkXgkM3mjZGesDPermg4WF
bethkYNsTSb6EuV79W75sCqp9RMeuBAp/vAPBsLNpTsygXISTMGd+rYy3bMpsghrsg5o1ggsYzXv
Pf0nS5LonKLz7dNsb12AvbFzwj/yP4imoVpFAi01sFl4Z7nY4WniaEp213rglxtco8WmZrslOPHQ
2ho0GsD59u1kArvMpxUOH+MvZCyZoEL+QxwEZtrpJzONE/oJ5bAxfYgGzwHoFdhjQ/LZdAfXCSc/
594ZtkS0GmJBGHF6BJh9T7/X1qM5ttnmi3R+wC0bajwQbPCBst1YDBQ8GD+XfFiWbMfrea7YVZpd
kLem9P9vI6ZkcLiSPEH40KeCgFz3PjbYYvgfyYpSChMtNY9WDHFnhC8VyV+nbkqsGjSK8zKVZ7Bu
27d/Lrc8oavi8/uFgM5OISFC7rmqn2vtIKd0dsUcwobHNLNXH+9CfFRYzvVhUfNz4Ua1hPhdOpnm
OmYnghnmmohoeQjN0Nd0o1gC7RMpNFf1J1k3h7/vfQ4ifPFIpwJihd3unInp1vQYiadZWf2YF6sK
l/579wvjI5WZAqqxWRkP0OsdRp1Za/U9Dv58Kw8wtAqLn00/PNw2MBLfhVe61loXKKBmtiOntLaQ
Aj0w5YSnNQzgpXFyimBdAVJ2OkGGilHj2lVCJQorE1Y2aanGTABrgXgY7cHolWB/xZx2cNGSP6H8
OxcBrNAUNlz8skHkXHAUlAbpRhZoUbBCiBq4e4JhWMo9Zx75BXBUblWsvEDIVSZ6X1SLkgaao/cM
BpkTQ8INNTt7pkqrQeXB/ZYyuy3Ph1pzbF+kMjgtpnX++2gBqxKqLxJ7wHDrTRHLGsUv/Mxhm9Vv
BRUyLgzcrjVxvt8Yu4KD3ycTvmZzmKrMiHdZJiGYURWs8EaTN6e36yyxwE+kqI0xCywNUMKd/Lh2
UD+t1ijLPzpzD3rYNkztUui1bxKiTh/X0bZoD4lyvS/y0RjQFhydZsW9c+zXtLp+iFYVVt41a4wD
QgYGx7srb29kLjcjMUDul6pdZSSxbaLdTwr70VAuKfioUEoPRFP/Q8Q992ZT3ttffS4Mxl0cJ5xC
L29Pi548N+XdQTSVMsZiFsYq5w6FnrQsXmsLXlPmuzwvbAeLST3DP7aMMYLvKJ06AEpnGn0ioVmL
dTbTk2Ul6dtubLcWgckRMu342WSWzyZwHsf4Va/h2aPszAVaBXDTIlw6BCwsp7edvIsamll0GCy7
uPgiLxSQXXYRi2e3+x3cLjCh0CcdOw+tc4Y4hxB5CWAXBFY/IqFdtXlIevNx1kkx5LSizPIyLMMW
O+meEX8Qu3RgFBFkbsaG1/dv7lwEboUAxnAv4MXFqUOmpXdIZDYNO2l9j+w9DcFrPTHQ6bucaBlO
CjvHDfaeek37vFUwxGPIeE+9nuhc7tKT4MBkYRgGAFS8NeoqoFk4G/yDlcSnPJK5RkjD8CJmjrRe
k6SRznYxYMoN1WZ253PMjRPTJdeLAjcjM0fX9kI1E7VNaLs8ILJq+jz2VKpNNzw0fBoaVXxBHqKM
eWXw57J2brNxm6GQ6wbV6W11l8LzZSwzrZjyaDY2d+y5y9HzrE8LCCW2Bnr0eDsffWkjFk6Z3/+E
3D7HH/URt7TueTCJoDNx6QFsYysG18tfGRCkAwkxvCFpnb2WmGyZMihy6Ay34scxrSPkyoNn6ZPS
qS0febjkczFPBXa65kh8DEfO5u9aZlj/GnI4LDzARGOG2Zfyw/dy4yblImtblfgAFpXtY4n5B+rN
zQJim/a38/mNRdtWxscK3EIFB6xQ/OK/cYOR1IuyHlHFpjYBCTBWEtom0VqnPer0gV4LdWbEDvfa
NGy1A/dukQiZ1dEvUzZAf8BDJbVO0EWg2bWXPVzTVdNI66VvL9ghcXP+I2a5BwUdxqGQc1yw0kBA
CfNokvk0R+IbBkjhlmUzvdZhGt63k0BGuf5TqslK8372gSG+fQl1WqcY/VuxQNY9KQ9UB3N+uB8g
QiIgnq/dVNnpyJIGmBqmGm6YFp60lXLIVng2Mluwvk1Q29g2+R6VzItaBSiWLXNYBLD9/nrhIgES
Xo2/ar9I3xsFcl3HWaIyTHERwz3QKHGLXCmBehRATYb8u5o6y5tzoUDBRcun2hRr70M2MeaTz9MA
Cm4nbp1/iQR/KFuSHQhJweiWMxZyjtNhoXYb8HpK/EryMCrwSb596qvX6xFtUhDIqGytfadF5gSk
OS/3v92TVZ2W+25k3rzsFkjJzxnSWRS2w38+UyA1AGlBwnPLTfH5aIrld1k30Pj1RuECUxHB4gFi
pYwiGOUvWn5J5VZz6Lz0p1JdTerjzQ1v9QwAPaty+kG/qJlZy613W8+SSXiLY4rWIWzWCOnXJ8wX
LG0PVFd3Q9NXv7XiemHeRJy4ZWE+2JTTe10uxBWXWfhf/Zzv6iM7tabpeNhUHqxBN70qX1UmRzBz
wF7b48VXKdHJji8uA1Io++TR51orpRCtL/h7yfSjlpMSKm7JtBv+uTsxMYEd4WvR1AvTx5E5hewj
51PxRQvLoVioNR2/nKAtpDl5mb8TbVxKqBAEJw/IZvUz6geHSjJ2lgG3p4eO/qFEZGvdmJJqEk1s
3zIixtTZ8sHkMjrXyqJT9PfnxiGD8SMuMubFag/haPfUclPgqH4PeYakPrU4pmGQ45vW6Tj5Ti5+
VfGw4w2MDxsbUCJa4IFr5oLPthtA5BUiIjYhEbXrtZPwJ2/qW0P7lS/f6YifUjvbgSHiwZiKM6g3
rwYuhFsmW3cnBtf8pbIGHg9WBV4y6meAzcaAieBFSMmDW60Z3Y4T1Qo6bq8kkY1V7Ldm38HHU1Qr
V9kJE77xkJIkRfNnQteOc+QzkMojBEdUNa9fG4Z5gQhXLxK0D5hxsvx2T4rKzUy57oZ3nqHPX1A+
/xFzslf+DarCNCfBa99nxSqCXY7kAwiFAJgHTiLHch/gTFAUGVVSKd7EOnKDrCXW3F3AYGHLlzSs
OacnRx+u9rPWQwugkROVIEcJkR9XoP/2C9NZl7UbWXJo14pFmIWyRYl3O4a/fRhPdFnVEoPkiaKV
swdy7nlVk0fRda9XJvwAxIDwiSFvMu0XGiZugOw2xtfu/i1RM+9hUEYcmjZkbAJ56+noPhr7+FsM
0bIix46UMA41J2wtfoOP9kngFLEXDqREiZKpMuJN+93mDSR43xndpC76+YB6hc0EyYwe2iA4nVxv
MnB+hyjHkSVlg0tDbb3WRi69MyrwWajAZbRCLnIikIFYHdhaW4nKqYP+FOWUPCg+F1zTzH/uHR7O
mOfgp0CSmKst6qBzAYwTafAM2+VRotz0qJtiQoiY/uBScQAWwqDeYkmIjBI6/b4RuIyf3SHc8rM0
yQnQPifourup4Ym8NGQ7Ef8uVNQwPTigitKRCbKbglLTBEfbZ+z4vM8IWrv4Rz2z5NQ4G+Cznv1j
AmYTLpuQK2Q1ToESbBCcaXDeRWMQXpfJgxJ9XP6C6JUENgaeSJJE4NhsAyIfi9uG5irXJWx3IjDp
XXypLu18vmRczjcmYgV4m2IRH8vy955xWDaC1oxr8O/BtKZ3WkSYT6Qe+cOBX/QQX6s5ntd9147t
9rgvbzxVB+oEji5JK7hzx89DOj92bDRvrmmZRweFSfMVlOGUm5rR7nEwBQO8gRZQGgSLVUORGaMT
ChD2KhZXHaLX3mLVRYtTgujh5pLuJULjFnNlXSkihURdLZ6qsyIjmUkVoNy7YsgPw6RgQ72c6umr
x4+qAnuP5tgHAzYcOYRruWhxdybCBvCS55M5xoKXx1MFpHaaQDYy6vUtAK4f0h0M8AQl3LS3rUgG
XigPplImqi2zH0TmdvX0j5jPCKPj3wrNriGK/SnKbwgKUhiPCjse2JiPo+3lqHXBr272gMOTcmvb
1fVDeBL4LZwvOc4K019WI/TgkRI3JoXEU5a9tgJKKGblqXARJqBOWw33gEad730s+hqzs162+wgP
BqI86bDUgsqkZr9xZY/9B35W2q8vhNtsbWRqN4SLIMJBddan7ZQNIOzMqyGi90Vdg+89wIy2VPEL
EMHbwo6Z1ukQZxlbTjHtWC53IJphSEV0uG5nMPIDkoO5OyT6B03b8kqq4HN12l+EW9zlQmjmMgvt
vhs9uOwbp9dXaL63hmw/HertbyelvFtkK+MtGXScH67fBR4vIIzDCQPAd+FpSD4UoEySeyvT0tL3
c7KPKBUZkW/RlBzqTQiVaW+8foZuXnwvQMLCJIUhcxodZbIJ4iaMugt8PHWcDbMVGw3tLz3/naEN
EnLNxJrZNps3+NqypPOPIDWWTu9nnoGoAC0QOpcRk8ufux1XVZDu+Xi70veJDBJr0TAxAgp0j/9l
FZRwowbp7UgI9wNTi03J878xkvlN25WjTX7uDZXdoO1Q8xbXSdQxYFlli8OCBKekBYbo0n1tXYbL
FJOC2qN5/v6zwLbuMWu0k4ZDLmb/M7t8Jch2TH54SenHD+NVcBMGv69R5yfL+KAps1cO/vJM7umZ
XmTus72fbfZL2L6ndF+uWoDeS5gz7FswlaC2OvlMxlOaiP0Nl2wN5Fo0uk9kmT/GzMmG4X+nwxiM
howPcaqqhHTs7OztsEE6SNK0X4KIxJ25+H4qhcnYheQlGA9IfgonRa/JfGYfxJ5D5dDkSjoMtxYj
VhORCW5Ekh1mQRL4w+RzZXSjgLWXPFWcE6VPen5LToj2SKWfTDvBEDJjzLKA/Wt8wfL4W4ajFYdS
nARRbR31AIBA/czHDgEIQBriUNk4Arvr/pGwHr/NVgFHIIKX9j1kjz4mL/yiE27ZO1WYl3fq0Y+X
fqvtYoe/S/BVR+GU3rxnikeKH7MA7I7nqX07zJLgb3Ykuk3T215Nii/AAIrjgYJzJxbOtT/2AZzG
YrV7dI3TBbMWhXpV3EnNSo4DlBSZVvaHSeyJafUj4QnA4HqMpybNxssfWsALImqLkkL3e8NXTa/m
khao5PeKYvd+oxtAU7fFE0iaG6ilj6ZMPz8nocSTeQZ0UGoF9C/T+vd4sEvo4d7QmP6FKJK3QBrU
M5UjCelz97aSRZyXAGQE/beciJoHRLp2HWk+GGgjvj4ME08vZCIJq7ngcsCkfIjd0HPL7Oln9shM
vLjy1KWzPZ9ZBF1R+jjpIpS18emKmxQhW6btSdpzF3iWQ3CNzNhU9iLgZUI3qzStU7w2XFxLxmNZ
JE3d0DTZVMh0kaRkPiq84iol1hCdxQj5k0SwhGjhvmztC0Kuy97hJnB/bJPKa/aHleFPMHNXFVs1
ndQgDOq3Eylv7j17AXa72ftY6fR7IxwlgjzPB0a4Xfw2fLJk7SH1e1uS6Xwy9bBv6XuM6bnozJlh
XUg5F4OB0i0P8mHkugi4BzZGocxa3iTvC9TW5v0lD7cTGrhCBAuTMaqojSF4VMs6lgvhvueL+Hff
5E04I6s3R7DSDQ33ogtXLZ9ya+T7I3g2vx+fecYKcr33yeUAICpmIqFAx1LVkkzn9CTE8QhGgO+C
QVlR9zbcYQ3PqYHuDeU6TZ/KrE+9vJKBCD8Vk69y4YHN/LvILfFEJrnaKbkkUoU/DH4p+y17cSpq
306gULbXgXGjODNnAQE0/Tu1QsfX2K5fIiakvKY6kppch4Fomr1qwos12kU8o3eO8CmxfnHHyFlF
LeaWCPZRjxPcv9ovI23K56MJCziBgT0fK7gej+ifcpp7JsH0iKt2IoCKs558ep/2U9D6k2uprnzI
sTxz0i3FRYDtwtNy1E3zWjHeFZrQC1gFlgc9fBHBYxpbFSEqvxDjsxm2pJ/LYBbK7pyG6AQ8HpMO
zMRrG0NbKMSYW+MVimXs/aU9n/+xT90EUQL4OaK9vqbT783d6Yr/RAJ1y9KP2LQqy6/rULuk17QL
vjWM9HvIayHzOlWiA/svjfW+P+Zjvzbxj0973p0VIL1QTkOmpaXT9vj+sYQg/Qi2EIeJSWT8GwgK
lutGnLc6DRBs41kyiEu8asrG5SQ9+PYAN/CqlZc/y+B6VbBjv4tVufcp6HdPwF4sXJfT0HB8ss2e
KSShIzZu2Ma5AGtKBR52e7e21/RvyllF/2z2Zfim0kCoS0FIf0xbh6kpnd7Pr+yootajCRXi9+wY
Vhe+gomPJSuEoE0ESWTfsPBLgLWlLZ42pW5GzmT8fEhmTjT0GH8MnWbvyxKTmu8ZGkXFF7+yJdoT
pC7XHXIgcZAN6JeAYhgqPxZVcArCCIY4etRvm4V06H8SbNmzP9v87dmoNskTmmjEsXul66j17FzN
W052QqCs1y5lfHCDHkthxx7EGt3XExSXumitv/mcM04d2aNo5a1leLcj5XCtpRDL/NhQbIuQA4SV
IwfqbAFtphsxdBfKs6Yxtp8uzGJysjfYx/lL7v74lNvGkYrUcDjGfowV2BuS//XMX8Zdq+0kRHUS
p3+iFjpOXkyPDEwhk8NE3JDSXwAqHwSwLzshkdc+R/9Y79Yy1vSetzKHjjFqTP7UDfxHT2nmN5h4
/0AlZVT4n0xQVIU8DD98krje/7IfWcxDUxbU1Sr44vmDRdZpsyQqkacKZqOofQMBnoLWlCKcYOer
Tzyvdawypo3BiUS1IKlsQKpaRwBWS8CT2ZkhlADUEATfgFZ9fxOQZub7o7gj9keGn0KtkSyZK0E6
aaw6eSJyEEa+3k/8UlLe2RqEEvnIrtn9bMlD6AiUaG8kfPReHE+AS0+fsXHoglxWWdKrSe6JnT3u
SSCIXeL1mDKZkCUbCnQYoszIEVRC3839jLyKVjGWOv1fWMhj+T9dthdAlQfPSdjSlI93R6H+tNxi
meUj2v2YKt6fQy1GU+8goSEDD2Jpz4BkTyZXkYAh+vw1pFqgvt7cZQkC4fsMZbNh/eCToWzUb4ni
gPEJXLuSOepeeMg2Qw24k39RqW9RowGcORnazuCO03NXpeFAYVZ8I5EXeZW+QDtGmqwhnv2SKWM7
VYTTHwtLqdCjjv/brWp2Bch3Uf/9PAdoV/HC6ynYTSIhp32TEo6xA+Z3MF/oz7Ij7FDKeAUgAqCW
qhFEVCZuqVeRY9nbjcFaNBO6tTm6Glf3oJcGBRVVwcRVcqa8/7N5NPx3Dw2MK7GDWxqC8a7+af3u
uxd8Xie5Pe8ZPDwf0McasrEfExBkZTTdyTYBnRZqTxywIsrXLCLsRRSESaoSdt4Sbm7/iLgMz0o+
LVJKV0YYa5rMvdxJ7yG53aYANtHf03++4F4yWpeDc1C4k8CbT25TEMncaSCF8WptgF4KD5249EXJ
jA6p3PozNwJm5FX1t55uYL+FSG6PsR6O5pBnBJyXAKKnBa15DWlD7SAxW53RIvh/EcOT/SFuQ5je
D1JATLKsdVVTyRKUkxMpLesOVkDF7ikSeHQetJdiPNvxO3Ma5Msm+9vCk0MKZ0dTi6xXFx/ElRbY
7WL8ysjyY2EAZqNQ0QER0rZkBxaNxhwEC17YihuAqhgbsZBLxK2wNq5nmxSmlET9VopVQWk5ZHnx
Ip7jNJgJTg8fCO4UBGRIrncFC5rar38B52nXCTC3qm1IcPAXzbLVNSqPnednEykIctA461J7ED5s
9349rmRgo+Ac+iPyJhBoa9SjXytNwliZWym1KHHU9a5s0ZsMyQlVfvdlzUmxYHfCf/DO50HQNfBE
35BWuHwkWMreqg4iTvkyZCqwgSpcExZTrML9xiAePRzvLTR76DdW5kXp0ZyesCTcExOr2R5zfhR8
rx+5IBao/4v0VNCATvPau9XRkdSzqrv5JK6XfpdU2kbsK8fhJnSb1EPdPvW2/H+nCzRr/P6LdJqK
xo9fOLN7FiTm0SIMvrDbV+1QVE9K5t2aQVnGkk+b3s8vyoHwfTUW7PmjtdviPmOs8CdVo72TdfCM
w5BJsPut0RsPKqw2UASD/y4C/K9hzl5BIX3fjgv7dNg1iWusBJP/Sq6jumF+LOO3gBXaIQ9ZmiHO
6nWOZStFUdOa/G6OqFa7pES1Dim9EmkAhFkHWl2iuIK28Puy5ufl2eJwBpvMGoH1LkCoiF7KeNah
U3vC1Hm13W9/6cQoGg5PYCTOPa4/t/cJU0r+FNkq1npDOyLg+jbB3bKXlgIUSZVZzqSAHoa4CnMe
BxjBQt3yLS/2LpdH3aU/yHct9a07OeylVp/zjxsh1PCZiWx/+4TlWhTXcpy8hAov7xBK3q0/Qjan
+XGrOrjyqmdVXettxnkbmlzNA3Lfwbx1MIbc8Zl0R75vCbHi0/biuIg+ZzNUM2K0wNhi4dP0G2v6
xjk5dp6LtlrfvyEaa+7YMwuau3E0DHvpnjQf6WFlhBFsVD/5lsRvFHQmxGEyfysB2cug7K90zR9s
ejzuQZ8ULQtA4GFpsw2Yu7WlEwxYFJq+hMKHerkIIyc6hrLcr10BRbXtaLuZGZRKb9hcMggCxzwg
VWgOvDM33r42Gx9MXkRuuvYd5F0W4QzlJoDyMwMhDTZ7SkfsguMbxwuNG5JmVP1Kp5Q4H5MtTmlg
2u9Io2ArdcPDps3SlIcBi/Y2MqI6m1hHLYpEhitIBRxKgFml3YXGRy0L6MuZpfun3l8IXl4sqKza
mvQKw8z+GzhFGGpp8hA+rvfg6EeVtrZh2Ht9AKhuHF7uaFq4kU5lDOzrdf4+UIYk1bB12Q6DpF8t
1Tcenp/mcZJAL2JhaOz8shNqz3OMPk40p67WmEh2J0gKUguh/9QNR3OXsc3KT/0I+NA0Q7OfP5EJ
YvC2uZIXatmE0i2BWaO39Lr8b9ag0SiTzsNIZLzbrVBilGiDwRXhNB97gnb19dPet8U/90DbysnA
1uQ2pSEVTBKUcxesbYbLOuKRxpImgQHMPZuUM0j1ppHGAhBRMDZtkHXTrz4hAF7j+JNzwKad0RGw
Cu31hSZrgdg8QpJLVxH9YZ/eVEhToiycw42JSpL8pYu5Y3VTMCP1HansEXP9RkTylh5AlpI6HGSS
OVmIMfQ5Qa3uxsYx61I14imPkyeCFNuNtOF6YoJzNS9sFLPb1lMz5szVrcY7v7tTVpaVw8NSXb7C
gxbHr47MpCMxNqC5bFSvwcP8okck+s6vz/qhulb20x4BdpOlllXM0vQCPdLPEkqzVSE3ZDXihS02
dxTlqpDqL7Q7hvby9v++tw3N79oRW3KrNxKzZw3anE+G+3CQM652/kPxi0cyqNTQ2h5SvRyrYGs8
FxGIY4sb62BUG+Ezpmp1qfZ1LS3k9llRBKjS3onF8UPXqB6HfQ3I+GiJUHp661fVjZz9QdU0Ja7H
tiTvTVHvVi5kWc175zMTt9OgeqH5l9X9HV/TDhSFegupIzjj7C6SKEO3POLwsit8A/M3ThTB3Udh
GxdZ8x8Fe0NOmleDmpTf8G1jvbjm7pl8bEsDvJI9I0e00PaC8Gzw5vt16bn71ffnnLTxfpYsLp5o
pCKhcRxBaiBr0VbzkJKHHOU4Zmfg/hQLR8qQscnPFjqYVV1vVPbl3M766+y5Aagg4Rh4tuRfi9Ky
ikrcYGuypsb1PHZY7xLkodH9tSDNfUnglkYPX4srojUgZpQo1GGciqeb1QMA/d/WkWba3h8FeOcx
W7DotuAd10naXYu4/ew/Ah4pkB9wkzBTEWKHRKP1zxE0ySpooS5wj7n3i+epWajDrERAWGquuf8T
JSVOqJKhG1NdzWRidKJyU2wTM046HjtInDfxbvJoinEsUBMQxnHL6JCyqnGv3iRF9uBnbdnDupI6
rE9TxZeNforOnn2vb33Qkpn1t/0ETSODhyZ4NgCVYBWCSNW0TTlkE9swtQkTGRmE5WJ14aB4Iemp
hLs9KNb5AhfCBtHVuEcy5QIOOBXVBp6RwLEJGf5WEjPUIb5DldXNZhtkXFrHaQBxf9qs6oOxwTLv
xTcqwZ8t7wXeYq6tOy2RHL1dktXDDwTlghd3aUIBepRZ2umg/7JO7AIq3YRq1WRqiVIvTUA0JRD8
olIRO8LPZddI0Ge61t5NdzKV7wNol0z215cZ8Z2JvHOUFYEdEVnyzMz9LdYqJGkstA0Nw367bRCu
UBJU8jDptCG3bbsYvxjJDfCWxGSoJN4SoxKQHZwSQ0ENLNDfKeBKCPzrKiz88Fx9591d2somPP/H
X5ntblsoQz27fEm0mIJfSDvGr//yEJkP99HotyMsJin7OY7CBrfyt/d9O48Ih7EvWVW2eB3pa9+x
K1Y9uRgfCvau223PM4BMK/0p/UcEWnhlV9eobvTCmJnamLsdykiTytNcyDs2Yn4pL1RYDJ7TJuA9
bkItbXJf487lv0PG69KZcj4TTOYdof0O/BHWsUZ9rOL8T1uF+ijPBrfh8PVNopFGWHwgdODQF/w8
A/tiBgAsMJkuPq7lDfPL5Yd5r8kSYpQbgMGWjOD51UmtkfO67rlyJ5BCcavHj6rFfEYRPDdSlu0H
z0ppN8atNQEQCIPlB7brGTay59P22YiD25SCJVX8Zu8Ix1aUBI8o9usbbNAJwwbC6/TvhX8QeGjH
rgZr+E94JN5UZmZPVVdrMRosaaU8V70J11yqTu3427RMhdiumsg7y1qTDCx372CWC3LsboTQiRVA
yVlFrWva1Fa4zufqp+xNlBwsSBIaZAeIr3q9P7ybcwP8akTX81BKqXdp9ksoa3ChcFM8wssLK6gD
djHchhhZMVONUDrd34ESWuGYVPJVz5wabjKMwIXd5ULDMoLrYfU9ULQ6rBoMN5/UZLfFXjPZsbmu
W1SXuipi2Skf3u5Co3qVdHhqawmmpz9RtsD9Ype9O37W4ROF+BW0kvVbCMDvmQNAOQjH356wKHIj
G/ljjWrEGWliENcgk/PSgIXwS3eZ9pkh+/qia/2cdWTFamKt/C33qotSMMlPrYdNmnH7di6O2gmk
hbCV7r2H/FwysYs9W8m/U2bjBLIkHkjNJi7tYAxArtOgnt2tNx6kvm9IruF0gK5piIXJ5b4/rDDk
S8S120Qnmzuk1oR96CgmUaHhMwmw6jfPovGVYjkzBRKDfwktqCg6C+FORWZD1dQRgWCMiugkvPpK
Z4geMrBFbx6rFPqID4YYY4MGNKxG46Hy4V5N7ahOzAORxdlJfWiSV9Pm0GaUgHnA7DRNbpmFJdqI
eUKdSyZvUDppIBdaQhSE4uELbNqHrn77i8l1YkYHKgzqyLAA15V0APmbz/KNPXA4JKP9arpkWgvY
daxWYwsiWlbcaP0p7bCh2/P4sDtCj7V/y2oNuKMxIuuct7xNZJ58DA0e6nSROwJbS4/SCFPxKFy0
gHyK3J2IuKmNwvWRu7ch9guaGrNvhK86OqoVi/cn4dnLsQ0SUg4qB5jNwJZq8BGgV80lboJ45ReM
AyN6q8h1De3AAdZGBfWhPqRi3xo+jElyQ5u744kw1Ll/W5RNhyDXo13cZhpz0reTerf7HBeRv/Oh
ShsmFklJz8FcZIp8CAMOh8yX4jKNidu3Y2RmwRxVWTm+1fcCiB22JtWDb9UipGpXGIbyjGKRO/uq
mdD6yTGDAPMyyYZv7dgm+lpad7VF3wGAlnGLtvP0HdCf0zJZOwqsjzyGYA6RdCa2XlgC7D1pbhRH
YjwRCj4LYuebwTlPkC11kkJN6nv0sDnZFTqATjffz/kPyQSnpyv8sfngfCFdvP/xU3YCH6z7l+iq
TKs9EnjnipG5zxyZvik1zDkQ6CdE0H+DkK0PHE/0mDDxUhAJXPAIrSHr7/cr2YJmryLrZdVbZ9JL
SezY3PACw+zwQr6niOs8AbIzWsQB0N3++abeiKHzmAiWJTf/CKYgD/bdw+tYJaNNbMewMKaeEQKi
3pK3aJEn/98pzUeqRVWmoGp82i3xRG9TXemC+6mrXkOQArZm/TRzRLEsQE+Io6VfpuWesZcwbNcP
6D0YC5do8jHeWID//aBeYOUvJYuBE7ep3jPHIiazz9Vx5GCH1OwIRg3ojY+WfU2cSYLuoEe2JGIl
CX0Ty2jUv/MwjWKESrTvTAxSPteN7qSbfwfReBVVbkBNtfhgIb8BtoxTvTdBMPGgrqru87py5qYE
tOj0x3SviKoR/zyAJ0rEmpOX6adk+GFqGkPJVGcfihVUl+hvmPxJDDxIRfHDpgCCxgUtRi/NuNr4
0GxRv9xIpeq1g3lPEyrxCF6FuI9St1I801nQRycqZnDWcx/OqWMJ8r1HT+1FLr5B7TVGgVbYZ5AE
f1DXTTk0rWAyI6Eju1akCkP7G+2Xk8rp/RWVNCEhw76FBOnltf9ya+lGuX14Vgcm1d+8tc1Z5rBM
ZDStSMbv8nwU8fV7gZwK+4/FaqanTUVnZt1JtQDuRZ5sMZYJACNlXmiF253/6gdqT6zVlyufmpcK
iV07GhFomeFEtTdEpAy7eC2N6Lwh6NGtuouk7emKofbLDEld/dUA3jsfN5mSJsVA7cztvH8dGYi4
u5P6IBS/chVIcgihmDVwu/z/zTtuNN0aGcYdC3OjcwklftT/IXjuS5/gaPzTZIZwR2DuGn/mUnL1
mhSs2t1Gf7UGRMXX0Hx9ARakaTNIJTU5uLG2OlvFrz5h2mJlY+1F1jrStDIymsvdPZ+HWXYIKoU6
km65SXeBlr91K+iVRGFuKx2yYQZC4vhH6FFm1eGzI3sKBeqDnUeg0tfLyq7QGxgoj3G5H6JwLSQc
ScPMuOfz1ZRH/i0RxeL/EetVnXJQRsMdQmUrqnwql3yP3UGtw4qZzBitCmsRBTyxRxVuAsHU9p+W
De5II9KOcwstpW3Cp+FL2O7AhxBX7IDUcNq4U3dva7vffoUOsqplTAhvO06x6LUsUf2YWz0QItOs
2a6VgC0evCVSxM4GyD64Ypr98Ka0GjGznDDI8u6I54ELBkmt7ohOiaODfZ2GvBMUv2+otzP/gYc0
jyf5cvB3JHYTYJMPiXk+eETVDfBDrIUmLAu05OMzFYVGtNeZDbMolsvzWcxelexloY4R2iOjy3zK
Nv/Ye2NuY+I8J0HAEiHVEW3Z7PzEvuy6LFEjyJ7OdZxv6ChHi1X45KotT8oXC1+Phkv4si8ulCPJ
RTkRV3igeMakzQ0G/Qb993m64fj5NmQO9uULc0gtiFVRnLACx0RIapr1BACwnqhKF/ZpfeggM7Do
kC/3DtTZJiRtvqNRY7GSGt06cnwsfv8VRnROkekpgnHbmY6MYKowXOXkq14QDUNeLqnzDU6sTXGJ
hLH9R4Iv4U/9VyQNkcynRFRui2XSsT1Z6GzUTP8ytG4s9k+9QLicVmR5XjyEwNXH94Gmp5WCbPpv
G0VWxKivfWA/s+zCxz1q1smNUarol39Ot1uq8uuk0e4lXV2PSyfOsrTE/OygnCi85Y51dIHH0K7u
s0K7yWdvg0/YfJB7OnrzxX+PUMhb6OKG5niFf4u5HS0bO/Ne8yAeNB+XnUKdkN0OSJEZ2kwQM8MD
T116Bd6DswZYxTNGDuwtYGEafMxFj+4VU/y5espk3kcVwhl9vhGmMb2NoVmXd04LOmtTsEgI9HRa
9a2rEJrdrxXJOaymPvfj5CP0Lof9vDQxJOiCMbbWUuQzUC462x+PRD+DMoDuvJ1wMiJbTJivjgD1
tYXXpcYYfY4GJd5VOCZXVAvjqLg9EiEVJUwBshrGxdD/BMg5Va9kdXSxGF01gvfV/jifLHat4TVH
/K1FaTbuY3rz4Q90w7FPEa0ZLT8lu2sPQdGlt7eDFz3bMdtIL8/we36WuMrVBoRdfSqENWsTVc9m
lxXhUR7ObURTUtm30AOxmEoIeP6id4CmqLg05Ad2iWv+JIMdY/IC1yqzlroE+nVnWLyI4nIoumMG
OMwgf75gfNx0ulc+C24XUlBWt4DeqOyyjIqgzPdtbss4ASLEnyz59Xl1+iYanuMF/m8SCUe+ogHe
Ck5vsRW/EfGcbUgnd+5wdQAlFNiGJGF/QnbCXdwK2VV1RNUY0bqfMBZYcWhXReEf3t8hDxmhztub
wuURz4P4mzXrtBB/QQe9GbdlENTfDPr2m33s/fnfLQ+15VpXUDtdqWdebdnb0oEgYy5Y+51iGlfu
nUNrVJFvVzfPafEjMEG7kSXJDbQFZNhd6qddSWt3M6U4oFhEofRDI64wrCkgMKPBvTb+q0rwZaKu
1+JwKWupCy7RDWR0FPegsd6oCPeRsUrGrFWGvxDRKoK9alJ9X5EFyjnfWFsg/XwNOe917sErqVNY
3LRd9UAj2Wp8oDvZs0QsNXLZUXAnCDij+Yolbf4bmEjhn613zLSDHRnV1Gyxx7EV7EZjEx7jMgEE
t71vy3ts64SA700LTb4geyNVu/8rIWz3qry0jo0/9S8roubnIe3x69C6aNn43aaelMbX8o+LdGGm
SfQLbvbjtnu/w6J1sb3ZWUwSgiJxCeeFK+Wj7G1MY7avk3xqUFUMxTPiDG3DhSknzjZQxt3oRcMo
BYPurgxWp/saKDR65jEuYcFt19EWkUvaRbzna+b3GUEvaIRLSj0zGI8rWIfl0ggSI81CMHF8MSnp
yVzoFMJUEQgx6mkaubAgSYBMZoso6xCmW7wggglrgLiVsvOq8itDNL8whAOu1BWDIvMmbOxgyGft
1J58iyXimQkd7n++g5Wx8N1DmFvKimNj+EjxqUvgm0EdCQdWsizUTHH0k6kG1Ds1LZwaU9BYQ3+o
RJenfHHNHs4YpUKlsEozIWvkEEQJXU5hgwdElGg4qbobiYfiWeF2JkAXM6ID21jQ2uNPH3ow1Syu
BZi0hBjqn2He5YQOHTZLZabafsEx03cYTNSqPH5E7Qffnam2DVfizSrZ+MaX0LACAQGjXqP+Mhbf
trUwMJlKnDFdojpQuCGV99wBWaDp5evvDEOf+mHYRXMVIfBr97FXFD5rbI/+mxgu0zrYWx60Ptw9
ZVV9kv3Hcv8fTb/B5ZjbkDgFylSOaA2UVxx1xNVZAje0882bnBVwIVPoz3xfvbVSWCfjPLAnwprm
WKBISGzeBq9lTRtSqC0XlCGN0ZgSymfJ1lElwXTJXukxqNrBT4/IPsME5TpCAk2JkodVI0wbQIXG
yvrIeVUzJEGiWzZOMWr5Y/tIdN+JpW23F5Oczdl0moyPeQQC0z29FzwnSOkTTv5KqxHCcdfJfsaX
GzXBv8JU0W1Rgoxb9IM2e0OD9OP7nLw/rF+idj1ssvIKCAE88gCzXBEmePM+FY3AWufleF+66CPH
1ruEWk/t+3czrT11fAUs3bQ5Xb3lggG0163F97slyV21vLgOXwJWBBmhaAMhJyYBX04Cag4a0HgL
4/JE+avwXKNp42B8es8+skmHBekcNn8yYYKWRwbqi126ddHsakDCsdYGdFhtZCZGlOUXBFpEzhy9
S3GsMH47nJru//TceSHM4mAY5qnHYVGRCzZO9Oeq8aD1mxcIVuK/8J0w3hw1mFzTBxRCS0UC+qQC
7bBv8Ocpuf7j3ZL6V+3vGLIEcF4Ko0sMxVtAJaCwzQQgkb7De9IMY14DuiYUCE5isvlh7Rp1IIOt
dCw/+z7t/bIG/9LNHyU+TrRfbjtuzklK4DypkN+pMbgpXfEgspRew4RgK0wIf9X3xp8bKnjj9t+Z
kWwDLLc8mVdjynCMa0suxu0HTWcPzMEKaUiGgz7Lrpe7vAljJRvDVV6/GzBmTaavV42oyvmGgIvt
avwGWTeh3lT4DlVKzolAwQa3JF2TESE41XCaSbOa2e3Qxnn0v/kX0NW/+WIYObvYk2LTyy7WmVaa
dBwCuiB+dpQkUXJyQlww9bVD/YhwwzvVSzC4J3pAA3oaDCXSwNS7g2NfWiBgXOUvxXYaa8C+osyH
RvNcx/PReb0ie5fPUx/fIRM1LdOBYA3WrrWgMcPJxlzAcyKTejQvQ9RKn9OlPTZV8msgfAUDVktT
I12PuFgulw7ZXftqNgy6fD0wgJrkFu3PpXe9ZEyGS0GgKEuLFuTtB8ubpoShgc+Bdb3UZIVgAui9
KtZAqxNgPX2b/OQ4/4xI+hjFTPOuN2fSvetR7CmhpjS9tOqwsXMZGdrDz1m59B0Pe6Hzt8eh8jtj
mfMjNCEAfv7iHzcIyesEgdLO94wpB0eE8Qq8RI+jBfG9Zd9orMW/2BqR1JZjpi58Sce9FyQGyWNd
YAIpkmslAmWjJ2L5qXWmhGHUxHLuO5Rh7CiGSg8stnxPgD4FW/9NmLWDRTPKUqU/h2DX9a1txE9A
Gk7FWVSXnKWUFJYRNPLUvbAl4FpnPcktZL/Hv3jfjLa2xcYcQFpa1S370PVYK8v1TmXvQoIXixyq
hzuz1AzRDX9DbWiTdXW0P5bBp4NeZ1ktNrwID+/Ck2UdXXJ6McSwkobwjljrGrB8MQR0lExu4+D4
JFyT4v8/CuwmjsYyTcmRVHNUPk8UQT/oRw0dYY8URb62OyczLyxyKv8iArQafo6myKkSHV58z4eY
TtDqGTXmWMG/AFSw/IrT2JuVQ8YfApyefCAlZwgRE7BxBCSnZdeRmyvkUUMVJ20QzUSJg5ral8Ts
4rgbFIR2CBxptaybXr7WzzowfRlw05hcvgzzjjttih03FYYimcQfXep443Epl5fdLJubdaQNE+yz
+7QvIGZ1880AAkkW/ugg/RpMF2YFzgH5k/tw3HW2I5ijjGtT8/FyinKdfdma5uV9g7D/ByK/flh6
9CNSH7Lx7KGYJw4WSW7hnjJiBX833ZqR1+k1d05I/9pl5LY7Q+0UaT9VrCfpWVnTADDcsLpgMuvO
qyi3Fu8JMSrAHnoSsDkAEq30GWQlAgxvIbVDFhz0NR87xc+couB1yRJTfKX00S3GCerjAcA9QfmP
3pOPc7JSutrybE26+xE48rwk2w0RORJWZmjGg96OlPP8vt50ajZdFvkhy6FhihWkuN5iam8YwlfZ
A3leFdA0rYUIl1vSOZz67bqympaqelcEmyt9QVeMbv39l+kICaiuLvLO4FBtpbdpCwcsDGFJ44Gt
N4e090AubeezzBBpPILNbz6vAPbXfHIzd71/FHdc+3CMHOTJg2d3oJE0W/ojDLZUNCQErunN2icL
CoyCwR5p1u4xIEHxjwGhCFNzlp8IZvJciuhkvCJhpN/+VqKse+02sD/BywLJ2wKlccx1IG4NRbjU
n2xLBK/zyuuPw4feVU0KwWjkqYJTl9as3OIwncxxhTkFtABAwviQ+zsT7CaOSVA7xUHuPpNahwoW
F0FOczzUrWQ457H9pxaPeSSbyXj1OwSiEHj0GFsqdb4kNMXh10kItz6C1nYi6z1ErhUVSRArr6sk
1S4vLbfVAP3yN7LGBgzjMI+mTrTS1IIJHsd0KUYf/qYRYIGy6sqLSmSAQBjjJwJcUSm4cHZAYYy9
j/g/1eBkf5SFVNDd2Qd1aBWoRrAmtAf+yEvmuZO+R3t7Dl2W8D0zwke63ZDZJjabE0vmwnw6H77u
RecECxxleSJN5FbFVAk4la0d8XLtILrHRJg6o8LLmTsTOZRSq9oKLzcy5QEuRHL36kzugEJdm8Z8
mMc8JCEG1PI2ZkRrRyPIu8/a4Buu69x0LZqobcMw40AQTT8V+IttbAaCibdMXFR9dpIdPpieGWPu
6HCI8Cjd3NvVGbZECLZFe/b8qB+2tWAhxbJHBPgEqxMJts73ZIKdMR7Gv5szLXugc6+oyqSX0FXX
i1lf3/P43j3VYNMOPLfcYtoby5MJEbtZ97M8Xq9WETFHVyW9IkMeX2pC15oGFpN2nCOTffjaQby5
OtTDbeCbEFAF41WnloJouPBLF0Bw3vvH+vXK62atiRBPD3nNZ6PSHCErOf7ela//IBsrdZzIKIRd
Qk/TkTh3pmp5O07Hh+vYHKn3U7NVPINjuR2DwIgVSB49D6tHPeJKevx7EKYcd3nF00HNOnC8sChZ
+G8eW1XUduV5eN+XfQTTHizXxNOgh8pOLYxZANCE5ADaVHcvAnBVCcJDw8b6WpuI8MrtA2OAGh/X
08NSOVXMaKGn9yV5OeF/J7mMi5uou/rN2afSvgUDs1NXkwNoYi76SbfRFL+RTj1aKqXTeqFaqYcy
4qsr9ZDtJzVrvdGBVLzof0tJzzJAOi4KlooG6LsmS6rGecavWRZaBgvVvX79FwLDdUSmQwk486R2
BHcwYxVowwiqO+Bu63XnrKPrUBmstupPfudoXBLJ5HN8zDr3ixWKrnbMbABOI/CNmf+nSuVFJ6Tk
ilHBxyuGAnFBB1t/2AK9NyUVUxD+1R7p1P84G2nVFp9ulc0pLehI5lmpHIVVSAyaq8FF/M1TZEf4
vHtVY3flqXmPTK20ML0f+RHtAnu/5sHdwTA82IdEFa9PNCgGgDzYlCBzpzQJeNaOS2RxPpYih2mL
ivzy28NT7os5xuf14cuZeMbNvc8ZMkdIFlWprlRgJZj4SaCoUNRjySfsDRjNcCxtUIVcVz1sd7WX
clVuhr8XzUDwYDvb2wQWLMSSXUvjRbUDMmeqCrsPazxYu2UVOmGaJaaaM1Jmzu4GvFmHTgkrusNR
47a8mXD1Sid+hTN+TTFsjQnX1rKnVD8SHx6ydtA+wyX6UISPrPtz7Gq1574BkMhKgve6AALbCnJh
k/EHrGf5pUuwpRCCTsfN3Wi9HW2Zz20NDeYl9XfX9ZBtlNdsBW6eVD3zwIcpFkN8ylXsc3kpZ+E+
vOgJt+pwfpS5hoJzcEfIA8zm5ZBWbwMq0vVL1qKY1frNgVnBjrMI5rbXB2nQh1tVCkju2Qhxhsoe
HoEV9VG8KQnYyTM5uvqBQrQTcBO12AcKDkz/ozJ7aTQcgWbKL+xvIr3fal72/Kxj+BiQ1M8mcY/q
5ZrVTdOVT9UPXSwGfL6RbSRNC5a9Bz2B3LOSKqjwGCepZa1Vzrybts2cwjAd25MFCWc9kocp2zJv
SHjsXfEPnjDtBKIR6N+Pwvu+tbwvjGnEHBk5fn8lpXAaGF8nCJwzR9CCumdgqblcsC7rQM/Bb36e
p2WQH19QBkwZPOtZo7GCZdDdSwr2R8JhYKBmHHxsHcWPW5kyJxhgf4awo0ORoUKPktc4Z9QZzIB9
JZGzaXdSSg2Vwdq+HqAB+T2SUS76rW/7b/L/GhJNuBMeNADP9Tv+YVw56o7KVf3LLGAPwzKFe4O6
SN12smhSMobF2N9oN5jj+OLfDE7EQLOS3vhPKTZeB4FLjGNkJMOWvuzXgO5mmftYGET+JNKQq12n
WDEMh6p4j2Clt5mk/KcW2nAEMdJ3EzuLTGSZ24VNOTtWbs6Lf8yW+EyHlvJOj3xQoQ2RA0xM6z7Z
rL0klTEZTtEE07IVgs0CuQltJHC+u5aWmsr0L8ThEbPhvwdxp6L7k1O2sMtOUixcR1ExKwNV4NNe
BgOYM1zrwJdKDbtkTaSXfBdKj5tEx1o4iYjphh5n6ndUhLLc69aLo9s9JWtGr12a3BnFajpLvYLG
P2RCm9qR2sG5gl7cDv6Z87BZ3ohIhRzsWiY6KAaTaTEEq0e7aM8MuCdq0CWVKisnIWTi5l8I3esA
wglBdPKAjfWHLWqNqJc1+JFe7Cp1pd4a+lVbuYcI6ZwbwEBXw6WhJgsnLEAcsjYcXIt4cH8ppM4u
Ku+WCEG1zoR6EsEnRZ3bGkOhSZuEhSoJWd+kFMvgPjqtHd7cW6SIzlRGRV5p1ppJhnSJWNDFYFv/
HYsiXhjWKVDSTsYzbyAnTqQSRPVFLq/QGB3ZHSdbelbYhOp8ceaszLYc0Pm6kb315Z8zLUB2ZSs1
sRSMSHUxoc4Lg6Npnl+DL/twUDbi6WstK8OahSuoTIWIH79gBewuU59F2XQAOXp7PWME+UqWyiRl
oY5kFET7Zue4xWxea3SHJVJ/Oko+kyx0gR6rdgHSfnHGeFZRStR9YLBqAJIVEiIP1f7TguwwEaWt
OsJwF8KBdBW1iaz+F4B07+CYn/iLRdefWUVR8hjvHaY7LUbRtqHd6tBXnHyk+Qo5GtuI5g/QZDQm
w9Uiu2WdYVT+1OsjNW9iKLxhPrXl8JQ9/S2vSqtrcvyaNuxMXug+7oiFB20Zw9B/2idhGMlhTEcR
3hlqzu+EusPhWdmQiZsqMID3Q8YdMPRQavx15DZFQ+UgY/vZhWcrSdwaNDKKFhqGCpF3UcDYcn0b
gW8gnPGgy1uMhBPgdAk1X/3HWHXZMiUI4lWuNw/mntDpcDtevBs8cR9xYnG3Uvn5/T2z9YtOqe8n
2Lj69zIGcTIMUAUlFr3xwquxS7x/7EJYqRyZt/FC7fcjlfgV0VmiJ4Sp8yiR/KFLGBmw3nWajmEV
jtF7n+jgjr/pR0RMd7Qsu37Z6SQzPSAYyZqtb212+gS2lcpRu+Wl7wsbi/ThhhORva8wrT56JlHl
ymJfpMdDixIxqLns4kTuj5a68ArtZElV52Q/7LchWytbjDpYzq+UT2mN6+9Um0bCLHmmXc2dCrjl
9Sve/CFL8eyORlYesprJFlsLhxPjIUMtNNtY3AA7LfSJsopnDq08rJOErtCCnK4UZufc4caHgr9A
GCN70CwJwCe6nOjK+XnUUFqDklCy4GcNdDZuaZhXE7zWhsvGr1S4llBkQfk8FTe0tE6QO7XN30QS
xToqyOTXas3sI57vnw+qi/e8D2JrrJr8+ZuR/vQGw8Nwm3Mbw4wjvEi+T6mubud6yxY/ItiS8XNe
bCJTpb7MdiekvNmsYu8jhdCiKtB7PwkJA+CMgyu8mx3zIlsWeTpnQvGWH0cCgEpmkLRoRrw1y/nh
cEV/deIlG86dTVVoL6G8JQENMxS08Fhvj+lfAm24Wo+MpWVKJrSuIz5MYxa7uKqK0ufyNjw1/wD5
0PcZsx99/7su/Bq120AAIqDiFaWMVcGKLXRAHauHLFHmdamAxD+zjZhglB+CheOzfWAX2/1UEx2b
EMGyfBWb4MdhibvCt2hxF2GWiut4Ie+Hcywz4UcJeGO0HkbcX2OMlAglsz9Uo8uwgJqj9vDX7A21
N4Hej4HhqgLS8amoWz0JkDqDfAl1/nNC/yU/1RACn5V8J/nlrjyfsQ7SWtR3BCOeFQA/7Grehgj8
b703HCmzATw5dc+1+JLxLtZd2xLKLa4iorS+OTwhfY1xbCi4EDGb/NEOjtP1O8dC2e93H9P7zyih
UN/q0zZwHGfsK6UtA3H23OWvSr2b+Cx0r7EDjgzOUXmlwyK18xsWquVlCQZzFydY2AayN85IF8ue
RgAc0p9gh8KXw4W5RXshQrfMKBZSIiuh4/ftewUD/y8Ne3ji5Eu/BuI0jOCnXQeJ+dnq6ImrirzI
1G62lgsAT6cLIGi4uUWm621ig9DRuXUwf/kPguNJDssdfvNe9OwjRb40trtKj0N4bcxlv/1vPIYI
CWlYvTdYmcIGhg1bn9h0QeKZJ2kPuCrpowM5ELkDCNBAtqe3FrNGjHSLnuV1BzoEBjb3ZtjnyxaY
pQsem/hRvJBxRkMd64vrbYL1Jm/LBLNMcmN9BTbodmGHA6wpvj2v29ScZiM85G4yebSho43/WcGB
cChMClJmIrRjtktsMr1vOitInTWaTmUXfpiAbV2khhN5h6vipu+unA3Sf/oXzjffTtXwV0SsNnhD
RdSoIBMnPUYv5aevmvI9tbZ0wh3H+cHFM7lSMeJYgUygzMiekmrc3kWhRzHtC+khbAElwEe9pSVz
33JrpMily1s7a3b7sKYj6OpL0dtr+XLRZAlCSmtaSkikIpSO3E13VyzNV3maGcvq62wtP3G+zyXg
OOdOd1JrMe788UUjl3VoiCjhfxLxgo9eVRClq3ruoDjsF+T479cUSw+qJKsOn3tH1TGFZkT5dBJH
dFW0mkOZ4PsGFcmDYRod9X3OnuntkR/DfiNpuvC0NiP0J81zpS2+rMCDMBOw1l2MBOznAf/4GtsM
ybnD7O9rN0RTmoiDInvlp2LJZc0I4h5+7E+O/q7nH63P663hiyfIRyv9zC3DgIQDaB/wep7ppXys
EAulitzVMg/JcZTq2FnvVOPFw8BOjNvwqy8gn4DIw/NPZRHXIliBqNfXkm1kPk2aXYlzxa21iocU
Eytyb6eLvVE3UcCbJaw8uTpC48VkHoWneE7+3oedOPGR3Oef1m7Ybpx7XITe/rrKiGJSLWmjPpwC
nmu5ca8XOIIHXou7+cTZi5unjsywFKHbp5ek8C2O+j7atlIHHNY8dmgfuVsCChPt+I/lAAG8RMEL
i7nVaHu9Fp80u64eeZN1DZhHK7N/7tg07gSC2xGnyH6alqZLI6nCgSwHNKRChe2ztn30JAticRCM
n59bEUhOaDWRnld1uEfTemtvC0QVZohBPZndd9A3K7FV89pGWJTPlqWtqT6PkWvIyoMj6B2W96hB
KVT3PdQOc0lx4ReCS9H7+frEjt0M3eXvLbiiuDYi89pPkpewwrf+uMsiPCOve3JVSYDyHsLBaKLi
Y2xDJo56UUzBREZ5uYERgHLCgppXe6DllbJudD/uUr/VXX1tcmuLZtvx4Np8Q/VbhLrHVPNGHAcG
rd2aiClqRBJ71nWhq5yS4J4ZIVSLVPpHpylD6sH7oq8ss7H5ZdiYLXagFJDx6tfLpe5L2z1SMJTJ
VOUF9VQOrpGNygmotYX0kJnGeYjsvTyJus5N4/lTdwl/I0eI/VUV1oZabxn+Ry9uSJ6yce4Cgr5V
vjQ9mr5YVL+HW6FCx1QbhF23B5PJooJuzA+EFm3VU2Iu9iTlbNvNA/PuLK7KJDA8LXmFpFE454Fc
sSb4KJ4t8HD1mQYOc98iK11/bh6hxJi+2WeILy+aw6kjZyoetTlnPMApN6ncoJnd0p6zsOL4sys0
vo9sAJ/YDGqVslzrwKqAwolUniANXSEq8yLAeVMnk0uGGgRaMDIZIfVEto4TFSay4A8AGJwJwPjO
YsTfGndgh7y52fAKhpMp6yt9gXhoa6V8yQigDxg4N3sFq4ekO/ldu81ItLaJ8ddVpHJSwCXEUqV8
Fr4W+3CHRWbrwet/sREb036TycXhtCC3SSOGLw8o03Zu9RzVAdI945hgqEASg/mOAUngoUV+bCeR
bwWe+aXxjBMMKa0kocG9yw9XNGm3mnIg7k7dlKQmnQGg8j5e9DcsaUtRnmTVi6bwxTssPNtTaPxC
R68yXs84JN44dQat+v/5cbpTrUpxGrMM8rMC0/ix1BFUnj5m0DY8zgvB+LCZk97hWP3O2SdjRcGU
mtKBp2vSmJ5jzqIak4PbMD/3xRXoJi1QK6KvpP6WKDmYa5FGNJ+8GWciaA1K/X5f+Qus7X2EPsOH
LT8WRIxEFsMBC7ZnhBlIyg+V9GPU5oArCu8yLPNcM2eP3KQt8Sjkuyfpt6zXkHOU1Lh28XE3Re/d
9b2pS0nugQei2w0T1yskAfxroKhqczESHcFk4CTUD7BvFhF4K7LpIAYD9e8WfnWpaEKIew9sGIq3
sQRJyBU/gQbj7YYMiu2OJk1FATe7I1mNWL0RAnkO7Xyx2TLVjfLYSXUI0Rb5M9WYhHDcRRZ9pw5C
2AXudYv+ZVfo+NLvC3V0AaVsbNWQq72vvgq5jtFciFKQYV7AEXtfHJtwV00dkWmiOMhrTTggZkPY
GXAQjttMo4lSVpJM2VFYmUlNKnchBdGJ1Tsuj+ZrDae469qbT2R02dGchgBQ6O4u6ITTOZm9PeX7
7NY7CBgdz1rF2uO09szo9hLD8XoQLcNH97o6JNfdIHnHqYs1Pi50kyadxzeCniEECh8TiREdbVrT
yKiVynE4jMRT38MIUh+cUQrWZL0UzL0E3x8ooH8jBXWWQRD3kgIawHR5L7H5rs8rFM0zFGudtzW/
/MKlUJjh56BXDDovqi3c/pdy2OrlnGMoGCHI2P9lcERGJuHP76M/Hp567Uw6p/+fgf0rY26hbdME
fqA1reLiGIM7IKhmomrXvU2yXbAmcLp4qWwYt/95f/TeG9ZjGFMls9LtXfxLFKOlELz2uee1GtER
u+5lGhYVoe0qryThY8HKJgzb+9ipWaDWdBs4zCVgwtnHNjKkUFtPFsIPR/ollyJKuqhQaVJRlw9P
uKu5J+lBvHZOxDFIKXkLsU/eVV+z7Mcpx+PIhnabdD+8BxwLS1CzURVc4ko6YSSFrNNSG7dJgOJv
QFWyPfhn0REEEzRLY5h5OgnWZ0rv0jZyOASoTKqFmcJ178KrM7l6vFMc6R+NKNfn0sPqdmFsF9M2
QnKx/wLpelk2jdbtolWCAL6pMlFWKkoGQSNLT/oOOiiCCc3KHPzHNEsOqU2ubuwaiRtwpC+bwzb7
iJNu11Wp3VsPRUNrIFu7zIf3MuOEkuUYnYsBcj3vLPrLnEOkxVtfVvWL8DFwE8IFpM5pKX+s/FyE
tDqrmgYu7xTFfcXzLPFhJlYhSdEcIohrOIdHn9qz6pjrpYqs+K7muNn8KQD+j1I4cqbQHAOMrAFi
VmzIQcezc/8IAS0SJm8RGVD375JkYu71oSoAZahE7DiCWdaXdzC8zbGF1s3fpBDE0vgB0kQXBJ2P
BN54ac3OhW9M+T+ApPCdy4waEl9CuYjR4I7qzAp+KWcwbPMDH37RgEjtFnON1qKqFwoSO+XiZ+Bj
AWg9YX327KYJwOOAVQDFDSuQE1PE0C7otI+cSsrGny9lQ9gt+MBL4v1MyIaqWizcF2XyiCGwxXBU
lEwL8lKa4LC4nNefh1ehQEyILOWn93NNsqWSEu5CfD0wvtQxu88NDJ/S6Vv4IT43ulAX44Q0z49n
ssXFc4UqvAte7i/rJjWZO72Rck0qRExkiTSs9BED1dASkJCeWSCxbQ53/Gt0wISa5c0U8CDaMvie
JFHADjHPuyyLaWk1N/6oCucZxXF6dkd3NmFFXcDDQET/KmkP27PG8l7DuoY8HEJk+m3GixUM23cv
zrubuSVaj1PzzHyV6DUjokhykWSKw1TOInFbxjiJwPgEvxdDS2lKYeo8N+tDqPGPHx9X6LhTwjef
1BcR6G13av5N7xd2CvTUxmmg4V+2ykOOvf0Q9K6K37rGkmB7p4oUdyw5NeozY3E4GPjTVW0vxZ63
AQYvIoQ3aCXqpeku1rL4euxttq+WNs3RJO0xQe89FVSXEkZC2Erb0D7ERWZKqv5FV0sHCfaYeOXK
oEMmyvMAdYSCN/xb4WWcccKqBQ1fNeVvF6aecP55dg0R7Ffu0ykKT6Ie9RK9jRvwsek19KsTLnxL
KK/yho8TKBQghDAoKYZoHryiMKNRH4aGAM3AXEJ2f1nSCC1WJEcqctWze2/Z5Umqv+LTAap5EAm/
taDeUS1GWVZxC0h7NWkrXZf4UvPKuF+k9twlOGxSv5mtwQMRjhOFJPEhCgGRMs3iv2Uo7ne3++aC
g8B733+/WOcCJuyKGCquOVJetzHBW6H6tofWpMHXkziK4dP2ZtiMzx8kEMAzHS6RCxB+3dh7ZnyC
WFtziUbpyCt1vQcC0IojCC5M7P71kAFl9TLeSpBRQnu0xeJkiqMSy/zqlRHfNK/uVh443ZUHuY7E
XMU8SmdD4u7EiIAdS/HvyWx7nHY+qxfVWQseNPHS8FNLmKCMpIVXNskhivOkhqFSMGaA3W5qWLPp
xoG1sEbBEvL/eTPmiwxoaBFGQCR0/h6/ikquS++zLKBYMrBb1gmwq3Zt6g4qPb2xvsMTNXCMTvAh
BxnKtw1KWTgGSmDDH2k06437+3aeWjJppZ6Vj7yUyou8zv78TDQqabwRN/PF8Vl4nGNvSCjr+anD
8UdQjfcCBZCayxU72oV3Nj+zWPctFjFK1bwzGFIdwPF6WeSQ+/07FFbKBna+7zBNJtQg4LzBCOG1
HKivPkzFbB56chY81HF/u/klqL2n0pa9UxizNOjUjEfddbJEkwvsd1VMAD77iKpxREiwzy23PE1B
hFBjAbwCR7aofmjSDUWfNM7DzrB+KZGWzaKgH9tMdFFiudT5rP2pj+KBmUjqtEd0kUO+64mOxrFb
xQRy2QAXGJDBZWN39AW+t6A9qeYV8DV5X7iP3xCJ8n8PNpP4/BQ2PD9G/NKD2CW7eXVr2bBeIsHO
NAHPDiB4ggKTRJS+sbERTabrEiS/b8D/onFYvLf9/AeLJt5wrwHrhBy6lzSuSoetaUfmZb6bGYas
3rgDWntF69Abx1YD03LUwHCBhDjx/KRXBRzWg8Quu6YzkjRxqkGm6AaRxbJRdf9I9JhVxTlquB6u
6VG7Q6oegumlGSjDJeL5VjERFICAxvxyZhgugyiP7yrylNEWQw64g5IYF5PdVlthXA/dYqjRRjdb
bYqj8aVygbQfa7Jm6GtVlZwAreAidf6TxXH6UIPMcOHnAKQbsixYCt/ScE52BaU6rXTdbZmzxOVQ
ophgOLp5+SBe2Gi6cDE9whXIKSqb5HPJvuF3hK8FboyBG3EDpInhMNhgd4lSBtkzesaDWOqYvWa5
oe9+HLfu5vrcinQDjki756tPkgOrWvwzKNgI/B9pQqYsjiKe5nmGVC8AtwxF1lRaTd5mrMVlggVB
U1eWIANlL8CmY7OfpWIz6VutkJ3D2vJGxko0xiCd+dblen1TzstqWXjZvtAtx83Rm0PvgD966GIK
MBYUe2Ra4lJufevX0uH1nXjnx+hM8Ef51k+uLjLDj3fBPzan1DL39heVQnPap3LUFXYwE8Hm0MiA
Bx/YpMyB0F5meBLwHKw2+27a8Tb+dJIH1M+U7KOLTbBSavKEro9oD5NmjXw0cXWl/mFUWbTzI9Iq
Cw0m1nw2jx87uYJV5U0fM9NaGEeg/KMPSp0cGTUmdbgV2WtDF8ZdUkh8oM4SWd5cGS2IrHEYRbOa
GzWfcoLLsyzMBh6R+w4hSEYigEttG2rZ7Y5D4eOpcu6Y96MGVAn6fxmS9narTxyR0448nHvELYI0
MR2NE/V08N2LscgDXkDiSvlnLE4vF1zvdw5z4CFvfqD/wDNqzYmRs6CNRNKlBkvEMkAzPjaxuVjm
H8ItOtQi3vKmA9ajoNglItd1+P3RIkDaXLOoVgn3O+DIqGgBWUxWAdMSlvKb5S8oG2txbK8okO8O
pmhSuLmObdjxdFruKWNqhvRmE4VL4kcajFfnATlO/a89wriB7+uukDtTw3bpnM3AjlGK37VKwKjY
YbgTF2docotr7U6m50BBmM6tRf9PffFen245U4+t1tF3G6pVJnt+TeFKmA6oPvwRCwCdMZezqMtt
vSo5tDSa5jzfeoXR3zra9VGhYyOTXnUfmHaRSh58gZPcUMkzJwfvZdNcRBdtNYEkbjihM5trNwCQ
Bft4EQo0RhUwE+JYFC9CCnF0zltkVSK3gCRwIylbCGhP58VpTYz5CJwuSaiaF2z7YAPmC9bzJ4dX
f7DLTnffnST5+HI86rs6n+5CPRf88mxiYvIvZ6p+k/LDnSx2KDE3H6SzxxD6heS6qFV+oTmiftfz
tKI7vqlCi1maq4IwT7anA8xd9T+FPgLfOuEHIu4MqvE5KWPOCMZ2BN2LXiBjUtL+mySrdsqhV3bw
A4viqXekqOlFaVkjqlbbPdGjQIhPYUZq93h21S4h/z0yVnXwjgKloV0fghoNFZjvVe/5VOsG7UWx
IN8I0xmZvUGHeQImwI4cmNSKq+zB/HCOTqRvu7/1tSg4eqAe+um3hE890thX+OLid+bkyXXUsVdp
9EQ4EK9KsfkdCSvGuMYfGbqPd/om+NGBiaZD2wvwcffqbfzh0kVNZy5S3YqZRWG9N85KS2jPDlXo
r6flAflUh6dgk3tdro6b8CTVZnfRx5ocIWkguh3QCUM8O9iCR10HHkhIlNmdXw1nnrLIsdU4U2ko
AZIVU8A3ahTbYOXDnbteW4/dpv4wvEv1SWoY1Nv8/DoWAGLf7SnTQpboEu3JopGtb0crvpOIjUM9
qrmYKrZ5vsyysYW9G4+kfaPodQeHqKLc6CFxG0Vj2vTxm2LdKwrwLdGiI3lYBrvIlhnwKMTqpFjB
opW+whRYC5Uc3LqRlkYjeGKiZXJKuhoVwLq/piabseV6zZrnIDbbcHc2rKSk/jf26LD740Anv5r0
HpPo2HIFKOnSoxDLY5KzihRDCbi4Kl3r5+vHeIqiHnR5OtNsAIo0fm5RREK8A1IxbYFd5+QCGJXF
4YNdEI9OyfvfCBf1UBJmHUfjT72Rsygtcf50j3qi+llR8hADn4wn6zT7X19grYvaRK4Qnu/6dB0M
3ON+F/5IEM8hWlSmfAWUWI04bXgQ0UHOnt6FPryK4p+VYC4i5mk3cHiB6taio8wfBKy8UY59ibqM
Du/JRVwNm38ouRYusL7pcd5oNRm9Bx4+ggFo6wfgZUZNvWdB/GpjKGfULvFIHNzScekHekR1V3BS
wlNAiZf6NgexuqJ6aW46CzAxJOAjvjYT6UjGf5TRsV2W0kzBxJ0yEJZejaq+jc3FOV0mRWqnF6f/
Lm5g4XZp2KdwrvB//bJsvH6k6pybHv5WuSZ6GkD6dqoiTZDIr7MrdJSnOlRXdOVo+Em4FlVew7QJ
dN4C1FOjNEG9uJoJDrArDz7TZmyfJRAdD414Kc4w2ZDLJdC57RSu9XdYuVovvZ9K6fE+zwQbpRCn
AhpA0iqPWSQ9ByubGlG1i/a30TR0OXzC1obrv26939/JxAVGIm07GN9S4SvONRRtbAmKKvbqYqDU
mVeQup+G0DOcteDzEnXFnodw86UTvuh2vK6JAvqTeFUZ68Qiyx35y7Uf3gaP82KJMQAapOjLEoHi
qdsskOItCDVxEB1J78yuD2XYwI8BN+2CheP6I+4RQgkO1h+VhNzE+AtrqLinKZoxVb2vt0MlWvdA
lK4ujEAHcmYg/HHSWZhQX1Z1KgMbs0LkymozjFlHDlQ3F8V6/MQQRuGgXKRtYSdPxZqAuRPw0+Vq
0RKVg3tWC+gTu41HH37QaVF1cVN1i5Io0QEbS9rD2eISwkOxH2KOuxoypo3OqIJJih+zCyxVZ0iN
YJq2v1920pXCM/wRfP41oPHEZDdzXR1KgESUd+sjYuiocS1sYiWbvXmNHgmxGaXBh2IR5y2MVbeU
jvlwguhgEREr4d8tnVb2hfO4plfQm/YI+5ZR4+Et24pHcW91FJ6d83j0Uh+7QKG/30nWOc5MocwU
KA9Qy/6KMPVjR3/P+V6/vm84dR5ooULxqA32k+cduLkIio3eyyoAHu8RWZ9UZtQD7NV980pbz01f
ind3I/f/Lmr8ErPKXqPLwRcPVjiPr2aACnRmQJxKlrZLgQ2RkXGTlopmzugKQiVaJcEvlJlhaKXV
w/WGthFFBIFNad7RnbtYdRhKMMqZw3+R/YII2CKruzSI1HJJHGkY606p3TZVbwyg8+xxqoc2TwMD
/TxUp1sOVSdU03dbdGOurY02I3o8rzefpfRyaFD764x1BKahcVYOn+oz0O5R9XRLP8JqI6kqEjFd
Mwrt5tlntXD1egaRnXkLA3pJ3wNJ0JjNu0f8yZqc/dqJD9ypdV9VP1wJw2LVqnDKy09GhmExRC8v
4krYalJeZriJLVqL+QEiGUw1cHU2+WePizZFHH0uzjhLGUP2Jo7IqFWIt0UoGEkcdyiP+ctwcoKg
kFY9peUGCgMulfKOMAqWozqvPv+BN2UVdhARJZlOPVBzq8r3QJlQsruAoXHnPsuct3OT2/+0h4FM
suqU74Xan2Ct6rM1+LeYekRj4pZDSfXHjuYn1n9wL5cm5mDTFNPRff6+meQpnJk0TFkqo4Ve+SKT
rEld7uJOYOxcT+eKsqVBtHHc7b/0EpbiYugVre8klKPA2pbTi4HsbCozpr9FkRYOS8KtctBZzFy8
9qHujimqrdxZn7eQ89l41Bwf7s2oS/lJWfE48Nncnl4DjZ/OG7NuiEJyj3czYUsvNKbtJ9duDUxL
lW0mvvYEzRBbzWr4AFFmcvYO79KxVRvXqw7kGHWlGokOZLjsD0ArwGdMImd4DOG4JngZw0DNnYkZ
jo9mefx5ESBye6d5F+2NSdiwg5BgLkgnm9TjW813wd5UxIXIgFrGtTknxqR0cLbMjfKMfPo9/Hgk
5mkaxlK5HBIAiRrJ9v40oDuGEvg5Ffve7nzpPnTa5W1rFQSUHLu3gzIUrHdCwpvWbNESOR9v1PrS
aWAtQKuTSJjiU2geuLF74/ZS117Igp/wDYdDs6eC+Mcb2sUPG17gvmhAD8tHO9OvWnNRPO4Cfm2g
59lrsziYgl52ccMtnvn0HwColMZPP06w8Bxcvd4Q0U2+GrKkgltqaPoLhjWaXWguYE7HpJvMIEcN
3LdI2f6pyI9LBqzlWC6xt430O8zCfG4OCSj/N27+Byginms1OU0yaga8aUnR+0K6BXxJN0mXEg/Y
HvV3iVScwASuWpvKr1K9JqCGUMZeqt2b9zH/5muyQ0FCfHY6K+v5m43Ho4x/0YCJR6XwKIihSlnQ
s9fH1try8UiYTBTH9K74EodH+d3ez+YphYNoLxpPwuKfr2OpDDjukR3BmvyPCZH5eJJ8ZpZ64NJ7
dukQC71saTo93UP21zn7P/eoaiIbPA0eTTyELsyYEbF2Zrm6aYrJF1qGWoKDOTKqGRvwV4vQptHJ
XH84oToDLFFvBBLfeuwnIo8tg7iB5WC4F+P6esEzTKS4dTao8C5WmM9wUFLHPFGDC+j/ZPBlQnf9
9vZMeT0bQLj7VwqH8DSY9VBLsaLX5TfgR4PwCPjjjuYci4RkALG/0KlxqlinHj6v0LUuQpQI1R1s
0SY3x/dWF9NslPg6dzAM9wfnsw8sQzrJIQPvLUOwfjAjXtLfh/7JfGH49ImJrDnUbfOs8/UIt6OV
TSnKNPEZT0X8ryg9eCFVjdynmGAjOBwjSBdCRMpgze4j41zEr1zEIiKN8aPty5lyzzY6eFX8mUuE
+rJnMPuQ5PZJPSoxZQVFDt+UmoR0du7TBaCcRaYyW2/flg3LmbKrP9Bg5Lx9pvbPfCpK6vDg9fIs
lDvcDkWW8ilM2O1+Ty1XnRIGZqIJT2H4hj9PZT6/HQ6cn4jgzm5j2R2oJSiZztMibuVaLRh9KJac
MrjGNrVQB4ANeetkNpv8BNupuy7afdC69ALvZrPB8l4Pbv5PSVKc5VSRQgGYHvImkEhJD5GUyhnv
pKyiY1nMjVv7hTtVghO0AvL07hoDAIr+iKnWESzKNrvgoadXRCXrSNkaZNxHPRIclnvk5BKGaxnF
aXn4PBjTZNoHbBq1yxxA6syVwyjz3OvXEeM6mbv3vX2diJpt7jw7ztqxXk34GBpkqgV+lxMYZIgC
Vnmii41hmfIB1PskWDhbrSfOwF3l2M2l4VzMXuMcw+g3o1xu82RxgYR9J2oDhyx75Q1iy5t/hf/C
Vso2paU3NdJX47IB18yGEjHb9l2qGolB5ZOu+rorg56SbWFZD4z44sKSutaeDIyPj6nBFi3cOvJU
qXI0gK+G5kZzsifdBUGKKSnyYhmwo5eBC65615iZMTxX+U24JSy11B/nqq33MXDgEwN2kNZ7ifkZ
CRK3+nON7slTPkC6wJGdZwnVQCPuxeCsOZFlsdi70j0Q9iOV622l3RmtXaPFIf2jIVDkERF+X2Va
j7Wkb6f19vrwsnr5Q/4NoP4JYh0O7XOWgnW98drcGLjJcg8ENYo58yQVFqzBcnZF5Zrj7oERdVWz
lpEqqIL1waMJqssYPskXXhor8Gszg5MGfNhqLgWtR1N37XtXsmziyiqYEDmPb/jBI3TvUjZa63kS
LU6+cS3mrboLe4CkyKRDMDnn+1m7OtuVzNVAqbx2GCYi4Rwz5MajWcfsYaWaXcdryUtjLPKvgOBA
RrPdfJdLLXYUtLJHRkUoAT9cySt2e7NVHObBLFMhFu71yeysJcY9EZQpegb3fnCQqYXsgRboCPMP
xLulepvhrIPHw7WomVFzzgyNVCALPyxJg4nqoXCdZfWxgvbictp/ymGqHApCzhy3zwrnfWpp/B4D
BO7g5bUgypZ7/8pzJR1QMjjmzUxwoR1uuCoQ9i6wVAZ/ezbd6kjjwOIAkZdBfsxJbJyE38HOwOav
ttfp9/kyIldB52qyxReysLrCqgN8vKsF1XZhBC+dFQcvYriY6BXs31FiV7Qsg7q7OaskhSgpGcB0
mCcR0ou+jHQuUbHbURulzXkum034Fb+pyHtWNaUDUd3KHvOABXXgi8I+oiLsC41mFJLRXiPZtGel
XPTRwHMpDyXqHcHrG864xeD1yy/U7FN06QZuirEwyoM609x8e4rlYEhHvHo16gP2iuug2xt11w4A
/vMDV63gsHIb8Plp0kfWGD8sHRXlDSGnFDHWKYiE/w+sD6tn6uME2NUeT/fzkY4yK0e9BWfbkIAj
7jEPTCACdYHRcXRhADdFuNkyyIX/H68aahBsG/kEW0y2j/iX49J4DqC76r8+tOHDKJCIXLwQdHrW
4R7gzVkwrH/UfqVzPLTqhvhzSEh00YcobJShGvSeYCjiVkvoOm49kqV5MJhd6NnlVVgkiodtSBjR
3vFF71oIQIfEZJsEs1MBbk55WjIE/oek6cCE7PprRS0WwOCUzpW6P9di+RmGyfMH8GbAWclI3uC/
dwNdcCxvqnK8Fh1Fpfe9EOKCG4yi/nAm+tB6oGF4TUXGx8JFHNTmgYb+KseFy4WYHGw3SKkArg86
8+f0gP7JiE/GPqMrGmULdZjqVpt0MB+P8MQkWTtAsLEVwtSBQp1REMcF/N8AAzfxWqIbNO/qPuRw
6BaRJWlABEse00mh7kEA2FWkirzfkuRcgZdqu+hNTSKGkVqPGw1MDE9KpRHxYO0tY/Z+ob0PIPX4
D3N8TyNKMXGd8pScKczjZHpHwjr+oNbJnzlixaaeAnboUYFgxQL5b8k4GS6n36GnrL87pTKnfcX+
nt8uZEspUO2rRgxbyGEOpA+XBkJEn2AcGCNic8I8PGsX4Ra/LBErZiHOpYIBvac7B5F+Q2nZB6Pg
7kARPGdKedjFmYq/hchMoyy0JVd1T8W592uIB43y3lKWgjDzENMMxZzkBL53zVac8V8AsH8HB8nX
Qz50YpsYKLdlqJqpqpvchHw525IqNEtFE64qjJwyJDSm5JOsjLS4vo2lHS+f8TEHF88m5JaslRju
MlLD74kEN6oqfB+pDuSL7ZjpxRisXe7xIXBas/qs0ll0VbDg7Myjac34kIkASh/EYvm6EUcS8qE8
fkqPzEVk7dWMfDmlcjC2xIriJHAqwKshXq9X182kYiA2tA2x6Uk1HO+F8fZhTXxcZQZD18ynOrP5
p46jEprEZo3W4P+sSqBhDT6b5UGC1rhbj+J7760qMs3bFtvWUL5jN8pD4y74U3bWEg6O9z9CPALI
fzWtanIIJJcLlPDim4bWl/7gJbLJAKGaMJYVmp98GOMsCt6aDUsXvyYoZ1TFCDee2w7MCcPVfLiT
a+2N59vuDHRJxrodRuid7EsPePgbZeu3qg+20hFQc71gA/m2G2j/zSRIEfMBqdfZxOxFep8s+sea
FsOOka3EWDlqhdn1L9inJ0NH7/XlZ5YEvLsHUpKMbEq36ZgEiEDvSeMPvTs2RzSozm0yKqYvP5KY
QmhdP2tNk/sH3PfPDTCrqLs1PN0GKhbYid3s4P89BijKXaMSp6c1rxFKQ+iJEeQ3uqlYadOTeK16
y8ECGj40Pn+2Y9YOXAPnQzsKD9OX2OBNhAFhHSV999gPnvjm2rMztfQICs+r8fwy9qVS0RoW89fJ
ltMx/N9UM5eItXzB/ygH5FWIotigeonGIri+cL0jgi84mPO5b49cDPvQwUaySPSS3GUhKN0syuFK
51LeYrGdtTl0fMAO17rWjsPoOUBhSnc6f0dBL+SyPJtMVQ+85JAdXa0Pd5/DR2+2NenxEoygRVU6
SP6NHcgJ2Dm1Qwqnep3V+ZaIGn88wI2xeYJJKWU+mng78C2VB3keI7IqJPOJgSc7cL86HOgtkk5Z
Gvn/rF5IFQMQcV0eNEBDBjWfdVnKpRvwIVm0uQmhtcnfVx+xqql66EiCr2P4MzCU97NOG6HQcXps
6iMOVCH8T31gjiqst/w6unwSZnJCpvZgzC7/62z3n2kmu1oJjDc7+V2YIT2jsjCCCPXIjo0dP30r
ZUhTx/sCWAo7biDAgmD999ghyryw1NtOS6Y9L5r6kA9drkvjYSFZ72VIjKMrdhZybPiTgTaIc5Oe
LD8JWJNoGv1kDwVXe0jEhnXoNlb+XqbVvfrLr94d0i/FiqOXL/zEvi6EPs5Evg22EM8QUP0URFYs
L0XBxwdsyyw1EOIiJOvjKyur6/N7MoSPTB/rEGTzSd1P0FsLwFFo9iKVpf4GD1869rlkdpBNStbl
1zK/m0RNVItqx0XiDFcjITLJKf6CoqWlO2lacaofHt4OJAETHbQDSGJ6ugYxQqMSrFWy0iJA/BTX
lHa6bt+2zTXYg48SfIx0z348gkQdh/qDfbU97BMLzTTqmllhxuzI7yCQNIqvnMZ5I+5aNI6Gm5+j
9yXFez8Us+pcWmHgx2cV+x9hnXJSM/PO1v247Gk+ltCT6Bd+HtB4497uDtoZDyfwreXkFo9nL3Rm
oVpWF7jDjk/EfV5kH8OCWLMqf3YD9qVZD6RmwValLCvH7r0Hy34gMPCwAnbLqkVhQPEG+YqQifNM
vn2UWkeoA/rY6QtgBtic3kjDpqEIqkiUupLVvtYWn927n5/FPDxtkswmPCx3MtZ7yTnRSYbMB0bm
uSlMjZYRbZFSE/4XqHiMU91SAlvw10p8aufN/BvsCJ/KmOFkSPJ6FJqw9+A6Gk60+GDPfunaxZBD
fdNm6WWOESyZabM5y98Vp/njpGOY3qNpfCycWr1HkRVXwo9pVoxSu/mxjaaj//FvngYmBz4Mmqbg
fLsEPjlA9t6kqgO6NPR2736UeG/CbGbztplD5J0A/08Actw8/+QniQCQfVdh49qLs4PRK4beeHnZ
evS+vGMxSQrJJKLuSKSrM/oa3OthHzVKqiYBkhbs5SsjlBatitJEUkHhWAwua2AP/UFuuFRi3sj+
lSVlrRmqGjYLZdtsCIWPxJKjB7w+IvQSbjhcTl8ERgS26DHWFNmURCrgbf7ImuWvjNd2EvCkit6L
F3RpwD4QHikMtnCuMDijDa/UoVKjgt4y5G+DKVQxH3rDVOeqllzm8fllP2LVj324cMVmap+zEokV
sy1yxyP6NzjZv+vzashtOD3Q8vraHzQYLuX9UudXR739jAzZdavwJ9jlAX5r3to1NQpMvnpqnKVp
MDmjbC2ysf3tFvwywGwW5+Ucpjijf6FK9HRvq2kfZBpVjOUIjeQng0gv3oK5WYau3bB+1abkMTSa
SMRrQ9gfVHX5Gmc2Tc8M//6FKgWvmvDd6oHccFCaKte60iDrnPaiiJSHOJ9kPT3Ez0qFy9DTCNLb
WhuWCJgv+V/tGhW5bDOWIeMw5Ugb9SgENGYvJSFfRUpMjQuJbdcn1XhBw+8a7Aw5/T5aXW2a+93n
V6uXaFe32lge/U2zrVbEiraErQ7OWnhnOe4Gscn/ogB0cL9xV8za4TaJaIbwJ2zW0N2WnwCpWI+C
wzNBeePLthE5u5Hl9w8gnTzglfoiMaAKXGT0ezjyXV7jmhej8uw600Vm+oGtpaAdFsYLBUMzY0JV
5aEhH1auK4mQzoBLVXKEqMJzcr8SjR7fLpmHRqvQXN9+nJ8krQRdtbrTwxqbK2h6evMlHEeWzBpu
onS4OozLRkKguTUE2el9GJo3uiy0a1HFfGioFWLIwBGWYIdjX0jHqplnE09NY8rbs8YC9yS1B2MV
dQBxuxU17z5Bvzh27Zo5pqBGuSYJvXInrI/ZtjBBMAsKnim+D0V8hJGisDtF3dMehufSBZBACKyx
SQdeBNs2d7CcSf65mSUQG+2Q8uF8lLro0wUWuabfD9gfnrVrCF2KGfQ+2En/IduRlu7ffguDv/io
d8nGObRwkTz4z4mSbnTPS4sI60yJEBU+21y6Q0O4W44S8RuHqmAnwmr7Uvg0dtcbAfdZj2ghgBDe
BAsm+WuTLIypmLKxERVuB9NjErUCD+RxBOYcs4keJZSL4jLJ7dVa7OaXmJ0VMRDyKajPUrOB0CDB
xoKu70Xcd2raN1tDZcGEWC6/VPOVAJ91lsjYmLKUhYsQdQ/aYdbxvgpE+3U56v8lg/iTMdnB1otu
z+yMZbPd+rQhqlmw++RZrhZYdrOWuqHjoibZa7vanu/yDcCqB6EruQgMumcLYsyY+B+xPLfBjTvB
Ar342SG0R/8lln6C6ABOt3cqaYw3E4osm3pJ372mVpX0IKU/jl1yLPGiUFiH6SRpcWEUcLT6b8v3
PVIUCshqSdaurq6V8iLj8/+BcP3Whgs1HrnWO7EkzsgDEHslp/K/5AewlnPoDS4hw3hkWRRkuCOd
vH3jSFCb0g14req3hLdNkHC0gcBpCP1T9MW1kJn4PEJjv87HorZD6Yn2fAC0GsS/jAh4PUGlLDUP
5gYI2pytLlXkTK9DBKInIfHKd8cn6ar9H93ORCdNdkHQxSQL8nqPuwNadvyXS64N+xk6HZ0EDCfJ
PAdDZOvVfxSRujJZHnFQZvM7QIoT3IzPxWcGxdeohgzGd0SvDc4nMyxrvBwEoNYbxu9OJ4DC59mN
3pN7qNaAlxWtlETekc4Jml/P3qYCId6SkBKmL5XmVgX5mw0A8Jdx1p8IOZpBqPblptP3nCD3G1xJ
IYkFrLh55RzJ9fPsyMajlL858ZKKukX5CoPL8rMPKRoFARY9TxA4ngeDhDOzMSQtiWy4UC7TIRU+
VTMcYhWIyO8EpYGRghlgNKXamfzKsEmMijvofLMGjq0oxvFW2jBXq1SpPbcjLcdaLLKtbdEEo+GW
zvA3PWW3L1E1j4bef5FdU/pksF5B3ZtOV2aE7btmIpsTFqIu2BZZQDm787LjgDIV1FSTpEXb0TCq
8RITR/d8UpQfsYE4UE+8mQ8sFivRNRRHPMRojWyt6pR9xS3U34wDULWx1+STgNEjPzx1HaIls0P1
uB0yvvv3Z1pwuH5v9CALFdgqMLtE9udJ3u3ykEV1y9xuHbh+wEcywrYZemZa/corZmYelQXDgC0Q
t9fXDl4mE10dm1ivOMthwFcf4nhQiiFJTx0tDaBbrjIBQv5+bVuAX2m/NwzL6BtFqfDP1ixLoZoG
TyhOqdBJKvPwEk/R8+A/nvQJkDHL8rNLORULsqmpqqmh7MCjzGke3qEYr9idQS8zz1werqo30rZ6
ee5B3TVse4UiLdy8p/xJsZ2w2zzDza/AeBChnDMaCSMnnHu1NUdgyeCoHLtZgLOAubu3X5OpkM4+
FDTtEpAjIbMZNiUbkdCg27Tyks0Y0dsIDEiu9o4rZeaeDzWMZrGJV9pe//E0NZ2x6WEk6do7Wp1a
ZvWHBrvSKmQylcnRHqgWArsg8eRl1eUpwg+Cez3E2HbKg7t/taSBYL26JEn2+R5JNtxM57vUq7zi
2Hc60ND8ci4t2MesAMvXjElL6B80Xi8SSR1tAiPltGCFGJRdUxrT452G4b1BX8ZvmsgfP/M6pOPR
/kqnGNA3Y/x5F4dkeE4eqr/H4QrPtiTJaYomHi59FgwIP4TeuXNafwFwFY/F7MWcIv2VvC4AyRWe
z9CrpezDAPP6m+1VlkCveElMrk6TcHq3X4hz5hklawlwm1N4pNY/R+RwQyWTcwLURxr4E9ogTUVU
gKf1gdBMEwh6L3r4TtOS61DU6ACiAvbAz4B0sV8R4hXcJUN2gOtpwpqClN1qc/ORWpg8OlXLdNRf
BEuZMn6p4lEJXlmS/uR/htUHaynqp0qMAmj/XirHwiwyVEMGm0uXViXJ7W64yI+xdb39MVgiSClF
65WJgOGcLnK0I+ybh+l5p9UtiNTdlpBW3KxwfW+rT1Fh8ukInjyGVruAni2S8+Z5Dn88tXoZ08hN
/PKHJZDoPC2or5eVaZHTRV2imzT29bmzS1eA5V5gtBKqOZqkVdZsbgePKIlZlDnxVl1JKQVEJqg/
kDUlHryZ3z8kG+YTClMfMu+B4yQ2x2f54o3yFOjrowRoGwEv90ggfBCv8TeY5iB98eVLu7OWLR3f
5BtLn515v/xdXHmwLrzUarWDb58UqKAJKnEUEN2AfDjMeHDA5Gbo9iR+zXlnxdY+1wA5S0OI8vhD
heaIZOXdoLHTAnW/M3fKJx1gfN1wbe/d3NB+WlQbMWsEVIZJSITFYYM/eofsgpd3qZYX9ivLXX9U
xURjAxH+B3qrFYGdFLDYAQFbEaXYQeoGLHslE/E2T6T8HzbzyK+ssgq1Adp8wvI4xNFeoQvkGPJX
+cFM6Nukv7hJs91ExvFjtVZobwJA9OuOfivbv1yzS0nR2XIAhuDaeIcx+Hpf6UjEolv3FkpX3p0w
eySNfN+CqnYfZq2AHvRpb1taDU3rCKASVgBLGPy9zyEd40yhH1yG1SkI5qKhlm6G8PfZ7uFjjyzX
+ROBo3clvYPnzyagdU8MP8is5JZU3fZTqFekY1aDdCnk04hJ8TNL/QbA7JgkYAAlK64HmIpxb6XK
PwKLpyGxFdncUNdtonJhXkpQTEeEn+yqi0LkUQeMOvc5BKkG+DpbLlwt27MPknJ09kisnj3pLFMf
rn0fquMa+D1S9DevN2eX1XqwMcen5nSwFZsfMcpcvjj6HJHO0YDte6HS+BWWjhtzh4eTI/DiOC+k
ZhLYq9QXIwCvnUnzp93zIuGvI51L4PElgR4vC5ppBuGjRTRayzUUQWeOQP5PNWJxgjoDaDunjhJD
xU1yub9sf4z7yHSxcOJzbG+nlk+Ma3kXBrQP8vUn2W+vf3p7J4sxTZGweo3A2gASZ7v8Ya8HKdlo
Yq46Df+J7w343VM6+JReWSl7NurKg7ScbdOR7ObqYHx6q3tg3Q0sq5O0yv8dE58HhQz2pjauhfHi
ZX58VNBW/tshvusPbYPL2pZmM918qJCMFMMFtBmRZPXpHuM8hIYP02L/yZEZ1fmJP4UeXwRsiR+J
Ji1Wny0T0goJ4fI/SgmXa5DN8cSDBeyLz8h2Wz4lxRp9xeUm+ihI/5fUq9Axw2a0rqel1/aTwgls
w3OFEDtAN2RpiSEafi/uFd86cBdJLbziKsw5QStAhAibXYaMFbjhbVqPFkR+fm6sjAWfcxgkNuAk
goPO+NsGJyUBJlhvH5epiQh0f12kOntQDQSZIOlf101KSfX+1HhNOEAUdxzEht/9HLptTRbvbKDF
r1hcOuybZoAegwj4Wi5hiLGqZPY/hAVXoG1bsu+S6ktDex/ZtEqdnT3ejDjRj/9qQFdhwLRAK9uL
4R6DDBlTysl1P5MnOM1JneUMpQK2+ImnLd49JU9YKZu3n5GpmXWVmLZuIb8aqRSUhBswGzo+CcQt
C/dCfm+YgcXE8zMppfJDBicHBdGtRW1KJUe9bhrEaLwrecTqQTpJT1LIuoBD7O60tXN+zPMyt3/k
tFoF/3PLcmu7WtkopxLyQ99BFfHh+dQTebovedFIfI+Iqqab4FGdHYKJGRXgKLuvbt76LW/oisxV
O3Vum/fZj0qW0bGaGHSpZchTDLtjBFQYS9NT8QLnn/y/IDaXmdWEu9x9Ai5HwMzZAWwSgc7pBXXd
RSuwEjZw1Wu8EroAJh8+zGUOx5Qm1zpN6Uvo5YXJ0+j23WH2GoqDQw5nrwMR8C9R04gHqnyRl/1s
1q9dXDCbOt+u3BTPGrK7MotZzWmCNg13fZpoEEejlnjebTPRJ1SP78D8RaX4SRbQujbSFPAY8g57
rodKhfDf2MxZEcUnRD9AVWlzgSDwIltSkq9Bw6sCG8uO8nsulmQSaENRp5rBV4sEwe/Hf3rhtcHD
818u9Fr5EUI7j3YhvPv/H/HylX7vOOaECrhmxvjwOnC667rA5Wmy8gUtKaEdwWmbc2F8N99HGxgn
+kwF5uK2+RzBvpINBVT28k6oF7f5Gci/DZR29IeDRhUR3Ks8RWac2X6qFSiUdSEnkouCTtpvQQAR
V1AhMLJgL42+LrYE3O7+Jlx9fTATOXarHlKBAdSPk9f/57jN2i95sl7XFEu108U6V7caXpm2So4R
16nK1YKEWcY+RxOR+rJZGL5haNvrba8FoLn3No+zvcl5ed/eG12qm+OWvFPtwrfogSQG82beoCCc
PBfOvU5wucKDw89AcWCE026biWePpPBwEGdlhT2X86UE345ARm/NE00qoCCX1b7Mdf151QgKo+DM
3esuSm/E+ax8gNb9l0GSUfjgQfv2lQPEhtPneOE7cabhE439TCaFJ0T2m6tAw7YIxqeN4TDJd3Gw
0EkXBjrVJOe/ctUAmGDbixwmy00W2nqIUP76EYxOrzMcWfmyc1Ln80H9+FZY8scbsLuhV5XJ05j+
ohuLW7jBPogOLUyMDuuFRqzw0HHIqVB7Kf0sIXK/PZ6T6qhuNQvV/HZ58azErm5gzxQtt4Kxgx9P
G7AzsekzdSJhpTuFhJE6PE1xjgvpk1BZkzU+K8fqbhI+SpX4svMP1kc7R3qTdrFVhemCQHkBBjUE
mhe4D0uWeIZb6o7mCbdJsIv8RVVtShKuIIIOyRyfPHdv+QPFAs0OXD2PuLYistdl5cICcOpgS08b
bI2sEYwVRP396wF8AVtV8kFsVD6I5uU/XiEA+zx8VcX3e+5YAmYAwhONrizI0XRT5Xfo8b0xWb8D
8dPoN2A1V1QnnOH/xzLgsXJdIhA4qj1X47X4x+/Jzxxpc3x+R2Wpz/t43Lu6+xplFxo+KzArYYWb
aejmO92ovrbuOrZ/OofYO35t28SJL6skocF0r4twyi91/EK5c979ndlw5dysrKl9u4mml9SuAMio
5fVDk1PRBXhBkVhSUro7A/LtELoypTX9eVuc+1YaFQvZ7oI0vlaTrWR+wn+uk4CRSoPOicwLcfvT
JMu5Bh4ZR+d4gck1wP57JCZLkggtM5HCVJqFW1BrOo30zBnKtKfdCQms9fu0TL8GnRRvOLrJKazn
eu5PS6UIhsgoGb9CldtLd6F+zQQ8iaoRfdj8KCenfsQKFyWFLQfkx7CBIGe1bO1fwqrbkx8EbOCD
kvxdYPd3sryZym1XTDLGSUg3pjy/L09jT68KcHl6T/fk03unAgS2Zl4uUIQfwbn4im5JWzHPsVu2
EqnT+Q8ti2J4EPQeX65FRloWTTKIQv/Fkbwvg+vBZMANI5QRoRMrEMgsEmyiyFAYQnWNwoyAkwvY
kdMTyUJgUxerVDpTdyHKbpzg5rFaUvvPV2r3ZRdZTjqg6h8ZNqIwbQRSlJbe5lafnQRp1TKR+PMd
eThIez9vja1kWz7zqVFR1G3qHWStEUFw/vYSlim6J0MqihbhQj4J9mH0xJwdm/dpT3EUhjiViuVf
1eTgFPMWMIRRC5zPRECOLnNsOAjRIBrsjCy0cDYV17jS6Nsi93BOruhe4Nb2Wznmdq2gpR4NwGp2
ZCqdDFm3FlrQpd8/ZKePEXG+QSGbnyaywezUpyxbUVdEsH0oJxHpoj/R3jsYNf5w0EW+qRoyywkC
MB2tajKXVE+Dy7s4qn9VEPieyeRdAJtYcUUW/CfFfG5PMFwe25O+JLlYHV8BL0yo8EJNrPxQ8kh1
l0mki47W71GyWaXArtR7QesuZl+zWzltHpW/V5kE7kMDZqbwwjDyT88N+kIKczWG43jsXP869JlF
cZYwYIJoz+olBx5LMJ1v+ENsYHUNgpTuwSu9tPuQSTIPMQ9Mj3wW2C6+oIHKEX9MtfIJ334Rayo2
eLAix8AQ4NudGYkeYNmAMDYOhIW+whO+Uo1+4QWDPejI79cuv19S4I4gbBMaMiSJcbb2hh/1ziqz
6LcwSBx8Ulq/B5uOs25G8shMyh/S9JYptlhk0LH1rUMK4DE/b2oRPg+7S7R5ZZUxalA/x6epc6w5
98kvPwCLXEOO1VXNpPCQ6D/1taerxed1EoxO5HkfHZZB3dk18mxCWjRMjfVIuJsfYoJ02h0hgkDO
wgdFRIi4tETGZ2Mm+e1DOB+MvArBWuar38H7Qgisxhb9vajzrAX2aFyqEh7N2xcB4cyCpm/k+5wW
NKEk6iDh45Urfe/nKwfVqmKiLDZ2cYgcsIFMldyos10ti8E8ux8U+8x+StkIRwVzlTTcBmfnkbSI
XCBHLyvwqHYCNn0LEdMNj86neYTELIm8UaLtIsHt+Pla9gnxCDRz+YeRW/MOTu7hBcEyzhrUtJs7
vWheZgEcxv5zs0HT8qangyQtQKTMq+enrJ9JWQ33bdZf+TJKQFmUBovSDbE7X58hHyYwMqWrpUs6
FnELOn+GgG3QlxZhvt4YIvEJcZtC0ZhjGcYQQScZkzGNBXXDv75LZpVzO47JICy6V4UYkAI07k0q
fUokxRbHd5ctTBIle49vUOw4i5fpmbFpFwyBsEnk9jlA7h8Khu1Xx5cqk0erKivReD00fd5Br7AN
dzB0dvVel623QBF2lBHH7P8pCul9rILcXNtPf0gKc1LivN96392wlNg87AThBdl9/sqQ6V902jiG
gs/wqBMQ9W07aftxEn5Hx67WVYwDzIHN3pFt67rhzmWeFMVZgael9pppzzpUaaROSE5QUXkgqav8
hKJxZ0s+NtVTe35FBgp4uC7+5I8FZMMm1izUuHpl5Ik/28MpwyCPPOr7KdmYvzh2/TeAGuUH8uAC
/0WIeK7ID2Zeub8uZnmzxmdLmKkA1AceEJlC549m1E0JXABAYanBdhf04S0VI/DWV/te3ZAYfmSX
Bb6HOsolouit7avL/RChOBDq80X1nA4H4IQvPIkN5qossZ4aZ6tD7gvjFAlC7RRO8vn5+OGGZSX7
bPHASHfO1RIlB+NADuhO2tJ2pVuJAo+4PZwdPwLEMwD6Qthj+evShD+A/iQlpWcXwACmVw7M+E+5
J/iO9XGL5PZ7ntf729JvAvmogrg8zUF7c1KKzYwO3ZHpfuK5xQk7uwe1dy8EdHMUC50lbikYa2FA
shgWFLfPHNZNgA72GKk7zaijsGvXFb/ygV8DX7HDTL/xE0RcBus2inEUM5LliLZylD7ZkdjK8sJI
rctmcrvwZoSxJDPD5q4QuF/0Iz25GUTJwEYDT5I/v+iixcJZCK8WCD3cudwx4GKWUbTRywp0OMzL
Yd6cHoOMAsibgMNlWu/wh7pOwYITBQnlRdmLgbbjbB+Twos4vtsR69QOO5OI4XmL6weJHJyB456F
llmFVJAvxb8TWeS8506/M0HeK+QjlVs3NpeiQ+LXPStUlOfID5r+oQUvvtfAABvjZFK0czlyV908
GsYPyqm0jfpH2x3S8QMO29a8QnvLSuCImyDv5thgXb2zpmW5uJXbhgNGmqhVu2T/Nv00EsELK7Mv
GJUYcvjT+gexV+h79T7QKlLooQkxVWErSnS8uxWCGteYIj6UCV9NIvXjmNcFRikA4xVSlvzADICS
HhMUSjvKXzO78PJXpec1h8X2IW9nLlJ0bfQDd+puLhD4Sz26sXzHVxvqb19eMdvoht0r+yburETr
zi7aDmPPAzG4zhTmFe7D55vsq/wspJWUSq7IOXMBbZ6VnR8B0aoESrfNf5YvlKy4ZnAyC17vfYJN
LYR83TBEW6ZP8DKb26PDSQ1s32DjVBJmuLEZUv6CrC9QrwIyMP21gXIL+8KTok/Oot0dMZ784dHa
30AdUg8bOyqfajLQJxQ8EvirHzsRj6vRWz4ryKcU+Oj3/53DiIJAjEaA7OJmXcpN1qvViwNcTXrq
5q+v8bJyJxhf0+QMo0xqUKo3HbOkmy1WgITBXAK4DObY0ixK8cR9TZ/fACmq0LnWknVd9s4RcaIf
ZpoDyhLsl4GCgVHKHlgpVyESuO600K7uBeKeogJ3xKSKlEgZwi41758w0IRfKfCeAG/BJ+KNaKJX
DYDDBSwLNOPHhFv+o7XdfsAVVMjhJEHJsLD85ouZk5tC6DfLAp9e1xIZHtP+bWvCO8bFeIu+yRLI
sFmuL/pfhOhO4a3/4f6Gp2zjn4k5UMACG5gQcUijsIwxzTbTPjmapYx6dYSusn9p4k+n6LYWOXkQ
6kPYrf7vSkcCYpT9LEXjY7rWwIAlOEDoKIxdZwlr8PUhEkaFphzlwQrDG3Wdl7IvefzlQIDzzjtV
BoL6y4nMONcECai+6hl94L/sT7yOyniwn8vQhzPZD0jugxb/Itq7YLF4/oCWX5dCGGtn6WqLL6rQ
1V077YNvbvbvPkBoBkX9XGZRETwawgLQP4uB+3am4zmWZ61MbapaPa2X5JdIJCeYXzahfxYsBnwB
ARp1HtPjywkys4wK9hCmZT7ed26xcms+w/T/g5VZnkdKoudmv1a1tTTWBY4LOHSPmM3E+1bblVrY
q8C8/ASwoDeKBtqbGVWgoeRt+M5zyx7IPtejs/lqf8mSnV57iik4qLBvvrBapoZxD3537mHDBREB
7MlhUok914vGkDZQ+LBaT0JwkaBB/hGf8+7ejpefQMf/n6zBbYTyWkIznl8FiOtgmZ3wz8jam6Rs
JHLAd3A76QqcGHjZd18V7iGQjqFiYqAxeB08GSi6xcBrlQ/QrsL/rMOR19NqkdDkn/oEBiJhxQ38
Te2y6uaYIVOe7QKGgUecRrVz1vEFwAq3LhKd/WCQCyrpTyl+bWJkLert8wkmL3fqZiq+Et9nRdHI
mWDgNokZiZhycuppL3QI6g3J46bq1+TjNRXnwcM7lQSsqlt6NgnvJz3g9zEe1QIuSz0aMUiCsYA6
hiY0YXptylXxuNtUroHrNvaAskCtmd/VK2gIoIND998vb6NpTuxm1D7KTRBrKRmUFdHi7Yiu/PPa
XGjHlaCuUlVQUaXigKJNACyDqUO5eketEmVZNdhKTpD/6/Zxb/xpnCKAP+9dOqWp0ro+MddIYTwi
lltIgueSQECVL2X5YpGrU0OH7uDtFTIYTzBLmqAy1hVwvjosIqN3YdFbh7WB4c3SkGkDmQBiM8Cv
vQbmPWCSMSufxSXNrhMBQXRQolF4IrRovh9rdqEbinAuKqMOFkF5qWZQMCgaLG9yGPVE6bG0zuad
hEQdzg8gx77z5GokI01HNuhOXzg1wpibYHvLZp0cKW7P3YpfdxSV6F41r/DPO6Ua8J4MygTC6Ia2
yEXyY0zZrcvvhV6sY7hSZJPiQquWCtvOYTkl+aM8nIqyNXcaXzZRlVycpHKiwbjjMMu0lvsBcWuA
/hJC5oEE4PasaFLvCr8JrTFY0EW4IK/Vg1+Obv/LKg+s9H8PW7+TKut0s+5ozGKY5zgIO9/RTgEK
ufPp8V70+dF/9XnxaFO3Oc4JUtQB46DnOFGw6pIFftCf9NjT+rGRsV4WzUDDHsFAclH/wghdoxbD
AIlLowECsQCpXW82u+zzMWvOoLtqhMZJEidI/9dCAFHk26EbHzSTW8BhnrqNx0NeogGR4X7qpQo2
xjjSMKRn9K11DjjizYELTuMPixwbjh+eE9FNUBnBsBOxyaDhScARMxhaYlHYUWWrOPlThVLm1+Jc
tNn/esuF22UlY8EJMVieZ/T6RglKyXxXEFdYBJefvf6YKMQeP1JlJWvY1r2Eqv3ZSEoXw73Pz7ab
h2kdceQ7/mVCyqxWmpLMqEUGY48nXvdIyRlSJbxImQ+8U+CGiFRBqYF8xpt9sgBQO0loNKO9Sj9u
66C8KNeyYWM68CV/DcnmHtUsDAHvl757aQ82k4oSGv6mNN9zslw4QMVEwzHU3K2U2YYkdSpcgSqE
qf9Sr6nw00hZg80oU3wDRR9Ww8BIoEnt0OOY86VixAI9XlCZOuTY7NcoSGqlrzZfQ/KJsUtmAV/T
xouNB3xoibVmpwhjgeBo8VHfy9In6wwrmU0M90qXePzZs/RaNct5X92lR17KzOkiTs0Zia/Ja5qm
wvJU3FitMnFgMJ081z4DAKh+5bL/TorH2gN/0JXqkz6344/BoL8WbYGFmP4/6ydi2ICwrnPBjGKF
CDUBGY2LWBORihTbKDuq7T/kxnuIm7WXu4BHefsUyIJGs0NgaTYC6dfIAI7pu9yi33grqC6cN+/8
EdRdqo46uZW1ucK/HHx8LSvFrsTUWY0Rgf5a1kE2VCtZiZLslAHH3jM9445RLcYuhldeKsWT4O4r
6CVPAtN4PbAu3Ig35dTdo4ny3UnF9EtNgfL8Q1gTlHGacC4Ow9RIpXED27SfSFpAaCHiApGcZ0Th
uruCvNCz/Wx/zzSiMmdDye23I+StOGIe317GKMxLb1LazZiJ35bZJW/jn0hPSVK997fE/JvXYbWP
OdNsSsYn1ZMPI608aQAXwUnnfZGeBq6DlZnqpcC8SWcf529iDahyBnbPP6Bs3IH34kmSP4axFBNp
0XJsMgoFgPQbk+BjFCA19vGx8CPf/7Gbj56hovfiOyWa2afYCR/Xlp/qPZc08zFwhjz3zLeZHD20
d5XnlEsyBrK8hs0HQBo1Y3cqI03OI7oq7ZwsjtgZLgT59ju25Ck9BpLBSORd4VcHlEd1NxdLYbw2
0BrwXcCDkS5D9x33tyOzjL0LGbw/6LPNoh81b20/YCeHOecV1DNmCBEYnBtmQ1YrM/7XMAzDG8P0
ABdEj2kYOZxN/XEojo1TNgPs6tH98xkpjjonPMp5JMixDxEiVqEiAHdW/6l59Loj3g0Zkx+RfYfQ
2znQitpcdCcCk6S/jW37W6f1u0BonPXW0YL4kWveWScJmu9acKSUboO8pg7on8elTjHYZBlyrWVJ
LeXcJ+2PHU6o1gPFlOzgqDgYH2pCtdSSDR4q8f5l2jEeZLCaupjvIirOVmfu9OqdQ0vClVNBf5L4
reDluwBlhsGJczTlGwMRkASjWiVoiVUC3anoXpDGOL56YcO0/TyG/T/XtSqe3EckKOi4RwMvUHBi
7zDebHL85RQra40D4w4/ri0DER8dfoAn/TBpFsai61zMjv2O+ijrmNEvFe6lCLv6OqEGtvAnsF5s
xnTOgt3MV6jz231oWPKpbvORSKBIt8XM7JEYbueiniKRb+640IW5MpXYYY7Ht8D4LyuuZlEtVOXm
l8hIEz82o0CtYIdjqcqSC+uk2hMUQhGDCJ0v2oT9LubMh7fwmhtYP8FRxOPPb6UU6MCeaxL/ClrV
whtKhxu3jMgAmhFAUhw6vvIJk7KUZ/p65QCv2h3LiCti0SyttvjtuwqRh0IxOefPXZ5VnmV1aLo1
w32itN1FCuCpNOCgqtKi6sLPRkP0DQIIR5xUlWbrmwRXDRZH1BKxUHICLWWL8UazcahtL1VIKrLJ
wxiHASX4ppldFmnByIabTShKI/lsgcBrWFjEdqX7qs29yu5TGIwfhKH84WYjEKntenIcgoc+Qdd9
3hW3np4R0q7CoGSHqejbUpuZNUJMUwt18kAuvdmCHrkb9JGQnKkv3uR77SjJa8iVD/qETlddruha
1HLQwURjAvvvsbtMk7YivpMBFW4B7LLSGEtgxDimn+blwCsX5TcC70/PANefDJpsxB6WzP3gbCDQ
qrHVfeNV4MnDApI4Y8LaT1dKY+ub7U3Wry8vE8RbHw2m/ebvxAnzNR6kLgKbQHgglpFrE+a2euAH
QcORuinUq3ZEHjJDQtvrrdmAIzpmOubXMFfW/tuE/uLemLdLd0kR5iDEWnHq4u7elGLup+mT5muw
sM5bif1z71DtRRmnvNzR+1YqA3vUGrG348dyfCE6pSNAc7NKAi9vPnnqhkEQtU8eAhot3IBVBcH8
2kmqO9hAmzSUQHONtdDHLug1sUg5jXkpdEQfLeNXPl6TwSZaB83If6J+VbOvbYDEGwOCkrpmvlG+
hKiyFdmbTbf5AgU/VpPJLyBFExWbstZWYFmNwDgNu9lFzcw/r6aDv6zVAz8vSq3z+jQZRNP1ozIS
CrTEM415TieKzVNbleaGh2Oo3I5re3CvmBEa3WErVyXllPgdH1JXqnOFcvaeStxQQ3G5FgErvB18
NkfEgYlpU1AyOqlPUlDR890nMbb1PbI8cRKlhFkTKMtpi5oKwEiDpfNuOhk7ing+8d73iGUmhLjC
WfcXqqkoFo1TwdNEpZBaqquaOQWV2jqBbtOdKoBruECfoKBFEee9DDWplO23Nkj1uRk0g7RCIzh/
dXv/RYvu814GFuo6Af8iBDFSX/FYNHLO6UVsCKYwgFyQz8+hslLDzegcXD0BYPwkOeWaAZbR1Nut
nLy422uELv50WQzGE5PaI7AtcGgmm5xmt34VUejqfzX8InjVKFZBID44AQqDMqVABUIq8ojHXUp1
DEI7LS8rvM3L21jYMISOWG1EwWGwIDADeXFc3Kbt4If4uj1BA8JwcEii3pLKrmgyZbZJvw/IZsqs
INxXWY7+4WoH9XQXm69ch7VdKlBh8ANhq3IqPaNXTJe/jApIAfX9KvReFuvuYydLhKWbUYEJQfgL
005unwN2gb9NL2Z4Cb4m3PQiw6uukbLxoyINLdmhQga1ZuEyaOH9biWu2X+avLTqDeC3CWf6v5TS
P1MJONEh8r2CTeMs2Q750k9J1V+WHhknk/1ZVfJHBChwynbQE8FG8vModxA/ZYCOorxjYpSmI9m2
Da8vDsCxct5JknzGPx2R6qlB2PvEG+j/FpLvkfZ9DMWUXtUAkeVbNyZlz4RQG8bpViz2SZDqH+s2
VZj/xSBRF3QxE174L9wKVqnlLBiChY0nM2Dr5FU2Pg0oBYDmul/9CFr5LQ8WOzaCM0uVlmxPkpg4
zqVcXs7j7CAmTsHsYtjMFkVipxpmXT5tqbyX6JX0PQ5vssXRTIXTF3ERk3qqWNKk62xEhkBz3VMt
y8G0HNbEbmtrXfBV5pyeGafXGlmyi7C5UzxUZp0KC1YfeE81ngvCrQGYvf7KheXwY8hdGDT/0JtK
ClLttFRDhJa9A7RzXRv04ERv9BNwiipmZ19akzycwijB1sW1MAWT4vhCNwjvUhncd6+aqJA4iHqv
wmFMj+PtnbEQhpuR5iRQ8uFH9eAlABdZIF+AKeo7KQ+YrBsWl/KcrMcvKyCknVUPC/bB1dvxg6m1
3IfG9UdYzNDKGxfpeyFRyRPZmyD2N1P5UPUrfusyZJNZe3XlxwHazyoFjLzNsd4IRTxzJd6HLRaA
Mnpv3GRIFWRqTwhELar4Az65RIId0vqHsReQwzgyHsZgn531RcYIiENS93CUcONsrxXLqEGvrDEM
lPzqf6sLPFy9l7C3jqPEebRj8d3HbCBDD/FTnRsxlHBE1tqSsK7VoTwY3g3H6xjGLc1ddqZT3u5b
yB1fNzNjMCCGX5R2RgzFEwxPoFeUGs2SegCXCHP554X82cHbSEtBbnshwgXPAl5DIFJFRg9RfVbj
lMEAgfbQgqSAO4QAQkx8crlbp1WHyycDUnBdlbejeqmLyvHrzgfVa6n9/ri9wWvoWI2J9bNe1K/z
lOCldBUZnvBBBZyGxsMeDVqcuBvdwfdakRHPCfbEWRSlOxSnn/zvtYiiHucZOs/ymVCVBC4osUsO
QynYoxnIOZ1FJ8zRVMsw3JIBa+SDUiohUUBzAaJ72QmbeWBvLY3xFwLN8PyAZXv9AGFnga01qTqy
nVGNU85KA7WbfvGU2k09oEuLaN47IsU5OWMq6oT9sHzKFm5KewF9AdCToFkK1SyLlDq9nRTgb6uG
Uj4FOqX/3u3v5RbB7ivPARbluW+AUXt64VCJEGr1R9vioQ8ac6H0tBKLOeIQqX/CrRoVAWCTSlB8
dW28UoMwU6hJx2y5/A+zNJ3i9ITlGQliJlMQdt12556Dc50Xa0jgzDj07xS1WLEKZkcxeqP/gZ87
FkdWlmPqLPINBR15uf07F2zjyr11JNWLOzeohPvyYEEHbUvLYnFS2rHUWogbr/HBYYecvXiVmUt5
Cev4AtN7JlNGc45zM2aIf5fdgFr0VZPWgqiaCfuFKAwaDw28sp+qraFqTPXXJqTaVI9vBhGUiybg
SJ/xcAlAl7Y26RjCsa/5VsHkzh4gzDCLXmWqTSC8c0pRJ45uQToiEGCScMwCIjE35A83Q9vpRrCe
V0FdNf8dww88zZQ8mE3l1uqmwL/cyaRsxKn6JLflPRr1j5rFOokXGwTeg+jKJlWekUCSA3zsTK+u
IAoYcC+0u14fhdLvWSq1FJUJzF2IJePJvEzdEj3CIDPtMyWkJ3mUjA0YKsMKiJEF8BqlGcZQNV9f
Iie+rrx/KbOH1cK7lzC4ecxVkObqT0JG9FCtHJW7wWFRNmIbOHqtKzRwGp3dUDLgXkh3ei0qhcA7
UJF1XwNGEb9jUToIbVNOa1PnT6jGA/4PSGVBZ+vZzy95854vL3Fg7pDvVoyNtloYjcwx4pblgUb/
G4YcLUDe9gtoPuvQkbbgEaO95PcrOjlDT6asisdgRWl4MytWjnwIE2qVG9zDTHdu3VPJbk0Bfyna
e/nO+8/GN0tMryCOMPD/nIwWgomvxYY5IVxA5f9oBvITGJpp1rbiNd/y8n9SOtFRkPB+ZuIS8cIw
+vncvwgGzrgVwIstn4m1aXIv3B6n+LmPQ0u801plMU2LU5dtbIflT1xR3JEGgYA3/iF7WA4sW6Qf
TwT5kmUzRGGUNDtAjM/lpW+B55K857Hi06tFC4w3Y3ldMckkeaDxubqeVSP/mb3b9J2xc8c/1sRP
UneLcs3EpdYEBfkOKXPzX0YLPG63hd/DBeH7Qkws6wytuQF25Awavmr7pUAq8m1/vtymnXKR/tbj
rNIfqcWYedDHHQiNWuZCZKHxEDe9OETmpTijLnJM4yHb/vUFIdCMWmqD5TnCq5OS7KRhNlWvpLfP
XzTtYPAI3f/mL+jbHshrtHQb1Z0pErF18WeYiMQ6rs0rpS3v+V4yzOEV2C2F1X2SgWhTPZNR7nPi
wOw03cRZwQSj7vRPGhik6NniIvcD4zK75YwH6sYEh/2DKGPODCltEmxwI58k1S7+snENqLoc3ISD
UwdZ8jEUxKIl7A5c9oNOTuA0dHTA0vY0hLAAEjXM7zqKurmjvXrVyZ6K40bnZGHS2z+5xcDc6rHK
xyH8wPmZOvGa9CD83llnBILQBs5X88f08vTNPenZvA6dgMUR0i3DHO1h2Bc1uSc/Cj8kvap0/0m9
P3vX4tapg934K9L3diiyhPy8tYtf2BdZUHL7wgP3eo4Eo7YEaB+uUm8Ko9Zi/HdhCt6B2c1NAozg
Hu+Gfm1IB6m7RTYniq5FX3DhrqtH5muQ74aORNUu8F9dJGed7TmK0ieNZlnQ7QThNh8MDVD+xU+X
athNWRUWfwgkeeJ69Sa8EhE3XlQ1XOnfBqtaXOi4akD8vgV/JNSrx28sKlky6OgzkwTvsEhIRsyu
jDmSDRGB0QyHm3SNHMPIR/5rlw1xy2tpmaKbGXOlPNZOQapmNy+DDFUswo0oLmurSM+jJs/NJq0G
jvldW8CbpYzivOT1M0/HIhmurXNl8JAJW1OLTShyZDSCxxTvoozQy2vjXcFO1mLUN14r0SA+eyi9
kM5Fy1B7zXon+2ZiyPFc0aWxlyau6L71ZF2lIg5BMfDO0+bwq/KT2eWDdmy1or77QRdaqZYblq26
jMybhdl3ryzTD/IZtJ33KkoUCxfSq732xk6ODosgwpX2YZlIbIVKdmMCmAlkLnRMMU4NJNKp7nP4
nMIdscyz3b40cYS8x6z0ozG3iVbMTVebzBJffDyxtVLVn0DvLE/AxKdt5otZmd9NKYI36MkTzJN9
zIYIukAKsQUqqPmgFb91qCjwbb+ezHDrt9WOOFltCNbIb1BMJ9GpRDvum8YUSTM6Y6ix4qRJ097Y
zn6UjuUMNFPjHuJJ4yDdfqGml/UbtcUPiZD14YJ4RFJCw4lrH2niyoLR11vpm97mRfLGrZRiJyt+
aSXA9jqPF8DZTj4zLkZe6/3/bsS6EvGNeinexOMhSsHrk9Hd+yD8NNB13aTOs7Jp7MrtBvmijIOy
ZwQGHAHi6pzAqzPoW4szV7JwUhE2yONVyGF35jfEE+fuyDMF2uAyhUL2XaLx5iCZWa+hRl/j2Ubv
wwQiMBuKEUSbA2nr6tFmhOpeq2SvgOI3sjpbib3uYgmj1fXh8e7S7rd/t9LTADmHnXBjoOorabsl
dmmE1wRiKe9GFQVvOJrQOAIW4x2Ezi1djnhztMVLtVEHIzrbD1GutQhBz4E8X2/tHrQQCVQBd4wp
JV2Hm/dpKE1YK7oSscbBWKqkXE30CCDKZXRXFvpVvf91oMScFsO4UNtvzh6JKKY/HSLdxMBgSTq+
ATu0RKY/mtnZEOaFVA/aadTwThB+rh6XqkQVgSd6KbVS8i9Yd5nZIVMv9bihdGzdHl/LPKTO/3nP
fNzecfVR29vglaPKVvyI5NgXeEsOI+mRGnXeCpywb1/hx5nsSt2D5Ihyd2b5jMdNp4B1vkBGAxe4
6dawLTRTFEEKeo8ja+afwvKRHfR6RsIHUQYxJX53+63MSmEJpcBawMy19b3WYnLefUuIuuIMixmW
106JzKfzRWrgRiwtL4bywfjyEZV7OseRe9owVxNfBEG1Kn8lBNfQu6I1rEiQ5A0r38UzZJTQc9VE
yolJpIzCfwhjxAgsEWm89yKpN6Yh7gPRDv6HUkmhjDDgprVEXBO6X7q0uyCwM9DQjS0j/AvG6m7z
IceVWR0MZOupyH8fGjTzba643Uws6t4U8Lg1iK/KzVWhc6zTm7yUszT9Mkp0eLUSBPkQrc9Yc40M
gZ4Iaipt5IvxDh3ykTKnQ9uMlGcZs7tRiviNa/p/vIAEmnMhojjnuKgcuBp+QLqctqejmbi3obc+
ngxvWH5EtHVBtJHYWXqZv3JaMNTT18fsRZiUsEtM6O5hGKdpaFdWqAzLR3rvoReltv9hYJwwV3bs
qsE9/huF8F0FKO0vcX0xulapevqvRh+rTMxB7gOME1oDhIBpIalSScvUBgiyDQ0eLzG3gAulo6u/
4fL0yjwyOCIfd5rl3xolacpaJpjjSaoJKRf2ZRRkAP33A+b28j0P1SEUte50eEBJKt4AQYuQcTAJ
JGYY6h7pfcht/zk4a09LoonuffHztXy+Crz4XCk8b6UwVqR8zVdfJD7cCBITK2Be87JZ7A5W35Bj
fJiFgoN3HyCEZpuvY+t95wqKi4M6txuiNkeSCRexTPo5mjgH4tFVVwH6Y2Y5xt0BNhH6xTar4Rty
ksmoYyEpBX4r4p3Rd5R+JSuG81JOTfJIh1/gSBrDdt4W3TWGnGkOYfC7nJTg3y1Up9VIRB/p5Z5V
OOAOoNNY2dm4RkBiiULaR/ho4hE7h7gb5Dl6CymxT35znqPo3hkliZYjVZwy42ml//G16D+VjSNI
up76zaEZTV/eMJgFFc/st9psTFFls1ZyBElPeRYKv6Sqo1S9mJ6gLlbge+/Mq08FSb21wM500RLe
oN8HGmRVcc5spH10piDXtGZPzrpMnrLViOGfPdEqvkq3QhEJhZCD7UiwE2uOABbdvyfUepe3Pi9q
g0g8AcFjhPsGHw45zvRsuK04sigsKo/N/Hi5BIv8yigrhKKjfwHeiQb9S/dlyCPAp6Y/zYXUy0gl
fQppEfBd7YmPiHRNDVT8wRALLj4Zs5mcjjDlcCF/xav46gPLZ13Tohynp71TB2jGZS7ir+Kwt/ny
LFykGzYrOdp57QsXsO16UNpIUHLJiwKluxeH//n+9mi7IcWXcq0wVy9BS5EMDiPAzs88D/Ikbzc9
tTXyQ+svmXut+GI6im5xAgMkTBmawfGSywLP+o4x/P3qddRCzphKVS16+yaH1o349jb7yGhoNAh0
bo5ffJZkSpx2tO9uhbax2iKApbsxtRknRS8rp1P3hdn4krVJlSiWbvjegkDPeLoFhI1fve1PoO3q
o9q6bOobuJ0Ol6Tb09pqcf9jwSFFlwV5349v8Nlfr82yIYVnkmibTktFTJaoptqqlghTdQ1o4cwB
hxUzK5wXNhOpTRkGZDc9ZcgKLQgGnzCt/wi9s8wWGtVCMYgWkoqoJvfmR/9pckTrYAaRIwwOQo7W
RZt/Xv9FYsm3RkG69G9f3Zpun1oBjli+jZM0ZogdET44hj7lnA2XxMLRBWFEbsUEvUpXDZIQjCG/
0/W4pvhyiJXqLIVxaZHLhwJWXPvJY/5QyF93O8Q19LbvG3M6y3xm2/5Tv0VresL9M4C8Q9pjOv0Y
9aMnv7H/6K5uVsKshxPP3Gylo4BfTArpi/HFH5jrLe9Wc/Ri3xM4e3Rgae1/i9s2+WI2sQZWUTh+
+R69x/M9j9FYd906/PIr/CZkE7Lib2Vsbz8MfWLk+0ONHk6VbWn+QUuvQmKV46tgSZi0LNvBP7mI
hNoDTe4NCV/KUjV6FtU0MpguzKJaZ9lmEz6uc1a3DOx4KpIuKze+DAJF7AEsJqmJ8O/1M1o7q1qf
FFe01fHTbwpLwUMSWsfuASOy4zpcp0qJDQtHK25ip190Jh/v7BTXCTE4JosyxQmT75HS2L2IBVFx
d5nBaQekMZbCbmclQ86sRejtu+MWuBUSq/AGL9tXX5RxPiepQ+5zIqT9L6ptRfKEQEac+FFb3ElH
zcfUvEyhcdwGHatZ2B18qk4Ln7urhEWlcmXTTB9iQNyTuoapG5UhuxGbaGzL1wcro02t/4T73L/9
CWJnbEKvMseoF0ppjBeLAMsw9KiridCi4Kfurge/mja5N8VI+XZxqV5CyTmBuylHSlrx8JSr8Yet
q+DKSsEie5PBAp02GNwUjojszPdaIpf87njjb3BuN3ikwP6ySCKr+XhZ2gG1RR7KmhdJF2lp+/Xx
LCnx+eow3Q876Csdzh1EjN1yRPsCcqjYoLsTKATkgnr3qth1beulIvHA7STgsu5odl8FHiaiCH6J
2iTTnlZGO3K0LI4uxgmp1edWrSRO2DkUNOl+aUYxqjpE80EpfIFwEbM3SwiIWECiEE8WDroQajlk
Mj6a6PXiB24PYw7G/hYZkNWDUtfFQybmUBvg0rPFScnIlxMOESsDWE2pJpcE9+nhPJRgx2Zau6iL
UlGOFHIBjShrYf2k4QkJVTKo4VoLpvMZwdaFCwsyoHxNbd0nvYu3/HjzFdJqneT7qbepDs2yNE9f
XUE7q0WSVC30JGK64lgrviUiLtP3kz/4zow0WvbuBWrOqLeYZhX5CulU4hxjcCaYkzq1d4pGPMwq
Tz0CtCTxdDDEH4Jx6pO6cEcBm1S9Hquz2PoCyTP04N42EyoOU8aYIi3cE5nDewTium37qnrrUfUb
sx5oqPCMErmS5Zbb4jTHYBJZdzAc2iyou6+xI8vvet3nDXzJQweJ/MxL+5H3ZziKmBHFojKXVN8n
nPsntW90ncffugU/7MwAB2JKtd17eCG8cqbXLgl7ABzJ2WddJi1mqYbgiQ6m6HcD2utW3Lzf3ZIn
bBWwLwUA/BmxPFFdR65bIOCiPCf3AznrLlBVIzSk16toxHREjVaIX4TVAzH8zSqMf5V7R5guOgKM
6VoE/HUz/4/fKZubMQbHNP9T0nBpPapvmZzzuDb9+/50OQK40/o9+qmP9YSTZD4HL4R6aQ1YA5aw
eC7EjKGLjOLNzwt6ylYTVoQQD8nBsvhkzw42nqhzBApcnHhSZ6WaMZGwUnFEetmFJ8Fz4uZznfrZ
5SRUoPux39Ey1EzZUIbyH+Idh7Lnw4pEwcMQ3aclrxRfG5XTi4mAk1QIrdWV/7Wemet5SNbXdnWE
lT7QPmVuyMDVPcy0azYYpAh2yimCA9VfxbtnXJDxyeETfuARATBQGdmG3LEWxhFJvscIn9P58tS4
cO5wGv42h6XErEvKhf2k2DyR9Gdgb0SXo94Thl+MREyT4VnGmails+KMxneBB/teMdCBi6JMndsI
hmjejNQNPcADu3nNbFtZgoB+OtKFr/IC9fpbPi75z8PYQEFyWyc59Ov0FsU56/mORh/BkH0PLn7H
v8p72RZUFoiUKnR75JaxW4TpYY1/1rGT80YZ1Zhep64U7zmLauREmYJjk0koL3TQ2tCgEtg8x7uU
l9tC6SjJ0UNlmNwdvgoY9hDTVwF7VcIPzdDzORJmn2sRAxB8/PaNR45oozffSSb+kI2XK1ivVOEK
e/f7y7Sk3VNLJltGyh8gwhk6bPeJ7uh6IQwj6BLJWl17LY77BE6Srlz5CtFbPTwZEqK0gUmIY9f8
X7C+ttnVqhRgP8nl6G+CDQqI4DTTefMRLgdElZMnMjMJsxSKL+EQKxygRLPE84ApTZifdVHqT7HE
Q5roJGzoRwzBkdkjym7dh6MdhQk6ooO/w3728itsYTjTNXHPTn5C/qsWo98Y+cQP2tTI5rv38Byb
7VlphEy27UjnVS8LGsUyQXXjGo4DL+hLyj3byQhvARupyYEQSgEh0MlGKX5q4UhBBh3qnkId+0t1
DgIBevAJzF9CwVQSu1RNIzkr7TXDJzn5HDRmJ5YEuu8lEokOGcfY+chjBNbnk/1hORjt1Kaacsh1
HsFtHe3RwWRlA94ISrD0FnTFAmoUNyZnoaKgpT/3gNTTi+Om/M5qbkAMQhUUke0L80pBFqTE9feL
4O9EklX61TdY/uvpGASSO9JJtYlK1FmdVgvQNQMQGT10KLltt4BK7gynX/yic6oEbh2DrR5Xd9mQ
bJaOY11vx9ApeZ8KPkBQKBYDih/IAl5b0lZ35i1qyGVOE89vhYKEKnKyQBCbgLizUfGZ/GuVN1O7
/WRQDxI09KhcA+stKiCEIcN2Zd87COHXUlymVSmH+hcR2jwDllI2xELjcTebLuhk1CagrNUaNViR
zyki4DIG9b6RBxeHG82wjQTjOlW3bUv0W0us+k1X6RriI7/iIZqx/TkiyYtCy2OWsW+FsIhunWNb
YPfjU7q176C1ot2R6baU6/KxNpYPkzRyg3mfVbIftmK5hzlWWtBR/b4a3hRuECdoJPzJsYOiJV9a
za+mujYm7cR7pfn8LExpat7junK6esGpBIZRLxYkafXWjzaZmzw2zgiGeNyQ9gcWD/Sgz5mqtHy0
pBjE185oNJ0IQHDCJQeOT0iyLi4/LCroSwkF0ns+M81bhXgiDjmKzpER2AvGjNGFuUp6Q2Q8rSx7
Hcous9PQhG94QhejZYFDShCUx9DJ2NHB5ssEJRhEu/CR4hVzDR9WerDg60gchNoroSEpYv1xoJky
mmcrjm8fQndJGjh86ppngP1fU6sCDemCfaF3yhwAhAh7HTVGSwsE0UAW8FUzO2yaDEBEl3cQqC8B
j04jECX5FMbmfJzxEHSEdgmtGYV4YM4WVgq4xsIBr+vPEZYqVK8AftxJJNMFTxeW9K1fcgzzzKvQ
knafMBz5rcbqeNTJFXOSoQK2pNLGNzHjkFUkGDtgIl+hnMREzxXm8YlRoZZWUNkT97y7fovs4vbq
GaFV6q+iCCr6xmudGuo2RiyggEJC6rUmWj6/mru9ePpvXRUuHSHxXmiyZgTAjAjWv0SaH326XM6X
qlwJruzBSC0stQmTlHuJz5+LloFdeFqvxjbZCSTAW/+CU38R3fSsrOMMfb0yGqAqaiOaJf+bqcEv
Y2EP7V3Waq7iN703dTs+Qu9obWBEbpowUfFwwaajLepDTbntzXIjzi2Go2hm5bu8DIUU7vW/2rU4
MFlwSTvd7MzebhrhyqsOxhgQu70hSoHPlNjPyTTzcZbS0Jdb+E6nxSDHGPszAfnW7pYStrq5cjj+
QNZRNC7FDiTxFgRXtAYmt2u5O3GOOt0o9+k1Jk7FT0RrJsvE3PZCxhwyNVgjdDwnNArGkeTiuky/
/2Qijh7OMV69HgZcThPPfJr5Z3pdQ9pHAVUH8eQWlIIYOmRydRwPvTayXP9BN/yfWHisMgOTYDFE
kNr+lJQqJVzKc4OsU0nXKQPrfCVA2t+0p8G/3m2aKKoTS09cCCu3ug5kphPdU5BY8Qerdzty+MVa
PXrIfoe6WUHVmdacUXcDNEApmMRT9zvTMvdKEUalNndJTm2ujdFP27clIQRuG07FOUBNw9MNEts6
9gO/E4zNgxWF+Gy8irWgFDlrnbDmtqNuud4VZDZB0J0ridM7YHa3nBR69Ap0aS8NhRGNFO5JA1qE
fB4tzdGjCR3RmCA2M2b4PaQzL/JK7x3Eu/twsYuZQIPoGrtXfA1zXPYr2CJWfHJc1bK2MYhlqXXW
UNkWXmlCQzhP1BvGOV/88cge4Vz4u+ES4Bpari1jl5Wgpz+mREXj0ss1CoL5JhZHw6g4WUowVhYR
q8j6iWvuv7DoXOyUkDVKTCEfj5KbFLFDXaGay+nUJu/e6hPK/NkyhfzBUFqQBoH6y5aPuDAEEHWF
4nd1g2LXAG8S6Aa0L5UnRIWc0hwWTv8N6tx6LrlHdxfzP12AVTnM/+mcyV9W00kqPkUrKrw617r6
a4eoL/Wf9/y/1nYCwVAySekGDXWAsGX0RUxV21i5JN72yNtTyFdDScW7THfMojvvXKTANd/V/Lpt
1heeYThZgeABGvESYZUmo5fT2ilE9ddgPEAmpii/CFzVacIGcdnteWKaPN4n8Am5jQ1oEnfbbqYZ
jtBLnYFzYj/LJGPJYXY3sWZXvt7XsDMDb5TYZmyNkx8u0RyXW4hJuwTStcppTQsun20vuL26kcNE
GtGiTG+DsDbxxwHjnMU5Ff+GRZ/5B9CKlvg8AletiCBpfCQWkV7r0Of6xNCM83TXOv5bFtc0phF6
iVSIx60/cjRvCL3qA7mJCv2eiUjU9D4pi9Qkd6gEJZLIr+bBB9ygQpbZfexmy1xy6g9sFpQ2KnR5
TzcQ2xXk23A41bmN0XQNCHIRQHB8pPb/nfwLo5MDRj+Q5s8JlHnzW1aXcEF6vQ5V+FHQpu++Jkn0
VrljnNruP7I65gbJ12N0teD9d00YsHRUqhwNKCYAKPnz2cu24ue3O5w9CXZLWIA5+Q4Laj7/X4/i
rNR3M6uBjDKNNgBqME66yGN+pcuYOSPMqdfGe0ukM0VGjOas13Eu2sV6fBKa2RdpTPvIXla1fSYa
rebSVCf8t2Mydn28kFruJT2Yq9B9wyvcOFmqT4LcBa8iYjk1KqcARuwvUEPlU2hunayZQD7PWXBu
Lg9yT9phV8S0AwnwVWuwA4vFDj2jXCaVH9pcqpC+vd8x3oQj1Ly2FUjwROoeQXzfXhCnB4diq3mo
ewpKif3uxMCrBIHHrNv107UhxbKRLp7dQiexUU0YF8jr83LHXtEaJiNd0AOOLTL12rnpHSNOACIY
9rm+UviISjLXxtpL1mqbovIid267K5tizQHFU3am4SU2758uZ0L/E+oAmhx6u27spODubyv4OHFP
2mP4Eq4nzzy7mzs5VtEoHALbQlsqnsLq15HpduROr8lXu409yLaq4OnwTgkOLBALogRrzt5UqqQb
nuofiCwX1AdBFqx4Hn74IiBqDnBMk5Asns8m8TdBqIp0GXDw9P7+mUpxr1FO7IGbXIN6aZQsF2wS
kpt1Gd5j9mGP9/ftlqQlKfXlNmZldoxaFt0oU3QKkxz9YtRB6Kzj3u0ptCmgc6n3iz5+ZNIddZ1P
/chc/KrX/2hwCjXFgYls4+Srv1HZAGLghzXPtcgxdvZI/HoHvNQbo4LwePfMgMbORmZ1gk+sKrD+
UGdamHvtHFzkL/2iU/VaWhoEj0kTTgoDlwRMuXMlfL7pT1KL90idIcu+WgGcZJDJSvQxz3AHPAnw
t+xMq6R2pWILJFTEX5zjE8GQMhyhonom4R2U8vtC+A41WvVDN8olKup1w945oqJf/p9IlqK7SGCQ
y+ImngLjcXlJeJYp7FW4S4eTDoT1Z/S5GwaUw3lUZf2Z6WLqxV9iK54/5IZwYtAb4eU+BvS2mHpz
pUaFtRqLHz2/oTv1D+k+w3Mmp2yu6co5V2P0d4WM43z6BaXlw11Hd21jebU7yXMd1a4Z9jxgkrTb
fZzN62gc0+8KPwzqiT0g33hyaoC/rD1n6QN9FFoaEdLrwSfyohJG5WkfXUKiYiojV5lEIJIyhyUu
DIcJtIFpgSdyMVzog30aVHmm4P7OZysmIP4QzPqkZ+G0IqULmVfGXEn6VePJfGn2NMfkzejdYibY
BhxPVP6RqlxFoRPCSsJ3zMAk8ixzkWzRDZZ/mD7udojVoUtMCjGBc6HzI1mp8FIUFDQca1dTafPp
iocLu3KW7IjtvZZz1BQApJEX1tTGa3jv9mMt1UOrOufVHtZkbr4OYi8dSLuCj/8tFlteVRPbvcxB
+kQ3Rt93N6JRI6wt/LPEX/hCsRbIw31pBP5ICRipQKxc+BWjMPutQSeaF8UJGTXwpSX3j7Ucy+u1
FpnFC03i5nhN1LN4i4DgVOjhkRlTDESyRFrT2ekvMaew62xYzsnaaUQX8oB61MMTksg67JiXxvJI
it7QrR2PyW3lSr5XNrvR4SqUt8LxzWotsg2V0JxtWDCY7+i678vLCCenzU/N42dxq5nRnhbo7fJj
3gMs7/eEj97zcqYW39wQ5N22BBgexJTQVTxPfDkuLu+sQoe9dLIjuhhkFfsPWn+8Nd7R3y1jz6VA
uXlntsLYYVUTSZn+ryBoJ/66cOKy+cg4Vfysf9u1JaxRksvKhDE00nhDuVVEOrHOjsFZW6c1UZY+
8FyfWpPPQZWC9T/tS7koioz7qyod+zxtSF5/6x+YeNNFI2kQ1qIJ0Mph+KD+I0tMfi8sgBeER7fF
tappNJiHAZQy/6r3kJbyfblorHTEHLlN9RzfLQAAwtqroSs9Aui18rCoAj/amZm9ArfGGFpo024h
vAmM1LANHEEA+RFsV5qt0yFfBdnRK9HYPIfYATsBOtWSu8qpQohxhORkNZ1UChJjB+EG4PIhvQJP
nbJlBJosc45ouPITYb9+NLwLQuVPReeExXdWqyZ5nr3yosFVdF1JHUkwJ5+Ols1cYXdmnuv/L3T9
lPlJSiy40NKmL3evn9pAsFZpZS88SzZTdOUB6pKwYKLoMDhGaWyQJ4AI+hdQa1rlWeWlgWWv9YGl
hO2w0OLGs30YSNL6ku3Pg5rF+HSgeqfgnNBQv6uC78js2tY2ow5ZgGYOPFRTwpwUSfssOeu3q8p6
Jl7reZxq3/vcOFz+2D2d5Q5nDNdIrVVyCsQG/QuMe3eLIkzDJ4XSmq1UsIVrrPnRwB7shJpNrzES
xUgvI5vtoeyYj7OEUM1Nd4ElO/psGvMwvqJSNuXVn98ad+2Jlo/ZisBVrrdIFRGKZqrVG0XRIwwC
LPuK2YbMEDLkHWA20Vi+LBe+aQWBSRGc8zoqQDGlsqtajn7IMekyi1cAH+hmUQGF6H+3TEEtuukF
NP7L93VT0CFEcJFeBrO8+WZ3+I26hzE2A9RLGaZdfkBsK7uLp9AE8QT6z/09v46FlOukfBwTgJqN
f4RpeRo9292c/jLKeVQVyiDU6PT/98zXLSXHMBKFrr1Thaz7tWOkuB+mDoQWQLfAnm7wR012VhZ8
NOUZaOaaE8N/Sx06YRcYJ0URh80TFq0L/S/qyP1oiMK7tDr4laZIeKDKJzv6hhWDgurZnxUolxYq
YIgPNZN4LfcPopDRmQL1spnYghLpP76v12fupYhUarEp4XIvc1X5eLAeZBbHf28G3yYubP/ypbQI
iSVDX3+8hKHvx7RD1UOkdZKtoFGO8OOe/u62yrVJHGUMGKtDIUDmosjx07afsBlZCTtZqnoop1iH
pRsBTlyZpDg/4DlHQGKbs3H+xM0YVKYjSwWaquCqwFJ6KGydBmrC9hylUMYoGPoKa5fG2LVfCUGj
DSM073wy4T6zoseNiDoUYpSRpVdxDdsfJD+u6lOOQVGiiJJiFQ/Q5J0UKTDERw/irQwmpv+uonzV
Z+ODwOyuv/eXbVJGoDR6HPGImy0JTW3RKchVPYGv02cKXOEde4QsHeMOPBHZ9MKYBK1TiJFOiM4y
dfNWUpgOxtCnkjNVsCANCFjcCnlPgibWDw9deTUOTCaph8dOmnm3lSnxFDxaWBCisqyikyA0+syB
Cjm7UJhRaj1zBWtGvzkh2kqPJd4gZK5kPOOMOgFp1i0YVHlMeOzfAJdD/ykJ9LwmpZ2QgN2Kq5AL
hcczQzMY0M6IHmUIg1ztAZ589SD22x18XkCCeaFoa6WgGR/LpEU9uWKUdMcRCYp1G2sStgRZ8jrb
697V5bNgOchM6Rh7EhqSWO/sd75ymYj9+KyPYBnW4rUoZ15JIAzqZ2G3n2T0L4kb51BE+LlfZs2u
WFJHxHtuDKgyb617HCpn5+e/MbIcNi0Q2y5BLdRIjgvSZYBlGePaG3ghEAfySpWu474/3hgVcsQF
RgyJPFx4P1tuGljDyy7YhZhLxOvZBFmbMjx5tmL3C+CL29rObLa71pjqleweHniyGdmV0PP10TVp
IpJGB7xz0SqXDGlAaedLOD1/M3vfjYNalsyqO/7CIEHS/4USDT56yFbkpJxuAGynfBnvTn8I28jT
2eWVs160CYkdkZ58deWUGasiDc+ogIQTaCeREAP1qA/Omq+EomAKwJxBeoOY6FZIX0tOSjNXH4t4
BueLQ1rH8OmsOiKDdH1PbNbQ9gEi/hNbiJo23wPq+8uqFb6CMBFzxABTrSgnVnJsffLFzTfBX5DU
wk7KvDZb73rW6bFTQZZ6lDKCAwIbTXT8mBS22PGs+r+SAwE7nXaLkA/ycOrObJvVKhpPL/QKSjnU
LdU5Qo2fm/rn8v+uQdSQ7jMZnH/TEtJsZRlX1Wsj+77xVI4bMDvVh/+j/uTtzaLGcPCMwvDfOmEL
FfYB157de7AhtrYnE2ox83l/C5S6yDzTHz9YY51J8XLIORJvEIMk8ixzFsQUyar6qaJSQVneV2w7
NbCIgVpxQJbpp2hpqQqB+RSxRZLASKbhPOXM9q/CUb87Iq/owuJ+Edbdg7s5TKfmDZCnAB9w+uc0
+5Fk4Rj+5OL0tzialQMjs0vJzu6d6hGfmhwd247AGULZaQrbGbqErUVg80DD3U/0J3yg2IiawmuZ
e2AvUjoEK8P+BycvFI2z4ghC9+nQDZjHQFPj9quhqCYwW5Vq+3WSXb8wFZbo02REavnI1Y+tWjta
g45ZGYK/bSc/5amqzlIeyhvCTpNU5fqOMv6Z0B1tZW1nKwLVrGZqvMB9tlGTvsyV0GXo63QQfLyC
E4GkXUFiHglSFHRh/8Ftm3L05XYMHICVUiYdRIuc2LAm4jSsDImi2EXdTZQmhAJsg4uB3WW82B/7
2RP34brJkJJ6ylf9PaNQDBbQzhj8itvUTlsxrFe3b3Opr9L2q7G/PToZnDPpyli3FkxJ7mNJwInl
6WBSS85+eBxyOr9NrdPRb1TMUzh2msQAfW4L+mtxygbD0JfMd4+J2P10N8g+qxNCPLTdsbEhs83B
RbjKsKKfG1JEVcplwlG98DYw6Ct5fJOPQ2PDENqnjrAAvDcLVWoR/Ww1g2OC4AbfX6BapIzJZKMK
di6reIhwt2PmsCRnzBEbBcKNgpnXU7SETpqw7GB8N6ZakzP9nWF5MgDlaeTRHheZf1LkN5aCszhF
6g9LyQUDy57NrwHI1LhFSFLBm9ws/hUIZNxtVztTwg/kqG5ig2q75fHt/w+uY5hXLis7j5pGq25n
TvzI1k0Sctc9lTXkeVgKxcX78SoNDMmpmvTCbg6UxOLkpsXPDc0N8P8KEZrNF3Q2A+9ywjxsXuta
ZkLp+1dEn/pLOZzwtYe+q+luN7QAbvgAjjnVCkC6phRUJ33axnDiCMaHWCD32s6hlA/KucfsMzQf
/6+JEyR3ax/55vKGjSnstx0qwxs1UofsyyajXeAAGGjA1VfMN5oT62qVq+DeB9rRNtXymETy2291
zFvjQWjwrTwnHu6ZqR4sHp/iOsU2WULTv6LE9FAnNRnQAqkG49ppSB3ejD8pSlAPAaix7DRyXrzt
ujNHK58xqy3+I38vbcmgAp9WKCBZ/qM41zXEoZRrhbEhNA5ICElvtiK9ng+Z2Tgp3VzKiV4GlPDU
X56ak6iFAqomYtbFGblXIH1nSkQuYJvaFzVLJQLy0g0eH1nB//jMtRjbV9cU7MqelBRRvLcbILEV
XLqhrqkO/ZGGqaL3Z7XOoLszufME86QX963LIN51CL7Q+Msr9P0MQnOO098yBiQLYatq2MvcT2cx
0agIpd0zGIyQBdHOHlITGgIH9aSeknsL3hzBg+gqqhE1gf/1bE9sj9ncr+JSKOvU6Bedm16qjPX+
fBCVKFenzIctk2pJeVmRTQwv9Y2QAW7HYy6lFVqvvIYhA9Qj3qCJ6vwr3qiSG5N1SwhLuOXVQdEi
auNMVhQF1dO4GjyEKRFcOHaOHL8Zb0kcSkcJ0s1pPPx/2CkYvk3veX2+CRKTwV9TaloZS1FY+nnn
mCS5NCG4naPQMNm4wCb+gcthgKC+yYS8+t533ktCUV/7hHDu6BQl+vFGDd5kVLccjVlJ4EvqYbSZ
BaKPTxIWseM4F0qAjbq1vJdc3ucPlr1jU4CszKNzihnjI3elV64kpiiFv6bgYc+mZkn4DXzJC4yg
R1AxZTJ902HZe9SANA+T3k6/dEF8X2qSObtZwUcvIObTg9HYFONE+TA4eF/2UX3JEK3+17XHLO04
7uwZ4lqzQDW8v+KiKhN8Y4s2dbjLxtcm5hY5FN/CQyFWyrqwKh3kZehIQ5MNxdFE+YM3bHCRsO+K
+bwlUcSjpwToxgsczDzUSqPwZldzHOZ5qT96g4ezXVNWrsfX/CPzxGIIRLefNTcaGnqWwBt3fC5/
Jp/Pyga+jc11tu9MYr4gKsdDjiNcoyZW2Nl0snqLGHU+mXxduQfR4oRQnAQ6r7nFkjjKoTBr2ogo
SMNpcBqlm6GkcctX+kyFpsTJ/OippWDzGb3OdMNG21Qlr95ICwSBMbRNOyf0RbXBn8dz9UuM7AmB
c6kSZa+NQcQ5CulBu7SLjVmg8iSaz/jukg/yceAGNhH2HqatWDrTcLmuvJaXKcPACWc/QxAPPoDR
RvaZERLRtX9O6ShtMx1AckN6ELHdqhw4HAxKYjMBrjdZ/MoQdCrNqODRmqMiIwlHjURK1JWWbCG7
vZpDnw8myMDhd6FMDqbAtGlAi0DQwdxud/znSwuvP7jBqu+QTFRJhW2ShRNRc/yRW5ofB+KiqycP
P3auAyfu1edrgk6lAIkhBJjp+uFAAS+7nuhkHuWViGhgKEmeD3lHIsbiVA/pJwo3LEnK8t3lFxn3
qYGmKm5+/SYIrVLTMBVEn8gsH3qNP+RvXha3/++CI2qVo+Xd9PpQVWIE08eMAjAxHYSKVzjyZFrQ
XjCWjlGoLF8ks5jPca36Quq+qlhevzV0YnDPKfi9HAAxCOhUjQetHfTdZFhOzb6PDKp14D6IqPg6
Oig59zsGqZC6YPWIE9Y+AYTAZtUK8GRTBSwMjwc95wjvxyufywRkAcnFUd6gxx6JUQTAbpjq+deC
htI4kDPuOw99fglLLDHlLnkO99ETW9/HWuzMfrIeUlA7teJaVZhdcKeynBKGrWkf990kjy52zG66
bs6xX189QcafikYAsEdR/2kzocLOGtj0C1jize/I3HDB4tUWKpSDHSD12lQ0zZRlb9OtcvgTs1GM
ENJ/VLIywLGjhLlB5ppFjkiG46GyxEaJkPeZAg0y4/jvLzcFSMN51LNkwoyaj//MfTo0IO5hBXHc
R+Cf0xcPXwKVxRgUcTLWFtLQhqPK2aHO6M8vW90u7WAVY16RZ+HIcTEN8LjR4F1bZopvNPTU8yxg
XL8v7yAjuSKgckcMUBprbZRmw/TCrvk5K8PDb0saoLbGIAc48GpRzWUfUWwrvtYDWjKQ9F/OARoQ
MsKNDJL9dvLWW68UEDwsvNsOe2hdH0RHNn/ZEEMhoClRRuawGnMh0kW7Bb/usVKohW9fl0eFiNGo
ZhQUhdkC/LkHUmg5ltV2kTJb7Qb+iw5u0d7Hc/c5lmyP+HM3gfKohKoKdYwGsHF1i2YXad226Pc3
uTtO0yp1J4wLw5BGAS6SMKmfZWW+iUUa6s+EpwXw+YYFnocy3UwMbFUFavhoedGpGcN5pcOTabvL
l5cC308Q95U9M7VZue3+8jCwqQr/XhbEThhDlCef/yLauHYX3nQirE3Fkt6y2LwzwK4ok5+EMm+1
UkHaUuMS82Bzm2TYolk9iQ4gFz85SEHrXdIHgDmDNofTkwqoQa4PriP1KdDncLLiIeC1ukI5VsY9
iWuKJbTymVYuMeDlCQhaRW4sHsGGalrU6DRSN5YT33KZej5dEsFXBS5yQBz+MFN3xDNCW8DOJ7c8
B+Cevw77v3ypi/s3Sx7T+KycMBBa/k6ZIUUBVFPz/nWaFBxAKFPjctRZfVLZh0H7gJZjJflJUEuW
ZBRHljaSxeysaL6KMoo8M3se++dhpIda5LRnsgVIPsRlKP+kK4NNlbRTZidJkwjv/orvEY9ay6lX
8yJzHQBbRzQnNNCT2SwoUg9Alg/ngd4i4boQU3av43TaHHGRUODq4gAyMVqTmhuSjlw3WFmdVwTf
B0AVGWS/NS5CPlMi9p4Nf6NOnr/RIW4V9bIGRwXsMzendfoDSjKvGQVAqF2UcomVgBBie5VI3eD0
VR+wP9SNJ4ujGHxYWvCW20yEYI10NiaUV4L7f8TOYy3XmmSU8UQKm7vuWyQtiejEBH308L5ctG3M
bZtCeEqp+L/5mOYxQ8UruLIy8y4IShVCgMNDCHeQpT9Jm+gTee7AaFnxu3qEuMdNoUWae96b1WXD
CBZEFC2enhrBL843CzzcP9vD5gyb339d/ksfGF0fKsPHsfHxDJ9dX2PKEiM/nIvzfQKGDuEXoYLx
Rih45qUaw0RJwF/OmOA5PyT0IgCf0V9vwipICMvz+hH/qpL80u0OiSp9gapc/nvv2wF5CEO2o/RV
zxUNwbKFd5ysiEMo7yD0X9/HPTY8n6SLYW16vh5D//+EV1GFCWwrCBMzrNBFWXRb1y+dXBV5KI8d
hZpj6paLBkfkY3Pi+w2kXj170XgAHLJ1zHt4spaFGMNlzMIfGbrsjStKdcu8w49tHDTlKWWDtK+x
IV3vRi7HI0BG5r4pwwMExiuEKpL469Ao3vNiqrHDahnSwB6AgCvbZhrvUj9UpWeiKZAuyegJyvWo
yw9Vo4kUNZXJ2gyncomxgrTZ2mKf38H3Pq3gUObwmsN2n0rn2gJTpctInsgZ8U6pKwPK+dTryCnS
p0LK6cvpfJFdWOJ6yhtCbKrYCDSR02iQGVxYIOI57Dx2JulusHNNs61J7hx7Mp5yRE43YmChMZzC
v/LVFH6zDPAxYRKiiGKyy7RBxRqFtYPRBAbBNNJGs5VP8YoOk4QEwusnB6YFXBYinKu8f62yWoAv
YalNJahLnr211rLz5DC/Cvv1UoTplZhpAHM5KEAwAkTn/s3WGT0QG9Z0xB+sWOGP5zbREMTZzfuq
mFDdcObP2TMc3h6YhaywgAkE4j5W0TasKpAzNtdqbp44AHw9LmGxys7iJjiELpvosaNa0u0VZSc8
SNJRPeg4JkcUqQWML6CEPOir9H02Frgtg2MNbc2ErkdXsyEWswaQVkg+Ol3lDj8aXp2TBQ+koXx+
TiVGBpSGMY8T7RQsixOkxvu9UpuPnhR0S+gZyllfG+K+Q2Wn3ncmgh/bn0Q279VIntSOiyHFBIt2
yjsc/uuTykcR7KaKeiupeVj/ucKPvzCdv7il6fhARyceRxIJDZQYI0FdGSWYXWOq1Z78W4e+Rh47
QTDI6kuVKHnoynMc6Lrke4HlkryIlAp60GvdNMhmvyIyGTIz8ZVH6/lP5iONUqDlNtayU6v7+fF0
yg/7a3OADNvUzkqHi0L4FXzihbjktgbMOD8tAkGj29uBk0BF7WMbn6YLBdt3A9OXcSgqgqu/ts1f
R/HWgqMtrI23GtCKTEor0wrexi5cL11dEgt9c8/shR6VFn5VXKYIlcC8UBuAE0JFjd4O97kSjARY
fzhL7kd0k7S9GXzNaAqayyb7FPCGQ5qYqOcihDSRTSl+YgDD3e57+W23j3gbbmottTYP9gOdKL6r
PGticcT5IljnNQOpXg8eoXDMBKxrh0Bs9Jj3feHloPPO8DM7j6QIS5XJsV1HiVXsON8UEkoTRAXW
n4XwSRVlZzhNhptVFX1SY7b7zGX5ul1IbxC2I7EhvuWI5aPhNOzOKtkqqKjqIAzD0JJ/VW281fJi
adzlmYcNdv6plsAzSYCJz4/sY54fdYK3ApanoZwcLg9SDl97nlAshZKUog2aechCLBser39M2VSd
xFN+VGYFKG6ujNLILPtnTRnLFvzzDlY92YUyvHGTJYnqRJZEA3ofgcSEOZX7Q485lsQ0fj0jc1sp
FoNSOEE+YVSJYVP07wODNMdhoIbf/4eKSu86WTR9vzXMlBvqtt/AStvgAF4AhurmuWmmNNMm9146
WCBXxLGfSBPWgaYFaQDEzPH+AxJY78fN5hBn4srBB4XtUUjlM/asoCxYYAGdShuNYiB3QTaKtpr6
Yw3/Xa9t4oiRoVND/3hIi8E6oOCPfwyfexHccWTGKZlQU8ihiyYrFCwhtR+vyYOgjDt8Lto8poh/
6rwxvbxKApkAXJISRiLJs0qo0HrAExP5LUdEX3GTI5NtDNg6ehpwHT8ba9kH6iEQueBdCWT+E6ps
QlaUFd/oMiP7HRJgoMK53KN72lTnScQAbGjdPo6op8qFElP6ya3JL/8373FjvQsMo1TMgxTCCn2z
nna1MPUrJQwpe76RvZLG0FoupFrvi07r8DXRq9OZPhATjbSNfrxIRIwx2TM5srl7wjbGwEr8NKLC
rxJNhFmpFk8MrqrFLTfoKtTtqzwUppoU0kBK0rGTce8AGv4tfnuRhEJtvCO/a++nVkQMKRdttPXH
yqiqqSn7cXHKY1scOXmf4mxv1hI3zvRv+uaLEGvroa31czm0kZQz0BdB6agB/zoEACFzPsjdb6KR
zivooE+M50py+BWBelE3gCx2vJFFKgRajAOT+ynDP9WTLb8n076rtfE296BBxziFjWxVvyBo69d0
rY8WLXlFu/kCTAypWYoCLtANWMKuu5K88LpHdNsifZzIepdQ1LcxwBeak+qYqQqZBGH7eCp+Exac
IbZb6LaKy2T4EP0zTBj34qGI8nsEIAMhlMSX9zcGKxjzUB+5o8nMhpG4NgsFDPGKYlcgyVPNjugL
H5VxTr0N1c8JRDfwE2L0bM6EjYE6br18hZIn0tjN1z62uMgN6+tUcFddqWHy3Z32rog+/i6VwQx7
NCNxlEqxz4l04sjNyhFzrkJWCQQIOVLInfEVKyY2X9jE+QJcY7ZqFOwFWFI8aNPGerBocYRBvs1/
b/NqmKaRcazJ9vggpSlJvpu5hpqoYiF38XxHgvlkUlKNOan56nBJzoflYZbiPvbWFbjDYbylHIcl
kQF2oYM0akum+cMKyb4OXKJhMvtX9dDyXxeQY0xA6ipt9Bxm5Z6dTM/9pMFm6EAuiYUKbL4a9iSH
DHHTH6ixTwg5wKldEXKzayrF/nCMVCDB3cZRVjfaJUDOfB6FvmV5FBt4FWEJHGVzdevfqBw6+0kP
P/hBtVpsMw1AX4SJrkOJ3NbQAuQhiI3jz1eoDJKtF3+aWkvuowL64/9OAEiHqXNmAhyCW8bDTj6k
O/J0s6EYJPagaBuPVudxqL/HkHO2vMhjWz7PXJy8/hiSHmAa1xesbd1+6fDGEoiNW0qxa0wm/Ug3
p0dppI4zL2e8A7EVKyfmd7M1MoGE98Gp5TeYxhuVQ8NhvYX568pR+kw0LLWOafBry/Amvenjo7xO
fj2Ht0zxSEVrV11gdbaYOEb6/YmPW9gYeazpK1mryEmlrutBHjp+/2Nm3VAp+Bo9lRKaG/ZWqqtz
uglM2tDh2d82k8tqtFg6A0AHV9KKX/QMk8Ajooi8uMHurDaH6qv04plvSnkqXzW64ivj7MCi/YjI
FbVof3w8uS6ZxdtGXIm5D/uJmKe3AH6Ozs88owUeZoGEmNMSZlXIpeTfB0+tRLJde263wHU/tsLX
9gRBmPIUr7Fj6BPg67gOYNp9nLDXbBVjzLRlr7ArxncYqs+hDCGKvqrS5WuF93r+4Od0tAv50w6f
NQAqw9vYq4vlL0go6/XLguSekN7W8Hlp0r8BoGNG6Zn1opmy8hECPJ5zXhUmmlecPo0LFxPyzTae
WJELOXdNQu+Uff7k5ipQeWzJtkar0NWtYCLRGNyocDrqJY4ZEyFdJn09iiqr8gzePK3rZlBPR4t0
UpqBNRAowxLASPp86l/FgMd5jWkszUNtiLy1eChoIR8ALm3f8G3xOgMsgd7qQ8hDOdkKnRChsowG
lKha6zIbRxg9j4aCK5Qt4E8HrjjKwtcFh/ypaHtWXMSVSUp4Ipf0pQ4c15kusNvWUjiAK72sENqI
vZ8bKdcwXASA+41Gd5AMeS6lnbZ+0JuE09c1z6kCjn4P0S1VGRUhEpd3AyCuIL4Y/mMeTAGfgH/y
5y5N19iRo3E2BvPukyii/Xh/mQ7tfosRONs3zeXNAfQ+hjNdN4nB/kFfzvjlPOcaeiBWfDSTEDzj
TbS5WUb1f1CFk0Xrc63AhDKPAUmv+Nf0PMrh8+SqdEJ1JTEJWPIopE21OO1SbEh87NRz085wk8Ok
YrWV+VprlY7HXbaZodjFwtFhuZ4Agx41y+nWTJgqy7mYll8uQqT27vIDM8vBFOEdi2b6d4821+ND
H54wvtbxj28+t3OucPCtaGy9yoio+rboKr0/kfaBS5K7NXPCwblMRvHZ5Y9S7F1wpCm3Y4APNnv/
/9MQZRCMe0ZDc2l5Dy0yfKlFLlwFlbBJ/fpkYdxFlym83GRf8lx3ZnfgE72RUMRbAzvh2b1PJGM8
DlQYvRaJ2F2fKjYAnWWWXcyR8TF2f42SmwN1R3cM0vy0/M0gxFxDjwI+24ZS/qQoK/qpgzg3wvX6
YEhm2smECQ+/C8INgdwoAL+tja/9TlOu1qG1vA9V1b6I+eJCtF5SWjbKXB6NfzsH+mCzrMwesCpO
IcCVQX7vqL98BXgk0uyaBZTVGsuGf4CYxnuUIDE4Rp/I8qDqaokOW2o+OJ3qfYhrdgwhYtyQD4VY
7jd0HbbKTCaU5u9zOFcGtVIvqWloQKqP8Zrq8mN7yBlsJtqmhV+ldyzXjj9XemsJ8gCdbQsswy5K
WFpt1ChTn3lZNTvlcFs/3FD124ApU/FGCC/tB04xLR/B5Oor8XjTaqtmjPOhblXmEyjqiUS+r+Eb
Ud+LaJYr3I83lhp+Dxo5FDYHRoMDnKUksiLN7XwNPVEd67s725x2QcJUk8UvC7RIkmygw5RnPjwu
SwNmxqQJZkWp9GjIA2bepN2BZUv3F5//LDXgD5/D8+tyXuZOLDygGOUTwD3eLBvUsvib19sacSdT
MYhtx6+rdxYxy9yRSdRoInfnX19HOrp3ToNixvyxt3l5rcR2EwTKBjEM0eBGo/BfQ+XLqNv4aGgQ
fNHplKI++UIRxu5bo8UX0y03sqsTuKInYKvwRl4hIgrDlV9MDy6hAFwwDUxRizFBDpc5F1WoFc1d
suW0Rq1WNNYKBB5F30NfYIgeCmo4fwaE4lcomJH2F84jGW/Cj8dy6JSZJ0ljgo2x1w9nj7m+O/VP
otz8vKeZwDHwgHHRemjsVFNV1UPKm+kUiM/9E5dQZFAKnB/1Q1b612/E/zZXYTEzAC7HdggfmymB
djmxYQTT1IMD34MelEmNiSGKfb2C0sFAtbvVl9uS0HT51lhRP4TkGrdKPHBSoQtWLpHPtSElmYRX
JaXUzl4tVJvHEdf2oXRhKtXMjQlrHpoBgqzlZHzu7be7f6oJ22/bRaBjwu+VVjronCqNw6yTXy2l
YA9ta/o7uWP7pibXXHPWxUE0KO6HrxyikMMI81LueNkb8D6Ak4jQDXGviifKGCtpHwrzbLlXG+Jj
z5pJiiER2AgJrg6+bpcFKVzlcbKw9fggJXj36sRUmW3QlmSzTsvf6GzCgtenncO7fHfQr/XslVdP
/MGcgTVv6b4A4mjdFbYiLJDFvJRKibpNTzXxuOPxD8Xbrw8iHOqeiR+uvmnyjevKf2osHXWlS7wS
9ta83vyArDVa8SdZxMoyPRddbMiTUq+mzdvb9YSsy1xTIQSIvQeg0bwAt4QGxv2QYStLwOnIdVkJ
7P6j/SM25z1LNMoMrFX+BdZgdv8jUhThqJKntQ18F34hprghIejKTCgMWzVFuJesWHUWoHQznZDk
CSa6hQ2JkRvnSVAnVRWAxPKRXIPxPosXkSdHT+SlaYVHTCI0ExO7UbDZNTecgyO/UVwxQ0xmmchc
yAhUeyukNKKKiwWOWCvWJXbVhMOAG7NuJu4BBJSEVyfpD/9ic7l4VT5ZF68OxMVNMs1b5kXGo5dC
pAiT6u8d5kHWgkTcy0SV4tLJQeEwZjCVnjj3Xh3OAHI2tu4wYqlhcSmiBSPpnTaiZRhrSU5m5/Dt
cNosGIHlxYNjwgo+MeaTC5VKCavP3OTuRDlQInuK+geCD9n1JaMnEambty6sZgHyhMieR1c6x+S7
dxnUmpQewFgeFS4nIlxJ+TWdwqtHNhqd4iHLSXNSIQQJ8zyaWl3NOrRL+R0EQUvAb17i8PWSQSfL
w5efnopj41hDgIr9fqPA/dT24a47kdTOwkS3hs75V8iHylRHoviKQYv4iLPPasDesJ3qOytAjpCK
0f6ZmhhkAXES2mYvfapj7NNVHHqxJX9O0OABKXGnvWQtU9C9Gk8pXS9cH709Byh3Rv/qyX8j26rI
TOIRTgTiYr14kwQQBj8WhO22mHtF3koT0SUtxsgMCIBz5c1IfuK73AT1/qtvH1Oo8RzSNGzfUbI1
CT7DjePQhBNG24zym8UzhUtht718hi73TEEO9TJw9HHhR1DL+oCcQdJIsDx8RZlvSoPhY9XnWSpf
1zSCVMFwBlRE5+2cwldw9KqvJVy7Br11W1SvG64ygyWSRBsYrODH2GAhiKfdVUPOYAb7UPn+8x5k
9G/gZTkd+STajPvCdL+pVOuQ1WB76ww9IuNtdyWgkCWRA8/KCMTw8/6JDXiByBbQvWi647yaAHGu
nTXDTP8oq2bGwJRyzvQqhXKSjKX8epsiymxlAkcf4onTGydygvWjohPheATbCkW1+0htXz/o3VMX
eoX+ORd1dF8y5murmH5yturLl2SYURJFPLfOtazAD/9bTkIpeOUkKKYiBVbP+xmwi7p2MPcCdKuJ
Ahp1j+ksijBeJ1dIqgXRNIbVWsmwSgnR53tJ3kU60UclXcd3CeqSTufR+j/A6Mr55TJOfDiZoswQ
MZRpaLAPnn2T+TiMBlVHHpUEgn7h5gx8qQQehgFUrKt6VH7Cggl7SgyIPvM4oYm7wvCgkcH1szbi
IJVIeOoMFFTieRvLfABKzvrUE7+Y12e9SjEfOnHevMXB2CJH1JvhQZJzHxXE870KA97R3balxuYI
h9FpbUnLg5orbrlHpHYMGWtf5cZJeOVupexZ2wOdnXF9xAU/7BOzbc4x4dE53HdZcN7aXivkRPIA
CouyZpV/BgwdieumgM/9x8Upg05PVg4fgjyxC1sohC8zZjrj5l+jmjG0arTzGLvY8cBJWk1Uy2OH
FoQpbVKyB1ysUfD0PzgNrsAWIQtmxJKC8/v+YKzYbM5TUXYROu89siI9cddwHQLzgNTMylv9Gtp1
kDaLk+Cnt/PJBGozDjDYiO5alTdAKFOt1u6NhLIE9hbMsSAY1v0J7rPMx+3bRc9v2PtJjMdUthuK
Im/GM4NqODmlwZmZN/hSRq/yIYNG6wthmKHaOenY1VQxBnMD6GdGGXVvrKGv448dC4GbjuDApgIx
7kBUtJKb+fz/RwLRacoqb9vGRKhQW1BBxf9HBOlwKmaWJ8YDpnCfQlYlYIXqDaBcUI97yod6EOrj
rYLOSq5I6B2nci4PRjQv8AwLOg0jRnIRJnnSjgW91wtzrzpFtRnaijVOxkY1xyld4yE6jVfFIuiR
ZVpQp2KIvg3q4HAqH8il7NiSE8VS/iHcVSOIoylDc5qPWHmkkSG8kf4X0aK3Ams5MOZwjBKcie56
iY+SNHzIjjZ6jrHjL4DRaiArkeJf5vzLQWdAWF8AKwoY976fSp2BMOJsfYeTY5q1Gq3A5xmmdsIr
MCLudYllqGXtgMUA9UV15Am8rWpy/xO0m2FlsHQ0Nn4KZa5hIV01mbmzChcOU3AMSb/SNQ+7MqYC
FkJy/ljU7S8leCggZBEoYy+pudtN+6v8h223ZVR5F97i4elyX8sV6JL2MPDx//Xx0KBUDC/Z0r7w
d4WCK7ADVExliKj0o+gNssnNJD+LMo89GwV7f9PKAtrrHrht9C9H3HsOIsKWXy2JUi9RaVgXdNT0
ANGJYqUm/TvYp246SEpSpb4JvAHzFhJ0Hv12Tu6fcKVP+4XCy0zudXuiR9ZHTVZzQajKWYRLAPK1
Jwq0OEERVIAX/ICjW2Dj+L3xVfmuw+nBoFMlsZWdtoKZekOLXq7AykY8F6NNq7g2xF9qaJHzIzHU
lJR2iuKcRxxg2zn3gJqtf9hseGDrEPqIBnW32MUt7nHPPG6TwPgtywp0ge5Sv2jO5gAG1tBMEL0y
Y3h2Xi1Q+WbyHAfj48oma5j/2CMEzu+6l2BbjP2pKcrGc9AKDv86bd+91BOF6Ww9bqujXI6ffvBJ
cZucpElmwucrSjOvTs1qNuXDMlAZ2YZxkpCInwRdLYVtbbfUyMS9YXFjbXmNWCnwRmqdU/WNkUS/
D0adn6Ysr22YeH7KMqo8gN8hiR09xm0oVkBEllYVBDm4khuWv1m3v0E9twaoc5XPPX58pZiQEnVI
NuJilgTTboMj1Kzyp3e5ZwlJSUb9AaVRA63cYku2PRjQN0ZKjlFVCpw3EU6jffvOYam4bd65BatT
9JDugNpt29qyQYgumNd/v/NyGyNwn7HytVfRr/Mv9373LNps2W+KLDgK3N4Xu1kqTNO6iz3CvG9T
oKCUghRniyLigTsDLzlxoUbPU9HbiRVeNyHRgPl+7+dTrBa7YtSsxrTcSRhJoP+oDkiRAOm4TdAD
FnfhAP2f9zrUGiAWVZ5uwgcuFG6lZVR9cNmDw3p34tn9Rh8CjQiqTDTUmzbeki8hfUMIYW7mej8J
rLKEE025Akgr8e59SmKdrnuxLTnbQQK0cQ70rrZs4EI7sap5woi9vSPz6cIrsbBnkq6ltqLKQ5v5
r2w3kbrDUmUkl6XkwGr+yots/ECnPCP32Kk9wPD4dMhwaxuo6pQgWDdJQB1/xvXoCpJy84h9uImb
JhYtUK3SR1E5ozSBa/p/6Upi4t7sd02Wdv2HJp/beYiU2afpHBDh9b4Dscxz8QEJ8yIS5YoMDkUv
6w/G47kcktu8GqLGdjDrJDhjeBi58sI0Wq7xXcRDJjRzns32vntRX0YshQhsagmZDFMPQf1f7uCb
9W5ofofLPiqljC2TMkRrm4L28BpVswXCfJeAc6g/NBGr3uXJPsd5yjNyAQ4YniUfZsA2ZrlHiVPR
HrhmlbFGM/Wx/aC8rcBi1J375HsgGkutVTXXRnp6YMv+R88ySgAfy2K6ayD7rf8xtLuDx1UPaz2K
ULyKRfj4hoU9jNP67/g0a1ZdLrCI2PMHnLh+vZyg1iCcx2toIdNN3l269Jv6Q+W1MH8yGWeqCh7h
gZAU2PiAg2NomD0SBIjIsQOuvsVeyb/Cv5K8HZJO9hSOnNPow/u0bkVlu9x0kZsPNx2RvcCYFmFc
HY0xTw2S89n3f7dHDqvHSqtjR2caIbX7+j+TVAGISRBSCSXDBt3GE6qKh4oSTss6MJHTyTRTpUqM
Nyt23e4HpEYAgTATIbcVyD90TwO7tHFuIymp3mdqk+QGvXSe5HoksgBLW3oQY495sGwLfrJqcQzl
XWjyS9pPhOUl57f20qRt2reEuYgOT6c4eYwTa61kegdUTu1veUjg++8ca1tZ7aw20xTlyRasKLkV
X4XGAwWrtFnxEeQHSGhsiUx0kvq0d49cqEXR0fMv9nci975s0q348WSdquCO8Afkte58INIZH7DK
CFc+h4C3yRvdV48o03KiKeG83zC5aDfKOADkItFTczfv7Z2ib1+L4sWvLmYTPknguMbwTACyFzhf
32NxCwKp5OjmOvEMNIYI+Pji8HqVbEbAMfw5bY1cBkphGce3RB578utbE2M+t8AG5EltaWWMVTWv
ioASuX5kjo5KIbVdor/6gzqoR78KABH5GiLpkI/N0sJtOgh4UFSfaEW8h3HowPlERbm6Ads+nQqA
PRIRZBH9RrlZZp16nFnfgI1sDEsmakOMf/7QV6AeOYrQOWLkcpCMFbT1/eQqDDGhI4q1K9q673O2
Y8xhtkaxHT+3izEWDlJPbJdtvDhxJLY1/USuU43rAYmQOsZCQhxmSc0Con3GbjC2LbLjNe48E12H
cj8Oyu2pOmlXMUh+AWbiiwKulqnrtG1ysVLEQ6aD2vIH4Sr8dlUFEVH6oY03cWpvyg4gN5nI75m8
prIPYMYZc6nByjMsvSCUHihO2Nhpp4yE92i22v2XHzFrxxbxVLwrLoGM6cvJKisTSO1tO2etbpGq
ljO6DoMBJuq52DTb8mz9mykp2d0Pzm2o7YynObaAV7poQ2e+c/Vsl12mwUieo7IqxgmYDVt3uAZz
hbXhc4L9hlsSnrrMEr+XFYv3KZaee2q0VctgcfZhNFeJxId0evebcRedQhY81fDeLi3Rd9rfSvHR
2MMt5oKG899rfqzftnMtK9jkdw/psR6tPzrnUJfChBU53xrhQSDsshQat4dMm1YM779T8rY4T+r8
LsbxQP8kwCcbrmst/pl8J0A5AlQQQ6Sa4E8GNqG6FN0u9cfmXTG8yAlpuecAgeeeNe1Y0KCrtsub
e/FjEP+ao4Xv+c2Cj+IyfPMU/zGd05K38Gj3FZB4mEFWuZ8xgCGMLoS62cKw+9iH1HQ7QxRup4fE
LeUiG0utTyaNKdQIehXjsJ8bcp+/TRN6B4tXyrDUfxuLLfQWshZOKg8B1CN44K+HxOk5Qwnz6C0h
4S1oOtdZSaIlKWE25zkylPvJ/nssn0e8y/wpmxK8R6RVpQAnOEfpFwkcPF/ZAa0D43gt1UYxh2LI
kLzyg4Qef6OdzHGXP69cY0yUkx5Cn2r350hYqrlCUI7K75+rvq+YYyit1GyfDClgZlL1bNH43Buy
h+K3jBDHlTHn/Lq91HDpCfRo996hmtJD5jkhSv98fuZEJDvbKIOh2k8NGS+A9WMAOOvlXzqJOZtF
3fZr23HkPNRau2uoIHvj+2wR6nqfqLwlqlCsz6R05A+4SU6mBsf67z2bBzcktHc+gIuCIqbPFaVF
9jeyY0GA6XGSBptsPawB+QAJRqDO6MmWvFKeg8wx0eAkQddkgKJEtOPAQT2MX9I1tm2rKv3jlQhb
pKgFAUAh81rqESxj1p7iUxc4tDCrSBzCsUWni6Oiq/dKzzxSeFkFI9dBOSvZX6PbZIV9A8/VSHrw
MJxIXvJsxsBSmie+wgWZ0tg417qfgRXutZbQ4cDeU4LjQu9eNcXRRNHnf7eqf0ggR/a4/4iJy7+0
Z03Iev5oVtvI1uhh4sbRWXvxTmkEGj8P0XPDiPXA9j4tnDljTXIetVSNMRvjXotnOZh2dJz43U/J
Ut+b++kwfhp7CTAt08f5OQGRM55c9mEXFhoJumhzFsl6OH7+gNJYdJiRkmN+J13tEiCVPeSZ+9BJ
+6BhS7PlYBSkkktKB1zovRt9wwr1GfYiDjXmHC4RjLgqu+CIws1k/4cziYrnZfdIWWWN9+fdnLGX
f6OGaRhz+BtbDZDYVCKn4vacA3qCZ/jTBYrcCIgHTJstqfrfhgrFeSR0jISMF01SoONFtclFf08E
GUVjt2QawVxozkL4rU9TDpCJIXpZuGKo7oxUlG0u0TgWEIf9TV9JP9GlEGOX4CvEqRMZEpv7gsog
Vf1ZRYdhlrLl1YWtNIOjlel8oCezQQNguMgYxArYMnJrbuV3bIPnUxbRZRBfUml5kOx34fsQaHMB
8+SkPLSvsgiKAJnaHB7/vSiJrXI9Ia0BDkKAJLqfi4RJTahYTs1JKnyIqursiZV71BVrGzs1hHbg
I3uxzOxnfRFv028BOifn0SpGdp/Sev5Ho5/HMuh8havUjkJctylAm302gY8/2sV/4m4eeBNqYyS6
cyP6Yj35BXaywCLEFQP+y3mSLBGuxkfQqeNwGQWoYenMdJtQ4NemTV68zHB6UR63Zq9Ad75qpYJL
Xu9y7CkcNiKXtytPR+bhguzu4EM9CPE2bGHilNkpNPjBpvI3USlUAoLUBnktJkgOj0i4bnJJN6fF
cKZrPsL8mArninnZcU4HBGo/VoG14hVGQsVDl4sg54DuJwZ6/5+vmHC67JysMVR/l65Q3FJMJGZI
nXVKNUYdofxDl4BHVUI6ZjZKh0zT/ZzznbVPyC/wGxtXFX/j+FNGqfuPFIb+kgie7Os5JocbK4gY
SSf4C3C8PTVGSLe2O08II8UQqihf2WFpHRlDVcnl/FrQa4VOWQfNN17Rfz0DuLndCbwFnaP8BzNF
r0BMhIjWDikQLF2/++UJh1viYsjjvXHvu5dMtwTxBFoNmx/2BKk+V9IabXSKfuZ2pZai2D3cDeIR
pFz2Jbgvxoax5zd/KTpT3FX9fs6/k+WYx1DAhJMJ67X6aWtxdkbT1N51ldwOSCbcPNGGnYZNNr1y
9n2PE2oEmohjj96MHpLA/M90+MRRPIxV6j//T70g/ThhBoqQlITbtxRiYuHcmj7YxFJsd0fay6yI
02f3b3OjfI1O9K647Ek/RWC4/czPQa3vjCnZfz83gx1mQ9k7QwQ8llrcel1c6UmNtLd+nWX+Z4o7
QpivTS6LhCJVkDytUh4V4P991wN2DizgpBtYfqC5Go3YOa5JijgGrkGIn1tbHEdBNuNkAeF5IoVt
HhytofctMMIIl0o0ilgxbYhtS0dsklqpLqDXhPWkYCYsYav0VvfcaFvf6ecWCNiVrclj7cOjziIl
v1Z+iHFKpE4dVFkC7+OToAMAf3jkpjvoTvuOwEm+qL5quwZ1FJuu8Ev1kZDVhdM3LjX/8BCA2Vcp
ypY2dfq+9ylFMjh4vPmW3n/nPMirkdlKJzwngIBvDv9ZHGhnslCSbWRhHOjQrAbqoLYryqG0RqkP
8nMQLeCCv5Xo9jYHdJNGpV85heFFGS/B3JYftctGfUhRZ/K3uNqnl0ISAHtY+qvAocehcFSBOI8n
0NEpxeTRAzTK1j1iERPWLH1zhlWXue9zGi8OpMw2UODFRsl83nzvC4PGmXXQPzGhEfQHGGW3bIOn
81OLtO74D6lQP7Za6Dz40ZFmBz9F1bQjcIzKEb4o98+lWE6C5l7LshpABvzao6MadmmQWDpRQNH1
e9UmrKzhIN5lceLvzhu8ihqLSvCZH5YI2xOmjFTSJZfVFoQ7gBvQzbK/k1K9QQcsJeD+VmCBijF3
rlkrAsd7b5ciVw0z/JEBX4nThlP+iuTo/zPilILIChQnO2UDpOsfhOjjS06y+4Lz88cnZcIKFq9s
8qQ/8AEBTs72FNxCEksrgUs0aVtsSALO0giMwMagGVw0rlJS3kq+6bRoC41ySumTpd3V/fmCOCMz
HY0PuWNm8c7b5Pf6i5yU85wMGf+2NIS2YKI2LgMVmTXvjbflBdzYqkmbqv+twjeguS8v1J0e/wXS
Y2pKd6dqZsUqesBw3gl7gC2gqwYdwXtPKiTh7SUOtKr6Ep2Hg24Q0oyTC99O6T0Pj/AfDRwQ2vg4
7TkF5APDUkvNmvtmR///OoKZE1vSDhwgIVyQVcyFNjx+xd9OpE+GODObPAa5SyOvn1aRxMYA7DPz
9KON9qvuGoU4OVRxtHZzaq3c8/kGXodYgXzug/wzG0lbtkhSp2Itb8fxJQ2zCuKx3OlcZ5k61nK3
UFgTUy7O4ex6PDx9FvUmB67RpPLIg2ijDzHO82WkFWNAZ1oRomlwgkEymumwOJR5IBCp8aXvKKw5
UpAFxCiZuevFn4U7QAMkvIWBJDBFopDX57Usd3mtX0hVAzCR9dVX0Q8C+qlGHsetWGNkASz1Dxu+
/OzyuQBmoK2hlRcxwP7uRQugaOz/lik8jJ21CwrFrW10sF/4JfWDHGiClaqBQGbA1tW/aijcUVbl
uRp0vC3cm2qGgift3WJ3aAbVDeZs3Qyq0bVnQTT3yoj9RhYgOnjWxI3FlTvMqr9FujqAafnLtJ2D
tWBMFd8VCVtM61Uz/TdWlQlB9mKw2KsPOGN58Vcw7YfN+TypFOX6dy5Dfv7/dSnK5UlP7w8FVhF9
oEJvWJ1tagSFmUPpAMf2lmyBPbKb5SQHBYKi8Q2r42G21UbSVVKMV6SGY/BnQK4+dGjClgibvyRV
8Vg2CY4n2RDk9dv7+n1YiKI3gbg2LuXUD+51TaWxhlnOU73IaUW3Te+MPGVqsQJCjJ+93DqHWk+k
RG+wnlUyjcbFGHhXF0vUmppdfoXefCSu233cwrEg+TXaSC+Z0lHSf+oKL5zdBVItTfDYEWN8MMVM
upUEYu26BZ8TlMUtcRvY2IbkzDAQz+fIadQ4RJtbOj2yDwvoxg1ELSYTtFuGtudYvwex8j83Bzc9
VGiOonj68HANTwVWyjT9R/ByxsdFW6W1x7sXULKYOGFCi2NSEv63KKP1L4OKl9cF7lJU0UZzK8kC
c4DYsXMb44e0YfiRQnXj78sQOf+aj5aYu3jPFZcCdiKVwidIfxzD/nIAVERlrciIYxjegdlO45mx
bIWUrN9n3OlO2sM6oB/1BHlIA5gVjuyv0iCvkqlnDb6pC0H6Un2urTIU7CF7XxdIau/hlTL9g14Z
vaJT/mOFRo2R9t2KYd/06hmOO+wZkB0aGNjGb5n+0RsGNYIx2qBVtUawlLN8Nhy5u6hRAAsoqlvd
tMNUJBs2HmBLh4utIoB8NKAUG/f5O/ahgWK3m02NvVdGxQCyrvbWJ4B5tLbRgojIllWY0mnuNE/h
xnafOnwasRsUByCU1XYFvh2+eEWrwElV9nXKyMjb8ehrS/RItxuK4DSJxW2qomwk+edc9lKDg9qA
B4O8oon2lUDI4a9xRHbxp0wAxwUc+Xabm/VDbu3ZSAgjfsoyFKgt5AvtetTNCI40lrEbdYZzQnB/
7DRjKr4AN71WQsRwpxXRWAIcwgXM6444k7Hyxf6k76NJstGkn1ZAkcMJch/SEnma8LVV8ftmGzog
0rrUPEFdZ4hU4ZexePLb2RRzkT5aQI3icGQVriFvARJCTL9xbfJXic9KAtr4iWKBoDXHQHPoxr4o
A5+GI8kmuWFi3I1JldCaJjLTgTUtwIAsH/gLsAPV7tWfqcdqWvxieUJBJS03ALxptXATwt6at2fh
qw5NMQQmmc5e/U9ArCUFldhLBAWpeijpjxd2dkqzkXN+ghCMlYC3bUJYqEhi5YPlBzH5qlQItqWc
Z6O2c64xL3pDL8ENd+0BThZywEcfghxWzryEo0uKTX8zrz8mFZgo/j+CZm78Cv/r6+uSTTjKe8/2
j0kK8EpQLOC6KTay+7eE7aTe+lKSqqxfliBoAcOxy4QEuhYxa/+BuX7jYSC5olKNnY+AGhC7tRqM
k8gWNrIDqYkKNFUqLzXiX6rTmyF3yOGI+gIJSY5ZXln2tF4qTlXWhhjgcSw1tX8sH6LR5GwIaIon
8fL2flRHrN08g3a8MCzQF7J3shGfQVyGIRXGrIlO31+KGKfK64czm8Upr9D2CBxK84oT0T/BC3Fg
7K+LPgqyzuZ8SsoowpA8FyiFhyrXJ+5rLdNXJ/zBY0TUGDRUE38G1wKmoNLX/0Fg6k9LeDERKWoU
zHPnf1MvurUMoSDuoY5Sq49Z0CMmmve1wYCskfeaUmpKOzmbl8tVqfLM/YawEKlTJt9CXcoh/JkM
tHBgcrmu5sdnUx/8nQNpUQHwgKmMSrmWjG+zVzmRdWJ7pOiXSq6FGG3+J1BpHqpYJchhYKWIji3A
n1EHumFlSbp9KlrxXY1UUB73o0/ZE5CIhdG0uWYf7bsGVaNlfX2rg4+TYDHfC9wYSRvSxjtOLlx6
uaMdZzTMmnE3W+yqYUCkLSQLu4rHYLtaGI2501sN3ofBCIiZOQtR7L58tD24fc3wen6sJlGBAdKg
87mCQ8RFWJKyzyYQoOLbK+9ev+rmh4TCqda02EQ5JhJk3JFilZ9TUbGVdw87FIl8P2iARjjkQdsa
6gsZ3VKoHA5iR5YyoT8F/UdlodTE+utXcKGpfTGahCD7ePXNlho70ybcO0HgqSMft5yzDUA4bFHw
101AOduSSPMum3LDv9HC3gTUCAEYZlFygY3rd+NAM73LbHC7pt1DwAZKOuisVSYptI3rkzOn/DDS
bUwBCejf/JFWLZgI1kaSAz23fbX3VGYf5GI9aSp4R39jX7ojnBn89pgQIh4ONYLsTuqxoirHhxjo
/0xICZ3eAN4DEu4KCxA7kfUbS/hpqB1HbrpGTELYWV9SuyZfHCHaEimFgMEafSLQI5KSsh/da8YI
FzT61GzIgV3D4t+7VthghY5xhGJUudIGVlilM9OEcEmx0qcB0EJlgC58vXGW6f1tZ0Ba514Dmsxc
pEhsRhwtbp7Un9eYFfLpDr6NJGj25NbngsTAiAajQgWUsK/WBCQvXiHko2KbnXidhfhQVO2SvERC
8lI2+LBYh8+lMwDqj8i90u74DMwcmxKejM8DmKCqUa93DBEjSEr13JBm7EXvJdUBJ3rFTrIVKOUb
HlG03weQIinhJMx6RHaFETfPXh3UX2EZ03CRtBX7HdfTi4gI2NZqalWxHfRs1kRFdDl1leCt7SGy
b2tmq5SaiiZ5oOVYJsSExRGRk9wGlxaWxF78M8L+irq6iP/ozw4feycIWHXaZheamsX7By3cZk3R
r3E/ONlKap3eNCi5xKi+8SxHVwlEcLSaZSHS3lfKvnypVdUtefuq8+ryVgSUFM/BUoHD9nPK1hvJ
1m0X2uGRW4nTWhVg2ecyZVe2uHVH1IoKiUclHNjmV5asnaHU5AWH5AwW/VVvYdxVDCi0GCSogLhz
2B9DJYODcH7OU3CJemSuYm67ik9FYYPHG3JcTQEZ7/q/biMSypKrdFOHASjTgp/EAin+72HzbhLz
mMxQ4zwCV2fE8r/hgKl++ZuvXmWvaOtzd9vCz1AAvWz78zcRlu5YFyYFhvDpPMVreXxw12W/LEKy
3PtLqQXpJL4pQv8ALqDHxQ/KxtxwyAhLOZK2kwaATrvBo7QA/5Y2FUSXI21piL2swZZqOaw36gQp
FFbsQ7gOq3DZgwhyRrYlvGR6zz0sPuDMjx1J9zXTwTKlG4i1ty0Zy3qSLtxgwODYrmDzJFpSV533
pFZ5/wR2/Z3Zs16EE1cqgKqDdWx2KRzosF1q6ffYpkERq+HNJ5nsWEjLCDlx1uz86PUIM7ZP29Kv
fBA7HpCXEEVYpc0FjOyoKMDhsGsRFOrBB3zxjhoroHyMayT3CM6x+WQVjMD5yQdvnt4Z+iL+yRD2
xn9jt7oRNnk5a3lC15Gnw9LWUJJv2SuKi1NQIfbbMckY/K+DGZqA6anaERnab5YeVrbVh4M4BKFs
DD7s1vsRDpmkYyYJZbHfFtkd2mlUWOs3xJtXzJQnH+mjCUmxaG7VfIsCQoFe1aRr8zzW872sOGXZ
BhmxivBXwS5KgKav/lhrvOCB3Vn0xSapwmoQ5D5hfYcXLW4SVRSulRY4jsAr9nJMJfXfsDud0lX+
GgZKw66zN5LJqqsBzsORjLaDoMEc2eBxNmBwkLp4JisG455r25HFftejqktmi5dniWyCCfc9r3Vq
XsuEHXYa4NhFSUNJJdawtwdiT8MhV2Cqu3tbgiBihAIDMzHFK/D+vC5b4tH6WOQhY2rMgywHStkr
fcJIduzdeiW9m+EtGTsqg3JoQkNdFouJKInbKufhmdCnGjUVxp319OwqDwXuG5LWkzDzD4f+HEdG
W2c8yrztfYNipmXcUoxQcS3RQ9D5wjrYVGiYXdjWpYGmUnocJa6E3DzcUaYkYfkMLsaXxKKm9Sgm
+iOKezJEeSw7/3ClrnVSeGM/+6+5SpEw12D1ygAwsbE0IWMNooV9vDkqrMhaeTSToM4RkcpECqIR
7xnP1hrM5by9BxX9mAS0xQbTWhoDLo4nRG2hUQbgnVzAGb+UdqlzDUm0PF9yqTiPcU4BHKGWfKYq
9CTg5bbFXjqm6ICRQEx0Lt6NSpPHNOLa4Jx6zPQ0awagwVVnP9UyV9YubX9gYPjLqnNwKuR4eZN8
/Qac4ky4o1xivITwyWYaWbQbl7WV+EMUSqX75R1iiS3kMNHxkxouseoxVN+2lZARdCuVKQ/pqf4p
NEQgqDwA4gg6XJ92RYV/CosFWe3ohyoPxNm9bsMGFS9QXbWHHB94UB0ByN86b/J9MHVQefpVmP3e
BldSxV7VbLocYccM/DV9t5Go+VXd4ENJ5r6Hi32vUaoYsDhjydT7NRuyq+04HwQcmvuB4uEH6sCa
PM83N3HFrobUJSOp1avzxXlEBYHDbojsydj88VscT9lwbMcAzzUcv5DH3o2tLLZpkhdYaFcMjMUG
AOx01U3K4/kdHD6mZWI5Gr32CpIZlZ722c5BYp3fLq7KAp+aY0atEMEmh4hqjozKbuFM6kBie4jb
Do4vwW3+vqKT8RYLaSi7+io7Qz8Cs168/865gbUD+tZu6+RVEo2Fw+gzoHcNQguroIw5yeBNaq8x
7MR2hWhg92GoAFeI/lt8hJ27wecdmE1qyeSN0ZzGFnD+z+Pc1ZI0VXdTL5g4wIyMH5F6dCNWxl/M
VXndEmrh4R9OBho2zw5wKhM2HuTigkckIf2ugeJJb/j4t0BOPCLohbvPm5i+TrTs/7CO7H+bS0yU
G7xLI8N1nEqFbBuAd62QVnJm6ML4ziGOX6ql46VmBulRKMwKbIKEe18opNve/eb+UBy8U47Gmfp4
Mqbbs6ioK5Cp+uP/TvWyACVUng7n9Iu7P4GfJFnNBQuP36x3Uu1EbFj/2BECbvNaWr2YOkkLdX3H
9iZ+qNXtc+vTqKyVFbzsThAUkd3q925cyJdqPyoSK5Jl+KtsjEUOUlha8z+B/whrGKYWoeSGmx7+
mbT629xfb6sg1MNJfAH91VCc9qz85bfCc64gtIMoLGmAyCMpKTxWvTAn/cYYxRstOpyb+mAfQtlp
DfurM4qiwyeIFrcitTwobN3HwVAUmdFLAzUPoYNx1uKgkaP46T1cD4wJnXrx+B9S1XpAfN2GCwRZ
hDbaYgtEziycw/ecGk18AvJxxmuMw3H7faSNjXkBLTR73esJd3KxgdzqLjbbQWUerjsVTTJ4d19E
zcYf8YRilQ8Jntuz2E2aMRrcXYUGPzGhwZb1OBnV3xJfAAtRWEW6frJAVK43KgybvpAYVVdWiwdg
L+XoCnUX/3WAC3YamBfl7zZeyomqjpYSS9V823ZWRHXIxo08xRXjtGoUyTQVSCt77ouBReamJnAR
sYVs6DPyeEe9ozmOH8TDQl8EWLmRE7NHO0gh236bnMrqxKnSNks9RcjMC0e22IdnacczMQaq8Di3
fsNS9T+AkMV7up1Crq/ju92M2JqdwqsyaDKVXa6J2sD1CNMlE6zvqNM2uxNCnVJGR6Hg/ZueGSQ7
zzYsYgejcpWfApBm4pWuvhZ27goHLS2UgT2FyO5xRwcin2Mhyl7j6T4lBhRwCwWCStPVcoxbjMPK
jTJADa+Fd2Me3BkrF6ag521V467qAZlTusAdXzOBGHe8fka89mdoqi24Um0+iJGlWAK5tn+DN+jG
Jt31KwKnIW0xV8//MQSEfnBltLSTBtJbmvHqc7kMh8qz+2qv/Txcc0H3O1gu+hrXo7UhFYD8MX72
uYx/3fHv0x07olBw452kbhjKV9Aggj5W7OAMr9kClfRq5+wXYwFaM1mVJz8ibAqC6E0eo6LpFvwa
qokgiSDrznT4yrm25L0DgzEVzeDvo3w2o4f52wOaRzilM1TkzkYRBXFVJQ1nhtW7ilIDoEh5sXdU
2ni/4GI0f4m5KG2VcH3zxU4Fxp0nZ6B1rne2GKFmW/EFOONIEnGCbwvkJFXu+8y8BcsAsGW6hf1v
hyXxiOqg99j8+y0yLDb0deJOzJWrR5AXy5Q4LgwURVnXwQ/stt6u/1JtvM9svMfc50sABjgyrUci
0SB46Is5zD3kfJEGl7BycTld2lrmWAjsbi+I2uHUVI4cHrLbQWMkxwMTgQWht0xlVXJuesiChb0O
NwB0NUaFGgCTBqh46yIhQrVmZCGI03AXgSx46L9MwngKgmfTztu+4rCsEBW18xsnxbiT+bgmsJFl
WeivO+hijuPOiDnZPTzzszrY8mRknIHzhj0GX4aQlnlykhFR35nOtHAPjNtW4FQ/+a8yCHgKuhPD
/PJfkfHyexTVxZQyPVJgxdzcoEea+0P8ktg/a138Hxm8ab3vCpCP1vpspzOIl9wTOeXYuPYDic+l
qUcdVYJKNuVl+fy8ahAeaHRN8xZc+iwjOxOTFNeBvIB1l0NQwUd6yEhQPIvJfTFd1vPhcZ7cq8AQ
e8bygrnS+g0U6txQuip2+wpB2V4r9la4afRDS989SEb+NKFCseWwb2CAuglCnXdkGJHbvY6zbN2X
q6YFnr6gjNIkYOXAV0zitiFoHwnm10RJCXBIanOOJ2s6W1kaCDjKii8vsvp620sIW3kmayz+yr8K
vmKEwhla0g+qxgVt5j5XRaPYCe+UrdPARmdgLfOP2jQiEuJezNTOEQw8OAcWorF8bMhKtxVnQ4SG
3EufqBF/sT7Mwmd3EmSnRLCR/Cgyh+truC3nHY/96upwK1L1J3JBDzmD5j63O7E4ZMrK0SQq35Z3
RIQR6Z+AMOM49lk1FwnXeO10JWOOA8CYV2HQYex24gpTZpLV/twDEsz7CJaMZg31sBWFgMccp0w2
LYhtjc7Juf8Rn2X1zh2cZQCUNGgoscvj8uiz8WIb9vD7I4rm02LhaHpwPBczgAGBrUZkPCeUuoRc
OWPo7KQVaWxTiFHHoZMkcT8fmZWKenVi7rAiVZpe+6QoXzPEibqzchErv16eGezobNtyIipnMjM1
UsXG/b67t8L/RsgW9tvnaddHf2y0iM9R6NUI35EiTi9yJ5/A/Bm6N6z+1dko3YeyJGO2OMQ1bM5s
8bKfoKvLnUyp/6QeuRBu7hZAFqehyDih8C1JIL9IRPxDlx5CCVA/YF/zZnSjbZdU962sOFbD/lUn
XlHIbWj99v/NubYmWcL4eJHoc8l+CKMjswgKoM7mQezfIoSJI5baZqNCrbKgD7WJ8A41izo5uqDM
VmW5DuMdFmTEOiO421ytW+azPyETnUT5JPTTIuayh/B/EctOs7od8H+ZG3VJdotAKEvglgknLlX7
iHH3rEu95sKpI25EeUXq3lNMewjNK32RkxaW7bC4DDjKYNq2yh5wFlQMER9w+LP+HV9EMMQSN0T/
/dTwMCCakU2JBNssM3Nt8StPW/iODuHnFVHK8xEoqKtqsn2sK8JtpZJOBUQTAUvpBGx5MZg96iHI
f65Ss11dtVlfvltt3Bv82S0dF8/ZtppQ2v5bz+xN35w2hzyhppoAIzx5EqcGS9u30YILnNnkdFmf
qsJJlAcRVaYtxxBYy25tMO6Yn+ccB38yVXglVX7LAkrgVGmfLx8hUX4TJPiLjhD+guYFCsozqJCF
CieA3uRIFVQ7wdkbs+H78Tn9QuC9in+xEAayIKnjjhJf3pRLACTJi7M01FwkZFYVI6sC++3J/r2p
MsqkpiKX/8jSvZTgIH0plMD/zOWSTMQvwH1MHo24SzTV84EPGvBz5VHm8ODryPtHjIf4nUWb7ZI3
7LbO0QNRuigTvD7qfi6vGImM0A9fHf+DuGl9CcJYledw/13KGBTUKAVK3X7iI7dCiezJ3Uak/9GS
WUKSQai9/pWAfDP+cZqVxLueljIY6og8fLTsGbAI/UbpOIdESzJPvE1/4JW/yCD2OBraY0+PGSnO
MYBUqK4bFg/GFuCoRZqM1hbDxelTzpqKtcS+qBXKY7yC3b0WOsMNcIJUN66UTmbBorp5Be09ANn1
dVY/Z/+y82MMthZkvbYo1PDKrgrs0tWNTyVzrn4CQdKGt8SSglOt1U2oY/fE3RlX3eh1ZSWYbz/p
tkKF7Ca+mGmkhA04RTZ/ut0+FdF72TMQzk1ZuK0zqeSd9GrXRKTf4X9L6ePsY0dlj7XUF/ZsWzuD
IjH6i9ph7dF52y73UZXURECw8so4M75O7X81YCh2l97qaxzbIcx1LKrjqkPYWPKB0/eV5tRwesqC
zRs/e6PViSfJjKoxzmukh9cfvuVaBNsAl2ByQx59pOqCsZQEoRAZS0TsoyosRUShwT+KLmDYRlrR
e3EZ3yTPovvXKO/pkyIOh1m56q8jrUJi90LWINo8271A+5BpECB2IStaQOzBRzKl1m6WAnJEhGe5
yxpZC151IL5JKi1/6cIDTS0qhZJceaqBiXsFC7s0ibT0DZC3U0ANrd+wV/QCaQs5a7qqtcSYFPUC
WtkncqJfW0m8EncqDZk2DFGeQ/ihrrqn/GVeeAXA4ecpN1UwOBj0ny2K3qfa3PkWZ1oKJXExGJ2s
RTp4dnKMMkYtzVCPPlpKvCWh0tQnS4yr9aSQvOezbPCdE+Y2zQ6iVbcxsbQ6bEsbBRnRIKsx/IgU
2wgaDnt8uMs5bVJTrZPRUTqimCbB+w/QIdmEo6P1hd58E1IQsSnBY+aN+ZMY/Pr05pkmWr0i/9dO
TVXNrk4dfjRZlm5xXuPYh0EaHtYacVp976NwfpzbLz+XJKgTDsAjVAy47Cri2yXjCq8HBzWswOyR
QgqM3fvu3OYYVKh+GThRIoedBbGMvl5L3DglHJPwfwEePgSdgj6hurgh3V3516/JkOKnyUXYJ+qA
ZJP1W03DAUcEQpYcoHTICh2pC9OgCI1aAH5Mq5VeVd1OxDkb03N2Kh0aEV+5lNbpQmobL4EUecQH
mgPRXo919SV6jg2V0LVT4FAH1wdNu6eUU9Id7pbdrYxnFDpy1hAJnrM163YAF1j7+MHBNpXxVC4Y
hLSpcZbyz8qliPBnqzle3Mv4hqUJy47GiT5M3piR43ZkY1OHXBdFPjTDyI0Z2x8v7JlnmkAbATlh
Ge+nxK5Zt74/6cS4B7gYEpMH9DkXEz1UOPihEVyDwn/6x6xWD4dM6lnRqZsUU00lLreSu9sMBxfa
Nzkkk8Bzy6Niu8R5kpIDNL6IV27uw8K9w7f+l6IjioTqwfPPyS3Zzrpp61iZepm7BVrufGfBEdbM
PmDLdWLtaMU3Q8u09F3hrjwd/we/HjeTaWZIwQbpI+Xd3kNaWBMjPYTQmJnefbpU4g92AXkw4lgj
+j+TcF06t2oeaYfBGaIb4buZ2bIzsjOggBPoqFTO71qr8GS3kj0prWQimMfb7+aXn6pTjgfQQp/P
kR+dLldCG8xJVFUKTKdPlvCrj+WVvLruIwt1JGFKsfCKZdUWhtNoUbGxXmdvQ4jfoDl1PGI3zjgm
kp5deqFoUNR2wLjQrutJqAQ4KjyODzGggewHg3CwtAqmX3TNVR8T5r2u1jXEUODhJ5L/owsbYT+C
hrJSRyxs/W4J9BBAKnTIupKXSjd/WX3Y5U5JFezrOHmE33oHKFg46yzQlL918IhBW9zyxQFJj7Rz
4j0q/IR/Zu2M6kOo24i96XqGjDJ/N1k9p/5pSSmy3UTLQ+wVCPnh0pjxtipTI88T9tPAhAK3UJmK
pGktcLk6KhQfshNn2TKw6sRzBY0ezlOWB4oDKr2v8wosf/GFtJeBKSl8yarBtceDFkQvNxHI0OAy
f2C2HY1ifZC9KZdkkq6XIcnBQVIzX0Gr+20RiMpGSv+g5wrwskmYiODYWhayL0TUdiPZsJ8NHmRn
U8DjdpNAVf4qbco3C35rQhgGj+X8M6SSs0v0HNoY847M/aamFapxH4mLDzhsWAToZwahhgUlNRFI
/bMYXb4l5rHPYYnX4ItH8CtBrQHXM+AoeRqmzN31/tZGweasxlIr7ZwsZp02ufLiymJvZDDRHQ2O
lRgj+3aS9F0IXhqJ/j7FYDzq7G/2HUmyz7ojWV5Fk4e+2pK1LmN8848hZubUEVnyauypW7hgDCXM
I44Fw5a0jnhsNVl/reIUwotGOZHfVetN35/c+gGV5Kl355/jI5A352Y6KBjqFB21vQn2KPc0vSUl
jM46o0nGOZp/bXV6xLtzj6qHUjLhZhwytcChUOQrIRu6GH/IA+9lmD40FnYHlIyBWZNDQzOS0VrU
lh73SdZyG0Of7v70+KI72g/FMO4/Sg/+wufiEyF8mP3eXO5UpU42FUNnAXWoExoY7eIdOwkpJXB8
9pIQRGziWczD3gZX9r+E6Tiwg+I2PzP+rUtKp2KDLjth29ANq1kWpw7mlDhUlCVuRTEYe/Ah+Pab
9bFUv+8ISmygC+gSZMyVVNNo2HOi4Q++3FAMIfJT54b/wCxD+69d2EI8MTed8SLdHsQ9ArxC4RlL
YHV3MVhNrgsmABJ02LCria/iU6sXSC4LD/imnTO+IILmSXFK/0ZFDwQ+SD69QVg+bU7j0SimnwiM
Fh/Qsjq5Sfkuu1G1zzGNzfQBLbdImVY+xB1i929N9anfCpHYiBVrbhWWreYmEbG4/S6a2LwzcQie
voHczzxCugd9Uu2cjP7Mmheyx8YUILvcYFCCgedU4r1NXQjbwNGg3LTQDxEAzzAwNRv/q7pZZTzm
mjHrsofnxF4akkqfBx6akPDZUpzR5OJhYOPuX21JRRI6DsmOcm8u7tRf9iQaKda1R9tWYuhXsKgZ
JrA1K9SXyRc3596PRO0ZP+U/SXDQwL914XA2Iy1rD7kOfMpMJh+XE0Qaz6a3n1xfiUs63jzhEqlX
1qUBt7eR/2RNQup7y6jngQppPOTdbfIwLLufnA2z7WH9riKOGx+Zapxvn6nL4z18v889hewyQHSa
7U0Un1ZMcLIeK3z9Dzmu89CwH0qe/GluAgewUQJcm+9VOthZlOp7ylV9k9RxkkoN1YZY2KljUE8z
L7RVEZMfg+O+Sz9e3Bi/BuJDv4fuAh6OhIla2lsSYepCumBhdCJpb3uzLSpS7rdckyxkyW3bfEgV
MS7nw4zpL/4krB7N9CvxSkNqYCI2d32TMfTxx9DY901X8zGz6UreQmBXmVtmajQMG0hIR7X3NILZ
5x15KWKckhr1Umg2O1119DlM3m+yDJb9hPCmqPbzCIXzPceuatJKgsK6scW6YMRREcYr26Hc+N+V
nNYfUhR/hMBoXjQwSDX8tg//4sR9FedAtQz9OzkrDUSaD2NG2/JHjCxTfc3jhHj2oSBBZs3bPo1H
CquTRDcxgYg65GnZljFAXNkPYAdhwotp2gp3oyvEWDTkZaIjD56J6sbIovLfzITyjHoGsn72cAdG
JTws73hYpZiKBax9fPkU8Cvhvg+aAE/6//Qj5xqZarKsspbXadTuQsGjvpiWGEN/aWQsykMrf5/7
+7VahO51qDmBFuyVbW0A+yAgkqRz/yal/QLngTxJaqOqdJL12RoOq+e1zIpgWCcw0betxapWDCx3
1c8P3pk/C07a6HxUgQEg5osxseNAeEiNbErMGmnK2DicHxashzk3fRd7MS5+sSiJahpBYbZmjHYA
ni0PDGmHdBgaYPrGDfca5kvgZgmLBQu6IYSFFDQoIHzqfOWosnbkO+aWKh87sUY/nOxUP9vBf5ZY
HaG5x0b4GgCj6Vsw0SDKFRbBRbJKQcutSeEgijHdVTrz3/iCOOgBJpc3Q7hEnu7mw9nNPnaIcueM
7E1u6UhXh35o9aGi0oSEVqp9s4N1dnAyeDQw8/ZavDqlASChL7rC0x5+FK7wq1NyZ0/XwQ+nkXEX
nz4gBvAsBVTjQbo2J0rAkvGqn1whrCcrbiH1QS/9vgGE9RyslHHDiq9INPUGnYz2MWB9JRyvF810
GwFozexfUywAfB0osUttS2oP3OE5EcgGQyd4KX05StohW4g0ioqUOuMczR+M6Jt2hui0Ub8XyKNd
eOmdC5v8ehxW35akmiWy2kBSKsBKZccud6z9WJrEwuwdSee2vzjPtkKB/nrhnwzf/0jaPT8qnXTA
IeBc3lkaEcGn75vNfL0lUOW8oDSxni2qBsNk+vcOw2TR9TYh982eQMwtwkmp43OOw0+SdOT5RdmC
ylQyWwbbhDx46yG/842yyXq3Pq5yyADRilcsOr+AjGNyhqTuctNL1RVTwqSlf1dgWK1j417GHWHm
p03ylimMHovGMduoN67TThRnqOgQuu9iCSJBZlu8/9W4kmxo8LJmP7IaRfujQq+WCOBFTOXrs8xJ
+AzS5yx6ARQX4gWt4c9RrwvMt6Km1g4yXDvWlUjsft+S0sGxUf60qR419C1CWsX+oNUl4a/CK+42
ZetCJIWeCdQRrq41VK/JKD7Vqm4d2LRlDuxRFly4aWy8JVi53psdkUHb7N41qFnC0x6YQ5afj/GX
cD8Ki5ywyhx05w94OI7o07VXccWPfej8AA9HWhbsJsiiKAK14ISxrFmXj7iSTDcYsGNwaA/Fb5Rs
e2e3xjCh/fbxxT+uQYSvBVM7+MPslweTpvciLmjo1T0DKv/oBluNCilHDRZKmVvzo5fb9nQVCXCv
rsamo+WrgosbeB3nXZtfvUvSJKKjKlg3kVSl7i9AjGLi/xAWkWIAJfp+TAypxKb9dhL1sIVlRN5J
PGRK6YYR7mMIpq5+raQqvsW/Vyt0PETsd42bcCo1RjdK+GPX4ZsSrlpgl4cDRfMeAEs9Jr4chrMe
oXLErkRIIziRQHX2wCcp+kWOa56dZsMXL+S2uRhUwPfOWGXZkcJzBT0Vrm+sTH95RBT1XsDGPOH6
N1xnKMtpSvXJ6vcNBoluit9NFao87CN5K+TJSNBiMdSLlUfDqrXsusXvn+M9S72S/75wsJkbc2te
kHo29Y6dm0h/Aw2h0yC5xfFDpXzwJxb8XXASoCIJlpfGr6d+fTWRRYShK88pIQKzu01atnpG3yaw
R7gg7NRHFACfgTeeLCdqjwVtm31sX0gaNEn9pFkByzDlvJNpXz+bYWhVucqrCNEVewQH9VbUO/BR
ywCdejYky6K8FWxN7cuPsuQDbTPHByBf+wd9fbPltZvxWyNtW11Uuu6M6kULtgjLZj3SIpr5kPGV
Y2ArJZNy/gmsO7IydvaIcgw2dHMgtvuxnYJT8IM8VVO9VOcjSAMnuMY1bSfDAdgQk2rGx+K9DTpl
N1cZz2vmWJXd6aEubEQ7pEARMsSVKK7L3r7VJFZQpNdmKWn5MstLevltdgcG1nK+jEPusAbAqp7z
2Fcz7En5H/Lj+2HSnnOEdToZmWWWLykf+usWGLRrRQDKEYN1f/kdP7PqNlnydlIThmIE3MdZgBs9
D7p79aAkoNjGySSAw984vUptUiwcmRZScfiSa63huQ4QWQ6U4vdvzkx6NMLZWJvcDHClpZZ7yQFW
4Vj5CcA/ft5QRU3X6OfWb+TKQO0kenc8kHgcMfrisgJ3ADtbjwFPQ+ym6j2ZLVmOKWgSGUmCvqH1
8UOdLsoqK+9McS8umucPRddJP2fQ6WAy0i6ZAL3sq5L8Rz+F6XqxvNfUXbHDCx+smO+d0IpJm5Li
rx3GHoxzNBckFsuu1/OFNbEjjtpPw2Gv/tQ5J6i8dzqN2/jv65AY55J0IlS2CehYFxOzoPhuY4ZW
SXlpKrA8ZIDj3+loyaeVCaxkLsDaSWcFJOLkB0j0DucPoJCOAbPQ7nZDAkf00aunSzwudJC/Et2C
IzIEnzgMi2caTq+hieeBQx9d1Jm0KJr9KEj7PIhDPtyRPIrmNjUxbhYFx7MaN1ImGccJBCUKT5bn
myj90elqcNSPAu521HsRHxwMlhCUS30AcJvyBblCw1eXXhS2EUFknw4NBaWfZ/dCbFczwrZz4Pa2
V+eRj2qJjFkZkqryBueXP94DM1vcJtT4kJ9ZjDZ9iJbHMcHqm4Q0eTj5Qe80D4J3jtLrZDcJuY8G
uN5kpyubuYxRSDWS3q0951KJoPRLn9NNNZB2eoaAL/wc7ZK90EsiN98NAtgTu9BKsW+YwRYCdeRP
1xFszHOf+b2d9w3Eyr4jgwlfAK3g/Z/ir1HDMGmGxYa9+AQB5OmMGvwueyiXqNLf1AbEXox0Pjwh
/s/5ZsPkzVXgcZlGj7BCzJDGidy5MzB4FqFSZ/w4esk6iqwxH3GGR+AvpA5JWDItknW0xWoksPLB
qa15Xd+K5lK3XPrMiJuOIh0CoY+Rv4+7og7OTMhKoMnpxmTxnIiOsfsk9hx9hqcDyE0GEh/6oR90
5m6UAiDem8d+B4kbWqrBAB82kY77D4+4y1Ded6Hq00qaQx5n8Q/l9g0El/9xQlwcwHx8HcufrtJA
F0OS2m0iYKcdOcZKDbybuKHtSupR6ff/RXDzeKkZn5wY/Cx3RexbZssnbMmprmFQxcCMPv8S28NZ
FXCupzRg30meQj5d1JJEv+jBjK3ZDayN1pZIqPOQWMs3d4agt3MLVzy1RpMWZ1pHf5Duyx5SPb2j
bpirie2rxSMG4WCbjE+yQOadb+D965t3LSLZ/1v1XNq7uDdEjBOXn6Ia7/qlOP2WADQ1zhXTQT+0
+AMB14PkuvX5va7/+BexhGnbMZoz56Anjw5MY7wwtSpBrFUU4lIVWy9SBrMyO0E63K3w6jvrw3ft
rxfCdmbeoziVyCTsZVsDpNx06zilpkwwKeDGepcL1yqZx9kjo1GX33I5j6NW2RuYCLPA39mAT6Am
bC0XqROuxTsCkUc2ie1ZuNRdi6uc1Udfai+82Qmq7TgrXzLwpSkaA66Lf9JHXG5m8jup4KwH9b0i
S4xVRoqO1bxB4I/L0TNgZFg7OnBPPC3dknT92FcGOG6+KxqWsS9UacqZgik2EckAdm9HgU0R04Dw
lwCIIblinlE7FILlfKJOzpNmKG1e08IkQ23376i1pW0wn9FPVk6fGx9rt4hh9f0vnwfmA7kyFi2N
sv9iqnLN5jKRQqaAsiC26o7+OsXxOAE0ugKZT+JAdNaLgfvH9sL/C0n2+qor0/fGMzu5Wn64N5KH
w6x6hMjfdNjtySxVOiZUE5F7sUu+7OdOb8lrCWIIpFQ2Y6r1rVqXuXnrDsUUWkEEc1kkXlTTtK+/
GTMwUeVugJFw9QtXogeA9SfUvKAheFN4rJ2krUF9Mncbh1koxOMSnK53scc8YrUQ1J9xMrJw75B9
e6ZLjZRjgBjuLiSnfVSJAky5vrCFQj9UPRg+LNcjfO1uJVOHf9SXsCT2mwbo8CjiyjT37YTgOwxZ
vah5L7+nmZ2gc1vARBK+uENS90AtdulnCk4GBh4hnSovenwP6/OSEMm1NhlCx/vsRG8xaRjtLQuu
0gOkaGuVbELxsja14F0JIsA0kVEBBsM/3PLuOD8M06hxS2T9dQkkSNjmJDoony6Kswv3GSKXnM5g
vCJ2VkGkI00NExxxYXOg6TfMOyV+JPngBm0I0/JWK7qtdy/adhHzPjlk2ark0Vh9IRkep3TVcqDR
KersOgw3MW4wwilsEFSIe7xxss71FyerfM9SmECn76potDPjL/AtIY9JDlsYFSXcI3CIGnYt2EA1
2olJvaMKb6p+oNTe5UhNm3ViYoyC+Zq4jSMTV7riYmw7IFCUU16O2Ef9ic45qZ54WbpDz5U83CKX
+XaIVcEH4IKYH8nx0UNwpgxBH0KaasrKHZLUVErwEU7Bg3PjaHoN7lNgzHf0ZZ2zTFC84F9qiyN/
LuU9jOmOyOWO7qNbmNii4aPGqndQOoQ8fYVWQRninD+3jdWDHzYXq6HDUkkFmYPmrfpVrFvu1yfv
J6CkrFnO0UUtAhc8QqMxfXiKxQvck3sWrMEdjMryC+Xv23M9LN4nRXfqAoGaTHFvWAVuLeJj2DqT
nFXO79OK33X8l6eHmM5NZqI+OC+tVFG/gD2NFPdS6vpFHE7MR8Mb4unEHxXGtIfuzsZWdCRqq4Bc
l3L9t30eoEYDRUlCssefN5+7iJcUD+V1rMyJhWK8/Fv7CXt7UBvBP2+scQ+ZibAoqm4NF0n5o9WV
SqqqKPSTGDyxlvrbH+kuxR6cteh2iDKF0kUnJtFBmlwPL26bWWJrdaT8BZV0otSAJbuTHMKkYvHe
MAmVE/ePjMSm+I2ZTHa+b3ydE3yxGzDxJ4p7Iq7z9fqF+osQYrnwoqmE+v9LWxenKA9Tx8VpjYU0
FqoHSq1tCX7m4syjo5t1WsRkU/75pGkmctykLJjCFg1Q87TAxj7sJU+/KXwwMuYLHollq40HUeRr
/Dt08+agYNQ0uaCKwYAMD/DqrPhovMVgaFYYyiIBETPO3Erx8ILv1fecYLQ3HUqQQ4Pm9Ui2uiX1
g94sjxyolMlbZLyNqsULy1HccxgoLcpBYow83L90vf2GzCglfpef3L7LhQZ349HskYqp9IRycsJV
0e5A1V41ccLFpJ9yNEiDbN6acHBhI68UNd9xC7GGykSZ+GAEO5OQYy1ujT3w0RSYbWnGGak6rr01
6OucXoH3yCRV3kANqK4wtHRrqAyzxEjqKkrQKXpwTfxzD4rjbQen+QfMYwMnmjhIxEtCgMVUPaRn
djkqTcRqK1diisSU/3xQTNIOtCPB9q+bitYxH39TjOU0Zw7NXDPNL/aiekZyD/WMyMct1KSYSmEm
jZwqwFq0vYWpvGcj5oIsPJabN89EsC6vpTtf14iMvUsLDg/VapEFbipwE15F3igj7gF/fuEY/zgx
0jXiBaQLHu2b3Ygb9D4SIz+w34Y6f4kUPXPOki+3PMakAZWG6IgoNsoWI/cSZQXCdEYEvAHbC6hh
dPyBaYXwiD4FdA58760qJUi/KrjWALaAwncOeCnXLlIUlJVkkwemI7R12mDnbfOgtkCMzbpL3zFh
rEqBVEKNPHvspachzhDHtMqChcjbM9UkQwMa12DdkKh9smbbnsrhTlIn80E5yXunPU91AkBVD7zs
rOjuJQ8sW99sX0TytQeEamIWNOZ9rt5lxlp3sqPm26t3mhIwH61isYYoDqaVDs82z73b6V8WsU3f
QsvI30iO3K5nmESSasT/ptMo3k/absFA20ltzTY7aq7ASl6CEIWKfP+7xeekDRzzVKVLPw/B7bRO
625Tw7aTQu4etUr5CwnEQbZf2KsO9im6JpEhWdGDgLIzc+S0NepgE53ATFw8rB/mYCQtcLFc52cq
vRceez+nGHFD9M+49dk8lMK1rjXPNBhTIGEWl93YjZuMtJD22ce8CsG1GwZx4Plkp++SgagOJ6cL
WklAUNERpx/y0OgnKwYD8plm3G2t6qgtLgVOOAvrxzIa0UzDxc/3inppXcB52hDO11LGDA5u4Yba
ss1ZEwpEjz/7B1DDLVbqbyAk8ZGnVuw80dlaaCCClcbEh2lOqOpjfe6yxy97kiUTspWTPUYW0G0j
Sqa7bCSvKHdXgRLwi7nSAK3AfLv0o9cdj1ApOPhZd/mZIxPo6aVM5Za3wI0eUOLk4f0DzQxnvX4L
2bW6mOlohY4s6/WacM3hWli2DhMe2tmDaQJhgi9fL0wmgidXNPO4+wWtp+rjm3Co1/TxomNQw9dR
tt8SDsVYHfSoHEmKFEgy60ZFxOx5xLVTgxgait3lpDq30TnRn//pF8c7jq70FEGif0Lrtxvm/tBq
kUdP27H+46F63t3gqpcIEXvMd9AlUo7Ivt2E//SkJgcsG2JPbFY2JlaPJr327lMVSW5MHmXq3TsU
8zIg+axMO2PwxrnqVWtT3slwvgMuS6WuNi3J8JoXk80eWobZ2uRuxHUf9efXYaMKiPmgkWLO60gP
XvXnH17kU6+U72GMBTtH3OxxcY6QuO/ugHYWoWNKxVLhoQsWnbcRnHq7ZG6dFAm5cdIrjQXB8cQP
UHuvxW5pyckY5VeBt4gL5jLop4OlvHkajRrnftL8M46UbRgHhwXFZDrmVaVfNQAmpD1osMljfvXF
TqmC6Dant+Wb2HHmcp86/ReA2RiVtgQXt0/TclHlYAj4ZzUG+wdoVmypx0d55pfBGGx989LfI3DG
MfsMqrmj0W11v/MMVV6IrYwiDZrypwGUlM6O5Ioa9GnCFl0Z2djpQubPuuTQ3rZ9jAg1wzqVmpkF
W/h+kj5nr9987eKXQfGXG0pQRO6XBFB3Dhc++ltenYMABpJ9G1+KN9u9j8spTsiVohcuX6D/X1AQ
eZ/lukAEmOTrvzXYSAM/726iHNCUc8aMsjrhqqZIpfTdE6TI+a08Jmv8Kr6mETYSWMmgO0RBBJZT
PFAWSpNC9gxuDhMFvNv1H9aJ4OSILZI2WNAaoSWP6YWW9SeKmSvLyWvfTnU7W6F4FWh+c9+97/ZE
Rzrc5ua39UsOqOdP9O88mkZ3Hq2Ym1n/tDbTt2gzzDkRick7yBcHzqRQYh9LQC3AOAXKi3Jr5AX+
OSP6Xx5UKPAkxWM5v83u00MrR6C9C7QQQELKgF6BcDE9xt4LLBcDDslJy6cOsc+jV6DNTKH1zBUn
aSvUq2AFWd/7sU6NWimMmb+YwKNdBU+mIyTX46f7wbk3LKgWkQL9HK3bVm3I++rSqW2s9Dk6er2D
Ybd7FW82BsCnPKG/x8sQbf7YtIQg5kkw1bTX1NrdrEYBJjoWvIXRGlKKPqaRiJ4uVVXA7dPudmqN
3eizJpReiiFzRY8oRfpagFfpiu4x3YKoDDON7yFmvAfs6dSJVzPvf8HeLETbFm+uQEFR575143Rs
c1/AH6hIdWzrfbuNRjnT51riNwJ4h2AAUKlG2+FyW6KjsKP1sKtMsoyIlSWxQAhxSxluQCHYC5zo
o+xYIMcYa4Zsgs/Ox+I0dhiBxvhoLzT7zhAjZD9LhPtnvzfL2muqPUaRRINer4i8l726KA9NabL/
v/MSFcPC/HTBS6gls4v16ghh+V/fqfMM5UMChQQsBlVt0VdeN5UN9SPj9RnHACsxV3dN4seGX3hc
N9yFIUCfR4xBzpu9lzhZTGywOLyotE4m+Updo808jRnBkBY36HOvItXW4Q1WROPrAUAyz2HMxCnT
fvF85vRupckKt+5HJhd6pygcQSlO+gSKix+/k+ofDieq7dQd/Vzqm38yj50DN6RJfjDgIQ0Q51w8
cCC1/swILH30/j2MVXnz68VLg2ddP2tRsw6dUcqeRtbLoAeoLwwdD3jVh+PV1rOMRoEKcas7qfHt
VSgJ4VW3UOVppop+dUgbdWkXL3ar061ZBk915CuZa+weLIs1O8jYr+QveuN+uO55zNqO9dgq971F
uiQvVb5E38JZiLKogawLtJK44ccenWY/NmBHeZUv6umgLq72LOYhK73sBuYHWU3OJgjyiXJXi8ry
14xqobOTBmByodl+0D4+q+4V+jnSIXEPg1SFg8x5T5z0+UvdhXUwYyGP/7zfoHJ4UqlGvpLu2Znp
p1XelcZ/E+zKm4p2wr1rs/v3ZvcJwi2U9BsX92jharP70qe4pACYFhMzNPwqrtaCgMUjuDW9X1Ai
VGzsjYQ0tM3ncSePP2rwNKu4gyyPoQgy/AKZEJd8hYtQ6vjTmTqZ7bZkK5E3mWpID2+SW7nfRu1m
1s58GbZT3A9Jlg3Wkgsvm60c5k/cvNA2NIYA9y19rLNofGbAHXh7gBIqoTOHe4La1ikOhMTg45t2
7o/D5HYb4q2wekBKu58tFqcgYNdRYSoz+U9fadvFpT+ezRNDf25fqxqvNEM637fXrXNbWs+JM8jY
ZGTFUGE32azlwT61taNyPpNVdBSNUodSU3I7znjBHCiyeBCY7kyanYD8jU6664X6OYyxnLdHOL8x
Fdh+3ZsPa2PBN1a8otvrrLETF/q1g72Zr61wX+/12Q2DawAuMToyxMo/o9tPtGpZ13QLU1YEKz8o
hAHz/MZO3f2QWJYRRY6oqGKaw7dp+XKZlIotVJ5MUQy/b2yq2mnUEKjnKZTVolK+Ujmv35+EcJ1k
pV32AfBDbtslArEp/UfsImJ9HjGZjWw7uSiW75x5niQmbSB5A5k3YxJZ7Ty9Vzy0/ILPo1yNp0z4
5U6yUfkWcBxzHecll8S+NNcOd3AX2aq5luW79Z8xmBgiWQDOd69wO9Ol1qZgwIPYUaT7M1AHs0gF
XRmt5PKMIi6IWKP5YMZXmF+fygc+T0fsyrOsMVHsofNKnGTfRbWJ2iNJVPVFxiinyPWLn2hFUYmB
Fjjj6Xm5Uu1VfK2qgGk/NkoM71n2QiAmUjzsjXC2N1PdDzGlzELIFhQi4Uq4vtaUUkG7A7yFCx2N
yHbOGOwF5V8KhY5ClkeOQJk6pPaDipmcdQBxyUjeD/fk4uaMXq63jSdq9OtcK/tpLcBUw1+guwU8
96RY6rvWgzrCP5ZQ5zwWBtajmmVzRZqiTlo3Dfjv3CdXlMTgB1tlveS6sDdq15uVkKdLVKZmoWT3
FvMr2P15tu6CjkwLAGZCNKrj53tmbmIa6LFwkeeeHWlPJ9eljC/wtUmzs+ZBxQNceCeiQ0ex0vA4
DNsdkRKB+Ieu6KxcEg2qpp3zzl82xFfziT9SmkPtX4XplXHqSfdD6FJvg5AK4P5Re9lZiDhbQrDh
AGho42G92a6WmoiqmecXiuaf2g/FgQYQU4c7Ed+fJAmDwXVVz1BijCyxWKteQfT4gq38KMS8tvFl
sETGYyNTKqRAF+lFT01/m2jkCqaBeb9O8bzzuVZajJnsRkW8AY9+1k/trGcL27q4tjN/tiC1BqTf
npoUWNBSEE83XSxs5lsYXvDjfekEkzYrwfoVflUp8j3zVJbIDmmDCLulPz894KVDJ0jQxtDDr/TF
OOi0KB/A53fP/f0NdrTqsYWF9kbHywXPgRhfYT0DVxofI8l2flL2mtvmZr3n3yIB9lEalGGdtiee
+cmd9HtiTYDznLAtysOidpVbOR0LKxl0hpHAruH2jLdivYFt3VRYsZIb8fOqcvgkPKA+R23WejEB
BRWBIfiVdIzgps2LOksbKyKQ+z9BOu8G8SRf9PbbLmf31mdPA5TQYTzXQ4+uKPDCNbZE98Lu3yVS
pTqn26jM+CSdAly2OmoND2PzXg12phWVYDOGrvHLFkzTnw9nzaaGX97f204KLI5Y3UKWCJY/dJbu
cKFIXODdvzm7g+S8XhczmeJhXTdL0KsZEKBM7pFMA/84+4R1IspNAgt1BmFz8BNBVxwSmu6hP8Nm
Zg8IJOsw5+ZPqTmjl7J+rr8AxzvNFSPfjdG85sc3kHkP9QwXdoRzu+jn2vZd/irFHAVRioE/XB+S
AgpkAfG2qHN4OnEjnzgG2j4imAE1PLCVax5velP7sLMhfmKOLC4Hbq8R5THqwS5nv+XnWHPoALtq
PRNpoXufNBeq1EDJlGG3HaXyGKErOKvavKtIYRzZfz78VyEwCJvKEvJ2Fs52Hq/dVcL5xIxKozwb
MCypmKZtjCmhHgbrIXgyBMIO2XOAjx66b1QIvwFweKKkUKAFUE+tSiZzVRSbxPgZwuZlltRdb0/p
JeOqLbuxZRCorcoSqxz4cpO6/Fiug6dQjdTvD+hJen/jUa7EhkbjCaC9cOgLvq5z9iPnBFZXTk5B
3UYkGSnq0K/uScg95p0We2YAlPEb73DifNUQGzD4IXdwQIgtrvxKZoRAI7WYg4YqOZykzUk3Ie1V
LZplK60IvHijpxOMKM4kyz2nGhDXWuv/+wpploCE/lPV4V8KVU1ofdYJr+4rRH7QDEJ+fuV4CgeY
qfnAFxZOjBJ7y6mO+sKgL0neMheO8pJ5tnhWrti7cKpB9YMsvIBpzYgr2eNu83ubrydSDCBJr0Oa
05tuszn4NpFqhoytzQwjPZJkdoNRubNzXupfbwnnvDeUikOxJxYH1cJOWly998yd9pY+hnNNUTgz
T6qz/gZyJm/1IaZFQfRO/mSTCl7HPT9cZrCnkEC0uCwcFpl5Uw1gZmnGaMX+SRdq2F8EcGFUefqL
hJwyHyYOaG5RIQC35gXRDSyufUP7ECDcqjuMNDDvn15jg2CvvQzD4orJ057uE37wwWe7kvZ/5TWE
crYZjpO9LDFh5vvtjTzkgXxLQFXwjejRGnsIXK8fkwq5ofy9esKQuIWSQ3B2Y79vO/e1bb0FCrzD
HYOgrBaZuMKWIFsaQxd3sVXNVRuSBSztVid8oei3uvXi3/N2MBD7F5RrxDulzoPIoOk+jI1yP7AE
QMi2YMPkqpmtrLDt7/4Nd1crqgDIwhE6+zZ1lI5ZuGD2e0aa09nx/VgsO7n7qeOh0Jl5KWWv0rPP
oiKiGDl5VaBwHXiOSBTT3mro4agjQ9+t6HW7kHBGBlVM0NCKARuNFUwaZreLNWnfR8S5yWVz8eG/
Lp+anbsW3vt4Z50by3DqqkJq+cglBgqeuGDcp54FURTLfuTtXLwjSPcIFco1VJ38v/kduNWeTVMr
RjUm6ZP0sC62V+uumn5pejzB0WF2xk25x15t7X52dWE0icMt97Zwtk6RyC+0LiyxY8aT0E/Y6HEv
r5zqunfm1wsPMYpnF73xgv/23Zk1g1RYj4ofYXBVa2Af4nv5KN9bVDJb8LrNbYyY6P49ZseO7a3k
C9Wpx5pWz1vhGzaaHIMwZJGp0uYYsc2ANF6Kgl4PwQBDRkl1CGtBaDBP2zFQrU74VZHrvAin53at
th8bUCyJy4rQafTWYoUQ6N5oBFJdDseiz9voYQwFu9jPzG7T40Th/42xSQyuYjVk9AC30jhPdWbe
C/qClOejwKjA+2NIhIcwooBinoSLaX2yhwxoF8eqUewNeLNq1Nm1jCn/8b4eXm3iMyFRd7f7vwPO
QVfZ+FWtzbtBbGDYnZg2iZivnfY73iwZ+xLXoTSKbUiN1IKut7NOfFNKv4PGY1cmyy/vBEL1Rqc8
Q6dwX+ovj+zYjN1ZBXp/8JEXDgBbS+ezmrQYWnyakRggl/LLQDMDhDL377DKB1alptDbkx9JizZT
kG/A7xtqdfS6XP8sd0uPojW6d5Vjfk9bvsQhYKOxFZriJd1pRON+iPRjAvk+ActRKOCbDKNwEzM+
MKIrbPxxKEeYQ6V5pjtgRNVkLRsFxUEZUssmPcafc8vSShBohqXt67lir+GYo6tbCkzT+jlflAoQ
94jHjIjbIosuWrir9aIUXgvrTwtpnNdMfDtFfrGUrK/wUNYsD8pxBuY5KrFjz4Ar4J8Q9/gDst51
vxAPpTWKJfEnoq82sAiyBKa9rsCjrHgFsQh+JTMa91mh+uxKrRNS6npMEkMaRc7c5vkj7DOL9VWR
Rhi86kfzt3bpfAop00vBpfXF1xzrNqX9kZewWM1dKmwNpaBcc/di5mrBTlQjLxc4hf/KHtAFUOrA
lgKUQN3qdnmNPTzxLHHYCWbtBsRu92vH98IqChR3HI03AUDD8ucGIXHzgkcvbsr/VRCIvnSISh2+
2hJQ13CycZ4CmuiXQAsML715knPUm4N+abj9KKl6Izzva2280BwYzRtgiYkQHOcqYaEWVFvVXfGx
cq49bXVf9GUoSpnj7TVfpczvOCFajS60vUE9QhL+ZTeFi4u7cEsnGOQNmZXaCb15B7+zF7Jl/OzU
O8NNJeCl4mSA+GxjX7r8UtZn+KCfXmvjbzhl3qhBXIsyg4peWqqyY/jDIvYBNYi7jUientzWN+Ja
omTLS3Yww6jWabhMUvqIGhwnxGg5oHZHxcfC6YRDWTI5KrU58CAJeJc7KRho0NO1fscqmxamPHMI
lDc/MOIPychz2kfNgEmmQSXJ/oACxz/+WLedyKnyeuMEQ49BS0+MwAyV+lqdvXukBcMnDqHQqt2I
+rmY1jJ9XmjmDJZCa5PAlil0sQhRDAURgLuaN/SRve/zbHfEYiGYFKK2LQuFky1OmTSwvfj/qZBi
8r108BYg7YY1OPgLybMYWG99nxxYZp2OoawrrjZFKaW1IOLMd9D9pWLBWeIYiMFandpNsBkRD1D4
j2t4YIerNPKJXLiur1nxrikbJMmqtH1eXBRsklG4MM5Vlw112Bl3bzhCdvr2N8Azzsg2Ncc9McCP
kvh/6UI5V8MkxxxZDT/D7ki7A9Wpzc3KOIr0Z8k7Xpz7GY7aP+fzUeqtdQ1GcQquuIYmCtjM10nC
kTKkFqX/a/V7bdet2hD3/qW+Jgh8vtOYKupbvCgqHJC8ykMP4SNo43nG7veNjPQItNOeqEcx9J71
BXfIejjT6WjMvcigi+7ADYdo1oTK+4mCBwcN7/fKNVNrWrH2UxKekE309nKnXgoWXTDzf4MFwcsa
3TGWYe0CfaWH+nv0+8/J0rHywIYi2vdnXxJK0Te5PPXM1nCawrkaIxjpxYXXZXo26RJ7BjKB4Jmp
7Z2dSKBdSs0EjqpHOjnebr5EdPQOemgaUy3S11T1WkhLk8SKclwuVd8ddeRvpj53we7+/OinBQiJ
9RbOtlzwLt5eizBpBVOvKnhpOkPRXcFKji4s4rhK2XIGwzK2u0AJi61zr1zUExIESaksnRtuyLN5
kOLzvTleoCc1jY/HzeUIrnevnrNq06UOxILuRIFVpTBEh3h73wIYKheMfVyt/qYuVq8eAqk457SR
FegcwHqehXJMQDQcw60zmrAGUMwl7RvG5Ivb6z8aoNUt8MnPGUrOi0rPMHeisZ9HDiX6bQ/BiMQl
YDNjnYdZJMrazkJqcetUd1DBIujFqNluUXEDZMRwXDia9/1G3S8MEtHeieZjQus7mhhETZob1i5n
Byf43Nt3ysKzp36bfL6QyzSM1IBQW3eJr9pqeS8PbA0+rtg8qL53V/YN96C2Usia5XDoX7Jb8rsp
ox2oVsS4xqqCCbIslwVTYjaOzGyZCzoa8FniRN7/z3SXBm81DoptQ7rrHjCIEaRY7YM7UPD0fpMo
O1aGCH3LDrFK0f/wZ9l0ZEthFH16w6hMMhDhIqLug4Q/IIK0w9ExLDa7671ySF8wUyznLquJtf+w
ordejJnkmvG6eaZN6Mm7t18DJNW9UYqRpdD3nJ3xl2JazoQqdd0m3SjV+L7EJ69cs9SmO0zjeSXb
jfB6JQ9uW6hmd6mLLxGrVux8ghIoiE+tJbMUwt5Kb8hn22ja7H7VsxgHSfG/5Gfggg1EOoChupA+
EliZBZuBZX053TeLQEhWIPdPflxJhuI8z3qIJkMnGJTDysasxdY/absYeRqf9XhVC5S7VJdRoWUa
oJAnbFrmHkI7zFc0a70SIHU0VAXcg6cB3BK3/bRakvq+sfMTI3LE7jy20ahYiZEvwtDPBtQ66IwU
4cMFOwMnzlE0BKGHK9FmBY3tfF/GRVbY6XLiDLBH41/+EeYnthrdlbTxQt5VBbmvNNPgnen/syaE
3DBg/Yd+BtDV6LyFgD5tSOMAEpde+mPV7xabA+cGR/rDmPoMZl6DwRudrjOVuYeJBNWc9R6hAgah
UKr2wKNWphgU+J+Q1hDbCkncVdsmMLvELDwdjHGtQOrjEifClU2a0Vd9CD4LY5bjUqYsS8rtVKPM
xmF3FiCxsYNz4hlwphOZC+RvZlp3HcCNDa6PNWlPZCFH3gLHIb0VyY8rCy/VQQFCGj2FbwHo3meR
a0tfJPLV/0H+Q6C3MK0inmIJPPLijNmW5RaN7I31YjHerOYJRDAyZauk2klqhGwE4f4docr92m+6
wt/2yQ/AYyO1jxEOCYajFWm6FyJzhcefhDmgIffljpRom3KtdxFAIhB6Q4u/tToFoQFF0H3e3ImF
nnmRgn5x+ts+5v5luXiqby9fMawFMthPDxfnhSAF63bBdxFBBFcFhQwH/+Wst+EIxLCYuNxT/8ap
i4BQsFaqKv4GRaXwAqqnnBzkZLLuUfr0P7vT705geFJ7IYdrDA4yq8EGn3Yhc7zLcVgsBxqLkw4+
cux7d6eDIs8O82dG39gU3rnCVgOJSJ4VgeyqrVgL8mGLYWMeD71qeJXQDg76ZFHPoS5Qu7vMMjTJ
IkRclVEhd36nDMGgvvavPNFjnAGbsjbh96VA/F6UJ4Mdz1Uh0eEamZFNGpRsiTtPxBjcdbXJ68XV
Yu0Nn9sCQaiY/JvNH/MKeWTEDEIGXT3pwQkG/WIg4GLfhEOR5TpQHRa1Cp30Wywso3Vn4GlXWmQE
uCAHc23Ei+nAdRnVpC5gXh1OdvXmLIsYdMKctvCYybrebj7n00M5A/zLgnEPkywumFvXO28Nyq9V
IC1NX5Af0PFqS4yUysoSpl6MQjBTIDo/i99iuxhtPo5uz82/T2ptAOQsf5OOGICshToVN/J5y5gX
BAMWFFrCNehuFQzLLe51f7kUJEZmSm2HHTjOU0XBVqv+r7GvYLRTu8Q2iG7AC8+AjgxT92wwaDwd
CC6BU9LmDte1QbeVAoaxmVIJM2nvn5tYF7dzn/0MRbJXOxv+K6a4VJA1+3Y85Dvz5gMDlvW2J+XB
lX8pi9XKWihL13MBUWpdCg6N/vMD+oSkuON0pW0Fkdg+tfxi9YLpo1EuJJ51XhQEI65LPnHEaR9q
fOHJPbTRnoQ9vV38bC/asHPPV37qxZCKFS9g6i6AEmYGFXqjsXHBVROpCUuIO5Gzi4LLTkwyUG1G
gtgip5SfmUisTxvVlsXe1CRBwnnUVjviH6bVxhuxTtfwSXi7KGW4bnnWLC0ql5yAyoA145hsFeVC
+TdokRrr97Z/ouxPwdUBlZmr40TruuYyDYayQ8ST38DEE+rCeLM1bQapm2G/qUUxLhJUrWD2GLzC
qNmxgCCjyx8mDp1qEoQm8VrV1C/YJy5U4c5Og5twu9m3uR92T2RzkJi4D6xVHQ3JTpaR14Rm2ijk
Q2/bFSYsqItDAeVo+jacQ+7hrV5LB57iV2EJUeWEud3iKOP+Gj/IkXdIpCkfSfL8VSBPyrB1HAgn
J27QGxo+fc6YXy9goT8/QfkGamUQ/gdWdM9a2GP1kW9oKm/DE8MptgUgHcNrjl5SrpFvb1Cqv/WW
V+BiA3+s8xBC+BzxqM+8SuZfif460ubTN50yqFePRq9ghHtAALifGscfh2zRREePpnm7LGIWD+NO
LDbh6lbUfa7CPXf94e4VSQ3e5FqPsVC6XkNw/zzCArjwxIZoObJO6a/XqotLcpwVHrhhJJse8kYO
k+TYt08ZwamE6aoY7PmLaTf1swnh3P3aG8Dos+GAtI1rZh6iRHcPA3A3NVWz4eFF5fASzricq0CI
LPlW0m9n+1PhIAi5uHnqOvdyiTghlTCbtAm0zeQ5+DmJnHsmT+lNAmJgKSc93uTcisMmgrd3EFLV
+q+aItjRU+SXrRV8zVluuGvTriziQemPD4F3l0o5tHzt1vWtmz3SFSj4YY4aYf0kF0SrTvjhvmUK
SyIoztKzoKpgR6bioZq4aJYVUcF3HsHoIZ0/IvTGg8MQXAPSl8+Py8ATyVZmBTGThzxdFu8HWbjO
C+OogFBoA9Tl1ferYCr9nJKf7wjA3Yd+xr9MaKIuj6d6ZfnmnPP6HbcaQK5LN8ftAuGzglzWTOgL
oed0o9YVHxPnFw5DsTKNhiPTSsYkCzPCRAvQbYmQP295/MIiP9D1gzxjbsrYfDfhwjkPHujqQI7j
yYqYvxwUmHkeQPJRGRa2LNaxQVHrYcXEtzCvE+CEYmE+wLHbNZUlUyr3K3fMWDqQ1KhLqNyO0yao
5G0XyvHJG9gecaFb3HeRSP8IHvF8wcHjt7jG1BLbfE2xHf5shAni2sY7+g+4oJhdxRxz8cxzVZIG
egadtY0shhhHCoF7ZDgZqSQytr4bLDw4exzreJuyMw8vUk4MLC4HEX0qS79EIG3/rKmGYIDidBNv
7N+WI+c+AJ0z1zy4L6MqPQLOOinxNAv5BJwM3UaFe3az4HIOpgNKejS4iMeF+Q6ulYEtjOZ/VOub
1yYWlXzi4VNZY6CsG47HkZ4WSjkGV8PbBM8y0uYE4hRHrHFHLBmJdvFeO5psE2gu0D7Bu2yc6MyP
ZyqDF8/vW7aaBo9lsze4Rb7TGNCkvFzUwNJH4Sx4vIq97Cge6/ci1ZRvhwUZC8qkHTuVDeHxfqqd
gFbUOXmEJMhBnuJ9Nbnw5AaYVSSgdp42CeTfqI2OZhtC34FTms71dr7EVG3/M80I+rnKWG1jhxWx
9qD3+EpoPf3/EhRFNe+qQkGPCwOl7inz15uMsqV4p1kA2FIIX+OGcyPKJo/yWKG7YOaNA3TKesJ9
/T2lmmOnMMTpZNHRA6Iu1zowis/ZSj4nYgiE68u9wksElzgKCxB179W1AfYiA0/Tc5Mw91KM4z8k
oghblQZgbxeL8Nm3zPMVWHhBqVl6RWVBK4o1hmgbFaRkvG7Ng5c7L1LdsCTzCFM//My01rb8xPQS
4ciFQtUwtezQWUnVTIwjPHbB/kzKuO55JgpVTHHc6XF3NQRDCefO53jjG95ZCsnKzeArLBKkna1X
DpQ/iHH1647v4bjWvc55P9BRPkfwN2HTEuHM7hAC82S0QbFooXbrBazvAHEb2cOkuBuLG607CgUK
vMmjocy+sIrC8KeKFsxPa+5b1nU6IPBU/KVd4u7vgfo1ReoZtBVWJFF+2w7OQx9kwhBPb0rmtoDv
nwze+EG77AcjVVaShpyAPB1KNHr8+frLrgsvORAxconx80iE4qNZH4vjEHsk0XkkyoF3G+IRYKT7
KugwLlRdVPOuIg7/l98jJiXICRcHn8eOMkF4kJYDi2bx6WxIpOUHX20YTUkvgrw2Sd3PxsZtpNx2
co+XdDIhf8gj+LLYRgQXQV83i+7UU/c0zys4C+JFdax67HTcum2Sdvs/GlOBYvaMMd9KfFJEx6F6
UMfF738dcmpqGgdUzUe0VrD3vdUr4cNGtt7XhW/+kh/DppfRaSdvSAAgZqKkflafSN0AhaYYrjHd
Kl8ftcnquSfhO0hCx+sQPqAUie2WHXeT5arQsitjgrQNQnmOspfyxAV6Pce547tKiYmArGMu9XmC
YVvurNx5YyrnCGEFUYkJjRyIl1Ikunb5OmE0H+oxt45hEwCSXWJBNRfqAQM5GP428V6M8dkxGOTR
3o+h/OtZIo1SZrRSUlrbU6B8YMViCIZmpkpI94tY0GrweYv4vVv49KM7Ng+Z4THHEG3VAxk/cipl
dd1RZ9G6v3p38KFlf9+vJ0Eo851VJZBXHfb5pwpPrRUtxGzW9ki224suZxtkyI5fswGicER22+sc
rxDY6ERSxpfgi9Hhr8QgficT5PLbG9leBiDhpQ1v8OnQl6CAcPmB7JrKbXAwYUSeGeDN+sX6e1/W
Au1PJGan4q5cEF9t4aCvrII7QUqMRJO6QDjbF+WcdmQfSzgdQjNnrJWVAsUbHF3IHE4Cqd/U/Y05
IKCt7xN1mMOBcK/3PJhar46XQsNuMtK93OI74s+CPErM776PM7VIjwyp1ye+GdAJQGEPXsfXVOHC
R+efNaJjM7KZpWmXHVV4d2LKWH0Buq4pdUcUQpDPs9sF+Zq0Dp4A3ijLKN96iTBkg5RjR3YLf/lH
uHgB1H+q14hFtaVERmCAUcQYgoN1xmXqisvfRLSuEUa+dAkfdJn5lzUwBwvO+bVsXKBjJN64J5tS
sgz5zPnKFgwmccA/KbinAxJgs1aZQlmXhql+GLpdEi2iFTUccB9vq+dDibkbi4kfPjAsPKnB35Sy
V9kyQZbIpHgRMxsdvyerrzp/Z8p+oVUrr7DFCR/eSdF9xiGEx2MV5/+Yw59LyWhIGn8B3B6Hlmqc
aRODr6U8T7S5oc3TB/PaR/l7fp4mmhfJf64Mko/K3N4i03tSVyQnoqRaJxhk9y07WuOqrfq1BOAA
vD0kKFCJbgxBdHFBzE36PqHyzh0PgUrpxKqlQNVDialId9R911AlYCtUo/vCHhDVBxh5T/PL1MKN
Gv3p4rEA3e9dx2+AFsj5TuHs0WpobwfQwRGqfZINIUNsqMHb12Ew0+FPXv7nNcbbIjjtb12oYEun
+zPKR3jCxmuaSu9np8CIQBL58o+qiw83c4IMUZlYSYbNmm4nOaUnMFFwsaBJ6vg3Ib80YFG+MzS4
gzMXSaXSI4tZrT+SMiDwWmvj82AB+l1+mvzCw7wY5CbUCCvAAIReP1KRDAnln0lmSbHd5eqaJM7B
piOp6/Yd8wbA5LfkXfR7DbPmDAo8BBFG3UZY8j2AP+Ik/5WPViSYrRtOFnx51ovAjX6Ojf5Fv+Nz
pDlg/Tz4idgp9aV82ypD06DaBQN04FlYTRU+Lz++Yfp84ODavjC+vxg+pi2K+0veRVSXUh8DaYS+
uewgUvwmMy5LzygiLymtQYA9eG+yeHTfOBeb5ufSSKlDtW9Clth5hGX/eFPhFtptYNzFEc6i6XPr
x81WlAOazddi9v9K3zdsnI5mxOp+o7WPwYkutiQGszURozvxBVw3vS4kIB8pQJ9cM5UOZ1xIYn9c
aKWD5Aj5EnQr8jZh9llMDvOrz3N4oJ3h7A7X9IVJEacE5bllBCjhDbP/LfklxWUr+qK/NOexfzTD
nDSB0/S/hg6iC8bmWZBV8kZVjsny2x0Fs6T4PzTQX2NVat4s/qDxdVuZq2jqf+HAqjMNdYJpGQZl
mfLSI4aOyA0BeOFy9dWECBQIg9rQeLOkpV5rusfOCpjvY1Ij9MOHn6WUSKArKP5ETr1Pw/4gcIuU
UMWAlMXZxij5v8S8NBsWQ7cX2djDtnyFyMXoTwfFbfdpiirXeR+ShI5G9YMUafzMfXfVOS7nDjmv
2wvleVWNgOxEsFL4nVU2KXOiMZ0XWmfxDyJP0wtHSXQ/4OC9ZIkE4qDqNjkg6dFkP8/cCW9JYiGd
OrYIRLvgWMlNb/dx8jY/wiF5iwKKqhrRKvyT8Mn2NyI6nxOWB3mYuA11Wt8RDQ3ghLRQN4CF+xVY
94mX6JK87dsqV7njJTkLXStZLehsZ4pCoXuV4N6pEj9WLavVAYA5cdMLD7IapXynMdy7RwY3Fls3
b5ZDrRI2QV7oBfW7vvVMWzGKuYPxi9EulUf5QBGa9dP0snH/Kop9Tq4UZLfU91Zx3rr6y+sEkqJm
LfdbcdGm96Pq0HIPrmlBir1ZXc6JgHy9whvcOsSVfQXLzNFDjmQS1Gb/mJd3Yo26gFQ2JsxvwKmC
gzUxJdNDUnKWX8L1mZina/xyYniyNNq91UpDUCrwrec3TnJF2UkYtFpzdKE1GmRkkVj3Y9xF7HIT
kwxWy6eg1xukBQ+t1/ZmLQR+qVfIYM99w+bKxCE9JgRDLA2UECAxcnoSnIfexksP1ILCYUubqKOT
tlGCxImyl5ntd946LQdDLbelJCFnl7ltVkpdY+x1NGI3OyztCYWLMpzcYPG2lEE8rTGQ7BmnGVZY
vT4R4VmH9tSfGHwrsy4PJuOyqizRAhKSpriq/fZpp6jZ80Wy4z67c1m2LyL28B8O/UU1rtLEG1vY
EIvUndUrKjSpU1ch0gXr1VrwjmaM3s4QqZSGp8I0JSWNz8HNgVeql94zEk6ynmle9U/PRJ7+hm7V
ipL2AcHyRVgCiQcFL6UKzCeaNmMViU890jplZqt4jUJ7QAFcOWMgn+n4VgXOrdOpaW9ss3aTrESU
Hpyn3DXqrUO1j8kKZDtUvd9BJ+LuBOyoB28ABXQOFpzfa8ZD39bpNXS+4LS8CtUKVii81pUG5Grj
lbrzxC7a4cbB38gT0IRfqrW1OY1AlJ2FjiGMtQmwvWcj8HC9m/wGhjAfE5UDbh3y6Pp02wDJWvfz
JDsjokrOO1NueWkYDqqE1/un9X8XYc88QqAUKLxNnYIC5My8pPmKt2OmDNPO8Q9Cb5vrMd7gkzRZ
Vihu7UsRpg2JjMe021fNXO1E+WTd08GlvxIIf6+Hj1tlWViMi10vIN7fLzD86APvcOnhT3gXzAJC
kfHgrJuizqLh4moAdkRRuQSH46Wyc1hrOeb4Hp5244H0aMunu2MvIIJXO05iSv7dslPZBdz3/ZXO
wX/75MRuMJKHAA1su1PG4mAHxvgqmlmAQsct5Y+Ptncx5f42lqFaX2lEPPV2n3Jy3Ynz7yHBmIO1
JWNqldPo1Hr1YRVCJCVU0RcZ6OakyAWT6AspzTyd/bjGuTEcFKNgzIb+5ICt5YoPE2rm+0MYEQzV
vde+ouuJqYehhOlXB5GovCLzA8Ih7T7DuItefZOe/Bu2UaQExwW+NTjeqT7Ee8fdwB7Oo3UjXTG+
LvrYDcT+Xj6bV56iI8jQ+iexzmkZfDyuE69Mf4yPyowmfRoBxEc5XMQZIQQ+4uUsNR3NZVWsN4M6
SfjEuSzE2D8kmDCK+9GHU7cZtL+Wrz9ghFgBcohOwFRmfutVWsqdBVGBqK4/1dz8EhJrZbNhgh5K
lcwbqPof8fGcMhFaEslK93fKN8ttNYuDHQeUc3VsWnX85fAVCQJtHjx6Qe8LSJ3KVSKUcldTz3xm
3g4OH5tF+oSMTclOyURlC5JF0kU+2aSWIqwCxK7Z2Y4YNlAU/J5JxtRz0/UUDG0Tu4IE1LNjW+/C
RZ3bjKlBl6zZGxKQW5dTBk4dlcWOREzL6tTIy/2AUBJ+dqwuMWPLogagP1Tz1EqV8IvOvAaVcWQP
T5JgdsM8t34g0J79JeAVqy27OXVDJygBk5huSYoaHOAPyKhpTGxM/OLXeUwpTmN4phxQ7ZuKRwFy
dEvmSpJczrrDcEa627JfopZoH+3AWvMCBhxJuWWXCQGx60UTn5ko/Tmgc4FCLBCOLdYgtOoD6Diy
3toB7/xCZFcOT11i1Y/Pea1symOpdOqPCEbt1kTml8yn43KqEGvDLoeG8avT1GnnyI9zlkuk8uQH
v3+SxQp6CVvFaeiEh5+YHUhFKlXBSYSN8phXvudktVQTclj1SSI+l7rwpuqclVmXHx4EOu3sCnK4
/d4nBLt/gktFD+3vmZXg9g6QZRWyPf+e84GP+JVnKa0L9N5hQkr2aLqPKc3ySZrlKNtDfn5dIIUk
o9UBhchhuTSMGcABK8A9VzRGaJSwbdvkn8DwHnl3rDaHhEo/brNpfJnehu1lYU672GjnyxI9VC6r
2KlZRyoODGfFO3O7SlaelENoJ9pU6pY399wCbO8BGB5fyqwTwvcuQyg/MpOe6R8k03jl2R8bzv1T
CIOyxWBW5yy2VVM97X1PCQ7koCse+lag1XJAITpRkjCMpuAaKhD4vXdTyGbQXFrI6CNkiLAUrxLd
SnKLPIoqwpRrVo5rpeiZ6zMwfiBJqz5beWbWu0JJiaMlMmjW64C0doznanth0TNlK13nRllXmnBf
0gwS/5mvtuf15pN8tpgbG0cN2+mYV1BA0mFDroAf5Styx66fQJygRLoeWvVg68qKYNfTyj0ZZ3Xx
DWQKhXJWz7nWI/T5RjwV9jVtkCsPw+KVEw4IbYRUGo+CXb6fRGHZH9rExKnRdbzTvhrWpPfLbDQh
+4glt8RVDp5VCjAw0fVTAJJyVvzUmPX4N+G9wS6Am93p4SWx/VoBxGisbfgzFi9Ld/7IwVFyM+Qu
wkD6qMzmS8JIlKqmsTyq8tY6jAmBYuikxzDuCRvR68bsJhTSGG3JntMQRly7DMBaeSo4d5s810Xr
FaHmLRsLIVwxuyems3SoAsCTV3anLc+A+aOGFIFEi+PDiBEx0HX+I+s+A1RzdcYgeO9XDxC7/BRr
kb7OeeamYtmnIKR4/kF4hfxaPyYTaPoNZGKQwkjDH7tniahjDefC/v8SNpb4vsjqZp8M7UccpA3Y
oCod6L0JjtzHCn95PfRCmO7VNdArJF01EUqtBsr/fYAQW74S9oN41SeN/RSxa5/8FhoBQv9jaYyJ
ZduhJEr0e8NcUOLPsOzz/mARDcxkZCzjjnTpOB2bSgKKS+Qkaf4tlvcrpjFG7rKjIusEIsyMtJNv
vaajwuFWHpZHS/ZB/GnbFuR4TLt2sCd2D/Dn6vmpzyv8R2JoTipe0Y0/+6fIqVhQnYhR9osvdTm9
ZEbyj2n88daW56s9CsqRWnoLhRo5KpV5UWz83M82D1yFnPemmzhO2fEt0USSLDrZdiIyPp4zIA90
qZgiDUrslNSBV49oY0j/SfxsYqr3HVKyuGkOqSkYErWNEc58kKOd+zBq/Ck+aZD43JfgM4B3LOO9
zz7bxRytuGFO9Heuoh6PFnh4H5l91eHPgwgfy+jTT6B9HNIBDdJ8i2BuBknLOWORhDQS3bK58Jby
ivFgkQM0uGDvtDvNHJ8UCIn3SpKaoI3SNwNh7/gDSus0AUQ7QzOuyiVyV7Gr5M92LI+lcGn9TGWb
i2vj5kVDwYqffVkVqbpNv3RYemZE46MTd/MEGmm+5Q2lCATnX5el7LQTbJJcvTH62PC7mMSwGUJi
Lyhd+t9NNdf/PWBzRUTZTU2aC6S0D0r00/p2yUa2ltpk7Td0rNWkVirIZKH6YGcHRgb+q2cfYfQB
hufDuXau/3YoLVh0u7dALcw+NpT+acE6XHv0p2Ti5zNLofCvSMJTjI234QJtE1YZ1KsvZXXEp7wU
sEUGTTZHlKWgJuSAxjh8wDU+3ZcL8lh7zqFqz8XQaLTXMKbzLZj4UjCskdh5XRHUgzDl2sBVoi8r
N70X+c4rEG2RrNe3/xT1cGeZPXM7n44XhFGCd91x8oM6UlIRvl+rETNKvHasRexT7WQq5FdrjZuk
lUPxdrHOWqO+cs6i1gb77rcoja4OHgbunr1P7KQV1vVTOtejOa4Jw0cdZL+4gLvB3elNLkdE3iku
b2a6ycnji3vwJRi5gSXlsSrdxSXtdB0m5lcmVnk8GLFV18nkRFxv7fCTEZzyyIZB1HLLH79Kx9KE
YQEBRKDUZYp5ygNoEGi5qhRhAsRKVcGH9M1NXpEVFMqHkyvijtBqZLBy2lS2SzKvvZGy1IdrFVVq
177T8cpxinmexvsO6UQqfl75zMlc8Kv6YmGX6CISlD4vLlQuezXjwz6fH4nlkK9ZrA3JRzSUaeLX
DFFLgu/U0YdesN/iapbqecIcwOyVl9wk5zD7dmxi8hyZLnZI/90i3FXTWHbTy8YRs5tZ688WQYdT
s1zKFPKLw7+lqUm4GDbwqaO+r3kK1Kxw/6gqO9FHw8c6dpY1vagsxLuXaSBI+kHmN7QCRKsMijAW
ZIRXM1xMrM8hXNVRYuYxWto04N+h8U1TYlnFaZ37geCOmZxd3JTkQ5Yt2LnWvTi5rUXksewzbOrv
xZyY9alTgWVCQ4g/qYGnjIpvofWXcY1ZYXgYGbVd3cMBCaHTS9dlsYxhT5/sOlzkgoffolM6u8DG
dpwSfXOSDx5IJ8gKZpXuhXmfqsHdVxMj1fxaWYbLEPqcDp5+Ta2qoMNzV8EAnh22d6axY3b4ymcC
gDbeR7WUqKPoauxqx0r4gGIcunl2txfFBQNmOv9gn4J5EitVN3dLcz2BYDrmdhUbu/9SgDJIHrKt
+MV8bqSzdoqP/oUSjVmInvabU98FC3InFBK2DSLBh/+wpFRaNOACnFkcj+AtSE+OFloqZ9m9nTTh
cmsNOMk5EJli/uP4xaS5WF5jILa92pz71ud4Op7VS8zQFVuf4XGFNzTIBBjTbGY9S+VN4+K2wxYI
nFxJdJSfeNH+QkdxFKOcTWX/BzfGI3QxHYub+KvpC2QvavaoU1lPCd3Ywgct64haEH8x6xsKC36V
bHyfQxYVnlR5Bs1sXY9JzL14VIf8N34avxcZWo8R+qE9vaH9q1EZCVjN15k/0hi25b7mlqOrLBuT
4WDjLSUqnsT1Ax30j+6MtjTIHuWbZ6eaCQ47uGLKuSxR3t93RMfhHIMDpUGOQsYbq1OLXC9w4SIB
2XtTez+u20PzbDwaooQAaogfZASUelq3Mym23kjpisTgwhc0QmhTh7ukBwMCxfUNk2A0c+0cpq3L
dMRHuLyD+5OZfn3J6/Q1b4rwB+pzLlJqwG97Q9Jxw2ZrcqvGF+y2SoUxVdHeZNjYjlf2Kyv9+tdq
LCYrC+kXtO3cj6oPrSFTaz5nKGUwqviEUyhA3Z5zuHlBq8HJ8/gOd9gRSfEamHTN2iexUeUInojK
/Vr0pngFTtYeYb7fMzzmbrbllgAarCPLNl3euSj2AMXezHnURe0IQcjTvvE85AWw/jCnoUNcaIRk
5fmx+j67gEri+dnsrw+Cbrwc4ZHova4x9buX1kNGlm5kufUhARLufP0c6SdJL+sQi/cvBTJpWCZy
SndQadWAJqUwm7EMZf5dwohdtUHeud0ha+m+BNwsM9OIiWTE+/NQhbfOHAN5uSngzLbDqTwJ+aEf
XeV1MQjhJUYvH55QYzyBlRJb3cOCNf1OGIAS1Ie0eYesH4ZVFvkR7U/6qJTrb0ywZ6YPxmrAmnoP
fRiQwTBNjpzt9r59iKNPs8nY18hhfVXVtzZkk3uMw6Ow3RgZ/UJFVFAwJi2ehwrcPq5qCrywNLYc
59c6odWZcug9386z8e04c1JIIOhsHUZdTIOcmkuACW22f1otC9XhGUGC1rgxbd33mJh8ggQZcJT5
O+BZKlX1vUitlUDx84EJQrH3ADLO296v4l4slQtaLqDrPPn9LyB2Bso8+VohoVrdueqNOn1r6eoE
P4k2CnynyatfNfX9DFIs9wzjkmYq+eXYyr2ve5vxv34qx1q/G9VKAcpuOgmHE+1Y13BWncSnQj9E
zvaxSi3tQYVNt5j8fHawCovxJUhc4nP07/xIL1dobFdjHhnwx0IFlQJh2weebKMNW9JZ8wVyWsNF
UXpMLgJbUOVzM9ECk5CzfmXWPEh2hybtkIsx8X0QgSiGmYxbH4w136SooDgyQdXPFPW66EiMqqr7
k244K0fkqolpTLJ0zB6BR/7BcXgfLyYex3SPttR0PGFSKT+HOnXjAce7IGgqWDW2J0kk61HzZgI1
bTIHoXn/rveffznExrGD26bOycn2P/k3TxbZP9w/v+h90PpGKyfaBTclKu10mAa3jesQnGqUoCMh
/lrVDqyVre4lkybeXEP3KBqXqPV/Q/OE1nCAlUwfNxmDisgIKG5c6p/LIv5dEoFE9HUY12hLllHy
gaDQa3QQsNKAgA3m8oqq+b+VwwadDteb0DeSAOIRSCRXvMDEHcXL23RgS/FLCDC6Aw6+RGsr+y/T
CBgQsezzemKZgPyMyDWmyyuVHiyMO7m1C0YpQ0BGB0C4/aZJDelfL2dxdgBjhdnoX8u+UB5bSTsQ
ytOGQb08g2HkdRgXGVehD+rQh0nvuUiZO3S2CRMZtDf247xdGMKNgPbEnkaWNF3DJIM/kpipDGEr
8uhd2qMqmK+RgQHNSMkbK77c4zVqCsxwnhREEoSZrAt6bmxyu3nCYfBkjwKaZaBpUMmc5XoKnus5
0q8fB7XT3un+Vjq4MOuvU+spE7HIW7r3+Yk/q7sCckgMQdggmiuL54r0/VEZJVNMv6CdhotIF3hU
niYFDetSEXQTf1YhhUBf73sRqCaijaCz4qjUaUEt4unSzetwdYOSkVL5cLNbz94p/NSAEoKdiTwn
Suu7KkMPohNO+BMWDEcaHHrNbOdTOd+a6h8XWER30y71m5fDVoUo9TCnkI+wNHPBdnYXiCxwaaC7
iNg2VI5EjCInNY5RjMUH+UgggPZYOcYl8RrMDSG/Fljq5MhxeE5sGlA1GfX/NDvD3sNmFicKpZ6g
aBqpnQqbi2+geL1YFwyMjEEeuYQnEHmA/nqobK85aXLe19LVEYnM+KfTc7IMWNzBXhltQ8rlDsxZ
+6m89y+A88zhVhHk49l+h6vUk7SweEkajCL8tE94E21T8Z/NvbwP+esS4j/Gu8MKr08NWov+cCUS
0lfmr5JKXPuvyXrECwU79EOQQRNFyXQth16UgqwOUAC1vhCi1blBS/MtPfSG3NayfDmxq6KKnCiB
lN6c5TcCkE1XtRNLlPXgTTieE1FpnEdMle2JOQkPeqiwyn1CPXVpjdKmS3vCFJ6H+bGSsqG1zmhN
V/l4R9b/x2073bVKw9BclLkPVtBzpyQYZZGA+zE+UvWcE1dbV72MotG4lZKGikpBpoN9gN4nq2ri
ChQU2kw0tz2Iv9hn8SdWhSXhndDYj4b2V1X9c7wH0UKlW048hlsG0yhyL55HrR0ucimnzdlxNTwQ
D6LJwz+kWBeKUTTfHIFbHIF28lvVVa1lo6zrcM9SKtWeG4K/E8oGz52q9cTm0ivzhzSnrlJ/Hx0Z
fXLCH5rIldv3EN+X4JB7iW6Nb4rxKcOi2Y79l2UbUYG3zX5xzsCB6JoY8+0dJ0oJpTTKBveSlvAv
5UufNwsyzbqQhMcMdNEFlhA1lcscwPDURIHcBqpjU4J2DU6nrq02PfrHQwrB31nCh0IcdUzn3TjZ
Ca/tyriiIJRgJgI1wNi+hsPc/L7SCakr127f4koLdSf1lY/S1NKQOLe5t/lt0MmPmXHBz3rSwDss
odt+T0MX9IW6uoiJWKJLpR7IKECitFFXc0WFnkg6BZmwtTGUzVRH0qTnSIVhg9erw1bgW1rvgAw2
vucz6NjMaVU4D0WMaJyaywBJ3I7b/0qy1c45SqklVeOQ9KfBbZeCNjOu42OUAxAiYrWoeX542K0s
UhnXpYHnmnAlUUiPPNauuJ0jCKRLso0RQY7/AKb/kml1dEK541XLQEWvfFV9tHFGriTcQyUE3Q7X
NUF9fnTj++DtL8YKlsQS7lhW66LvRlbDl0eyB+YdO6CSoqUECjgC+EbVkdzpKzgAMFvvdgIydyq3
3rtGtX2CEBatpQ6fm/VpuiVsudrfbQdjoP9ODlHU+mnnpFl6TxMcHvD5011kL4WBtj4Nm7JOCKPD
i3ywqV2mjHha3wyH0naPOieG+X9C5GkPx4qQAw9NbI8o3z/7gDzSe7gHfusRGxyK7lUEz0RgCGJh
SiSoW7/K2t518u2AuapV3rU4hBKPQe+6hvdunmTRGdRCXknQ4vEUeP3Qs3YxOO5Pcpkahe2tf2H0
cKJsStnaGbO1jm6MDhF/37K8oBUIDaT6543xBgBJk04pJwo9k6POkPvXEouBI+XW+AKXB2/0sz6z
9PuG3m3PsqfAhXSHeLXKFgHwJp1pd6ChteoLN0Zsil43pbiMett2vCEFFQJAKazJLl/Ulh3avsbL
mjrUtKSE8vSU0oakYp7nKusi1fsP8lxsAoVIamscO/z6XtpZK3hgWHpUMNx9Rz5jSw4ntzdg26br
kPLjNSww2X08skl41aypBWk4ZoJ/vbTcVgfeGibnL7d452qEmIa7vwwLtJqlWaqdr0bgZMzXq9tk
0rSEz6GJqgpQ2/ZTIrcu/0VszcxGfH9coDpbY+hpjehEa6n5I9qG/YvartqhA9XCpu37MilZ48qK
vNr48RJACLnf1QmoNYDpC6PsGRxo71y62Jah+hJHrqEwEXUD1GhKvpiHXT93CSxolkl5KkSXUT+z
v0TxvOmY9R7SiGhzHjE6ItVhXjLmY0++NLtl0jVnZYfLCm8EQYG/J5mM26O6VYeIQJ2iKvq8sq0x
slwvHH5YiErxYUsCeKhAaJ+khgmcCCeUgQryK6lAzk6hXJeKAZGJd4tvTUHBq39IOmv7CIwlWmWB
xgzVflFqGES2oKOVE4t/xnrwisfgXuXySx547MyaF2g0lfu8VmSiYXKfkxzo1P66gBPWa8FzEXuc
D7Aw3DSS4FpfbD3AUKato7DJSifJZQ9nyZytNbcv3QK5OYA5yKdx/HLum/sKbXwP0dNRuylCqAVf
gNl7egOlB9uBxSalJq1J0E/BI8fDrKk/8y3F6yUTvBcwBy2MY3vjdNXcrz3fOUzAPjDv1N2MaKEx
E6UmBSvIC2oWVb+qu9orZcKHD38mmnR5cHnefJT6rmK5RUgAxMLxFPHX63iikyntWI2S1I2NgnMr
iBrqgv2NpIooBtiicSkvrr+kMJCtrSOfvV3yJr+WjJv9CEo6grOX6wPH9RLHtphNWYkoLqJeKjTm
1DLhE+90Kx0kfJ8mcUqkjguTDK6z4XlL2uiXzH3Z20dvGgJej4pGa9UBIxUhfYDrQtm2Vymphgwt
nGrbS1zQ2keYBhxaLC7DF3CfM8p+lFZHfGX5WH5xA7eCKa8rMQbwTn1+jydfOnWQausPnOwek4YC
1fxyPItoh+wRbuVzLsNvAC33ZQo0Iq5sXHH0NHuKILYcRDoj//KmHagSI6dBOuwPlxA4MaexZJdf
Onbtq9CE6iLCwhwsUf0y0CDxAQifpp4JQwtoQstTzaSmjvl4rMGeO2wDyeXbal5B/HwV0G3yizdF
miPFgYY3/4B9fOjonPat/MPXeHkx7FRdR4hs7BIsMx0ZQ+wNk8Bjj2j/T7eiia2E94OoGb4HulLO
zcYaJBBnllgJXkPNJTz2AriWOzl6KlPFXgOwhMD2NSc1M7Z37Dkzo/kGWJm/vBhP30GEEcRsvXMH
7E361KaTTZCxnrvBtrTp8Oo5F0MD7htLzwYs0/jG83gKkcJDq9eJ9r2BYfNqHxAoZXu/+FvpmWTW
cQk1ManLZfjRAfMvsgaijVtAU3RgTWpXfAfNAOEhsMjylCwcikQ76HY0EBG4YuxBftPBleuoDc3A
xd3yraOO/xBLlMOpRqbn5YGUT0ybzR1MRk0bMptuo+x7i9D/dJH58v1rQCnXJbTCSJHu3L08hIyq
yu2rmAhfCMJ94hFXnzAmtrxvujW+IsVxhFObd7HjVMKGGGKSN8N0wm8sRKaxFJf1AzBiUAkOGSO+
bwcNvLoDhalbTd2/VvXYqBxWF8OcD8E94neFa8MdAQnh52mdU+Ceq8VvdxkLohsg+hSsafoAwjCk
cYdYv6b7ltIJABySS/RB6CvsMVihzgcbcMWHkE+4FqUjc6uyIKuMrltcY0ZIK4A2igq74rKPa5z3
uHSBhQybOQ4EO7cjnh40mUUewo1X2iAjgpA6ceKSH7ua0CRbAB1W7iHMTu/QY4TTvMdbuop7Mt/P
0mU1D2K2735HqQNXYxzGVa6LAMQR5N6PCxhFGFapmBgC1J/t03BLgAa4VK8uLv0zMTyeVssV5pNf
bkzKJ8siVOTvWoNd2mpQFVdMdbZU+SWKadzdTA/5bp7QSgebTDc0LMsD0bfynvEkvwrpaUp1+rc6
xrwG+7gP8zhRJEmz45K/y+O9fH2PbISJRovVcvIXz1WrcPIPBSHJXwHgK0ioQePjheQ5pkE+/TdJ
YJSDsugpsbQsnHg4KS6/ONeLuNb1jplm7rPyeGpO+DQQM11K6NgH34ldvur+WHSPDTvd58KYvByW
E09oF27i9yOHUdCqi0vZ3fBalrV1IBMujFpaXNssBatFjOeyHdzBJJpyOH9at3HOdWXUxJoi+CYT
SB4OA1p8qyNW80tL7TdNy5s8do64+78zARLooo8FypDKQVkZLZCIbLH48VnjbvUADKrjyqgMS5vC
XYrrqBOsd00jsKQfKM9MpaR19K+8SZF4TgocUkmaxNx+7NErpv8zqL4FfyarouvIP4I+6WwvINJS
P9KJ6sZu7yBgCqvDliVBRQAv36QZHSoI1GgEvNGnZ6Lbf78uBdUAAzpe0vp4GyoWw8epkyZuGGk3
L0aJEOlVIOS0F/5cOmv5JZl8j2fy7HmqUHDX/PV3hsnfHDL/XCAB5yCGJe+HAG0j9lg8Z/yI2kJc
FAOxyYem0PK5rQtdMrr3TBDGdoSx3L22GnIkUq5Q7zJzbe/LI4NlBEI7JHNAd1fAiyibnABJZeKX
vnx+DjzjJolPlU4oH+g3kD2tRikLXC9jGFev5kzk637jq++hoLjjqPnFsOrC6LncpYrVdOu9MKOZ
V/13o4y4Y8Wk4NEra5HhLqbEYehRyxkhALDEQh/MS+PzP3KSY3dH1FIXZEcMQ9wKoJMnjjGHzEvR
+7NRG6pAL7NlanC9O3hdfDlPLaK/EHyuBO8oPGEvAMgiCeepUF9gqDo0h1AifuqJ7C+eLUaSNyfW
U+M3Mq07fu7DDXfEwHy53BcIPgWS8bRE2YKW5ngi1jQ9qqoydk6xKTFMfKSnpz3uIKWijz8C66lC
nn72SlybyM0inrZsSL9I+9Z2t5zaOeGrhtM+yTYFII5dQBfOU2lBGlSuKpAO7SisXJaRB8mJdebc
G29mmhI/1JGv7xqiTPrA9UXHSWAayOsMRPvsLkSIcOO8EvOoxfkl3MC5bPMGYSxbCga88r0Oljzj
sa8PVREL4nBITwHuR+AV+H7Dhc/otb+9lsJ7s+Bcta630VCqsXVRdc3LjFb3jBAwUN6Z6hkIWkkr
WNdtDcxxEUtRjpD+Tf6yILhQr0+uhODNCWEC4fR7zGwIXqFBYeCePvvYHcreoZalgInA6Tb6Yyih
cJbGAl5JKIvgDENnBx1Dw5X2P+Hm0HXkNazdrCyp0qwepypr4XUzmdX4QomWgrYk5Qvuhka0JPVD
vi2Q98YBSbj+snHil7zz/wOCOH+g66v8IK8wt64ip5u/EOjDCCoQ/xfJCY6LdUnO6BtYlDr9esB9
cRN4pRFJv4z3xUFFiEi8J7qZNe3gvrBjttDMrUMIsXpgRaz3X0tjjnlyFH4UDq09Bk3PMHoo1Kff
3jLJ9CH6zWqrd3YtFHLenxRsLKTiXppqkzZTHDv6T6mCRSOl3wQYSqEQ9uXZsn3Dk5ayFu4nmIpr
i7ShxH0v1pM+rSQFzfkYyQMl/PmZqkR1knG3mqHS7/y0mYwU5fgI8Hwxf4XJMy5DTB2Rq/nvgr36
V+nDECb+uNdvyohBYPkk74a0g6I8fEHKjYPtzK619EAD7n5lZqHXjOnCjE6VprdE6fYzGg8xOLis
lT3IF8iHyrZyJa6nP7tRYBj0WJ1oJRONX6zB6hYmMbOTzUQaX2iyTVCoCoGD9RV2U04cZmkzu4KF
/Bi3m+BjdgULBQ4kcsEgNlHnl6nNxrmEDxespvReu3/68vbCRCoQeb0KtglTDOFqNXeG12WOAYnH
dfnvnGSqBmgOP8jtDWMtZHAAm/UxCeOZP6ZQ7GFlIGZ77LHxrcCZweM8ryA3UxJfVG+erqBdy5Q+
zD7uyn1tKdRs9E4xOR4NYvjy6sWtYVK9ECMftwSQ4FgBLtMRKTd9r5OcVvxiXwzxJES2fpWWgwyP
pl2ZAXsYL2kU2SSaaFN/XGuaIbkdgqGVpEH5HZM5yUyMFh9YNi6Ew0P/vio10keuGhAo/96fExIV
akKkovclbsi4MYyHdyHu7fpf9jQOJBs09vNjlMLv5mZjX/vpDW1l/hlVujdFCl10XxllOuZvnAHE
U6VDikq4wFKPKXdNYpZy1lxcj7mrk8zH1LE1fxykWAk8Zw20tq9ulJsXV4heeVjGmHXfDkCTvsOZ
EOZ6xdWTZ1UtdkUHnyzf0nrxrBqo6bfFurcAkuNM0BSGZU8tOa2ECd0OSxj7sMaF1e1MhKdVYv5K
mVimdu3nq4YhdxLT3oqHOcZDhxl2f/gRPyYdoAfXVEooLZPzPqUZMzoR7Y3/H9c1q3Cmx/quE3KV
Sh84bReXbg2mrgRRD3OxVeDWtLZIxggNRihu36DSTa0hFLIL9ov6caUzmTUTKPABKm2iG3lhux0o
ugB+ls1m8Ak5YVMjK2yVSvTx/wD/8SPqyOZaFtUPvfcajdCb5jC6W6PnvgLlJOXAl6VvlJT463Vm
Gs0s0fXsF/vVmWDor/B6BWmxnry8r0A5CT8SXYETl70ZTw5iTygI/IYZ9Taep1UiTdYC6TxMe4TQ
cCJLfVpCe4LZQ4UsSkKh18Lnrp4CkRghS4OZd7BpydEUvJv9ppdibQi0ib75JX9Mat1p72hU3m5k
koWhRsVcwaB9dYLXpSWvf4oJawTb3AYqwHsOR/cn18A5XLENgCtx8CaFIjyuXwrAH3Z6X1Ysn6Uk
jOg8vAbTAfUxheFdX2uPk3XipavsM85tbFmZKXK6uJNbdsrb4o7U+9ONHjeOWmWJ/QpBOMjJ1zPz
SrLHrHmGnqp/1Getw/w9OTHsVHTtOp8OUsjl7woY5OMEicEF1qKHma/x9zN2dP+ehRQ5iGH9rgmb
Q9pbMJOijg2aCnzjjf73iSXGQzT7PDr8ORMdqxXFDCa/8JwqMRcYaw9GiEYOOHY0K+lrajMELq9S
+tLnBbNpORfbwX4PAKagU/zyP3ygoK6XFfH8gNBSzYA5ccBRegvxRm1pDbLORGHy5sXFmDP7bS4p
3WHoktwVFssRYJbNl+IbwOXHGAoJ2F9auXXcu7sY0lFwbZ88246d6x88Jh2RUSWxxiEOpIT/xNyX
AIH9/+IzxkfG5YFU7qM/1x/XaFVvpLD7JwowBtcva9+7ps+wt2V5+fTfeNJOfLxn6yFwuK33eGMI
Zfi+NoYpFRDv4NLtmt5dGDl+QC2FWuHzfOtVFst0I5Yxrnx5NsOjtXHnTlh3wqPzcKEMR3mQ64EF
n5Af+mavopmcfoS4MpqfkRER1jBHVf0vXZoryvFW2jfvG+Ilqq3pZrty7Wb7Xz+CCXBmKPFC/xRr
IGx2rujYZZAf4joFarBSpaEbxbzqWciWSflyv4hzQXsRzHx/+gzEaqm3ccRMrjClmKQTj9c4K7PV
R81UDeOVdqoc4RvMDzQq4r4K6Azdt8BuhNbrqFWfM1+kCRjeFmA3cl3W1oKF0+KO2qpeY3Twk7F1
MwDSxog6j3PV70/kJcibkf5fdyzuiAjOFECCoyKG8QxtuJEJNkCWZs235HXy9LiakCZawxsQvmlK
mb1aw2xJnHfvGMF599v+4DykjGoVq0Dx1632VvIc6+5a8DWCO0+SeR7AcvmKspGCWUMCUtTvi7Vh
RvtiHmOW2WmGTLVAEJOCTEn9ghWqhbDGSMY+a8NF1j2UqFPH16lwKWw2vp5dkZZQPH75SkzOeYtm
qr632CGK/3Q8nG9nVD7+w5uT/oEPE0vuUqmxjuXYb7VTG9Mjw5GYksFvdxkxFtHHRlPYxT6vlz/J
WOsEEssfq7nozrEtKWoqM7EJdQ0n9z54eg9kc3RTmJgigdWiqoQspPQv60B9O2kp39UAFdPi22Bp
HjygryPb3HRsockCSywhLlDCibUzG422osp3+AGCdWCxrrZ0trNsvTAE6rbKoPljQ464xIzKYR7F
B/TYai2IE169owH5TTGqRva8FSbOzXRpeDNbtG2gYEnFHqQv8TMKzMjl2iR5+pmteacx1nowjIF2
55TotcvQOi3R0ahV5Cmta+tPk6wf8K2S9JJcDn55/oyvKxjbwNBRLg+hB6mIdMdF8mhz4V9ktu4Q
JEP4YvMzKU3uef1GqeQjYzSjEJzFvvKIb7JUjaebmG4QPAObvkoL5mf6VtN1qpW/5c/rXs6XFy7K
IwvyVKG40ZWW/iojmeyM1IJ9Dj0wMjbYt3OH/aa5s4e/WDqb4K8IAOzK9KupvmbJVos1GwVl/gsd
ryvIrU1HAlzWzI37kgs0bH9rmRrcb0AIqCiR1EnVe/gVwaR52AgVXkaYWeuAMIN78tcKwaI+VhYe
TowZYMB3gFkb/+Ja0BcUt7mT1eBGrjMtXe0Wa80JT8Q5sD0u8KhQ/bZ09GKse+m5JLws4i6zte71
glkqHjSJAOzIH5f7GFILSYKkDmxpXSRpGJOV3LHgWngQ90WIdK193RZjia/NxnbttC5/7Id65Nnh
FPqX7AjZzJrZpeC04bLUfDQG9OXEN8N+Mfxws9WHU2jeAInDL3Wr25D3xRodsgbq+7ishLb/4RBG
jgmOLcEd/RzpBYAVz025iSxsXnBWP47alSdiTbOQEGzkZnonpZQ7L2sytU2Eu9ESVt3XZG4Z+/nR
0hFDlY70FsXr1/PQnXZyT2PmoNqhca222sDyMS9OOXikC1WJjEKO8ByEUZh3oA8Iszf0W3vO9466
Y0ZDOtgbxsYvQkyUeCdtxqR3R0GLLBqMM+WkcmcCjnorWNR8qcmTJpfHHu92e86Koxoto56kc1IE
X+F4JfRFEKsqxTf5zOzB0mr9jhDQY6hMABCsFtTPX71V7Kt7oKmKYVQWsvVip+SbF192S9s8xrx5
IvgLG2WDYcz/r8RQp6nQ25a5UAg6/bvECBmg2aCP1BOHCreewBdb/MAm8RU0EmQA7Ws97A6rkckP
n07/nNNewpyyTLiMQELnIksmc2E0ZmrgPs+/kUictZu4btl1QIE+HS8dPfyv7L5Y5LSdIm6RrIDV
/we0H5phXnakOfmOtbIczaomWE7PVYOP3F5G5nKNBL2Uw29fQP00bH6+A3H41itEAkKZfW9T9a7C
55lEVfeSn+HPyj3mKcsNfpWeAYO2mx+Wznp3q2EVX/k83bnhGixuYAU84bgKduFzG11yNdx5uH+N
b0ox6hiwX/ciqnMJWNAciWtkg9AtQ2FVMJ+mcuPyb5qb6g+6KlI1//DLQUGg4Do66dQcnJ+L6ps0
IerGJzb4if3fj9h4IFYjS9ZvXczQfYU5u9z1wWEEnSU6AJLkiJDL1KuIjD8TyahuIuPrTjHtYgpT
HaFlyDosEvFX/Z1Bk+LzbjGzYiVub/sSRCguhHUUv8lLjD9nfmJgVfCvUPURYoFuTucitFCoNbSP
TiW6EDrrKzFed5JDZBINi/lSB34HyzSrg9I+gGa+DLH1ggGHrCLgUx6b1AKV+FzDxrhqBU5ECY1D
/6FAuuDIUIVZFI/ubAEdJrWnM6AECoSxXU5cRUhKzpgAsxAtB/9y6bgE5Av0IWTj11DPHmUfXZoh
FNc0/Ubjz4ORtwsCkTUq5zzuL3ErnUwexh1YMZiv/shgmEEKpecMGrboQxbqmz2gr8oGALt6jzYR
i+p+mtuVb5CDLlTpPt8D77k2uEbzNQxvHzNGKSpXvIeoaHd3M+DZjWiJTFpFjm0zoyYs6Au8wRee
FwJhCH/qh8itw6tDWo9e3Nwmrbh+K1KHivodwo88pp1XQAGI7GvzmA7HUdcTP3q38+gU00a2EtkG
RcKde1OLARc1NgEfhWcbnmoacJHxi0N/FUHCRltOz2OWGXltKwiJX6eHtc4wpswYmeVYuVnPcMVG
IGS/jYWvJUitY1IB0zb/p3XpzvSAnMh88etE7MHcvtt2Gwyik50vsyEGc/nmKdknqmhfuf/Q4q6h
vBZ2wiIi/nvM9KybKPSH85qHtx8mJUVvI8J5U2h1yvkQuP9hoyH7oGSDkHYuJt6DIMqqS0BLMkZ9
6CTfi/OoJID9jISh9ZvEFQYMTiwOQSIHe7UqeRIWFU/8JIIg4Eq1l8JbeEnpKBoapaF0TAknNF13
OVabW5zApgtpUXdUWvliWjz7gFPOBZ8xrFpa18NBh6Tsov4PJAo9WBw1LqZdKt2MpHFuG313AmgW
pGaETDZt5WpQ8+lDiZeKsWiN6HeD9HBLVJWOhrFfwqqVZM6S2bISO4pB9W5NbZoTWyk8I0X91WXY
C7C+ZjSmfKuzMcfU/zys0tGv9aRpHUI0ykyP31KASeAqDEHaZwLFE/QFL2kHzEZRwBltX/LN/DzE
xVDTp+DomvrnIKzGBTa+QyG+G4ICSe9zaG0Ci8wYH/BJK37WGZnsDHmXRQzpuVwO72Z60pmz8lRq
xkhAyCFPRz28Vo2u2Aj57nBZRtT88WYPexwMip8FAqLG45mnl1Ec+ITrNLPJ5LLQU/QUn5K4hqxS
gjpizTlGCxa9tIF7N05CPyxFn5IxBcFM1O73KpLbguiNGX8evx8SX8Fc8QDFh2nTFEKSCZiBzvpJ
ZwUTmsaclp337cnVPRxGEQk4TWzF8yvP223y9wN+M3LyLMz8qAx/7GnJLq03kTkMYkadKbL7BL8Q
qvG15WVE42z+T5tHL8tP2tVkywHSTdBQ6J7TQYjoa4OICo5LVtmw4F6rltSQS5JqL1SiFe98uC3X
UV34uLhKr6wnCMtDcBtkYVee0AaUVT6vMrZnHqh1KupHBKli5FAKy5gbyjq08289TBH/gGaOnGl+
kyh0bMjOSWtC129uROPdpV5ia38I6IeQ1Go8ybspDHruYJlxBlXsF1qrCvkcUKT7SQN82kQj8Dr7
cu6QMu052oSVxqXOM4ceqtrAnz93ikJOGYXIUuzma+2NRsuUnayMp2DqnU5irOWei4Z62hN6wzNx
c9xD+iLIhX8OzSqY9GUZGbyKP3dKfdXXWXhU4nVt+raMPxpC//LeriyLxZZeUEz5FogEYh1PQXK/
W3lAAj6errsj0IV3SlsgXLLsvm+5bZj2PawqlCm38I5gmRYgXZFkCvaPcGx+h49gG3Dncx1Lm8sO
gmZyFwgB3rItU8p31eZroHqCOIB0NQ2WLTea3epZv98DehDHLKenfS7VK+/f3zaAFqu5pO3k3Dvc
lvCNxbDUnuqJ+jwUP4uiqm3QI6xrsLM9S26z89EHD2b6oOrGrUHMZ/TaknXicYrkIB+383dpI7Uu
SmvDtn/UTZw/RjjzJ10uxfA7MKUfOJwRihuFanqO93wURGCP1v2DMhPKhcaT3f8R1On47+RrtSji
R5TCBhlLJtArbtNFzge1eYVPloIpLkzLphjb+XIrldozJFt/Mv4EcBLcglipSMtXKdNkGN9CRTp5
FNhuBNJpBVOMxWoTNw4G/YSFuLeoS6Qu1dH0TwFgT73yMrMAu5uuHM2kXEz01MB08OL7VuarzPPs
4k+u99urCS/Ov2qIe7a6GBLfOkX5QtL5EUzQm3A6uqrH+DS/ldXbZ71+PPEyUprCOLOVeFWOjKmw
RJsIlPD+KF3xNCeMCc5XQkHBv9VtfR3P01saNYz0lewbodx39e5k08gWTqBE+urMp0m3Ty1hgjXb
+Fm73/Ta3Vm8Z3yYbd+flpOOS4tuTi2nBV/PH1retddtA20TyYjqlj3B3Zd+56j3Bj54x/mi88Dl
Tt2lN/AteMvrSslYrC0D6oKTuOfrR0MB7ZTM94rscXnnrVfHaO7QILqhcP79d4mSQKbVTbX42W+1
9XNGL2L3h1avqi3kAeERjeh8M5z2gWNU77AIV/Uuelte/kTDZnvAQ0DPfHR+ukYetSmEPuFNMqHX
i6pRTgbuYAUHnVloQZcw8Dpt5X7SaFY5h2e7hRoM2C8yZDbJZHRYfX523BNgzQoVu2kEg51DTdC7
XCSPDQCei7xtIGlHPTci9OSkMs2sNVFKfcm/5VZbAyj3x+BBhwlGr7uV6ANOKSQ+HNQPT1qfCOn5
Xe+i4G5jM7zXKgpShV/h/geN2j7R63qp46pfEfXrUVKauBEDDdO65noDAdib77DJF1B97PjP5SOi
TvXtQNF3OJbMujAKbTc9hSv2jVWw6n03Vf4E6tBmK94lLXdQumRPiJqQEa+7mMrTFoH337k0I36N
ySTJB7zta4b4AFIomptVCiNglLC52ysMyM9XFD90/Jq6jWPRaNOeU18K4J5R81j94rQOI8KQS8/t
Lf+ThtizIO+NXN1ogtVpzX4NZqF0QY5hDUKP8BJYF06VMQPiH7O+LxpBwv6MXLGm1oPamtYzdqbE
NzOvPrpbi7PAdjRsOnD0qZls0sGgnPoOJU99MEkRl4Dmt+SD2xK65RYLm1KJsUTLzP+PHTJXm0xm
gotFlCN5rRBC+uAhb2P/6jScAtAGuIjM/m35GNLqoaG7PuJvfvCk8WzrxNlEJ0wQBmJgWqTKZaew
FuX8KKQfTcVwb7YMxgORE/eBQbRLp/vYNbEiijiSlAEisBBbXTF/KDy1fy2F+0qTDBmLQq5+sGBg
zPC3UzlSah+hH3lwlbeF/kG0MxrRKJVYLWsg7Ii2t9ESqHBislaaFvNIV5Er09vvr8yz1wXBKoDH
oZUTs57mLosO+pSa47tjBUV+xQeatagtCLYJzDmm/qoc5JB1NhA4p1AIyNCwE80g/aBbj4alRIJF
3kp3QkwRe0MsVsmyi1taD5jmd7iGmTuWPqxeI0cz92gaxfHFSMXOuqo4GJ+XVOhH08gy5M2OEwIm
G7GwFyqLjPtMZQre2ozdyWlPhFW3/+vmn1UdsMKImXRwC+/FBZxrlpk9vUyO+QWRIQAZzoblT+4p
jdLr2sCwSfD2i+aI3ZNj9oE3xilMTXfX9kvfSli4+wlNzVhWXewkpNcd2zR+svWXP0dtYoJIOs3n
uxtWMO0ibJbzmZ5syBnDdkuzKiasDT4MBAHk29/OJ3KKkV3pfIemTV6A+yX0db4h4m4ffkmNIuho
3eW9onUCRbs3RC7ICrv1LUbu++xvZRXde7aF/7XCkpm4itlIRoYpJ7hXkzWX8BBkYLQIU+ronRqR
rtVsPQ9y+5g27QAoT5zpmjO9fH00+08Q5nXVEEw9s9t940Bof3GgLrmofExOce/FIR0Zg/rHDe0Y
qOQg0wzJLxcZl8KNLxbdNR1t9C0lXQsssGNjn/nk01HwKa3X2plcvB2lorb2quncjPc/HbyzYo/S
vfWP9+OR2SuMYB2E85Qoyr0JigbCI7grVzjfXh22cB05jqzlS3XJe/ltdMdAmWv+f6UTSdPZyN9C
SrBb3V3gPNSINVbKhCgt1ws582zDr0jMGJVjZRwMUo0f9ity0rsbcI9VGcr1tW/qhhUsauy4PFwb
L8gNDNdl4jQdq6LwPQH8h646PFnpc7YCh3HG4YgicYeyrpbALKN2II9i7/dmPAACylsO0/s1xH56
mehxuQS+0rrpgMEwSr4T1CqN0lxOdXwSWWqVN2DHIREe6HdgMYzwn2eNB9KXtRk8gqKzCJ2j0wFq
kkOtStjvyheLmasjkXO5Rw5kGNsRLOynhia0zN9Uy+AfOvqMX1ktRjz88AC+kq9onVg5GyySQdDn
cnnd2SqCXJrgAO47sDXYR6x6d30xvZ0BBWGoVWDbo6ShMW6Y4TWheOb/o5QvUk182IjQ4G73B20a
QRnDsJ9TbM7FeJCYfXb11dKIuYU4iA/E7NXp53MdTq4Mxekx0ZXOLN7CBDOsHNzJhbTGEoGupzuF
drNuODtxdC/F2RvZjpXdxJgfmnE+RQq8JPu64sF+iDWdruNZ32Kshs2nWKUgAtSDonrsi+daN0Lc
hr3sclmG+j2hR8bxBIU1AAdfbwyebPG9lRol+agHDw56W3Z4f1Xnb3YMneL6ukhUAHq4UiNvVzsy
DymD7TR+7V3mc6M5Y6jy2CbBEkjc+EgJruPDHHUMxZ99/q9p29b6uka5JKFYqDZZyUaKhy1icuUg
Twf6Z7bjgATg87z/2sl2687QoNp1kvCpncS2RpPceU9UJmdut00rHLc7BAaeo4hD7ahlkrd3zMCi
X7P1rbBi4TMEDRKoDD93ibC4uG5vLH8HsjlLJvdxhVr8ljM8t0XC+Fu2KIigSZYeH40pqwqWcMga
OUZs6li0h1a+8BHEMkmi4KgLkV/tonhWEJLcADg9Dx1ZK5Ea18ImFOlCrHLFpiG4INnEkf90Zf2y
tec6HVgoMNMYS1g4D0r35YVNT47yseFhvY2VkU2HOJFtr13SfYpcyDMkNTaE3lNH/l21y0Eq84vK
hA4aqhxf8WxnFq84gn5KDzIvXM9JikqvHiC3rNo4lBjtnpNtM2fH0l/w1VfVlWudNxmf9YvNeNX7
XD5AH2F3bWK6Eh8hcTRuSjaY1ZRefhOrU1efe8Ox3u6UU0O+Ck1vZyf/rOIu9Quq+8n2gsyW1kkL
Pt1L4pQvR45ShHsZbheALymXYfgmJQvPPtQQYneX+CyReUC/LhwMAg1bkpm3OLbqVEUWG7dav2Ft
X4Ds7HEzQqL/qY6cOCPlLBBaJQ4UayBSJXKhW5M6Hz29udzizmYQkYu+7iAVhcpjS+PrLHcYrzT6
tawoeTkDSTBxyU8kv+puutesIn7I/N5VPGzFFdCk7IwthCIWwAPEWqBh0N0KuPf2ewqEbG3wSlW2
6uJ0onZsueRBYRkJEkZRwn/o5MZUpbW8BFiZ3gh6m8Ikq4FIQ0hEEUIVxmaJr5waixMe2orfmkvQ
6CHMzMryQQmkHCMNzCmsJQfEa4EzEZ0PfND1TJ9p2j2CCkYSynyIdZY8pk83Gd0lJ/V0bm3GiZnv
a8y0QsXZHQPY/RwX2psKY2zDAYU3uAuw1oH4R4JZTTM7TGwa2P7Dmg8VDeSndZM6ecwcEdndZXfv
CltIJ54wj7lCOnxVtifeSYjiyoBpowRcde4S8qm9l/TsVw+CvtK2sS6hRvmL7UBYfv/YxjhcgI/d
DLEu6gP17OFQGPNvPs5ILoca55lTEDB3E2YqjWtpIc0vjWqLj/lSNen2zroNGN01FHcM99dpfdsc
2peb8WxYrvdgt56bIxO5eFCeqTaEkwFLITDz+EMlr8wp3+6KE/dO5koN3iT2kFTc3FCL2XeukFVe
5ZjGg3f9n1vtTZ5ARERteK/bTaZYQjy6FtswoN8njKarsVRAvXSWABs2J1dB2q3yCePdJEyQsGfo
anSI8aDUCsWjZXmp/Ymm9Ao9vJUoV1slOTAyu3dAe+9YtF6J3+a3cAk/mj6Ihz8foDGXs2SGWztk
zJFjemQfYcul5dmsW9DLTEhBRGSoqP1noK8kcTGd/pbP3UwgyYhjCl3t3K6IBNB5+v4Gl6qYTTSX
j3Zh4PU3hS+wfHpOLzTs6GYAaKCu1XWLiRTtMmx/9HbJhASczRssvbpwuun5DrjSzFzhm4jMZX4D
vcWkSoN/wtZrjFdVA9cU+wcQIdj1G/pHIlOMKwEYe3OGAbFuo4F8SSGJeRqwxlSNrkWsXisLMooE
7lB0FRd2a6xRS2LmowwLt7ogVAMNPEMazsHmNPTZCLp6bowLMsszElSUyySZY4abZUsP48wCwoq6
4BIx6q6L2JmMchc3rwZsZNEG8hHE0O6SfYOoiqf+l4t/FGjdH3Dn7UHAcFWkd67OGRL25+MMciVF
k7w3bL5D+KhhYlA7iQfR9yM8I34MC9egpog5MDvR826wLpcy5cSSD5V94BNcNAdEb4dyEqbiF6bQ
tzQtPjasZsZFEGRca0kVzqkf/yotv8XLhh3SS1ZIvcwPiqMvBwssTQjEDA8yjKmi5kqGLMiEWUZE
MY03U+kfMs2NdG8B+sGjEnj0YT7Yk+stkwdAv+R3UziVMfCXWOp05UvAkKHkD7iT6rEEl+bB+Qxh
T+2VEopXLSUglm+LhddFsvrF/LTRzchai0i4HO0jQILYjWNwOjeJkpTbOF7EmP2s8AFb5H5WouqQ
vz+bb7fSmort9dm0SEGR+hPTs2MVA1jWbE5SX4Gg2JpMn4lRciC4hWNm6L6dNEYvwcini3vO6Cjr
D42ojMUuoDSGyJqJw9mOybsrjzD0s6iUSMjrhY1nVQ+/sPBD8Begh4BBk22esOR39ioJTHeBpzHz
jo1x0bb0BZg89Huwps+LPWEnv+Iiqjp4syiCUmPa92muQW8QDzrLoRUxP/HkqBWYVq0r4Hj5BYHU
TTnxQoM4SGWn3GU0v101LieRSBaIIA/FkfZxQyR7ZYgOdirGGbiLuII+tB1l5yY6VnyDZhcJPb2a
FR/sqI7WMZdnP0kfUzDOJRBZmLFMV7K8bl4zJlhngaeoCsm5Idoh8BFK5L31YO2j8sRTCD2p5hAU
Q7/cOISy1PIQEcTE5bsYiukukxA+oB9VSlytcPQSvcJlAUYRZ96shhgcdsyMpCRxWOQ2waeXa9EX
aA2eX4UJ91UTRVCGMr7OPuRo6OHl0ejMiHjSUtSIRQDs4NmdmB5DbbDzhfQEI1VNRKUPGdXDvAG0
R6wb4quYg3sABYKKPt8TrnjZB46djOG9cbGpDMRpu0kZUs0+BsZk+OWRvzuo8PMUObvmKhTz2KT2
9HhZ9aT9lZ1ZcsmUiVtSuM4RyrjRjV44R9wlK/+r1Ptl1VPdkMjPsJnvYTAvjEZNOqDd394uM0QD
mWbozehxpU7geIf6oB8zOBw3XEUuE1/xkTlWdAo1uWIQKRZ0VWQ3nhEI6WqWqVjNmNl3e8eNPF7z
oIepm+QhhR7k/+vJ/w0+bICzq4eLjxwzdr5jK9kGdvt19nfMAOXMy0CSBx3tFx/Frdh+5S6YsiIF
hOwlmRx8XnMMd3OMmSY+30C86HspAhulPeGCbSJ1IF9VfCLYaYhWaN8FnbEAkfDDDq0U8bcUJHB5
GdIgsa/5CNICXpZIA4VKpODxe2LOWpTRjm2Nr0Ik5AQJy26Nl8RLxgb39b1LEBt8Bc7wGXa90nXs
5+ZTQJnGfauYFHTVwxkuxzp8c1eGjR+euUQ8UaNsh70f5UgQdBiRAglo9bxeJ+VoiIjQ6Q6vICzt
ClfUNazrbgf/Lfm+cTHT3BnBM3uR99MIN9CRdKz71zbR9UVkppqkoSefKA1svVzfXUj4pT1uq3Xs
iU1wJBwzBemfKMBiiRsd4qWdfuYuEibfpuPU9r1yzf7B6G8reCW0JSL7SOdNiVapq+PBKUbq1jrH
vReykAqkHBV9cTz12dtzSPdNN8/dhcZhNzv4xvrc9eGYHRO5j7PCBr1LZoeOJjIGB79ClGLvChvo
whefD0k8zRTSGs1uh7/UFAWGH2CRCiNVITGF7WiktJ361URIOdYpOmLBkgj4Y4mjueU/KbkxB6fl
hw4+8UA5CfHJa63dxOGPrPcaUOcpHj1p4jMKHbHL1PVyNolKVPxBrHrWJO7rfF6lGn5FThEhI/9q
SAatnagokQGkwQuxaF2vMj55F2SwW9T6TuiimJVaPcNgViZeTtzkC/5iaRKreKnB2RbHftj4Uoc8
Zcv+/pitE2PFIYqFtrR5JL80CFprc+mvDTlAZs4XIubips8XxkmElVErmurj2PAX8L/QwVERqiEU
BxD7Ni/5HwlopRiJDSM9/gVsBUnHpZbtnC0fl2SEgwJ7UkU4dTKGWRyBh8y7djJiWyQwmRw4dXNF
1MUh7+5opb2ETEPzORDGcGtQa5463zn3yRJ2ldGoap4hJw4qkX6Y9Xy9B81AAN4uvRjUnzSWU+Qf
KhMVfQHM3fcBGFedhtscIydcKuafwXMesyOHoimqNeAq3viluPxEFLb+cHkZenkVCsQWcDDJWE3Q
bZub9FcLAhngzpMNKMPbQ5uMYinx+ajFdRFR5MnLzX7UXxMA6c13qRNaMxBHzQvfTJ9UebDYivZX
AhB2pmAsSJ4arzBsh7vu2+LYfQa3EWUzSbEzISXhGEz6I29h2oltdymvm5ZWKvSR87IF753y0ZMk
sVS2gN69JVV3RAn90erkZ+zCjIKOs/l5wtIbISNoLxlfF+1o4mADvbVFCCEnELPDbx8J71mxFS53
RKMcRpHEfCw47H6DiyU2jGdIdQhdaoK+8Fhi7X9biaw7pfsi8ouWfpcUHcq7OmSkRTzvbaHBKhKy
s/5jT7CIUISh/pMRaq58yZGhyiEBemfc6KyHeI86O+jalfqqvuGL6GgblYIWegnoAdM9DcTwr58b
JrP0bNV8fVwxtXMDXDbBhBROD/3NF/CfoSS5PFPEay0wDEwP1HxiD7IGZ5i+6FihpcEWA9oMuXIP
YcX7X9JZZaN92P6Mc+d84jMt2fL+nyfI2RMhLkeGRCHUcbOBpZjM3fzx+31hhL7wHKfhaE8t6xBr
LwUlU8ibeUckJqVAcwLyuPuQqzKzm4BFzsk5grPZChj5P3sdOgqhwI5egbEzrdog4GJledidONL3
v3nyRQsA+DizU7cgIC2C8CBbkaSZpr9hRHuzMdb4J6jrnmQ+HjqY74JB97UrKjOkIf1621gCV5V/
DBTiPELBYZrg2ygPQ488ADkB52WJVE1QkOcDCeoksSwSVl1mKjkwIHiDgzXfIAk9IaSmo98dEhyM
dlCfxXQUX+CuiAbIFWXQruBiFerKvd5Zdyhkz+pLM6YQabx1s1UVW37iAcIiN04uUcxr6XGXTupd
7SozY2SqSI+C0V40KlxB4e5Pw33nElxx+7U/NTekEYjey0hAGiaHG/KCRGJGDD4YESKwZVR+7qqz
bw2fEFwtlQaZXp+AM0Xi++YVIykbl10lJKffSUULm/8kH5YFwVT/sXLnzof2SuhmzmvXd9/svd2m
Ao9rM3pIXlnBGfPNj7w2zqNJAsnvunrnWh2r6WLXjoOXCbgL/iRdp/Q/AtYPm/0Xvh40C+cloYA1
c3zVCGh/OofeRsfB+oP0u2QR3XIm5HLjrZQqHZ/5pfAMz/OcQGBy5ASBugh+ZefegEAP9vp2IpBj
UQetVqDCrgFGLH6vH+lwBY93jXUBxSH7I+Z88LcpjKkQspURgQkD0fXvy/GKBr3hv20tLwWE2UDt
vcxIy43os9aFa4SWw36Pv36KStW/p4y2JMG4H5qfHM6PdhJfzvNSt0OVO8Czq207xVnX60gD5mkP
PXud0f/4RQj+6JDTKbGWdKgpu+ZbZp9u7MXIcj7xtemndVYnCOlJZIvpa5tT9lvwc0eKHS0TYr/F
dh1nfNidzabN7vF6Pg//Fej6emS6ISB+6SSMZqYyW8lRdN43AchZ9dp5kG1fooI5ghfzEYOr7YUj
aKHAI4B7Fidq0Jc44xpIdgfw4vW/eEDGwS2LIJz3QoRGsnuYLGAzkDnXIxBLQQYYL3Vi4iOmXiN+
eHnvPgsB/KqLPnsdY8vYKCuP/QJirbBdo4oQQPfrfgC0VrOcPprQe/PR/T/u9dGVdpyu+Pt5uvhA
1qDBjjy1jFLK7EqrfB9Xi+mX87xmRFeaKeP8B1DdDFlMYgsbI5Hc/1JNXgGy3FhmSyA2gDUh4p64
F5/wGWFU/eE80RtVzJ/HDm7NQNFVCiIT8EKlq03OPyMa3kF+nGozVJXH8lMRD0qamjdHD3o8Y+nq
Id1/wekGeyBXZ26vSG3RY6EsgSogKXO6ykMYalydZDgBUujvD9KjUWCUsBJuDZuwInxsZ7iS08io
nyX6TEmy+HI9XjFygjcwby5/gz1ECthJTaZ2y8pIg4WofaCeHPqz2uesQDgWEFKedLKzBilCZlGj
JYIbqLgQ+j5Uz6O0APEQe8j4LpNAW0KkKbdcO3pgivaJfYKpJFe5YnM05wFFWjfm/xbsaZBSIC1A
m3JhR7RXot2FP3QtyPjaqjMxJ0fpctdqV8yge5pxKuIujH+7nuxQfytBOMFFhBe2SVYBP3RAq4BK
WvOHOWgbYfNQ+9/+RqvORXFkau/Ea8Png/LhYjMNCUzwGn32QtJQIXIVNrKi7zGNe7xDen7Xd9G3
ATwj2ETqBfBMKxGmJUQ7dPdcDSVqKAJVxVprCj4SZ99ARU3VLtTYD5Yvr7Veycp7i13iTUZhGOQV
CPQq6tUAwrOAVOsCWTR934H6QTfHnN7Qi42hp9UDjbrvdrQWFku3TP1L7EOcFVhnW/p69RlqiBvx
Tt5zbvVvjPSQF6/ZiXeB30KAAAlBS4uTw3v4ctb62iNrqOKWPHPNeyoEYEksYdmEMXhzAwu1SNeK
9FOtIcu7D8C23e1Dk+yir68kA7s/M3lkna9e/+YZEegHXFa6bXdYuq79qpCvE8BTUpY3gNa+H3sC
9XLZ6v0CriyE8GY099jSl782rcmh1Kw5y8l24DtT8/WoKfcY/tN7dW4ePIN3HylDTvPnxaXKShTn
9yZuFZ7oEwmMOczQBDRwmsAd3RFaV4Jp75T2eltT4OBDb5Eo26si2t/XxoEGevdMhwC8ExWATVHf
qbOkl47WCM0UOAq2ORoSpAAYK7pzZbNb2ZVLYpD4A3uKSZwzNDmsYBO2K5f9DZ/GNLciae3f1Y0q
CJhSGO8N677jrWY/UoG+NFHelwi3L9yIm1t0sQWp47N9ZdYSs9dfexIjR6EIGtwaBwc8y+swWzwC
g0UBbqt0p783yrtPJW2AXcEYfwijAhwgXefv9IoLOTv1Pt52jokv3RTLvQAXei217KsuSW6PkgPN
LoRQw/LtgBKB9N72zfMsqSis5OpxYTbADvBV2hqVoVzJn3LM195tDgbYJXz6CMifV5fefFk/ohPS
uXU0rAzieSbBRJsMkotdvh+Q5A2dUpCvWsqC/kNw70o+5D8tmssHPczEZeVyxF305uYHsSDMJCvv
NBZhTZiJtY09QpI4KacEtU5ewr3ybtzTMOTxzT5K2dHwNJDn/eirTD85Otvv2bS/bnzKjvoTH80R
ge9jZjR/HufpIo2vrBwpdZ/wRdCrkS0zWl9gkyEOfxA6ZA+nRn6IGkUY9vB2pNt3vJIIjYdPQaSy
Z4n5R+XYQkZ24EjJ/x+Z6M3fJE2qFujSjDrWrcWiyuZDOU7HjjdBQHiitRWnPi2r7WSArLtUG0y0
lEvcwKVfxC42oZA92L5XlLF/ejg1gFi/IQRSeB/wNzUfK+AJFNO+0JCoGiObproBc9C8VJ2T6ha2
7BTonXHk9VhTtb32wli5iYxAMIPGEZYoi/0JbVpoBQ0tEngKTr2G9onoawtFyBWHHeZae7cXhZ4b
9Raaoy9Gc/wy3JP/7uq6XjpSqdiBxn0zIDZByNQLXw+kHTiJQzg8V2GNrZou6OUftdhiGNVCR04W
w1ac+65vnoZKtPQ8bH4+SdXXBe0W7x1TZxJcthD2DvkUI/nQpM/e6odOT0eVLakDnmNZEMo2OIDE
uzBu9c0N+ivz/Qkw2/f7choo3BDZlpfQVoelGiwVVfr5lIzJWUpuL0HzUeqdkW7VUxddi3s5uh/b
TjcNuAIGV5K4TLOHoVMsecQkLeD/JjIj3L8iN4i8Fiv0i79b8iUsOCfXzai+IGB3VtVyV3p0Jdfw
+VXq1GP5+59YsYcODDK02gPtG7vceV1WP8YrYpCYtCrumSh4Hxm645PEIYeV+22Ic6xDEwPPTjZ1
jrvs7+JlB1Zr4o+rpqQNqAjpoN18XS4HVX/iTvkYbZGpArEMNcCN9rB51PoIMm3jtoHWhGMITHwr
gKQeCJXQhDIWhlHFR2CKrH7FTX82kKXtksMpMzivoxY2J15q0h1RayRlq9rMfGKi6I9u6qWyJmia
RfKmSM/1WOnXsSvOgFwi5V0nq8k6F82L5wO7NHlBsodhjBp0ewDWLm8kCXayJN1tBVN6DuWS2DaD
QbEi5hKWyWmcQ519QedgupK8kAcZbH1SwF2KIY1kG5UqyXs+nJsKF7m95CClVZF3ZziUr2abSkbe
/s2zn04hBaz6188ybIcr12Zc6E/N0Ck84F4XoXD1N79vD8G1uRcPtJLJYcjNWEDRVwXtMCdspuqs
NzhPVN4Y1sMkGb3x+3h5/zQ83es35T5nDfaKPzJuHJoIkwW21SC8AQywsuJToaUSEnc0j7Y8fyAQ
uQ2PWt/vLMsEFdOLzzeHSPxxc6BOmEMKlhXfG0Sb1o8Yt+F0A8DMXkXEphhoe+FVFcABjT5ed9SY
IdSqnAcNWT9H3iN7xAmB0frZxj2Hwg4W3bGS90221U/Wt6J7I8lMRuoqkWkcWafJ4J0CpQU543e0
/FOouTXJZPwrmCP2q+r/vOYy11QoEk06NHpJwHtpNTbUsCLEPRlW0yiYZWoeWiJzPR8V+DOA4Pvn
8bDlnOxrQLNfpyejILQ5m9tV3aVd0GmpHbcz3VPhF+hVSmDxXNpmQ3lvQTY5LM3rTQJ0+uUNEVKL
DO3nfIT8yl2KZ0Q0e5/JS3cbyp3g/YQ9V5xahURyh2Cgszx04VwzocPCvs5Y0ixjEd/aRPMoImgq
mZStoBvgINtwFGaPsKmPzvXpLdG31uYq2+XZzUJ+wHtuUsaF8Xw4m1kV4waekpRX3Pspr7he0Brb
NHCVr/ikM4+TMBP+eEZXbE1XGXfHssHo50NW02nPGlGKIeWs2pkHdR+/kML23leJ+YquYmcDgr5F
9/Lcwo9Nt2qer1L/9SgVsJfLErii0VCg95YoI3Y3WV1rp48s2E/Hjzjgxrj9++8Qjmq2ZX4KakmF
greynwTUMxFnObQO97Qmb6I7gqXQjXkAoJ6CujBPgku8UbJ/NwJbCSh24eP20zBHFb0zjCNwsDpq
Ouz0BFXstd/+WXkZ6jM2T6DW1rB8twt+L2oKHmGRl39fy6+CVgB6KLTLaWSTicZYTItNXnehTXQ3
TUso3lS6Ud26knbQuxgZNXJ9xID8d5NeAcaNn2AAKusPN3/a1Vk11XfkUnypC/mZvqvWcdDuj4b1
CKE0gyBou5QBqjPWXDfrGZU09SrCwusGOlqudGdJ8JE/NM4v0y73E+kDSZ/GqwkPzJ3C2Z/RIu/y
6sNx9PRG3XSb1t4ujeJq/ZBtVx9gQRNLUZWgpSjBrPa0Wfo2nuc7TFsMgZx68Gl7IMDKaFi6QPik
DtOSW4rVlA4WdhtJIZr1T3gJTf0ybMRAClOhlD4xtM+1664hCbCRb1M5T+kT210yMTyrDGVysTuV
KYNsnfidiY9r/J6p49KyV4wzErwIVOzJnW8DpXs0MEqARod4svGtjA4iDg6sZ3vF2hw3VyTStflI
xvAJBjupCkN3dX08i7JCDBWPsI+jBAqnUpP/uHgwexHb9DVQn6cPXRn+iBXOauqAB9n8hZ1WXIu3
0BwbjcW4alub+lWUBaXcTyLl6H7R1A6KSmKTa+s9X/ntgNQ3zUaW3aTFc1zqfSlfh1l2sUVGYJd2
8xs9PDh2FkesbnF95en3LsegsuRRyJCh6M/7JIB0tkCBLXIe73V6QPqnEWOBq7k5gCZBXN/Y5Zie
bKNLsr5NMdTVspI/IUjm91hDN4ZA300+jbMWeTYD7cQN4yeyFTFrz2vKYEtuHmySzEyZJiBiXZ96
v77g88yJpzmJhWJ1V0Azp4zgyKJDeniTzS83QVIvGFMmodqkZXUUAEfQHO4ADmBKlVtVVfuNHRLs
RjDBG7FyTLfudBVeDt9nLbf3MtizE0wmTep8x6xRUv1vx7bESZTpd1vweslZKAuEMhiYeClxCqcO
60icETURGW8Ozq27Pjdl6K50SNUC6Swzvr2VpM8TAsR+WMu743n3AIXGZekHL1sT3F15v6aC2zgp
YaV31R/MJ9e5tEsJjSHr51yDiDzLKLy4BwLybRUf0hHwQxzUw8+l/walI4hkqoMQ5PLLsI1Ltj/C
qPPrIrR1sULgBcgAHRwXevOpTK90CwnWYHdgyn8ZMSnXbSbiCLw3yJtQBEd70vZWZq6QCOTiqo7C
8MuzM+T7xSJGcaVxdjuZOOZP+wHjxz+bXUKVgos3ktDFOPuE9CiAdgUleBZDnVy3FFu2fDOvsgII
JFxu4Piy37FjcOsFC6CcveMXzXTam1YQF3JUNNVApM9lPdgG232sXjChhChjgQdaSW5Lj3eJbS1+
hn1FkGfERMsXwaDOde6Q4kPJhyoOKW5EMRlh7Cm1bnMoP494ONn5vbk3rEZnseIlV/gVf7XPt1Kq
QOFACEvtyBetsmhdRyBJK4m9sttX1xnYEfA0p8kinMtGu+H5ifpo8thVNx7Thf7j1VTtFSFhtjAH
Cq1zgpquMdGGbFmTgNNBFYfjaZUC3b9haP8sr84CdDZif3YuNarxF2Y+dzcGofu74X7KN7SxOQC6
hETkEWOrsfz0jqDSbn6MfwZj0dd4ex4aefh2envuVTlEBiGm8N8uutA6R1hoE+8hEWvW6FDAt6zT
2/fPRYwkpOX63Wj5bs7G7fM9LFu9sIphBzo15JtAyXOJsDyQBPr7jM11li3nHAi/C0sB/AO+HS7/
7mtEMObHv2oB9GM+RNEPxKm0OrZ0HIDthvIYGAi45LOIuqu40PFBkU9lEt2ArQHJ0w9wi2ZFdecE
qGqicB12XMEddpSPfBlyPU1BhzTi/JpxIBlFxvDqHHqP2JCqIidxPOzmIa6SLFXYA0FpPLmkbe/1
5ZIo4ZzfdKT9d72r+IEEVOEmUxOcAhoae/sHl2AYYIaEwG4TgwK80IRhcT5brAFYaRE3AMlGdOEr
PyyxlLSR9xmyx51jBzaW3X/WZI9n11JzApXsWSwbNs5XhL1vPsaxa0+dNtAluwW3zElUmTK/OMRD
/DGsVOGs70sMt4gDffP8OeF8iqe2HVQzYKCiSl8tJFozqq6ANZb4R59rXN7RVrDAAhagv4Nf5CEh
a6kSUraUb3SKIwfVh5Yful44AKJWPMUWqPioWfiPt7IYsGNB878sSvhyIYEfeqCu12FCqKNv9Nzp
NsfCHYuQiByQbGNB0ohEAzCTeE0/6d2t0XAMmMn+b+JtikdGTsPtBtShg5wQzVjCHJiz7CGX5Y3i
3H6kxCyVEvFHl++4TTydejq0HlaVz/6Z6U2rqGWW+T6U6aC/FJT3BFPS9rrZdXWksku2t0VRqOAs
lI/eHCD0SlMlhU5OplTFQ+YDpeX9+2j/GWxYtaLq5/6j7Msl9ra4D1HjtgZnRbDpTGLnzQSMxY15
MuO9+vhOHrzYKpzoGUKIXO+YDLD2UbYjk+d4e1V34Lwt8V4Xyprg9KfyMDAwSyBMqyo+4tuTKpyf
Q478iaswSLqQDweihGdyDErFJum/lptTRK0mQBaN6sXyn7ZPYu7lSQ3i3NT47WD4D/hEmrn2gRWg
N4sFTPSref6xYkXDgHQ3TecI7jV4L/ZRlM1UQGM09ITZwwlMX5OlZJSoOOXu/zgiujpxs1xNdagv
Tvqsrg9ym1lee7vt8h7w6ANXett4EqOeVZgSbaOliclq9HQ61vGzj5MI8A/UwrKlFyHjpLVhqJLO
eA/gwLbXXLxmTKeMP8IjuXStv6s9OKjv384v/2WE8uEg/F1kOOeSxnsq3Loy3w6jAX5yKf5KPHxq
pcqPasNPSnztNvy5yQBWqujge0sLThprow/ESBF1SEOvXSQRZJY9bqOjl1jp7fv1ojD3y/BTS38b
5KBFYGOTUVHLEoplc2znAs3xblsCIjgrQ1ej/LuPAiO8pWWZ7Xg8wnYGvf8J7xqBmBMe/FRNmmn1
+NE2bUiXodvGLGTjA9tRGg2NeV6G0lJi3vVB+EnduI1tD/nd0crwHu7u+Gbg7JPF9fuWuhKBXrT3
2B/kyZ3Ybnd3WjA4d8bGeHx654L+cNqZ7ZK3VvMCTLYgeOcJ5cKBJpw51WbRhtu3QvCgozFptizZ
Dc8r9yOFdaIAz5TtduBF8gBtHJ03EGqPoRH7a1kGnbmGp1uvkOc80vl2tPzilsfPJ2WEcedNUHK4
Dx+/uivrpa+ehD2qdBqLhXAfbY/8NBHqy++VT6GADLWDHxIm55ZeY3N+QxCJvfjXByHZW0/JtE5F
WPsTUpUl6dkHijNqDcMKwR+7B3dIeMnpYcUCX9TcwY2S6Gzfg/ZW3sF6s5rIv+8Bj1h7mYEsky51
jDMs5plcci83naXBBXB3CCb+BS/mc4+8BsHUgKc75hSdAaT2PCfSY8P6aj9e3+66rMO6AkNUKatF
6/rx/YYBSKad0KcgyTRKkqEBzo12+/NFjMILXfFZyXT3eJc2ue722FGK6UzWQcP0A8uUHxY8pJic
XvKwgGc/utRJa4aMLyPzV21/y6ULBz63X14a/u/p/vfDH4JhDzab45t4FjqSx/nr8ArdMYe15IXD
+iQyUNdLw1hop2hex5egg9ZwBupJjqbGLXXGlVQDtSXH3ibhQP1dkVZvHgghOGOPFV4Px3yXWqA7
a/ipaxW17g0ttteWFN6UgYWNr6P7NMjdw0VJ2V6gPt+RMjydQh+Ts8F3w29e1TrQKeSBCWzF1qWO
We6dDgbKOK9i2lNWwEMCiaqBWd0EjsDan5BT7TSmcwv7C8dq0vrEMx/YYSq0wVLYszmV8unPCogw
ulZM+n2p0pyx9XhWf4ccsizawuSGJWr1zdyNNdYssZgnLkdeKlvkrvSKzK6MrkPbhAVHtdGB9RLe
MJ+EcdC6uO10zpF//v3voDymml55w+KI6CeVq/wKu059njR3LWYMSevCcHEDnnrGXr6t953TWHiz
GvMw12v/O6RuDTdDbPcUu2TTPKi8SlhhiCYJr6tsSQWWEaydtnVAb4azvUY8IlW6gdEqwnGmP/Kl
DqK0Z97OwZo/yhue8DlupV+iBM5uGSMaYNxVLtk7qqCUF4dk0kZd4zu5NkbFdew/uSB8qVfWsKJd
XuwBSWqC7wDXjDuCHJ4z56TC9M5fEkiWL4hDxlOxkBDGcEfnMNu9UzirltuqMn92lKTgVtjJJ69k
ZMI/5bygMkrKAzb0BdFCQsy1g7BpzRgXIuNeIAn2qb4zWAntHK/imwwwo3CWw2dXco+ObAua0gIS
P7JCKD6VcJFIHIYtFic5zsdkM7w5UEaNZQpeDeKe3YVmnDNa67zBLmnbAxeAA/yRuJ55o0QmRbrG
fazQgKT2tQ8/BF0lm2XLCke0XAeBf7OJSOYoeowj4BUyb2V4Xron8CKp1XpBH7P4Ha1zCVbjiNxV
TGKd9/19S1czyPk2aIsC4iwu5B/mKIAMRv47sDhcrm5xKdtq71qOBV2PKh9oYzKJene8yicQJ1b0
MvpuAhMOgYKsoZZ+a7/3tp7qyZ0+wCh+8cDvN+twP7QRcxD1yspWYe+vVFHrYZ98IV2MoBS5Vvbi
SSAw+5tI2GbccLfVBo2QvH4eDD5+soOnGLiCzpfN4/fzod1ILil5Ncmvtyw7/Vh9vUpdYnW340u6
vqiWMbx+suBlSoGO0qV2y2Qx2MGGCSO6QtUAp7LbESOjqkoYL+15R/eYCekVdi+JzSTwg3DpvM4B
7NbHaprrmBo9Rq2WZ59MR3ylCfDtW5hApixnPx8jmTu6J8uT51ByWOdBdtX3hckmrStDOMsbiPVD
MMLdL/uy3Nf5P6bDrP9KN3ubOfQQ8Pk9gI/VYcJvKRxhgY2wfXRFF++ZAFP6LcXA/hbWbsy00EK/
iM2weGtBDAwa3jbZP5HKLSQTXoRG6v4MZNaNKxgUuPUTb2kGJPpBANI93CAxvvUvbl1j8hZo+7//
gO1N0zg+g+u4TxzOsdHXVmtuXx8Onq8H4sD/b7X+UU2kgiJ88h6WNZFqp/SyQIgX/j7pP9qvivde
zHfbLjKRAAowKtw10AcfjTCkJXpNs8F1iDv3gmnkw6DuIIsXMLr6fp9CWZAck09GMKZPMSXnz8Q3
OBDC2h+nSehU9Un8kx5atnRa+qHshGQiY/cpOVTjzd/1PzjZHJ2KqgV3jO4P3MjnaUdYEIC17TFR
2poCSydEoLkblU9Wy6Qe2S1q2UWHrEpMlA8mKOdjc5uM1F+Z+f5SF6Dk7R4P6xA4/u+WBCud8Cb+
GSLHO2En+CpgCAu8FmfRu0Sn2rpmhR3ZKFvuc6uhEgThlXu2cnBkx12wRgq8Fnj7OTW3Ini5uhPL
7t0OPfYYsWschsQjQurwWEoSgfr7BdzrceQwKdDOyuIevNpId3aDuNppk6pU7XTg3lgBcgARbAyV
DnP67cSC95cD6vypWRj7fJ/Pba+D6JVQldaPX2F3rb3uRwIqS2OTYzTL0Kogp5ZatFZtoHI8jdRu
H4DeCFytCA8tM8ZnrVqXWgtjMO4dzxZ99B/AzGnt/ubEDECE7J0iFbNTsMXZ3wuIMTdMBW0XwG7C
Eg0TLLaca5RWg8/IRQKAhZs8cqmjohlQVFxDOvN5I1TwASMlY30S5CGxGmYvMHFIh7wezRY/2n2a
vhQC72E+7PKr2bpo9itdJnQLyQSJkQMFK6L0XOerfDk5VJWBbi74a9rDG3+XZvgmlAQuUMv6ulMA
dHBnrDiL9eufK0kQ79+7oVWycuCS28Bpn1H14mq6eLSH1BfKNuoYPphUzvge5BQecsNiBMqDNVN4
fb3DG6x8mabn9Q1irXoyll+iBgH+lIJShW60X171XOZWV/GpxWpvrkcTyWF1OfHX1dRyJnvrPhDg
a/EGwsRzrq7CJhTWd3Mwcgsv+AhQx4gNHxEqbXo+QEZn9g3Ywsjp0BvivBIyqfGv8Dlr9WRzqZkn
CNsxbnmApL76GnR+wvI9quu1gs4IMQBZWGltKBL3BkSo2CaEOJ+7GZ+lYYd594e86KLhwKZ+iN08
XcfvawUfeQ7iq7F/QGmj3NRQS2M45B3Dzyu6hrvNTNCe2Q7QuPGizyUoViytJZJcLVqHkpfGh4em
GbFXfq099FV+pU8ScYLI4PVEaO1NQquPWstlnlcc/oCjbqgS8G4RM+gs4yMW+QmDF02dDSz3TNXq
Qa8UQ/4lZ/qE70LA+I7IVOS49ioJIxhXD3TX4ubRaVRbxlASki+VRaM4i16ZwFO9ZSdmWI0SBgZl
OSSFDWEmKRdApt1hJDVVJiUeuCLs0Hop+rP181lCZl+eoSP7KCi8ZMrVXXQyFG2fbmWfazwN68nC
LOB7Hf/MK1fPKQiD2dT0pOLOS5egvsX3sOj5cVAxbBdKjJoseWnxZviP+CZ0jHBmdahY/2LmVPMN
5DlPahsm67/d9zZIfuW2o4nmRkFsZaZdddfCxv7aLXNDw/T5tOj1kFf2DvZxGtc/WMp1pZALq2kg
kiB4baeRcqr6DGx3rCysr8fhsGvyJzvuRUh8xQJ2ukrmc9eAzGAHTmQXzNIwgVMf4nG7pEjgjg2R
jKVTUC/f1GyGA4qR71vyGDfCNrHq+coglgVBo1IFjEZGhhU4XbrYlqCeg3RTWYpNZ6sBmpaxV7fg
BQ30eXyyX1OSN/R3e5Jva0HN2lNI0YozyDbpPJcOjvTNEbnnoUI211SlVwCkNggD7fTHabuEYO10
Q4Xm+2VuAMvqTp/934UvyFSomEgVGfJ+0nt3dMzf3GkSAyzHj2SjAzRxjxL0al+Z1SGmAh3JpjBR
4jtEJVmDkrhkwLoLOdztjVEmqvalCmfuuGmkmJp5F0KO3amSEzKkDhTWiT8w02Egb/KsSOO7xuKe
h2TDeXAZtEAE7EqaQmOVHa/m3WgBxBeKui6A097qKC6q5hwTgt3h7uCq4DJmzqhELlZbQoawlV4w
00iDKRaDUK8mlFK/0buKmTfk1rorgNl5owWgYmBtbG6MfG7m5J5rCztf6c5aOEFarsPwzsYMlydb
/n5ACiLwsAt91MpLa2xpLUIu0LVVSzQr4L1zFNKDYZwvutgEfuDuwc4Xgp6SiVCpVjbnle+t48g9
oGLUQeSqPjtL513mnKeKXrg/zcwYMYsCZd7S95q8gafSocNoqPCMBakzYgnDheDjUqwxT+jbRBwE
wkBlFfttfxWRT31d0ybrBrnh9CP9neMGwJPtlmKDKXo+R3aeBBr12uXTgQTZmt6DGa2cNLWRHa7Z
SVmL1BL5sfbK9gV7fOern/jJp3tqUATwznHgL+SCT0yPvn1fh52ztAr39JRJFqrd5CPXDa5ObxnN
AN75wiEfT/9AzQw0B8uBhRmTVNy4vH0w3WIQbhZLc3BwENRu7/en9qrb7iyPvvD6kSBwjOo5qhPJ
9PAreupmGpKVHI3b8rIBb0ePjmxrSodv+wxsYoRRDZuH0+lLnTCxfUDLITPHgpwLOsp1NvZ0NsMZ
YR96cbRSSRZbSqcKsZgj3dxHQBiIFcHL8LY4BBr5pYPcPHf62CXlzrZ7Q7PWS48C2ReEpDAXNMGi
qO+XIAKnV4A3lskwmDkkUk0Ii0fC0OIFUCUC6W7XuPghu1lGY8mtEgWW4g/rvsDXFAPrB8+UUtzC
KxpITZxroQJdPfdBL/8hhH4vi5qF1CMCqqkrvTjcFWYW+8iVImb1hLvK1TgylsGPUG46hLIz+qGY
sfeMq/1pD2im/HA5yhsfBaAfF7JAIRTXuxSzwZI2KKVl9bcYmxZd1CFz7XBWz8s5Jm/qr900Q04l
St2xTyaMtYJffA5s6yB9tn6MrRjaPmo800BSPzMA3hG58n/NKy1lWAwF7Gzw7CX/Mt+crVPZZxW6
QthpRYJrfaZNaKQtMsdSysoD1UVGce1XnIlXHu/ao5CsMZ/Pf27lSPp2o04TFVLzvjYPW28IKvXE
zJYAP54/gq1jhhofLYIeBmUIM93lDRKhVw+dFfOSUPmejYHdpWxGcDKLvLiksqA0fQERxsPLQ7u8
v6r0jplbsUTzdnaWuUbF8RiawRWQ93SWmzsQn0ZnBNc0Z4RZUsv2f5gGrA5Bq+LecS/3MNUORp+w
TH4b58nQX3EB8w+rCmO+GW9Hv19lYcPoceSeftw2w8fnJzp4K50YzUv21qbYNNC71k/p4haoh2Gn
vnn+uOl6iHbB3Ep99BN4YU+z2OlmJczOfMuK/u94Iq5GlQ5o1dCa+YT4GvUulNNdnP0li7QeA+6L
o2rje/3eGOY0pZZtdcGKpuv/EE8xcdOdAeFMFoazhGb0isu99OmpRkt91rKiHjwKAu05hnqULea5
rul12cJBhhQdt1/afdGYe8vAl6t01mUNYM2hep4E40sCQD82rD5sMpUmREeFDIZ51I0TOsXw7lFw
SAohu9u54SK26s9BElOS8dRc2B4u6AiXpmCyQtGdKYXygCV82GOORS9q2LsXeGlQKYV3X/19ljrG
hip3M70uPWreqZJNKwwIJjD02fdZMefgLXdTrWpg42mAGMgaoUQuEGjkWQNMFDqPUQD+oCHQkgAp
chv9O+p+TvYiEZdCogg5IRmRSSSmlRRpsP1/qPAzRaR/H94UiZMx1Uoi6/GHZt6nnHDxq+yFbDIu
4GD+NsDrIK7gEeBW6ayc+dOphJXnXM+1PWQd+e3U9koYjVEa6BxRdIFKK6LreJVTVAedZDAmsKUy
r8mQtVWF3RDWhxFSETxfrQ7liF2FObk/VAg3oTCs9YaAcR7wfnJsG0Bgj5JmVRVcoTXcqfPLaq9O
Bz/5n7nbctGlNAe1DwThpoSYHK7l0Nla+yoOyEAwz6gUwbeNfl3gKHo1FbilGOkgBY2kIi5W9lPG
uOrfTLzR8eCcFafrAJGsdpEw1w9LVbb5RbhFYXgHQWcgTIYC9eFggKLyUWosp6Rg1wG7on5/CT/w
k0eVpvvR7a/oFFlyoGMTWK1ocaIj5oJ6vn6QMgWUgz4J3+6SKJj/ZJeaNuz58sacs7yk4GVe0j8p
1fONJcv4IkgHIAf3j1N6zVMKYnmhQZcHHgdp6Wqiqq7xovD6z6vHJr/euEJvF0eXA/1oxdJ/qfG4
ZnwTlQyi/P79efb6dIydhkwOO7Kov0HZWfU0ipxmQRX/gdBXBBgwb6nd/wZlhBIM4ORF6MoeLeqH
X0WhkUDuUpHt6nZ14q0QaU59k8ac2K0Xob1DA7zXPnWgaJcEk4NctB0Mfe2vYg1C0sI0Dy0/7twt
CByH3elCJey7Pjs1E4+irD17g1OXUOqyVDAKpb8/X7DTIgLuxi8KX5na0Pzs/k2xsq9AuLhD3pzn
tGdIv+Rq6SWLZEa4ylnpyTwFqUT/FYzbxE98wAK20d3TURhQTjCCkiJTvjybFEySvl1pOSPUGQqG
j6vjOIWCTvk3dbYmEe83QT+pBTSK7tbfUHdZPj7g5Lgk0xZUwXe2CNMHusH3JJnqA4kyE0hmx0Kp
Gx9Nvg3w9MCtteQE5zwHLyHKhvl/B5dRPBNz9i+ak/na/O595Y0nbAnmMjblmwbx5lK574LQytL3
85DAbJ8CF57tWcu4EEgX3a8fbYK5Cuno77VLatM54SrjoCRsDtObDouBNBQLgh+amYtm3kDeLMti
8zdu29WKnuu+cbObSHrfQPefDzaHjS99OBUCh4jyzSOZUFNr4xjQiUEVONDUiouTEHVNlxgcb0ZX
ZmA3du9GOwFYXsDA3tOkjE6gEZFwmGzJV0LyeL5IQA6/I0Mo856GNRYbW8NQWf46qBcUebnfBnbx
7IzmfZDAaHVfC2+07iDFSg7FzVX2HYykHmVaukVPoySZZQnXxGZomoLu64fyPxlGhPWVLpmY5/N6
qHsRcIxAiSmWcIDrsXQkqj3H4C0Qj8h1L3m/OnTU8gejLR4Eonz8gpGvg/mI5WkRRS9qqvn7D6nA
pFvSphWmHUdNJTqvb1CBrILF2UwUPRRMlbtybNDf9es2TtfjyIDhKNdyzlVAV6QDHIj2xflYvEsw
IlLnsZnPYdxC61iJPjEw6ztPRZVJnfX/qqn/nH05RtZ2ThGboBBKfsQXZFA80zGIN/ivamOy2ve8
RPm10BU7y2gyqoov9YbQ2gNEJvy8bf6LaXxX1VB9xouy7gcqLof8UdDwQcwiixI3DZE1+IDs9Jsv
/tsi0b/BXZYwaTr/kCgrklOHZ6iQSP5f/HpMrsh7qUBKxBeeP5riN0GoXMHi7T9jBywYkrjMdbAs
a+PbZobXJhNbaWyTePHHEY8BXo0L3K4q2cQ7u540O7/v3+pnIgg9GAcZFreKh32IeWR3Mj1zcHCt
ST47PzDGBYI8WA6Hb7CgOciWXolcRMpsbnU13hGRjvh4FSg05BWqqiY5cmAj0oO+7FGpCcRuocMT
KvpAX8jTxEQj/nedmCzFZWMR85gzxPnhYun3uvEHpRe7xk02/BYRDj0gFkDU1O4tv2LRzGNU80M8
GI+yVJ0Ywp2Ot+drKtjz2IyWjYZSL9is+P1BTk4xSmQtw8Q5haa0a/CeYBqWTYxf6eygynh+oBJn
lzUabEmHJrZFOZUirubP5JzOeFQE62IqUt/1Vs0pGjOJjq4Aa/somsBM2ijWb/ckUi2RD/KU/bFY
45W2jLwIg7G+6J69KBMoBPDAFWSlY3sNngEFM4kxUouxfHktjyOKUmZv19w/pVTvMO8gsB9Tmbdd
4/0bwtoVX4N+cHaRQumEQ3pvckicREgPjzg4p7ZBTDPFm7GrSAs97Nwvuhp47UAWO4dbPTu1TAy5
YI7qp2Hi+sa0jEyZ1wFoYS/CHouZDrDNzfqNYR32foojBotQnLGge2RsNvoWDcqi29f4yTutso5N
QBpB9ENJaf/YjLO5DSbtzMTt6C2EW60M0U6ZzeKmPV1gdVFN8hN5WWyG/LCIz5ntZUmFsKRc4/XD
yBo1ThY2ImSgEa+HPuMn0hwtqBUtnuSsr6pbYoviyWCSxU3M9qHXhhaBGk5FdFw4QJ0Vp1S2bc7K
GzKr/UR9WFbL5+nxHdQ80uVoSq4Psek1HZ+4hEdhtkguw+2KQepQ+aVxq2WCDcLdkC87M+EgokTW
n62zdnXulMK1BPzLwdXKXB2wEOIusw/N8ZusO2JeFoOMzjsMcbitnUlACWqV66izAeQozL+Cxaza
rT2tWVcBgIkgqEMfaLcE4kcXcv6vRhZO14lcMAchuHY5g+W/Kdg09zbOeYDg3npN3ukZCP64g7jT
Ol1OL097CfL34oBx4Zyhy7ZG3XUC+0Xx97kHA59lhyr9M5dLoeg98UZcQsPgYqJn2yAjeYjIwVM2
NONMwI2ZQ+vU3kK+Oi7dEIQWUA9RW0yZhJU1euvq6uusb4H9n6N0PlNvuEFzRNMAaA2pithB/02t
WXoyMEodZfcpCkAohyCX0sLVIybW8mjoqXOzD8I4pRfzY3iIN0pmbs71Z6uac8ggyj7Y5Xx+xajN
RKo6op5BBZvGd4uge2Juz99Az0ulXWV3bMxvd/AAm4o1+Nat7HdiTaZ4FhSUicqYkqTzRwHiiKnu
bbeX5pKfYaoxzgAo1IR+pcS/siDro0YrQYL8i5G8BJMuMoNU8IPyiYzvGLR9w6QRUZQYy3C5syfS
pmgiGjgS/X0xt9bq9M1Zm/OwaH5he+X9jovxYs32R+rY1fD1Kq3HuQtnzd7Ybfy3LZU9FaZgNSrX
JiQFY1QxgIuw77Ut/uWJ8xbFQrZhQ+2b/WA1Cw7sfnRdvQAvzwdapRQuFtOhMjTBNXgOBb3//l1S
qO6JTPmg6C968mmcCIHisG7M9Sy/nFcgFqN6+gLDkK6ACYr2X19XykCL/y3ojXvM7MtL5NwraySX
3OibxP7ImiiKg/95V0OmOjg4HiNFqHEZeCXwKzxfYs2kPfpGex4/7UF2DLPCRrUsBBYqL6y1yrWl
/nRskyZRuK03qZ/An+BKkVpkqeB6rPeEi7V6ae/Wr5fDeIYwofi9nE5GO/0SqNaR+oK3YcPIWWQU
Qy5JX5e7c4uJ0ola699CYwr/FUzz5SFcW0lFLLalATeAUWBJXHXVSIkgZWrZejsXyhCap3k1/1DT
niKjlX7eOK44CMGGa/wXLpaHxKg25buW1ou0pXo+IixAQx4k+7mJpfyWAChiMcMPn0+NFZR+PoOS
5D2iLfNd3rnliko2MNIdE9lIT9JoBDxFRjDNy2zEYBYPCMcJ+vWr9DzOcqDT01PeLpwIoTAXKOGO
XN+SRhT9QV4pjB899DqT3i84WQH5+XkkEfr/dkrJ71eSTkBsHV9s6LorQ3b5RO+AxgX9uNP+Br2n
qI4XpNf6nYSjzQE2DY8GmBYfyuwZxj3QthPP/eUnpdqYPL6K1amRT1pUFBNpwKtQc6gdNG070Qor
7XaZPAadFk+7r7rBj3T4wuWvqBYRK20WXOboEh8uU4sPM4GeUL8ZX24x7shOH0SzO6C22tcfsXWV
fgszxDRGsWMztMbKuFOz0ydDCh9LWLBLGobDsvOe4bdQluNFCP6ewzAeEK0wPKiQH8mk5L/5eDKH
U8tASJY2CVTE8cd5xTUc3xrF7nhbkqM7VhIAkDBrBfb6yBR6/sNGHM7UWUBzqpSokKFU1iCCEsH/
gFEJ8wFZsHvlV3wbMZ3rx574qYjcj5I/osaq9O0Sy9v60cmMyE+emJ1Yo+gD6bzb5HhhdJRn74m9
eHmVjbiaLsG1X7caRddDR105uyD3JSEcTV2iTLFwN9dowFUeSPL/0o7sJt994Wpmbzx7fvve3NEi
ifjFmWP8rfkY1A3+gVs0NcKXAK+Tlkyzz1ErI19lKPBlGPxP8bSxP6K+qxTGWMgeli3GymeFD5cv
Gda97dxIRJkmKYHIRCsZr5p1M6THgwoqQd9tJIeC9+gMxt1WaBh2UlTTnBus60JytbzsFxhyIBBr
GZCQuyr2PUGVCdxUxM2b8hvTzaTuBQ/SkXk7lCK8E8vj4QVr7xktyXPg/lYIow463ff/kbOu4eQc
DgYyGcgs7AIP71Yj9IikD+MhLDIf/lxFdr0ufnEp/LK8h9MMmC/YJfgoOubsl0FiLz2ZL2I4D0tg
O1Xs2A9BM6/oJCqNf+4JUTU0JzWSV0vjdQRAz4UOeolGAQGxmA5M0l7v/uwWKxYRdyW0WLfm3dps
vT8zRKZKFqBBK/32JMPXBtOR2RKemC8yrSFWS0f59cri/Uw6kzl2Th1llRmkEX9K+ut9oKy0MndM
iw8Tt04xFuISKnI+jHWJ6G4v2t+cTYylge54DHaT73OhgF+1Ec+TGHU9rdciUz+JGcAiUYFMjB8K
B/UOult8Z53DFusyTvhnrDPeda3Nq2zQn7pzdWCYKWCRoLAu9lWXQtFLtKd15+PSC83gW/WP5CWd
E+K8PSxwIIG8PUAB5wiAZddkUjZqDIIhDztbQZrBHTL0h/XcKHzBxAm556V8RZsmOgU7if4Z0eEL
JeD1vQQTJnPj96qY4oWXx3uYP+0faalqWwNtgUzA3iUi/AM7oWJMaaPn9Dwbs/s/F6ojVF4QdZXA
IwHOmn+BkMEG4j4OtfI+8owXMkcT6fX1/MVs9ZUzACrvRQfxDIiQEch4mMPddXjiKfWU1lDRfn1+
QD3zncxUuZzjQ3star5EkJvsB9S2BYHJlYuLjbrI8dIdE9s2bTjNYR9TV0u7kA7IEW8H5RAsSubR
lLApm+/xga/p86ssokkSRPUV1+OhZhXXKBUZbqjWSXA9RWPSis477VMeDtfOiCcqdde4mB6fh7vz
fiY/+C+S5xChKHS3tL7O5edVXHdn6MWHw46R84FZpehsi55VV8qBS1qqMMqL8zLMxeTMn4u+51bW
s660ON/sXjBmS2QV0Epd122hnFjUmwe7LZN/rEKyksl21RYEWRvxd9Ya51dJUSeC71CqnvW9yb1X
NotHPE5XPcJltTfYFWBBeGQWgR9TtvkuLVWVjD4AziTOxWJrisM1hXGR901wRTQ9CyjDUOnO85Ko
IM5GErNhxDYJJEDkG8qcaOJ1a1fmQgAGXzHfXp1dF7HnD9DEYXOvEzWYTOw+ZpYV2rnllGdtr9cX
/XBQjZPVGV6tYJeKZDSqdfGZUjhtY5Fu8pu42tHf8m1HIGMliaMm63ngnRSPk0xx85whUK7zv6Zc
sjfYgbnXzYiAIKdt0gmC3zfVphE/b5iGO+bot4+93Tl7Rvdiv97XJsqqDRQpUXz76HnQTpN7/5gL
FEYMh1LfY4pUoxhvsfY17jZHcd7fteLcQx611DAEwXAtpuX35cxyktRqdPm/yRNTu3EgvBt/isib
/THazydcEbs=
`protect end_protected

