

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fPF16TcpNgM9dNC6nyb4WjUK+7bY8P+I62AEEiiM/KOMhIKuPOHBoWeWL2UjxSNO68WLeYIZp8lA
I7rHN/CieA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E6OKJxjnDRUVVFwAhrQMAtoyRVVpuMKsXlca4m9CcIt6QI8vnYN0tf7gH3uVuxZ90322B7kUeFw5
Pu0UeqAoBaSyysHuDqXazxHy7oyk4BIWChvcrp7LULlVLcL76obtSwsXi1ORVmpdTi5b+AcD+WUo
OP1PSFj5jpodG+LwXm4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x+agogSsgbiI6PGyBpMY8RQCDzLctIr3EaG23mH5kJHlNmNKNolnP54yJ8Y7nIFi6yl6tlyOLMoF
/kxU0pyFmIj8QM0/MArMxPTiemXbDLS2VKtonyK9dDH7VbjFnRWwzK0Ngkas0+nbW3TqGPAY98x3
251QPjQoZCw3A7W9PDc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KNs7hA49BKKrboRSEkqIGldOa3ndCnhjRkSn8lL1xFfKUn+p+Wbc09ogKV6YYnPU/RaF1LbzyoE4
udPSNea4bST+08IjO5GAxXqUugcig44J+hzpGKmh7oO0TuyNbYq1CnYcsZXaD9vsmNYz8fBDoW2S
VK/mYa21mBKTOuTdQ1yp3wi73aJ1G9N6Ngt7ovDUrjyd5oNxxNlvWU8JkJDinbEnci0qjZ3Wu9Wg
y44pHUXf6xqwFYJpZ1ZcGRKl83P8p74+pLzt19lw9TPlTfKI++IowVjb6wo36ztNDJS0QjQE5Riv
hwbPU/Bt3S82MVCY5NAA6bKC/8NnoWMbmX8Wiw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QaRubtGbYrmCghuFdQuTgTEtoVYYLcPnD5z0C7mo18fwCG17qy0y8mj8xWiwE6bo49IP1/JXSIw7
rTBwHFOVrmbm926sWNrF1r3IHB83C5cstprQ1om7vnkw9XX87SjkscphhkrHmi08jjzW4qX96m61
/ymclz5TlAocMQJGz/jwscvIMOrrbuH4SkWQOLQnRfx9GIOv5Y7PM+w/wuDSeFXsAXz7Ahq3/qmU
cylNfSufW7/zfN4RZB4u+d28AXsuFe03aSF1dpW+uBK1xtNZccvj9h9NMN0cuwxt8ZUlLJw8l6e2
hqRfTTZl1F4qnnrJu6w8h8uEGrmgnQG1AW0epg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XXj6Nc59BeA5Kznlx14IKravf7ohERw7h0fbO7pT7/HsiPDCWh2DlTGpFUcnbNZslPN2RfE0nJNX
WMzLQtaHK4Bm6kxY71OsXEKm7MAIjEdLwOMtJTtlZrbm7chBbSxcW6sjWvI36jk5De3Yct9Ao1py
DpQ9NICUtRTwGG8SAiRkAXRh2Jv3rKvnookQrlVxIkNRSBMSgbwuTbq1ze/KMUZebBWwJNUVIC9r
RV/i9wjYXBOeCCUk+cGDC5uSpwdLXYV9ZxhQUU6C1ufAaK2m4OIUeBqPc2ski2O0qQYQ67c35k50
ynO8H9PTEROPEOn5c37S7feU+36OcOOAsVBTBA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
QdGxYUSiWvN1mzXojHT6B9BSHgsclxT9rty+sSaCM49qL0PUAJTO2e5GMe5UhWHncxIQsh7KK+kY
BpesTyVW3SncOu3vc/BAC+WBvX8TLX+ZCJ/85qy9SDCwEyPuMVHrUADK9QZP513sLO1ZvvrRbBXs
i6QD4M9f/wh+YC7wm7nWB/7ptwjaYWKfM4s1GwzDULKEacYE3m8v+ssqOgzlFd4BNxdvy08a4RH5
0/1UL9sly0f3hFCeWWUx4lv4zDtS0JmP+mRFBxsCNwCDqpfdmy3U0zTP0/Hh/8MPul9UP2jzI4po
4OBHgX+rNgC6WBqoT2J1jE14/p6GzR1G8dQfMYo5vg2UrH1BX8MzOmrNoe31j6p8WxR9U47fxC5w
HyGH9g4GBUOJ/qQ0fgK4xLKQnuFoQcpm9QWEhA1LIxOOCYEu1ETvsJwyENDnaFQ+9p98/dYe3HuJ
kQycxi5Z3vHZRBREFgls0nDGs2wwggpMbFKzVhVaMf5kMXaepJkVZfiwbfm5u7SvGRcsvJt+TZaq
XXWvIDiWeBv6MC9d4Ugf/KMeganlZxKKQESAjajVG4cTZ1bh7XI6lbB5vHlm9x3OR2MTmTZ+lCx6
eRnhISihrANaulFhp3HVLNafmNWxtjjFjFP2qy8hqC59xXOD0jM8KIeU0HQ+IAHq050SEmON6HQh
lvnu+EIxRu8qLFvoByrkfuUBDf9pTtyhiUtPifveAMAYSsKQrvs5ZFYetkG10ovcaMEOPZF8j9ag
hVXbjq6KEb5jIzq/3gGmO/+XD+YPsqMgCHWcy3PpEyb4IOc/aSRCXN89dhui63/8JrkLwvWDidJP
r8huPVYaNEBisEfkVnehrQf98uXUfyV5AVmNmspCFf6FcC/Q+SPOY7cK9D8pWAn9dCGt4KzkMCQV
m8ZEHBZjLSGeQ6W5Su3vzsxxSGkHtHsDNOexYmmlu8MR8mS5v2BpSl3dJ32nPX0mVvnkgQD+ublA
RgRYl6lYLAR/ZJaqp8JhIdpdKzrkzFU/1+6uFH48Wb2JWJwFxzFbaAsJCvkLUVGkqAe7GusaePrV
KyDk1pSqXiYLxQabVv4odXBnwk3//4CCz/14ONV6T0QmG+vI3mc3mSJ2BdeVGzgNLPkPSVyYD5Sb
o354wIc/EOSvTYxJHLOAxMF5mNwKuzh+fY7e60g5GsEEEjYrmkSyIO/wbn++IpV2JirKkFGNXeuB
7YaXXWBrMZBGLisQSc9hUzbvFQ+3bYpucyjCR/4KkOrzL5YZNVca154zjJTcARrB6MwyvEqhMaTT
LuVOAzaP+N2uMrqLLyF3IPhJ9WoJOiUImt43DwDBkXlEEVQHpn+wlza9vQT/Or3Otsznx+sR+Y+g
EzpbKRIfc94zxHXuDS4celXv/nAmqeNVNHRxpZVs8CbEMdloq16lKo+DrI6uXawdXaADIAnu27hj
KEpfGQhxG1jEedp+mWiz63uns600zhAdvdnE9nnlwJ6Ym1pjQf9fR57vI0O7OcwY5ZyAgw3eWmA/
oO3cKFU0lpH7O1IA3SRwPjoSoJS4LOZtM1lTSS6LyWDiVw3qBMLhKY1cjIC/7Wq+XQoDDFtDNGMC
0f7yyt60hYzTXged9AkaWjljl/bMzvIgq4FqHDu3xuEagndqEWj5XyGjaFN0ksL0oO6zbEEj/c1E
JEUpA8orNOFqVVGrXPweRHm8FKpAe7sKrrMq+vcN6CdNvnClY0pj7oljyPB68Vn16wIL/Bs6RH2l
GH4Lf5ceyc+FUo+18i8tiLwfRjbmrNoh+9OlqlSFkM794uQNbhl9hsiuYch9F127OaqQbG5ZIIUM
836/QNicJkKB8SvVCfNRIkIejg9vKnmfvUGYERxPvZ9KDPtgA4rgTaH4UOzVafzEyRK523ESJ1/r
B6naCrMWi+igknJ6Q+Aly0IHQHdufJP8Xkv5qBO/lfqXOfQHDD9gRr/WtLLI4WtaAcTwDSA1/VxN
JudJGs/rNSZns4r09q7gqd3fAuxSIAiMrbeK8UuOAFqIsQ9lWNCasb5kZnrRniyqS9da2j3rNM2k
u8mID2e4ryoVKumMX3kThZBn0nRI6uJPlbEk/L1e9XDc9en97ak1ppc/BTC8HrKzA/JhtqfUEMaD
aY/dtcp/48PA0FUYJHtBjhPMSaCSZ3OBvKzL2Qx2dCbQ9TK5X7FlgjOc0cm21pAQPevD78f1VJpf
Y2LH97e+rOxVYE2EssfowwgIdcCwxbTkl5xx5LPOpwPtgkp2HegwhIRbFCzJouTiiy4Rw0bFzlbT
PBqFdV/Iu8W69eW+qhjq5hVIudzFfzi+kOoCoTsKw+HfRC1ag57cnfPuRjK45VQjJ/2F/We47miu
6QvCTxdahff2ro4WOqx7H7mT2jMGeKHNQg5g2ZNLS1lf4A1BLqBqtTZRCZ1OXPuQNHvfWPHpZxnF
Do0J0lwBkfIEEQLDYuCOJXYriU+3s54y68arrVOfYyhl/TwxvsEAp5xTP9Q34A7NzB2SvppoFqa0
3C/5XyZcIqJeAl0m4nM3u4PscfXSWABedJMPuQ+6WQKAOMasdPIo0K+A3g3EKxgmHUVZRXqEVzRu
MhHXVlMGPduMs+mdJYmztf0k/gKnwOfR7BqFblLxz/F0w9GgnEuaEATQzroEYgXjbJqF/Z8i6D81
Knds8d4bk3P2vvy30NVAtLwFeYQJdM6hTYPFBSkUium8rZutJBh5fvd84AazvyJ9+hyynN4Sjnt0
J53ulLZFEODKg/wkk9cT/t24yiXOmGJglkYR4OJhmP+r1vIJ94gcaHhjHNfN6qCr9w2uuWyJ8xLt
A25AmZvsHiA7sh2MOfVc3TOn9nxP2T0jr54zOuyZYqzgwmh1jAn1sEyO/JSjVdkUgioXvLoJhmTN
kW4caEAu0TFyG6AbhlSNVmr6Fn668yQZBLcVwV7OId4ZbQFcCNtGF8JxW95GF/9mwOqfTDAzQDe4
Y12strck2qhBkXCXbVv9120kt6ZzM7EOpLBobVq8+6XRFzbg7wiR+2eTax9yiXFSilVpbhRdjr5C
XSG4IEzSYOXv+gEZCpdStZJ/nug/DNxjUa/m08U1EVpI1yyjtNUO4ZgHBBd3b/w/VK6mxbs1AXl7
bDcD2F8Qparrl+R9kVv3oL0iPbiyZ32OuKuCqpBhUqKpFjFIaMe5f5P6PqtUnLsyh+vKb2blWSAv
aU21s4bOuypjr09tzAboDFr7uSMvSUzxm0ykQ9Q/I+sTJQk1QLTmdZQrhVb+ePUW90hlSBWe0V7b
MUphCcUH2+uj+s9xpVsAapfmtWoqo60Qkin6rRuMTSqirXPIqpz0KoLYXsGS8T5dO+qEsln5nKvO
wqrAqlB5xKvaSvahsvV9/JDu4I14eG69rRzVNebbiH/Dc2HBridjjXPf9OhxyR9T5KnFpDUu6m/b
xMRkoc7w6wueK/Jj3eap/5wPy2D4bo6WTAcrL+uaVct4WsiDskNe8UBu3vCJjZKzSi9cMJkDia70
YR2aZQgtorP0VXPAewIDJqk8CuAElKOtuHQN5xGw7bpA8V7bc383fQJ+6ecHe+CyCfTb/C/Xok9t
wfoEeqGOQc/MtZqUn5Bh29kRZowMBl38VxRIMWu3WYFD8KggpVeR0aSFdELTG9stxh4b1EnkFkSk
Jn0+NAXpMDIS3JwlAw2+k2st35ewqMVHz/eYBfuvp5HMqarCwNcf6c/3fvbHbehba8mV8rO/UpSi
tZzZnrNhpHyQbbIIGmnhiOn5cb9Hq1lyhyBlnLYB88/64Xu7JVdmr79ruofJOZIllVwWfGHrHCho
dvDAd0qQEReumyeABCGzXicLnlIy7Gy6rtL1st19DK/u/S79LZDe4b2IB7GvWkFSut5Lcbvptwt3
Oi8USpgLpvqiqlO3Na22lB4aOhs/Vz8uBbKQoV9kDNP/XkFxrBbJrYjQ5JtaznNK4Cjx9DlDEN48
d3IXmUGBNKOHEHi/38gnbHhjP0N0cKNVckw1kmPRxNV2rRiv82KXcCKHDUhgOS9GZdzByO7G0Jyf
e/DwpuD2bcv0twMpkYDUhhwEFprI6SUbenmTpEqYjJ3nXBk29daVe7N94t71t0J+icc0OJ/XXViH
+OSW4DCFedbiEINN1n3NpFZys5onKuK2ANxIcWLVzvsqujfi+iOx0TOrD3u7vdX1fIZM3P2hCz+q
6LdFc2wVQZBZ0B+0IgNj2chxyEs7yFru6l3EY/d0upwkL4aSpS1Jnd8dietQvDd+OLZ45AnWMnYq
xOe3+vaPWx3b5SGhj+eXBqrguCd+9Tpu+zL2X8rDKEYGcqj5qO4DeoTGAsYYHI/q7oSrC/aOJfZ5
54FKt2dbWSGxbxXhbcx1I59SSvjdJyI0z3iSLD8bGi3MqkbqyN3va/nzaQsyLkd+KTw+gcUS+H9j
G3CfbONhmD/Elo8iMN1CZSgQ9zTtLflj6q0z7mqwH5+NXwmypAa4931iSVG9M6apmoBe57qV9tBJ
oWi65wIDJd0MUR755Bxarewdwm1NXUCWMX5lz9ytlwW5CZq5TdPwj3YFldE1gcp/CAs/WYbmgxWo
+1UkAVdnwpOaRlmG/JzfhUD0ApECZbpTBcChGcZl2yl4qEljjhTVG5nrP4D6QVFphDwpHZ7nZJgN
FLBTCXzzpltXFdyGM20IVnK/6F2vHe8R4Z1Xk4NHKSlXOTkojggpke0feCwmwhRAFtL2D3V8531o
/unWCq7qomvAZ+RjTB+mBOK0L1N/z+sDgLy2dEK1zOIEwk0Oyg9QHJC4v1aE4+ME3YAWZnAaEh2O
Uk21SAtmeARuoWXKMfWDZr+5q7JKFzC58HNgcK9wiJxvcS77i7Uh1X2bc9B0m5o0pNjNj8kOzBWo
BuiVANlN+6Ah3AuapomQw9APXi5jrdCEFs4bPCGzXQBDNJ+u2pCKgrKDV15sp+fIiMGNrSjN7oYo
m8VxjDlGS+mjEBIBjqwK2Rs7UqU/pP/nRk57hS5kU1SjklSIj+eO8IS0nnW4F1QJ6n84bb58HY4y
Zb2FyIO0U+jpyVj8Pzu80P0SyouScmKEDoIe8bMlzrH1zRlrhtT7VDa/0hMxJDU0ql/JcE6ybkiu
QSU28sJi/lRllQeupJKPXnXOxSUUixsFeuq6sxOQrRuFDyHvT8DEXiZc4/fT2dKNdj75aG9e8hN3
z+9SWZqYJn9f85DD9rA49oJTWpi+U1Re/4VEp8EBu6RSM2xCMPIB6CRjwYw+RxjUeXldZ4lvyzNq
nz38a6ewjXBcjhs5mo52bT4Fm3OcOEef6pnGedhyJ0SsX+hH9bmH7yblG1pw4iMiPg1+lA+OPHBa
iJIo+xUwwvHcXdXOPpB79qfiw4tzue75SqDofliM3dFmUqhosqtEiF8ax2+V67FRvhEK1n42Wg2s
Mtp00n2By7Z62f8klkRslD3DYcqjJG77z1fVgcc4rFvJde1ImgSQpW3gZAltI/FHBLnZ/7b9tZ9+
D4i2jsemTu2eUjO0y9IYceHaJDjglM/q0xCCm7NXUV5eQZKXxanpx6kOeOf4Zx7zK2xs/Uq6Y/b+
Ngd/Ui0V52lsYwaamLV3bgujFTrDfR4mla1YArsgaJqmuCl1mxKYjHc2M0Em+TSkPEgMRORpTPcF
1CVz/eV7o79LrOmO5qIcrPKDf6MssacFwNKwdpRPRqVTrHnw4z8p424HETsA+AWG+rZZU77X9M15
q9z5leQYApRxX8ce05HTzXXoYzD64N4s/iWQrjcV2prD7XZ+mwEOlFOLiuIrxLxL20aMIZOMLhZn
tDt9ULr/D+Niylvnztx7E2n0PIGGq7Z9lRrpUyBBJv278xHHP6Ap3P4sFwQYdx2GTlRCGO7TRZq8
cWi/wn0SLJzvyuhl8hjgZkHuIunHnSwCALC5Pop8bVCH3L6JWSBd+DNeCwnErFE0H8d0C3H6Kw+O
eN7j4EXu+waOwb91/tXu6TA3EcXyTqrEktaehlEQ/jt3zJsO3IvGAiaAKj6BtHoed/9ShCMyfyX7
pfS0Cac769djH1uaspD8IvpBlKoHw7UqZyROfKnAdEstgfGHcciHyl3DwUG3aJt/Tv+5X6DnzxZF
dW5KLu6zq0yBSWzAuy5yaHkOk1m1HOWA6GbSKtXwRBO6pRAGX6jypn7JSXfHgSAPQNhmCcoZpzp6
SPgBB19Z0b81nWZ+QMBYg5gS3vrPmHaVwvjUP6VwGypC6ema0ZlSOFelByLOoOOJL0sG996FiTOn
6jU4DyJcKqC4oba44L7n9J90Qh+dqLB1aXoMzrpS6E+eNRzgQVldOSV9HJx8z11O2ZrXOCmDNLrE
PSXOV9J/5b6cyopNWiVH+v5YOGVCbRQTmQv2q+4lnbEzOvK7pp7yswLzwZugWp98mKrYj3GUtAPv
50OtIZUB2Z+6o+vN6jwgkMkOy9sOPoc+HYdIOe8oL9lBUd0rWHGsKksD9l2YJM3cUo+5iwZnbH75
jOsWNlItwupZ7POFBm9AuWQz9KT/NwbniZYs4l6/z/6IHKSu+7O4m+MCqzEocFrx24j18dngdjkW
4VtU9HANcnayTTfWoGezbDhHGmsZBtQhMvE/R3gBdAbKi+/VUm++Bqn3n1ctSR0dSpywjtcHcvwY
vvXduXxCaQwUrTlWdU7v1+q7sKogbOICNBTTWdTocm/r5AL00VLaNjMFluerZ9cZdy+m1W/aSL/o
C/lXxV8MnN4gkkoBgzrtXQeaj2jRI5f4PNFukzK3cDP08Blj6I/5J9otG4htmpU4LOnfDAmsHP4e
Kia84esiyQDf55ixug+Z3eGt0YElC09+cZq/aP0RAbsou2omu5fAP2adwcvIP2GvcRzlj0kejR8j
8BMf415oqg0hJknRFl16PSLCuL+UhvRmbVj0rez3S29S0Ryl7BHvvm/+PyV7JYhnbIKCeCW7Bt85
Grf6hkJgTcVCDs3QdYxYxjaNB1tkaC5PtIMP+WCc0s0r2DUMtHuRZxqK3bjfP/fp2IoceboYymtC
9AvS9o5uLksa92LXXqTwZxyyDggy2gQPY/Iu2uaDToyOtl8kDejzJfUU5DvmnCtOAfvk2kvyE8A9
3vnzPn7KkxBiVxJX/26jH013U1ZB09Ikb+BEJBLZ8F8Ycymxj3c7lZTmBKnayv6OBho/lhArGgGn
PnNXllzKrc8hJuW33jHr3fGnqCaUwq4xQGE/J4SWta3BFJDLNhcUgUIotqu5gLL85jvJ8W5g2opU
LeN0Llh2OOUCfsy63Qhfd35hyCMp2XR6Kc2AmNiTfTvaDNG6YxYkbuQMCb5Wi508FQglXDuxXyoN
5rLsQx4wZkNnQTHfy3osA6+hN9PnPGist55jsZ6luwPYbWLUMG2CWgA2fwfEo1sLAH1jHVUwiKHS
Z2wbbcvQ8oWvXiRwqKyOtTkqhx6CrRLrcFtEyXugclaZsydA1m9OFNiXZIMcVbZOUNFdnvii+4dr
EW6XUo0LScEbp/YbDYNGl7SsFNzA9X3jgIwUj8reYp9n6kSJn7NvjFElbVK5SS6RZG8Uq5ZzBDdf
dvUVZrLedZ7AB1UEQNlIautlrna1XKEDlTXYgyTGMTlSozWewTrSwzTlUnGlgSJoAf8hYdR2c9Lk
uxSDw1x6z5OIfpsbKehrvvh+sAZ7j0dQKk5oYef7ehjyoz54pbo6vJPtdmZu4K2rQwTrwpVDTiEf
GipmT13h6MhE6XAOAMWoPgmRlqfsA69j3OTrP0xaCQQ3CuTDHR8sc70tpD6D3PZ8+CzNUv0wQLVv
W9sMD6agiDZtXJyYE6Pqf7EjUAT+9kjiZRoQCm8SoLmDJUIcDVqvUHtLOrxrvWtWWYYVjyizXBhO
Y4rJzmCMp/FijM0eMzKZ/S7YijNtkb1d8NCZHoKPwnj7QLm0PF26y9B/mseyfU9MmvYIE8X+wrsq
wUcyPl6yTZEaE1FlPKlExSLF8BpaxW44nq6uzyIgH3McCCQqvJBvjQbTF3eUHBgsLT4cQZ9zDjgw
RPWblqQgPp71o2PFyPPUE5/NKi2pcIlu3hEH1gJlX9V2u/e/Mh6+fGAgqD7tSKCvW5mkLdmJvc1K
owQCVT2pmTurPslcSae8AnGnt/cJqYkpfVR/34pyvJaTrkiAtYcKnTLEj34QNHAzQF6JgFRByz4T
CTHFIm0fq/FNO33sDPUaHaiifTEoI5eKxWBv+5pJVztuOa6N1J3txVNiSjJ/pMXh159jsjqW3yuI
Y0dRY4S9akFTWr6EjvpNz1AtRzgW7CD412w6O3CC2TEC8MGEl2qtlz4/HyALtkfwtFbtWCCq4Qsu
EgPYS8vl1k5D0TtfXw6yUFSB+5+7Z0YrZ0O4ujzb/jzU+Wbszk/jPj49BSYuF5wCsE8nt0OUG5Bt
yvv+K8MtseLjNpc2piAOLxBpHOTeil3/YIe+s40zuWFGlujN/xIxXy+rbLT6UBt4+BDKZCyBfBIU
mpBS69JMIz+iUPOyeloDLDNUETU8QuzhbqOB+EpNJSGvlgUCUhERyTpBTd+sud2oLInP6T/JYNBs
NBcVmvWfEBhEmlbD+IPLRHkmk7v+8h0NOxIINF1b59Q6Nr9T5Ur628ocU8I+9SLhL5WoQaGPF1EA
mXo/PvLrnscWhtN1c8140ujFppfzGkLkdtDNc46SWaG240HxkdtoVm0Xo/wc8A/JkKFtOuB4MRL3
gRqvy5cFsy+W//k1A62nJ3AGPuL4IyzzFYTwheDKLdrzShOC2aB2TZilbCJxnnpLkwKQz6oLTFss
yat/ETo9OSEMGmSreSd6UEk4aB0X7onoKPcyGaJI+TZrJIZuEM0tJtBH7rZhbqPQXMymmAeLcBUc
MFscLDzJqaRHEPNKtgTeJKOMqM1ffbnfhBVukKwz0RtbseqRF2zaPwVhv8kkjnJiDS+yOcN/Tk7Y
A/CEh7q0VCAjFFABcfaTRXgPAvKEpyj8oUTiPqLA43N4IM6APlSLeYLb974CLD3Z8/eCDAqPQnDp
vkKQyx7kwBuqDwDXttL98aE2/tWPpmIx/MnQgHXoAQoqiFy7+oRadSEFTaPEizwlI22qOV72s4yA
ywoJRDw8Hhzqh8b7yANINRNPqPemEi84c3LLdIOpP7E9hAeVSgqvpe2Yva/rs43N4bptxP5OmxHV
knNpE0/GzS4fS1e48keq8p25MDFsPx5MCfnwuFA2U6ua/hoT/YISQSfJR77RHToUpv95azjS3Y6M
GhGsrdxbw3HeV483j0oEn3+gMoqGc5UrvTbXtQfXUUhbATolbx2emx/0wvELQaAQH2PDvJu6zQ1D
AlYJfDKKROhdD7cV3dtQU5yd450W1CzLXQbfd+ZwJST6MyLipflCYSg7oErIylydK2fDFUPCmlOb
3NB6gTd3hqbi00WzGEklcQc1cCKmyIgmcpKiotn4xl25rzb98v4wpxbB+JPO2a+twnsDsuTJhIGU
yuK9TjDlFQ5B0Y4LO7av9K4w6777MQXtJ1O2vpsgyruKoXWUz8eYnLSdkzZdUPgeiQiWpIgzhSz/
8/CYUXCzlqjM0o+SfEr7oYe8/zd3ZWk/bFkyPLBHFCJ60MKyEzfU+ufS7gBLh3epxqI8pAbru1l/
qDfzRRS+mfMQW+O7L/tQ2NMlFpqoOKonkmDnnQJgbuZtfZevo7QxbFqA8tOJDafefpIyOkTEVcdR
ViomFZmb68KOXyhOjWWQ2V0DnVqJAzIIH2w8qaqSHY3v3jMtY5UyVcDipHypCCnGec08AlyrglXo
w7IU3XQ4cre2AGAjE6bUON9MEGKoqJPLNW/iJW3GYxEOUvEOx9vdZYUfyZylh8RezRR5qrAW31yj
3vpEmGr0S9Lu7NdyuVW/rmA38LRX6fN7DDk6er87AmI/iutgqThFdoy6wqohpR/YaHdABojFVAQB
B/aS/LYIcvlSFf2kzKvxcvGWJhdefvIAg5/LuYH2bTxKYr7gnROVBW95pBS2OYZwpJ1c/EUv2tKh
8pc16AEN3WmZOlGR1+oMpSZeGwV31IpzQb3F7F8VZo33WBnR64eNk05GKivnX92V9esYzPiqyC7V
PscwN0Y3AahA9KMs3GPHx1VZQpiD6u3roS6L9utagoFXNTNCAIv+8wbj7hCTaL92cTy8Qf2E9kN7
YqsaF/epJsWyuj0WxdK5rE1UHMzMF2+Grf/fXeHN59E4Bh69TpIYsGWIXK1a75oQ9Kou5HiI5NXq
DewU6Hmv/UeYJiybQ0yHA+wxBC71Ktvi7r96Otdiq2la+d7r3zY8lC2thlnYvzz8ggzhX/6jVKAP
EHYxU1Yf9Y+qqAdN9kUxETjECMmF9cM46mle2AKAfmKtlIYs7cKG/JkvtJ4z9KUWubtJszFqNzwy
SKYdRVY9nrwpR+AEJ2aUJlBCxYPHfgpsI1EixsTnO4RB3PIXiV7MD+P47wZWFYGjBc2FmUDWgkcy
vGf+pH/jMYhReKnNgrK2PZn3o1TfBP/WO/zlGnCAFy9SrgGObpjlnDN6LmwmIjYcgfi28a4Mcqfr
NE6kWB6XuMCtFvLwiJTkvcWbRzJffYeQz2j0zTfsMgVrZda0p3/S66o5gyIM8c7dlD1uuyO8eOhO
XII3iLSfrpkYRPqLmD3vON+eDMf2Yzx51t1KHxE/vl/Up/BIrJZ9WQYcGXMIAEu8Hks2Rf1hl+8h
y73k3sG8dk1Ot83e1pCTH0dORmHg2zf4XtqnnpUXZX2vjjWKwdrUn0cz9vZnaQJKqyIaYeYdUqzy
aRpXP0G67IoWqyWXg5d4iGQsFhKyQKbGy04r0ueOGxyv961PC+4nJ3akLKQCeSqOiGk7HqrG9jfy
qxlsbkXud4VAmI6pDYsvhdTyf1XKZQB1ht/YvoJ2seU/46aqbBORJ9EfR+UeXdYaq435pRLLmu4l
lQ7H2zkebtCko0r/hJH/qTlBwiew4OVg8GsPej8oU7uzmqwIhGcMBwIiDJKqvrLiLdA16gQOUR19
/ShQ/5sIau8l2UqnVz5ff2AMwACMBpTHOCXjjmWQ4HUGtoOI/objg27XwS8XPBRGoP/6lv1xV/Qm
y+jt8QJrG2Hrk21GpYQCsaWByt/yIx3pMFQMMXjYVacvNk4rILLXQzD41LZYbL1kDwv3LZsIhErh
gDANADaSktm/NSqt2wcWREKyxQMcqsQ1WiaubhVfXLIaRTMcbzo14/cviC5FWInQKyiPwXCZSykR
hQDJIO+sNSRB4yWsl58CtaTLm5GGmrZ3Suugyk1COmPkDNn5AxadXlyZHjpYmlYcUiwKL4DVfNjp
D+lB6CVcR65OMPn+kcpbZWemAcYJ19+8r9Gw5Tgnx1a64uLlJ7eyC3OehFkCP5FhULb7Zo1EGAVd
etuA2M8nKfcjyfapR8bw6FjGWKP2pShGSO45X9S62mRqoW7O8QCJmnrG9fFUZWfX8PDElh1lp5lj
WVn3I5PUhycbRvnqkg+q/iCg+8fkStBGcUkjos8VvA16BixpDTuZmvBULtFEeCeNzv/ggASrjtrj
LKk3O8fIT7WcJLUgqAACwKoLGyQGSVR/+VJQPN3imT2nH7sIQp57PJG97lG63cqFEzjTFdgLqbCC
1qYlRMi7kej2Hk70g4cX7eHXll1gpEAtr7xiLi28oh33yO+EeflQpy+lmIfS8ieTmtncya32ux4B
ysabTzHFg4CdrX7L4fCIsk16LLDnCF9ga6Abzwd5a5TtNd8w71Fhiy2OC8nj+nmEl9wuWOq1Wpn6
Y2/pswICGKXeJmB4HmdpKLnkni9PD1YCg35DWAn+LCME4HFgDQ8VXanA0XPXrSp30H1vvNMqEKsc
wpahP14pb61r0S9Ja8ws5+H85bXD8D9ysIx+FaAFjlpyDeN8ajWkdlUwDShHmr7Q95Lb9e4VLHdI
GA0ECKW/VzXLsEnTmrTuG++xLgMdUoqP96xqJ8JY9em1P5+qm68j2H0ScrC+lMXwzuCP2oPcj18i
iRId52eLhUrxG/5Tuf6R9QlJYmxxn7juiNoT9stABlMhDDsXj/PumV0iKK+DcTkUFtM45i0wYJkf
7+gEJC9rkSTaogHcQ2PLMDSegASrMHXnatbfRi1xizxLDTReA4fKCGyZCLHmNuYXJJeM4elYcPnW
Wtb8GW33F6Tr+XWI7BdTiEJQMrAHcK/v9gAhpYiic5GK+fOEOztOGlInbH4cspYR+CgxWdiwmTpX
BPzAeaEd+jRgDKBRhThA9MaaJP0yRao5fh8u7aad8EnE5o24fAfMH0EX5Pqlu2rEQNAquIN2jA+/
XjHSWyZ5rr32UX+80I7gqiRCZoJBtKVarsLBNGcyQEKID5UzCx1/WaYaOvApvcSgB2xOOM+EWhAe
1xJ5t+AVHo6FNgNCoqH28rMHfskF8GPDfabiL9dg4y36Yfr3hNFc5wWIqe7O7+m5NRXPEEUOknzO
QsIxaS3SRgbU20zc8e2bpggNT+lcLoZaIM5yGjvG5K39dNg6Dx4XLvQ0uvouCywTYIOyMw42u4Zn
jdeZc5ZtCi+cfO48u3Fq8A6GrR+lNdoalEmtT2Q4GVwJDdgWTiaiSam9fgMkP3bb7WiqG1LrJsSZ
iF2fZjNiEASIFty9Db46Hxz32/c+WHD7rvH6+Liv/ELaPNQVZxiZmCrXlRFHKXV7gZ3/HThIs2VM
AlG4yk45TPSELkcisyJoYchXmcAKuXNpEfbsLjZ0tnYxfJ9XXoKNmH8OLVBqAj+Bm2FXbvSofNBO
PBFp2nL7QwfAvXJ8yFmkCWG394wBicRkENmOakO5a3E+TzsL6HZsQNK2x/MlPF+iLPLLgndxBHNi
Gi6q6Z3lpRMDfjfSyZfUQWkG7nt6YsyG0I5W4D6PDUsq4rYhNE0vGsadCM9W9pZe1Ub2JKM5zVdB
50zVQmVdxf/v92xPLAqVKwNBjJU1nyTlMjR3X6bI2KoBFY99i3RGOZyehaKEzzjidnnHLok2NfNy
DkkxzC5a2j6qvV6cM4sKhi+r7FDOL3BzNmo70b3PW0llqicP2bBWJZR598CldXdNf4kN3iLM5nXw
or3JGBtB4pkj+a052DsNwiC0vRpYLj/s5QTnkX2Iuzy5OrHVHlNNNW4/zggJVQaaHMpJJK9cISwL
iyTiWzNbFvN8jigHMF2+8+7jvdBby6vbzpfUG+yNijXeMVoFnhLgeivHst3fIz81XZaxVFMLwYdf
CY1t9y6Pqu2r1hx8SP+vJ/G7w6vIqWWlu+3P9IBgw8V1MoTHlBtxDoaLC5tunG4ZHplcEeABNnYr
6NjuoHcBbybwNyO3friP0GLaebEgD8cSLbws2HhnGCbP5n43cK5bksiaDw10QNpXPFm4mMLF1NpP
Pnqw++tMkiBXjCX+Mil71Jwx00umjW7youQtIM5fZ2edJ6XtY1h2tQdEnxns/uvwNYHNApgdVb7o
kXPoX1dlr2dtyoz9e7/v3Ht3bZgIGDUIsSPwOZuGLYZMRooL5KDyKgKlDJDEO3rG2BOo1tfzPRsO
cLY/f8xv8U+fojMz3WvyOnaEcc+2QPvCaMgdO4QJjnt1xfLC/BoWEEFaKK1Cc6hNKYi2gUMlt1Hz
aPd0bpnwNJCoIfGPF/WyQWDNKtN0QQxyTIoejQE6LYKjMXX0n/JTCHjcOnYN31NKZh5oUBPPobBX
96EE2NWgkxUqe3ho7q3XLEVT2QBKqec2IVigvnNFp7wPLCjpvdH4MHKiemGDI2fXJzYa3v/y1DIb
9s3xVE/kDS+rtTF6TB9pdpnXfg/jBqWx+93ipyGXa6ubJsvqEJHEL3RtxCROEe1eFSmLHNbVcDgM
gkJdUGPFsfDmkGSVbghphciMNmuqHjhebrJ0h4AlBbEG1EKw0Hubjmv7+419PXl/fkFpARzTljNB
RidYRAma08q/ew1HzegugnPX1vYz3ZySWjLJZKWb50d5pnxoLfizIgq8TVs5T4+zYJ34wpNYaMN0
TZFJ5iN2H/DsGsZPo0fiGKrxF3eIpCl2yZ1uGvTba6hZOfxmySeEVU9gRIEvmTHALzyJbS6Aw1s0
68h81gUPP1bDq7A33VxzKCcG3gbsJ7st4w9sy2ZHxgsoQ4UhaNAkxBn2RMlltDBThpSEWrxVAHt5
gahyiaA2X/UpTLtIRgfh464g1fToW+yxAFvPq8DHE1oDflY7HWlB7XWkcmz586ZGKmSTAtJPTr8R
841HO463N4bqTnXF4FPaixNI+Cc01wXZUrrvQFzwAGs6foOUvDMqgKDD6wFayzdLEcmoCxQieNZS
RskKNm9bTr1PS2RXRaHotwS1W/nZjVjFAgyClsPKNChn94MOQKChHtuLRlUTTxDTqdPQhFNlAfQV
UYNSINHqcMpn5P9We5LXdj/aJ9tit2aamqOxhXAsCerd4CsM6z0t7r41/flxyVp7CUirtWcmlZ6M
gfRTXmoFQ807PxzcH9N3AkPT10abafAUFGSYQjxou3YF/e7fs/i7Rz1Tvqr9L8aSwKTMA2hdmX5D
KNz3P1+hw2Iyp9N+91sMBpwqPgQk2AIkZ6k/fgkuZNq3S+FiIsGEbGCgMovmuHcS/88NF172EFP2
N/lgPRtVkmlEyopk1uaHQnfgmYOndU5FNySoaLOBpVSVpRS/mxV1talTT/Drm8w3I3/8AWMhj2/i
PFw2PnVwRUp+ENCjcCSczQu8vUyXEYlsslafSJ63ka7LnPLPjSLfVTo7ElrlmdlY7U/tY0CmIfj3
9LURfQNgu+uZqMEI1FPbnAF6AbfeL6UF0AICJ1How+yFivzPCu8spTPOJCbAtkmq03I8SqJ57nSX
ZnURZbw3hm9iNLyXvEKSBRcoVqDZ+gWaIie093S1KCpVDD2VpCcqzGMi/OyaPlV8iPSpd/UeVUfO
qSOYbttOAqSLpi4p/FPxiHX4oP2lQV09XG3KfwYKhrsF7sCxbUuuA06KajnbpseSkFcwUlEWr2iB
+DDzHEzFsBVwEzZ6ijqBPLmdMMDgkMpnq27FsbtgFgJ//y724SFwMmjHQfpJT7oEywePT+aeCwEy
DYNoPGccDQ7vrtk75V0vx6m8FQrVk8ca7BS91p5Cy/51zSrDjUd0EiRr71rtPbLali+Yn9aCJDrP
QXMQhAtQWqnPDkbCZ2AMFYZSFCYzpfeEoDh7+t+V6pGMZCWHLTLvQ5Gv9kS9qGcl2k4iD2S46XH3
trCv/OdIocTr7xtlLVDeXrWxHAj47KMyfnmV4Baor/3uCzadXyHH9vkAlY53W3bzf9UdD2w+Q93r
rXWXpVTFx+MLW+Ghs7gLqMqSSN3vm0oOHg1CybFHueqfDvwk/3n2rHvateiKXBKjG2cJHC5rFbai
I+xkGbZEju0u4tA8JjoQFAQYT8/zKHJH5nJjCz2P5VTyh+/2+5llxBTkz7BM9QeJCzLwsm5BdXdT
ZLXbkyFiBxr1fOZYeo+1HW+9ixA7FD8apGObxq7LnKTTjx6SX2ykKPsttZM9kirFaTAuMWbAmmSS
nb3vdhn454rpADtIleq7/b/zI1xMc0lIJJg/iAY0t+507k7pZK9abxC5mvO48WKjQ7WhykpKSsAb
mncbkUcQWxK4BwECSE8snGh3R8DHAMtO32Q+QhtNTbZ/lSlhEmEVRD2twEm02dcyFw1craFPrUp9
ClfiPQR985MHibLydpdWglLIZ+gAPo3drMpTaiQv9bWTMohKbN9r1KwfKyETq5Mp1ycvmKoUFDFG
Fnu/j7YR/G5Vpaf9WwcqnE7r/F52p1gSYXkosk+Bck7Jv6iqJemuPIqzYeIIpHcyPKU6P8Z4HB0/
ZcsC4yvH3DflZysGGgvuR4TK8N1cDDf8qpyowwfGou6fTltoL1bNNKgwyDEmR1mlnn+hfOZGjnqX
5+a29LUvdbQcWUlKkqR9xm7eRd4UuXw0pFzLOYqnmYu4xVYiPOFoGXtx1+0mmVeIOLE5BZIWhJj6
mDA4kSnzM7Beg7kMDbrE1cEgZJBIRzq3EpKRVUTR4oGrZ/LsZsOLoAFefYOTxaA8ICqGrgDJz2K1
opmdNB5GffOAocP+VPp/lfCzMe18Rpicl3QlJzg3VlX2Qt6V+A4J3B4S5hC4hwYVTm9jqlRWpe73
IQbyDKi6YBsv6iNVsXLzgYzBEUPxG8nfHVKL1zxjy2wX7NZg8xLIsmJ36truZw7fruBKJm8fziY+
60Ym+y81p5DuSiYBx/10szO5W1ZP+U6OH5ruKzHhZ396vtyDaW9dIz4wkcm1WSVhHwsKfcYce8io
lKiIvuWjXfcoIhixFWsnaoWwxx+1dGVMhF+QceNJa+OFsizELK3wBKkEk2pP3PBv9WsCiurXz+ZM
9aEe024SFsATkclJh2yXcNiWAAMd5GYCtEt/+WBnIz116he3gvstPEl5nOxCU6xi1vQjACIxP3RA
zxeznkuq17p1M3xx1/yNUvPJOwnuKBtmXOtqe8swCRqXq0IQ/2O3J9QZHjfBNyOCJl2bXPhkTMDz
4i84uKM6XraHUjlCFDO5GRyuuWlNf4JCCt5H6YYq3/aC8VQEGF1TwIjRlgpTgAszbVCzeeecugU7
ZxjXKowfDu3PvGgFAf5qKH8yON26YJi2DbJi8FwOONR1rCGIMNUgC/V/o2qgY8BHny+MDf9mj9zN
A7A5Bt8g6sc9wDjaz9bmt7ttvBraZDhA5YrNLtffDurDEJ6tBJoJfYjyi4R4x1gjHU64RqrLP4h2
REWB9rar17iFCIuqbErge9icJ0UtyY/d7NO/4H49NHdAWSdl46UYKqU7y7Uc4hDnN5fTcObMDEON
O5MZZwq60cod8DLtOMy4fXmfj6TrvyAj2ymd5SwoO0p7VPVZBj1ZP1jw/x8lP9jgnpLXvBLEuS2v
QjrO0Z81Suzs0KK5vVN1YjWtLHwCfuaZck+RdJbqSiOUjp3tgdQ4y2xzD1YIupbyfI6ErF1Jtqkd
08ifVm/5vUAT94bSk3b5qqfDm9LSW78dTG3kAuUsbDuySl6CqLel252i2mAyuH/qOoYOO0ItdZZM
1OtUZvo0FlMKwPSklZPhP997bIdGrFWHtfGK7Gfk7o0kvIruJ7ZQCPrtdpl4vHKEOOv7SxOx86qj
UoTfYiZnTz23d1HMwfV3z2b7FFb1tTkj702qLOy9az3pp6uP8Ig+4IBtyZyrgeb4Ii01gBhbLOMo
/ZJMSFKjTxsx+VKFHQvjmWB1OcV8wrvOg/WpSDWSXTRmqZYA+YWQDZhTMb3XlfznK6o+xQeXplOR
yNmSOWAQ/3cPGvBKq/9GJZSTR/syeo5z0etcgZ4Cge9LLMq4NWtj8MyENm62Hpq9eLARG1J3gtnj
WRCDxp3QT/Mtl4I7j6TUUAmUzs+AfxOJXHQEcBOV01mJcXVEctuPcYzguN+Xa4jpiFpkaPdKvK8F
LIemQQXw79GHUqFBCTZ9gFErMDOXqXDojXN/FCAJP0WzVonhYgSuhKk3jdfzlv5w7TFkS/Z5F3vh
W4ZvozFn4ddnoCd5v1l18arBdsiztg6Vlw1RYOgiTnnCnl35aVCR4K4VIxCc4qqVerxRdoX6e+7G
D619NgQri0AsAr0oJuooM7MSnKoX+StmjZ3x7FyikpCxYF7W3uv19UfNbyzse6iISw8YJAkgYdzL
tNDpht822uvJP1GjGSqZXiPVVv55hC//flkgQAFSzJYJt4RDrz14GYhFHSUc5Yd3nfGJUl2oWSMg
38vk+BHJpqAber4DvhKYW+4uD4QL91FlvLK1BTOIQ53hRqXx1jafi6KHFjNgQ1K3BkIcnZOs0sgQ
Q1G7SmIEevdR/g5ZZfeX87sZJcD80N9SSjNqOxBq3b5cBoTWDQxdo+Hu5tsTajP8blaErOimqLqw
TG6B0//MfY1uKm4ajzA4oPMyJzJb0Ma7E6AYz+Uk5v1zaAMUCu1Hglef62djb6snQTIHuZp/Q9QV
InAxvS6Kps9wgStWCFeqEayMdxQ5Q/YFP9RN86Cczu3npyJiNxBn3zzyQBsk2xD8d5FweCThbiHh
thnEMscK7DbnP0r9m/mg6cld+iyPSAKJ5qp59pdPqxb8/LX6HcIrEuNZOkSVf4T6evllpJm7/Z/T
cH6OPdoO49+MrdBcCnYHTHIbeGiOL0qAvZM+/yrzQ+Ppldl44xB4yzStlXDKdTUUzMtfMxamU2lt
M2bDwZPC230WXWO8TI43kQ3s7WIXiuMNYhJNKDoeS8aZDJieKzai/pm4H+jRI90DZInHNhhe5+jb
Z1WjpYwp6w2yCqY8ducVGezipRZUwOTFfWzI50vpwon+C+L3fO2KXDQg39BsCj1Jk6Q/FHF/OdJF
/uWfrIbS1oe6vPNZANmnlACNEzk29LYNx4PocHPmd6QtVwe7jgZ+i/cppor8FfLknkRna3ZAB6IC
BU5KktJeusMtwrlXhN2572vkmu7v5ZT2iU9COuqSsb/8+fK9bahtyxQbvxQLyowNcyJRJd/ScEuA
a2KdL9G/fCvq60gWWdMtJy2rwdeLghNl/40qwY+MQHi7vKy7BsLpWJLGKbEEsXlsW1MF5fzdfWj9
CpdrzrYb2LuvwtA3YjrIQuOQwM5Df/H4MFfMw0fBpGkwTF8nfLR89N+RZ5A3Q5m8QcUYGo+LYgqc
kkCutxSAOyxSuI93spmMgjt4RLCR+qErVX+U/DhwRZhYyjFsSBUMSpPbMBOtGE9aUsCWFFGQlxSU
GFX8h0gnXrO83xSj36P5M6kl6lNacPLXrrrvMB/Ygtg6F7PV78t/w+VJ46Q9zv/6F27Rpz1InupC
PGuiJg7KmsOT1E7Ou20ISsMUczqxJDMVnMwB7W3hjYbOGWaiMYXEIxPdHFux9ikbBrkR9tqDlWyz
kfiEuWHafwp7CHOBvQQRHVd5Qlt/6uDqywmwocdswY8a1fBPzk7hMgxxDYluxJdcXPTlAKHcKBVv
4ovWTvPsrzj2nNb2KiQzsfayH/cNm9clPLMkJbrPMxrhX4GJM5/Rdx1ki4OiOrgGqPUC2nMW5maB
Kkrp3HXt+u8ys6JhH/fkt01dV+78m8b87bivQZuhV1nYRuHWuoZEOhc0F3W/ZjJwUP54VHHOxGk8
Oik5kDz6nltUoaar+wUC4a4BCXsM0QEHQlc+eFTSVQakSsxalC3C7Pjmbo7TiYr5y64beY3GlHOi
oUDI5CZ4fYRVAPlgWrlkZ3UZv64y83jHPxPlNx47xrFuCVA02uJthtrbOKGMZv+Lu0Q6/A31PQLq
FMRy5tDZZoA0QPuIG7Ek8KQdLbc8SksGJxMs5aSbO2qilBF9j602f9BJAkQrn7DzK1ty/bDBP6m+
5Qzuyiv/MEggLC2oc797qH5HwOs7NePhPtJ3tDtFSWgH196F60nj0ifToAHirC29DAnK1WaLHh4L
420zYEB8uv9HaNzxDgY6mWyuQg02QPU3cxGskoKnu4uUL9ZHaA/x9fphvxHHokAWmOOPq5LeeAFw
bf2cRfrDSzw4HVMf06PvvmpLfqCpL9nICZJfIIyt4CgjMDz3gukyhpdaSc5RlUlWaunpeGkLhA4C
1KqUD9q9YO5L1CMRB/2tOATG+/F6WpAswbVQ8eHiLsk+V2DQ7vjkQLwl0CdyGG1TCs2Q0jChGzjP
ORb/1fRqAHBQ2j6dagcReZeFfgVwScmVJzkmBmBnuHgIfyS2a8pA+zRdJVbNg44UnAMVm3i1Gdzg
nr3+zoYT3Kyn6wFYEuLjbSdLOxjUPQEmsvmgJZ2vnDUeAkb1pcUe9P61ZOZFSPXBTJmVvv7/o0Tb
Lgeo9TL9KGuui043p0nl8QnSEGJWyU3B5ivh1tDVMRZ81tZwezKNF+rzF9CIqYsIOK5o9IYspe5f
SbccIQ+0Oe0WgIx2f/vw8Q0jTFibcGICJkDQup6IiY8t1/9MdZo4Jf1eQpal38U2MwQfmg5Yb2jX
DQUPbXERweIHHdA32RPLnNioxjDwP3cFM/rVygwSTrOAdA1uIfFzCRRVInjilI2eBcFW6aagZFGi
SYB2CuIAXIemyFcHZvUKVRZA0cx9D+7Dg8dsSEQuMiCADsKtzqoFWyM6yalK9sL1ycoBo6gCfbRK
Kc3ufF7X+gSkij7lIK2c6/JaMVuVZPwH8cC/RuC5z9scCTy0PjJa+++aGsNPpvg0t7JW/oHV9jrI
VxKTyKoIk4QNx5zGEQ35MMdV/WaLce5gzBu6MOcpd3eXIWMTYFxIfesJverq/BpJYB0eFwLdLR+E
mcul9GaN53BvzlikeQdY0M4lHqAMIICRQAltEGxTQcKzN5lLso/DNZrLcE6/w7ZMJw8lcWXoxrjw
klUEgfKxyJWRUoVhi8hT32pAu2HrdFaJkXiMNldJ83z5e3/nvqQoStIrkDfLNixEQYF8rDBCrAM8
nP2BCvQnAweztWxbj5sGb1bnCZ16jzSFT5BR+Jcb1ht01jFEDII/0vmNL/f0Sg32wZ3T6qJG5d90
/5P1gkyoje5nNre/Lm8NWDIOqHP5yvn+3N0nT5kZLv7O+Bae+PmZ3XGmcoBhMu8VG0zzQCF69evB
BGWQNeZQyklTZgckfg+x9EEtvc3OL3ze6iET+Q26W6pLCM6A3GUJTk1lRgWe43jrXt3XdBuqkTlM
1Ef4hHF5/HNOFumbPXPGqBni7j5K5C9G0tEfcfPC3Yk4os8wzVbzwn4ohBLvGeA9HWS51eywR6QG
1C718FFuxgTBs9CBYzfyAruOwnCHD5sEUzGqe2N9I0mRPaEX4gvxcMzJlbcvrQx40HQGxSE1jkqz
bxbB1gL3F6rwMBtb0fvmPZjLxCdNIXtGhdp8+2qQm0SoGNVR5BDateUcWezXf1pFqOzStSQP3biD
w/CcVb/C/eHZvYKecZ69LeYiSzu0ebSDP1X4JvKMVz0qLp7/NVtg6sGASuJfzYsNFWDxvVCwwaZP
4gGWXxpbtij0WYQtH/0JG5NZbdlYeeTa4RR+/rWhVEG/CfVKNNnaYh9G8Ogm1KMaVrOASJ11t1Na
+oGouDmeMkdFpZuv+u5weHt33+9XM0RgkLn9aLshKl45+UiXgalbRAfKHlJFLUtrPe8mDl0AeoQN
KuUevwDIr8HQCq7anRCU0GChE0MKVPUz2OD3WAfLwhbMgGtf2fVvlhpLKp3OpYBni/7Fl4pEBBZe
tzkIBMBh7Y8tgLNDNRt6t1KoOTwb78c9TJgD/RlzPRI3D5P0jzeRXZULxfNOMSQe9KjuJiOarL+i
LemEF82H/hMEWnjOZBZolUlXkKE5fhgjKwYzUAyqEtGu7YRgxi41j+4y1BGXLKVsmLRcl5UT6Lbm
F6V0WBhFpOpL5AfacqOaP9feQydXaL8u9ledtJ4kbIK1Yq3giI/2plYUwIqOCeJ1QvLTVivMkxei
Ov4w5A1S+N7rrMRBp7qGGScnhczqSEfCHQxwvkbmDiFF+pltNpe2scFAw6U5BWSf0riqhNwwSFRo
aPyP8rDfebi63lC3OLr9mSPv6iVOLDMeSl1+QbhwV0u+kJjPCRhuIToe9DpSv8npwQl157XRbftB
xoEKnug2LUNrWKfEkgzLuNFZYhFLu75X2zSpsohA4HGUSHkqkdye3uJMRP7yIwRhdqdyvx3GBxQu
5r28X6Sgv/P+GqJs1P3yQOuknGhcR+BFiqJe5Xi3UdfYDJVcQE2IecRps2iRRPGpFphlz1xjkSUR
r6KFRSY9gYBOXa1OfAPXYOn++3oJC/AkDaBIN0DOz/KjUhpsyEmbOfPKocqJjlU37cU1dQM0ghoO
rg8vqzKO/++fIVlDL1RIk3B0Vf5Epvi+7IF/KK4TOHC7d13R1jRvaIGNQc2uvMf0WL+UvHKCyAvV
xQkvIu89cPhXh6h5BEpZNfXv23gkQyV+456NKGkAiAeIF4SNc35SxINpdkcKRHv67l8z/MTfnQmd
1o4oXpwU9y7RZfPMNroh0FbpeGh70/lIztz1vsVdj2fgshKKWhPhoWUqp5UNcwnd2Sin8VP12eWm
cO5BK4PbBL1T/Cqv+pQv3sa/PK/ht6BCNV6GBxdStbdXuxK/GwTmXO3SuyLYG/dnbVgVYP6NL3p/
UK8uXw/AYHpxE5P/WaPzdhi0C5gtDeTIyn4ohnllXTLOhMZaG3ykyHWnhokGnrCKMunM/SBqTpiy
aFAiemTagMRirFDbzdW/+fUkb5ZtnaibyETm7jdHVm0X7NEb0lTK1dIz8Kb0tpc/gABmqu+LgqDy
bwgm5np3X0WQBojeC9XaMyQv0BC/cBdAbe7PNysk1LS4CyrFlht9+u28TcU0wAufrOuTC26ijneu
TY1YaEGdcdi8Y643wxG4h36btRc3EI4v2DYvL3J45qxhhc89AzggpnsI+FPUSDLE8i8FNcrH7Eb+
f12CCiesow18UEBhq6YXlvSzZA4L7onfaebHJixu0Q6zqIqv2qhRFy0qo5202PNH14mAqx+IQImy
VyZB+rO6TA6oc5gsheVc+2SOmd7XVQz2LaOfdKNEcytOuTLu5pgxaz+Ql+zmIgN4WFnw7KBixAXD
1N93R1f48GmQ48zbVKV1xgBJsLOEe1Il2mcsiwcQmYqOWdyt38PuWV5gvfmmc+NhwUkIl2hx7qm7
p+OLvThLuHWyOPW/7CmWl2VTBvGm/uNbPFt+eVUNeiRTxGXrM2IwmjwsOojq7dkbtewqxdhVXRFY
QYs6AitDanGRzJosYYSc49iF7gNLuK+jIdNHJbjFOCgsRh5oIxPbtnIKNJM7gq6KzJlOcT+sNGjf
fCLF3W5+NQCST6P+Kc57uWw22dPDd3p0AGLkdnqpdG0ew7LgCscHoJUqCx8ZRsj3G/BWBva/uiZe
cxT9Ki5C3BHWh3HICftVeEC+k8wxmkyqGhp4TXACaJCzUc8abRIp941RFgcxWCadLOjRnFQlqe3c
1Hzqq5uyoxIHUK5wM1rlT0/Ad9XBG1SSC/e/NQcUl6BbpiBooXh1vuxkR34IhL73lH4ic3aLi7aK
NMPowxDSoTuxpHqW9gwoTH71ksAGfMXPCngye+PKcMlJytQfIC0Hli2wekzR56KSOQ7G3rDQ0d57
b7WW91lVw6pi6sZjH5lQaxFmNojI3wEq8hkh+O69ua7sC3u99yiTg+qX42k+445OfNdf/nxC0KTw
WaPZr9q4XJg2K4IkZlRuR0Se3h8a7VD6voBEd0Jsea0kVT6QCU6wEV5VRLUTenMWXOOQ1MMZCDXk
piKCGdOOqDPOTwu5Sa6jy1dpt2fMkjLT0lsrH8kqRQ1n/mMPMDTarWHKPTgTHUDhW38e+x1dnhly
4kpYXtdwiJ+LGaKftpXThXfqbWYNcLJpHmUSUHRleNKhK1yF4JSYobZip2dWY3xH776QXIXcM4Lg
lD3o5B315YTg8BwygSeEoEBGF633UlQPnP951oOcxWeDWakiGohLA+W/dfH6e+MytQVbOx5zeoSu
iG4+R8Tch0XkOPcv36dCCA+/hfE3JjkBqqsgtmKnou/HCOUXsVxP8HUtqhGCN22suuvNud9UI1Es
aDPAnK4HwpiYhfPcunIni8G+78VLZOqzIfcfKI/Yx6h+5VhVcNNUc4WexK7rmP4FQn1eNGSp880I
sJ+Y4Y8LIDEfjGMbwdAByPD5eVfcG7JPhOzY9xKpAts31n00pPdAPzzbR0uXNZS+vMquDq5KX4Sj
Uj/VEhITqpJuOhsqHPk0svoK+RMiYeOuiVLbmgmdMaQAdEVzVN/lwOh3qFx8SrxXeQiR0KtpBPK5
4uPW1V0KTdUrQiTzP8VrhVAc7a6E/9le76cHOcHM/gdZ26tEuYNVXbvbzmDlK0N01SsTNKWeXueq
x9e3rhPsasHUNPos3Qpmt/ZgrauC0YQEuXbbna3n/xy5kBmXVv4WmX0n4nZJPsNPrBLfxOHC8qoz
vzIoy6jOoBxfmg1psNP58frMglCuobU0zSuduze3onAlAT3qz7tphKWwK9/RFphmj2H/Cr05xj0W
ji0RvyMuWhxJcMxV9KnapaIsBC2GJ2LhETTRNnTTwXqmHapHesaHqakZ/q7JC3+4fvfhiAx5wJWk
IMWmv1SRg9jROzYKM51h5ZsBEpRV2J0lT/ORADotUH/Ld1RXhX3CYygXqvociEPJqXxpObhHA506
qmVif08jemSI92MWsZswPhgnbSB6IwBk/j2ZpaHLEJIc7sPbPEhkZ+/y6LiHUJ8usf8RM1lqywaj
liwUc99Z/LEiRTaqkbbU2xcpcQvE6K/5SiZNmqJVPNd0Hc3J7MKz7AjobHRG8vSapbXIIpIdr84L
r1S4Tq42kGnY659TFYBvlUZm1LAvqyOP1TLdgZrEgz50T7xZet5/E0f3CUSoYqL0FgdOfiQgSDkH
2YCwT6+RHyN+NG5eHSJxlRJkI91foe5dLYi8+I/6Gu+uJ5kNUZ2zCUdBcm7Of1z4fCzzMqE3LiYK
FKO4rczTBsfTrhHDZLdt/QsPq3XSj7zteNzRALy2acifXdEdKjPRjzMGKUAOUuyc1Q32rb6Oh9Ea
mKNAwOA+Oi4d/eXknEJ1o9Hwu+Dq1YNfObn7iuRgtHBePwaecdGpKDI4kQxmYHCeQTSvOqZ1scVY
YTR6TsWQQsMAJEPeeBZOyti3PyastaB6bDxrnoaDt6ju0CLYwAssVMPZwBelBFzoMP93N7E9+ksW
OQHbi1GxjoQnl78Ynlp3gvTW1wYEnT97529iKwsyZLGIhfz8uhAs5yOn8FTInD1t8xbgqyKHO89S
/tLoiWFUl9Hj5o+f8rIo2splkCqUq4Lc4so2xlMiNiC0bolSOCu91v82EIFJ61j3aXdmBLqwO5Cx
2klSupMAfD4NrdJooscYidaF0g6oEh7q/tm9zYAsLcKe8SvInt0btAKkj65VJp2gK9NbD1lk17b/
8qEUZc4TggIUFeFr6ar/oVm3KpuKnT0bMlXFU3+++EhjYt1WL9YCnAbb2pRHE/GccE/hRtxoMUmR
mvFpEXt0cmIxAYlwOvLnZLWOwOhwJqtFwkbSDsDfAMpGFUdxGPJgzdLjFN3O5mKq0ukv1wM276FR
ytBgMt3jqSHxY/3nGPZURxibqZvGRNY79taLaJhtc7cYe6a5uW19exd8yl15aocxNGgTSrSpmexy
2EidY+AemzpUU92pONmArx/7FwsxbKeQLoJgs7ucRZf2X7gNdDScLt6FUESuXMDdxru8m8mRuaXK
m7xTTGWH/ofbCphieuQaD2GcYLxrT56o8e+CguyD8UvmHEMLv6u4gvK2GOtz9WcYvI8gBeifVOAF
MHTUoImb/AP5zGQQlnf3tv5OMVzfmWqLSyMH/+V1kmBDQhX/0xz3JH4SyuVMvjjSb0gJ8WAomKux
y/x7jfmh8dZ7pSnH/usGmytRwWpH6syP7hdZKdZJ+vCCDNIeE8eYcajQ7oIJ5TFmL+c6r7EYLDMr
N/57uOarorXhEft6liAWbVnliu14sPf0XLjGdQO/VP2zxrxjZOjo91DoNDLeXHzX8UA7Sf/HkTDA
GOMWWvJbP0xJ/taXV0c7IMQcUDfWc1GxdPyJXR5G/HCfDGT2L+GjNRbUc7VE0DXa9lmZlk3tDIQx
pMJpKp61Xz1DkQSE6Arc9CGM1RQiftueNwEVg6CfI2QFzi3qXQueA6QQodfbN6rJ/YIDvgZ6Ty4N
6iXaPP4YrvIowJl2ODsdwI2xRq1fac7JVtujdT4CHf2EiSMtTr6oTugrQCGCMsLGCcu+s7FStekI
4sYpHEcWgFeGcXA34ffkdlbGoxasG3sLe08x3xLtQppiGDW5ldWNW0ca7sSrC5fdmZ/hWVQPYzZx
fzjqviTxewBWcdmNkuJpvfAp5UWQtVSP3bWeecK/9siz5URrsz5wl9/cJWfpzJUkHXR0UmrE5ozY
UJIVqlM3FLyp096iPydIRdA0XRfiKhDi+3Wb+WQziUxqdqLjD0kfqcUUWBiXw2CbSFX/rVB7LBEX
XkamOTFmzx3kNtJro2b/Ran30yISttuWOB/SBsgg2g/GfzYJl15AtlnkmptcAVxyjNKecDexxfcL
vCkZ1/F3cQJdOqxm+Ml7lxWZtLDIt5c/8fRtjd1xcPeDVPoexhP3U+khhfJuZGbSqoxd3VDpN/st
bUTVnk6tLjOABXyNWr1VgeWVr+9HqKlFIJd0PUfONfrdVgHlrkvNu+yh9Bb26zc6xF7qZOH3l42x
5PjJz9bJxn1LMiUPDtZ80itfzouuZjFleT/ZStg/IpILDBmd+Q/fHwEc1sUq1YydkbtDmLIsshlo
pwGZWxAmdvKk60V4hgGHEfT2OrZwCfBJmyQSvGZbO7mfmFX9NGuI8IhkDxIIyta0gQdfSv5pN5OC
2F4EGmQtxCK5Jj091XTwxBVVsp6qUXFYpVd8KWdAsQl7ORx7yhU66y5cG/50EvcS3XND38smvmSI
13395AtbDRsDSVukmd7GeF9kSN6mEutyljtdyLsg7UOVI6rQbZ94DDknD97GaEfr0z1nmvumhAlF
h6/G2wszGrIu4NVPG3brLdWeE9D9zA4zQ1j7ynmDSTYGfu1ctL36vPzISBLzEc01jIwN4kOtBP4f
69iqn7zESv0DqcvLfmSN0YMXmJs+UDbWBAEe7fPhyBwLWWl2Wo5lhoW6Suq/+BLpu2UKyfO0f1Kq
JChKG7cugP2L/ycQ5gI5mKLFyxaEghYD3R/0sk/HuSzOdzPj+yTb3X7dB2yffJ5/jnk80QslMe8R
h0WrD8CVtwZfczNhh+vMktCrrmEhnj/iuyULCpQpJahaINc5lngGjezHEvkwNn85FFv/qYX3sv/w
rA4jG+LPxPeNV4PzGXbEzv3Bn5lFO1FSSw8/L+GZzvuTDT+0lso3HiAfHn2v1R4DCBDO6r5Ws3K4
gKUbg01JYRQJrufXtvikg1nyYW7l3TA0nL/Z5ZHNmJqZOUm+gD2lTkKpDDIRi4suV6rWrM31vc9F
idjBq0ps1O/+BLqRFCXUJe0DvbUvufTZ/LvT+t+3auqk6Y4tlqVXHd6Lli4/0WLaMVGrUfhTQNm7
clvVtT2FgfPCaJIZc1lYexF0IZUS46uwv5oso3yUnR/mxnueFQb4x60ILNnDCz2Swsn0JOe11MHO
G8SN2TZIMqPEDsSrlh10Xos9T90Gkrf4S/n9r7TrDnFYvT16PklPI1QHvkbwAjKD18Bo8I5McWAO
BlfKSb5TOGhAxkhq5F8QUcjkPAZc+25rrUi3dfjqLuFXNai3VdO17KFOnnxwghEi0FA+bwrsmOCR
MV3xEh/TOARxncAfhzyGnrc4jrR2qLqidp/scsBVst1OW9CYKJz/DrGMutLbb465h6k24d26VS1t
79a/mpWntxp2grvv2ylBhzTywzCGtI8rsqeXVlsOZSnNpgkvMCPXriJzaym0qnQuiIRqFNL8XILP
FWCRvst0Wrgxt1uOpqELq8aAxe7k8XUCspJoQLj/ff1VJcTq4l8Zoab/N/spHTfUHmkPm5Iv1Uzu
N432R9ZsAa1VLL5jR+sEKvAsWI2vG9UDKYhTdV5KnV4WVEKWU1eK/x+uXfvZHvQI6zP/emCws25E
1prn5id7wniJqQWcrrtmhXFUW29j8wYL3NJB7bVlbWMnhdZz6QRmwqa0/HpcCJwfdayXoda60SsR
l70AnRNd4WIOyTh23jPWOJUGegrMHH/F7Mhu/f53O2oZO6yB9vG/XmwYRaVBy7ypslNlLUzahHjO
r69KMAthVZiVLGaNLTjBDb703ip/XkSJrSjuDBAPM+xoKJVNQTyXWktjqaz/bNw42UtkzPJOEyTf
2u9zVIuBnvPfJN+uOHGpqCkK9Z2e5Xl6ibDY1ioVWRorF1vCX8kG/SH5YXRK5a32740v58f2ReMT
nhRPx5xXnHh2miO87nasz0B5LYTUyJtW2I7P7zDNVbTqFzv0zhoSMIohsoxyaJScVChyoF3zowaO
qMNWZOq1wKv0rwFXzeJ06MT+3xo8vWB3wT8SesJikgQmVd/ldq8mDVR+sZaFFEVa9j/MbuQKDXgg
vne1DRK5d3Mx7qvwky9AbKfV2ubbsClgaGWUUoYSAMMYNAh5NM8FgUa2PUgfvNGmwXu54toPD9HD
j/PleP94AqE55cCM8fML14B7QFZYGdlCmVUVyYUVEJttX7dqdTtCIIHNCqlZKnrN87NtzcwzlOFY
os6M6BKbsRv/1mN2badGUmgM8+9w5U4cp+9Rvx9012B3auydXDRkcnZmnK43P6yyKlR659+c8btj
P14NRG2XvB7n6T4d5LUns8h/STB7Gn6PjqKjALmpo8IL0wif/KRXS4kvoOJu5u+i3ln8ErjUxwP9
QeghEBMOYiC9wr3dPvwwjatAx7scSyF/Eaec55WsZ/lDHLdZ893X8JaH08genW1Asz1E0G+tDffY
zwVXM0bY+daO3Zq8lyoTCuIG5mBrcWKiHH/yewMhMYAbwSnVef/4cOtE9XY0peME9WWerNGpugp/
8MNXpFjfGlI1nGOyghlNLCzHUhNu0r6YP26aRn2Y5asn5Bne+runhvXI5dyysLCHDrj+Ew9XxD61
u5Ne01SUnptuggRtbPJhbIRD//NXPbSTpu5M8YSX29G/411SjZIkmjTyB+PjdzCIWdJlyKNMVcde
AEtUwf5bj6aMtxo+k/CZcpnaiq0ZWAYOqL8/8Nr3cXxeMWguWu3MDX7Th2QHXIxUvM6Kd6HHUakb
Phs+DFjvREcW7e8OTGSlfZ++XfvMrVFmgOkeyTcqshs+pxXrGhnKZK6PJY4wJH2mrCVvhGXxGXq3
qjRx8T7HvgeIquebweoeeD+JuLM1nydCb9Q7Kx2iDKJsWCYTE1+Tjmp9biZnEQfcG7uTAQJiJYTV
u0ARGqfGlPgWdhhn2iZmluOS3u4mQem9XekfSTX84uq0jddsbYGVOcrsh01BCgApBI/w8zljq/bt
uvcHnsDr53as3bL4USzb0EVgINZDbAgbDQzo8EvdHdBtRdWE21dcggEHoI4jcLcAAEXJHeOAdjqz
AXuTA149CkKg1yWiDdlEIoSA2vooPpr9BHbXbLQVe2Ff1gQx6dJzgtnO3IwKwLKmFKqZ/HUlK6Ze
1yt/YLMbaONumpZZ94JErWYcXJfKWpAH5njrJmmCAodAGEil7Qkb09pfD3q01ns8FCIOh+oKhED3
Teuq52I9QxirHVfYd7dTPTfUyKc+pv21moY0wR6Er7UFTsZqbn5OFZMmQ4oxrhsn7pABn/EQ6EqD
afh/WLHxOlZP5Fq97q0kSeA7OhBNuEXlMrfhakbhy44xXELTc+IzvVCCHzziQbrA6lYHFmK2qiuA
lrxP6bbGutkVTwtExcxg+527CB/7mt/hafds2mJzrK7jArZdCRb/1JfkYDB8gYmYGGq38jvHbtK7
YBYvXBnq54qHLsxoIvx7NmRE0BJaO/9qcR6lBcFTNEdETyIj5xS1JfdRVNq61wEcmzKQf+4I2dL4
Bfmq+WNo+C5p09gBqqAqbBjBka5jDMAJ7KR0qOoWw/C7m+E9KtZIrGnh5y4oiqN+g2dKDyb02mUn
KRVnCFS+97oVBAHrE0blBIT8AZCyMJkqPllCN49LBXswE5IiipOsA8HVc1m/qlldTfWbB8bE1kzm
wDf0HiW+d+EktgJHiwrm4cn3EJIiQs7Bnu4YEThiPoG4//MiqJbFKKgIz1PShVBAww+3uNz9hH3n
feXZw0j6QUBgimohQ/kSrv/7+IPRG0j26NdKHoyUflG0Z0zZKmifoqQK+i3n8MRg4sq2QvqVKcCy
XGb4M+WyoJa7djYsipC5l2EEl3qU9EVv0hk5hxSnr4GXciOX6ukTBihBBMaCQ0hJwiMCrZAHXVBJ
cWmSm9YO0yTrUNMgMpOxbGWGGtCTtojuEoHR75Xk8PknnHA7YYPMiFdzRl1SpIHlBNR8Hb6ckalY
817c7EZPk85TMuEoTO/4jbwL/3INyKR1HNr7+MlFe98koS7JVNl72rbRNcSSmPWDyND+3CcDH8OU
BYdG8gYwFan70yshl/+twuKEPKRXgiF4EDukm5bLubowXrgcuYky3+nbQteUD5WVPMMHu8QQh+nw
KFyrfmS2Nu8I+3faHR5nrpgXBhI8BvWIwg0i2tV8/gyzQ74LE6WPPSHanrCJeOGQKUaj5eTuVg+k
+wBTgIQqxrNsvDsgRQW6up+x8dW4l0SwzCEIxbwSfqca+KmQyKKEIwSx+EY6nDD4Abia9AWc4vc+
C9yTSQWiCBd3UT9Uum08BBiloyAbhHZGXoSyKamT3+oDlKltYbp3St3f2HDnP66q91qcYonYi642
Y+l5F+g5/meQBRTGVm//S3k7nGPYPUCXHmsJK0A4O9XErzMpXKrq2g+0MmKzFQhaLDghc/wE/FT/
10+n84dd3H144qDkLzpeoSLq2e6Q8OQT+uUu6cNOAwcAQGRC62ym+M+QjUoczevaOLHJH94CbSfR
w8p8w1ILo8cE8RDykbm+A/oAr7CWS5GwXYA3dyGkgDm6JKatZlqDhfXG8q949eJjjYIWwC9v4Jaw
ZobgK69hgc4BTc1Jy4938BLmaGO5sk0uXxB36rDh/fh/mDY5eLHqoBDbE85q2zwFyz9oDJceG6yZ
sAgT44kZI3bvQrmLT/1qr3/OFgVZzwEzzzBz7Q10qpir/DLnYGsBAQaAkvch2LXPGmj+ILZiEAId
V6vuMh/Sy36dH5TQlVAeNO3Gnd3cCYwZqb+dnzzw+IPmYi56f0i7dMXm00GOVnLOrdCjRDG5M4FO
lP2/F0eD/qgvSxsZEbMOSn6zpK3QyaHJ4UJz+9KRKxFlGkaFMil9ApBIlJ3KALc9+ayr80yFHiZl
JKixloqk7F2jl3jtEOe/K3vtlSrsfMadJufgQQjGxGePmnvFkScKcSbf3MTgMk5myDZ8Gjzoabi1
NuvnBxHbBRyJR9EAnSsi05ItkVlMOHE1WPdoXC1FsQTwSAzLYzDS39V9AgXyo0fVbggOEACzgg7x
n/x8XxthmT3lK3dOgCsm75+HWF0NF82Ed9qJlDW4xxdbMhJRs1/C5wNIeV4TeSzbDIR/s36lBP+D
57g1DsTUaEKZLAaOx3Lxj8kbNvpe4TSUKEAlscMcw3HZgQa3Qez0PoU/5BcTt6S+eU9HM6mDfqop
T3hvMV3Jz/y7r39g4mB/skVD2D9aGq2KGC9BYODEjKPs0kvTB42afD8b8dmqno8FWR00yWOZXP8E
g2QW/18Z/BuxM36RJyQVTkXZmqK6JszKA9tX0kLJwx37EZaMbSpbbI7AcMQ3wveWvBszpd3maQb0
qb5eCw7GBzzAFT2kdAllhE/9Vn5kkNqNYuah/gS5HIcx4ZaqrPQ+CZrrQCHXYtwA4biLb7kwO8H9
XDR+4SMFSpsnzi/mWYZZ4lz5Ioju/oDFiLm8L2io6jVB2+sFHp2Gc+IMsk5pQuPEeZENqvMz8sIn
uTq5bfzXvc/iBYahKB+F0mGIMbz5CVZw68UnF8NLB3UVtgCKU4v/t+TSgpmi0cTfl6z9s8iNgMEy
xT5BPAqGKjXL4mlwr1MDH74ZZM/AiP3eIgO9WV6mP+FijePt/aPoKXvb99IseV4pnwSvUj7fcrTO
Jb9dAag35lOmOZUSKOSkzX5j1P6HTqlhWKZ+8uUwafhNhmcZF+T9TWK9UcHaE4jwXeiZyXFVWbvr
fPxw8yuPFDNc6tINldl3l5TZBeRAyenNM2HfL010wXKQVZd9MiXs0c1LajmEwQ8D7+AU0L+DdZQ3
vkMRH3ENkCviYWK4gwSbVYvPqPvlzUVBnxgZvvtxiOCdT8CKP/Yi3VPE9kzzYP8mF7r3IoxWvFK/
i6MpfoMd5Dx/gMfEku0sGSzoZ8X4VC6EeFz4efXUaPI6Pupyf6vq/BGPZb1AxMH1J7vQYGwyrzry
8RFb8XXyx6SMcfaX1ZiM2pqZvAQ9+spOakLf/hATvMBlUARC6PF+YpU5JvRVlsWcQseRhrohr6pf
BJBUR5GlAf2pPKfk1GvGA52+nR7oNpdW1VmMqCd4brVI2sCYToqTJvRG2YP8+XPzLTZTAIyd8nhc
4gVMglrKxBwrUEzKcXGCppx62Qvr99FirKiB4bQxOi2RowgKFk61UT2CgdCAN6H9BcnjWq9TGXd5
uzm4gU17Y2/MpcsdozZL71Lag0k0rqsF2kIsb8I5YCyMi4fcbZyTBT/Im5YONH4UzswT7KNphiGv
zQDLL3m7XBsOsxupecRBRWZxkgRhscY7lnn7fUz4YMEQzednAy1wQOk+wFHYWt8MBzrdHLmdDw7n
5tqQahCSu+B6aeB7YFjblPflE05R4p0YoYR4qJ7ReO25dS7gEZGRvquKWa9rSya4qG5QsB6TbxoL
tIt13fxoNXH0AbMchS/trSIunGtb/xUQ4IQNhxwqeomEjqNffNPs6OyO94Nfkv87PIs/kr9sU9Ah
xqxa9ZdtlbkagFgDYDgP7vZY9rnq34OdhN2SInxxMbCTWLb3aqT4FgCWvGl+4KR1WxhEsGWtrUUQ
Xbr/qfKgo5DHY0X9W2RhX90Mq81wQKfNJejKWcUCbRyHa26jYmenXZhqbeTj5ANUsqi+YHEwVIx/
6zaUYOwS86ENmfGmmTR56vNfVTEaiPPeSrdpB9LNNHzbo7ZRvHC5jPpsH+248x3y7CeLH0QmPq+H
0esS/UsoWhhvCQ57GNe4ixNKbh7Z0oMa4B7Pt4+sKscgMkvcmg34devY3Mylnwqtj/k42wt6NTLv
2BpbEqJ35cQ+JeNArgKnwQ8b/nLMyZpXH8v1LhQTrZdwAP29nYihnowaH4Zbq2lCfdEroz5Fp3xi
pP73Ib9AnNcdPs5BKLUnd13uM0miOH4xe+NJ8v+Y1hDVEkM7F8vPrIJDtfNctQKGsxH18PnblYyA
xcU/iKlspesLQ+5SVGsQxinL9KDTZ12wEq9SMk8HuTnox81GU8Wc5M5M/5s/Za82d2T0LmXtPRd8
P+SnxQ8N9ZQBDDnw+Py8CntTKIzn3piK/g3/QBfgU3MCz9dUv6gE3UJRNkx1JsXrGU+vHL/5huqb
FwiriXoUeffCK9yntal1wiBdIJivsXYjszlHTGFpoyaLvV+bqe9TRJgz8yFOhqERsmHu/qfsrMHM
5x5NrK29fH0xI1eeqZxdHkeKq+sClh2sh7nCOTUhofheK9mGwK+HOrEJE8TMyuMSWetPrTXYU7Ax
e022Ee/4S0ibockkXQIjfIl5f71dn6NjiTl0A999b0daAoxjVzFEQJ1U7CKeO7BAVUoAzbgKRJck
R8zBFEQERssDNqiVtF7hmJa9dnGuWMatd0vigvJRMj/s6Oz4itPj+Rfg7qAUYwAFnU4eKKJkOxz8
j/Zm+9wx24g0Hznb9OqqQFZQPT0b4A9t0elznwudaOp/ml4Iip79EChfxE4z/ZQHNxwLuTFVv9jJ
gGFeIWFGcoV2BHqDsC68/kD+sBUr9ALEg1vEc6Yz/vXIlbFRlnh4Lh5wCUYrJWKq0LS7TsihomOL
KFH1gZbhK07O6zBG3pvG/EiQjXF1eDZELXkseXN/sVxw3KN6zoXwa6wzbyuOusWOqGIUl8Oqho4i
4l8wrNgj6gIeEJQMYdCiP8a3molHjrnmRx2Nrg+22s2CKZF2gyN6f88MF0h8QTMG54J7Fr+eqH3h
Q7TKym9gWD8DdM3smEvupQbJlbs4yqfWiPEenghcMScgk1u5hMqT5gaJY3Th0mXuFRTFXbeXFg3V
XLA95vY0OBrrdhlrLMBdQBkn2WH+ZCPRSpXlzfpLNrGzGFmyVhfz13oAWSsC62gDfeXEchDI9TkY
uCEzBWsFZF2n0A5f7YMkPrS4Xcuiq8fjfvMXCePDA7fJnoR/aq5zS+5KshMdnY3no/L+wsuvFpOi
AOhMkkshQIed686YmqsazmTdK0wF21Vs85R7mv+DLcHI83HyHTrR30EsBrpwBi/JSfFgxgCBjHy/
VBbG743RbM7M48WjhdvyFznYWP1gvfLQ7Xz2B0cnNCtAwZRfIlHZ5gaOknvCp7yiyX3Z8RkMKECt
ec+T5MjREKCg6h9O5ZK6DKdSLUjbdlHarw5J0V8aUcr4Xd9smW1jfAVUnuhH4x+G0bMzMdkQ3EDN
gRwefxMS/Z55SGa/UWbgjtRCUK4wDPm4HRcm1ie14+KODOHCEpg/lNcgcjd628gi5KgFRnvYnusO
TdNW5Uk9EzJ2vdwpzEjLH3wZDZjJEqftt5WvA1sYdwqWIuohmif/oHY25jckqUcU4T+IFQFgrFZk
A8Wj/eQudmV6ptqs6VrrPNiYT4E+xO/Uhkn+u9ZDIdbDaV9Gn1RVGQclonEhFb0f67izuZoEFEAo
dNc9r9h6tWfLadno999SprLLyLDpY+Bc6DDhO9URYhNvQexrwR3kWnkXEVJYK0TJIhEmc5j/rc+M
XXoROeOqTBDRGm51q3vbmGt7TuccXYrMAHQU01xcNhvHRDNvdUqnvlMH++VvzTXaWV/D81ygZwi0
tVP05jb6nWtclD1Bcn71eTeDSgjJ2JoC+RvX8AZwTyxK4gvpIoNiG7vt4/ZRwt4XdFDnmG9Y7d3d
BUYMddU2IFRLKTV6iAHf7pPXmpJHzifpMaqYoTar6QKhZ4PMPUEq1R+vovnLuLdF3CmF2QrYk/pV
75SndlUD/ty6tyU9fmmEUyGDB/on1gyCzLfrQ+Ar52M9fc9ohqIilzROBipjGLE6pl0GPbnP23Wb
bsWEMl7sEfKi1c8nN4WGgKTT+mRaUzSy32gffoW91SkG+IJrHVs1KqdPxgs63uiwTtcZK/iVK9kY
kIStWcIyBKukxUM+9BFapyFA/w5jYBjiw/iTOfwO0s9jAiHiF4cwshY2HErPRznL8WvWn63B3YtX
IoWgLxLpnwKCWvhftB9no43X4Rihj4BUqZwMDfZiI09fBqs9NcmHEgW/tCORsaUe4Zg73E+GZlWN
LZtbSnP5Rq8fpCAZfyxcOuJpaKMkDHVst44Zk1WmA24vn4sDEu9LxPgYbnRmwfIyqpBVGCBMCnr5
Jz/OLI1tm1tMM+328LWe6I/np7qYwNPECdTHelXEsgL6jLs+8WlJnooMBWfYOgj2slvFELcgiYL0
o/6nFn27YmEtth5MquMdaOJdS6potE3aWIPO6v4rrPDRRkntnU1Q2g3AiBD486jvqEPjZYXQW731
n51EyB/7Q86cyoJr2P9Jz3MsTc5OGrk96qVCvYZOJe2Oxz9sskNR5Z3S4IUIn2KZsd4TAXSs/CuS
zpl5RAEnudwQPKn0j/svvYax6uAUW3IoGVT1Zg/HHmMkObsbnT9WyYpF0LauCE/iiHq2F4/fQC3V
BZo8PdNmKtpfNJyLhybWdEL0CB9od1X50WSOQFEt4lG0QvUxriA9jDfrGJEdydIh7HdAoWIfj87m
4neqZT+aRTv9OB6VagRljaeQJ4Ymw8zRh/Vh3TWnv3LFZoUoPWLock9iv8NAXZN5LFIbq33JTcJS
tMgZFMn7BgN7lcgRtKFILxWh99GkSuWUzqt0ldUnKA3eCluCwgK/ncnIXxrsHu6TgOMbFL97Q9g2
3geUtECN71H7rJriFGu0uUzPy4mRxKx3J9tQBWxdpARWXBONYIgJViztzDLJrzHdhgOkrVXJsyXh
DeeWYQH9qKUMFSBlt23typ44Rf0ai5HEL40HKmeS2dqJh1nOtErOkSd7cLiUNoOGC2AjMyzULGOo
Att7HR5WFllCpnc8fQp99y4hfdQim6NggXTeETVsdBTM15AhawjO8yEBfkro3EbwkGKfoGgBvlCe
V6RzCXRFJOB1yDUglSRm/pBU4p1mVdTyijSbc0aTTViXDNlBQNjYMQ9g2yAl8Bzv7kqQ8usoHdrQ
dULqKy7eGwdFrMZRjL2FBAfcC+VWhlTxTiRs/22Esu3SDgI5aKB7GXZFdKAmqRN4nRJCeaz8gQTn
95exv+dkbeEOvQ9Fw8CCEiKANfF99lREhTMr5S1hASywBqV5IUkEVDj/tPqA8CQRZCKWEShwsICM
E2BLrnB1GCgxALSpTeYtHtG1Dkrr6XtQ00iVsCPPbLJ7MEjxgMe3YdmedoBv++FR/e3HAt0BlRi2
8jgwAl3FuKr9GtfBqQuMq4nBd3p+wYZpKuMTEFD7FgAtRd3aHQkwDjrzsG0HDP/SdfDykk1w8PTn
6Q0GLGrx0xhBW8JzxPZgaRy/qgkN/NMD2Fo+M653NvhCjut4Za/+5RUacow4VCEswU0kJ5dEX8RO
rX7JWK5nuVTeJ3P/NYfkenTrwmJATST6v06TGsmM/H/G+h26uiyrLo8PsnVY4GFaKksG/U/Hei8o
EW+KFE5Jf/VNwlHGt9AQZ7OtTGOR77cLGyQjKi1y67Y9xR7Su6jKHrIXI1lAu/h//DoPZ54RIlrk
kCVmCJiNtjK3o54mQP54RhIvKjJhezpmaPBjktrPGNFcJnoCVprzArDCIg9uZrUk4TXaHaGG9F7S
YCoSAx52MCxIGTVjXhOVXeNGHPmqoPTuljcwt0OsZ133S2jbjuny9Cl2mS+/opS9JwljsHZsZ4Jv
IjKE25WMslJhanZhAFI9rBu7BYGxc3pXEVril94AWrI9O5rBnMbL63wzsCS0NEpCIcFagBXcAsZ4
2ng3U6ko6D4trhtJxLiUOIXhv5QqZeL/lXEeHQ6L3K0cIwMP31vu9ztZ35GKTC/jesx5XYdQKeJC
DrkHj1TJEoGD9R8WBA+DEwmFuNN/b6qVkJEW/LdUln09H6mWtgvxdR31V1tojSLN+TyPCEvREHEg
ztkSX14l3M5VF1DAVF3NtmNiptiAW54UTGCOBgi2D2hRgf7UT/q80XBYGIyVZEg6HNa8M2LPe/PF
YJ4fxQhyte1+IyI2VgAMsfA7pWAhyLSPTxo4l1uYY11k4toN5LMLmDf7eiw1Bz9NZRYs/RyZCYnV
Mk5HdLaA6buLK/3Ve0gG1HXQc7WQslW3MuJCD1W7jdQVhzdKHU9fydvRWccmfiq15Khs6SHFgomF
EMKaNWO6h9oTaTm+am+29QiIL/mG+O0yc5P+ZEfzircYDRnQz2x1FaeR/eWNzE0rNvI+k7DI+S5/
jlJ8joUGZgDJBAKUvPZ75BboLPzOS3MXS9GoBUBqwr4pmM9NFouY4X9ndJe/K9VQ5wmur2HITEwb
piIu3iPAlO5mnRA8FgFP+56f1h7IDp9NsTD/814KpBzsutAVybl8en4xovXLu+KvX7Uqd3hBQuIZ
si2b922R45zS4dLLYrVxghxJYDJhC2vi0YL47V1HO6NduBEnktEQhr2MkYCKElMPSMM5Ot3OXSbr
LleDPcE27LoUDFpewuQfwLp+6Zx1D0Ctv+WP6Hqaz24yjsFBIUCgyAF+Ht/lIdnACiy+D8jHMf1n
N/IaYvF0YqyjZT4Y7d66HQCofy4cux+D6Nv57uxAUIoc/oOYmCIjRM1ECysU8AqeEQqkVe3rwD+J
pYiuvHU+8vLxo/+EmTmKaiyFVd3iEyp5jOcw5ByDc91oRHbFGqrrVG4aqz+1IR4H28ZsBTr2U++Q
pE4SzDZ4MGfFnbI3wf0/S7zQzieuEfidxRsGfgIJcrcbxdp+XggWYCBPl4qneejL8+bQL9wnSxCv
9YdX219U4wmrnBuZ+wRZQDgs+p6lCXRKG7HI7wihOw/6XmlceVdjWenYUXOuqP0miXSew3PsWJYN
OWJzlrd2tQ8GwOLw8RYZqS10y1qjUZ6rFcrFgJmmQvMTPaeRfMzBEJLL+2YhkDien8P67WjXWJc4
YEnANgHXVc/ZNcbxJ++h88UKzDjL5xN8vQSC8YF2xrqGbMUpI1cWdicxkkhv5Q1za/PEjWzuMok2
h9cdGDlAv5yX3KCcVV0J4idEfXpPufoTelnB4Dvt2H9BULgHfRHKiEmZO2DH4RcdnlnakHlWXZhl
B5MUgS2AJaWr9b7xeViyv6tXgBGY9OIEopnV21ba/+NXTTifGcLf81FzLhr+6fai+iFnyUSEwgbY
dzQPn04oyNictcYOzpmWzIqotE0gsiU4CpweHDwPhEq3m0FxM+Fl2I+5h3gkqpoNKp7qSRhTYCs6
y2e69KXmkBs0aMxqdiFiNEUfVYpW7cYLXeN/YsScJgRFpnLjXNwPDL02wZOkxZgf+p3d9mp7jrX9
i8EELba0/x/BLR0OYh6LpP4DrRgeJ+utktk977DAzu1OU4yrr8MmUI3JaJUQzzwcjPdgUwJJIlzE
51IW23Pec0niagE7d5eROm6iB5hXpBOE9kPjx/WEO0dqcYxwAzg0yd6s0QLDGrDfj65BFdV7ufU8
RB7JNLRXy0QjnzSuVsNohN7gMpJrEThG6qely1KLrY46d4/nXgjG3yYgm0yxxZ3z0z3RET1X0Cfj
7iLGUzXLc1lShUA4zboP8UutPT/pxOxjwBHeFdEqO9sLMbfFBhoPZ9Zzg6CCjECn+sxGGtAhgsMe
HoNTJIsJNoxK7q38jV7zIA2Xl8O8DTElOHWngrn0Mgrf3dKFM/TNRXhnQ5QVaBI61rt/cLG0xVtL
6KkzP4KMeuXTjR8RTpIlJpvx1jQeYwmm0A9JZtXZzySn7KpXI9Mq4Ky+FPouCPc7/E3Ta0Wf1yxf
LoktWSFGrxCy2hJZ8h6OPTCL/F64xhW+0VA/t2gwExgSo5U94JUe3Q2KqtU/pCzOrCQvp0joqQ82
/SRCvrvV9KogNJSXvn1k5Y70p5vrHAFCiozegfmi0KzchCvqux6QOi8rGJcgM+QmBPrzU8qaWNo7
zmbwo6O2WQJM562sKdu8/7qbDlgnKIbO9U+B+7lGhKm9yyjTgc918QClOaEjhN4iHtqFph9xjuDn
roErZNaIglAFZYYbi1sdaQ7/iFJLhmuawAo3lMk/Xe1hBxpsMOeZ+mvfJ7GaRsCXQi+HBhh/dCty
SdGr2nMp9CYpEm5zfyRUarACc+6L4HJiRtlkO6y1Prktyb0ucyV2VVXlhynbAr3qZJ0cikXvW4oc
5WNQYHWUcO7WwH2FQeeYVPxxO8trSN3dKs9aSWQwL+KUeMHGLcv9kByiXTM1DjljiHJ5OBdu8K5U
lxpwLvSrSKKDQeWwl4OzHaa2o0T2lNtcBi4Dfr401zU5BZL/5JXLK2O67OPN9axlH4qsa9P3w0EA
LzD/Bfh4MqWWuWCgHywYS3rrZncDh5JTYd9ym8qGmytWcpB9Tv4963mJs8QNWh2lMV3y+8Ryc6tj
TnXqXL/YOmFnE0Fjvr9qaLKGiXYhFhArMSZfzqpl0si/m8S7Eland7t+EpQfyjZuYUXQp9VouEdn
mUleXYJTpF6LDkhwGlZ0uy55r9rVkLoj+jzrxiK/zh6aPXWZykAuh3IFOUGNfuUXJecrgxEjX0TI
LwiLH6I9aoJMK+AVyAM9FlpciygwgaBci9MJtNqI8rVLOFGhNaD58QA6VMU4M7twqY6ImO9GFYFx
U1vqksHgYcR5xx9ACKMgAGBNA0pPipygBF3qzNV/jQe202Hzm8uNgeUg5V7uLN/cZ/YijXIWn1nm
eoRJ08Dq+r2jHRqdJo6zfdk6GEW/dF5oimGZUVYFuUugCVGpVC9aJc7uLz1lW6wMXrhqCOjyqRq/
MjqW4ve+tWiybdeSpWBtIfcw6qi2/0Hvq8QDsU//FGVG05jXGuR00LyLOT9DoW3Rtox8Tov/Ke8W
PAFO4/lLCA/FzTsNPcLhxR70ytG8mLc1vDSiGBJ/bCYuCbiWn7RHstEmTmUgx+zGD4j+JrNUSPnp
deUBbkCf0dHCC+nmC0TeYJovhAC0jZZXEgBRrLhp6MX0R6LPTA1KaruVeQZjRWf3ksSzLGVpueHd
uv9YSPRE2NEHthkaMJHpkRE59skyZzRXrC1THyMMlbzFNIHWTftFXO037nBOtYRudyTmFYdMxc1J
OnSkfJPnO1I1Oq9gIVkyPfP602aFqrAwl+lbiycRyfvE6By+5etL/IDtCTwH1T+HPtC0BiKBodFD
HMOmw17Zl3U6CX1oyoHKUSnKxDDx9x5c9MaQu6QJdEs/wTQ59d1aD3+YOM0oo9xCsNYctkL7Gc0C
IXA4UwJ6V57BVcFX3MVTEYPB7z0ozvXOvZ5GcUcH/lWsnH7IlCMt58jDgz0fPrn1NIFro9s5LLn0
uPjh89hdVZXF4YAa9s5UrY9dkXzWxMwO+UvtbbIjfLiZUl15LWtrmS8Adb2hI4bZasrwWPVobRv7
F/wMBZ3MeTRnS0ASlPljf1cJiyhU5i+VBH8AE+4Ixwbk86vOGx/u3ajrru7XMUUWRLHW7xdKDNti
QdREqDn0i3XchgCXjQB0nZqUZPwzDR7LMLRdY+vaE/CLWEZ/teHN2Enus69Hm3UWvsw7JRgxoEwX
npkyG2j3pJj83PwVF7mTHTlTAGYHQonI8aHA+ALsjSbCEUT4INJz7DvsW6oHIS+4dRDCkB7vD2l4
jf+8qqO1H4X8fiwVnHXVZUeSy4k46HFGr1E3wncCC86sr3ifOVrmFu44Vkac0VTzvTgwvdSSINyy
pSPkaKwtdwqF5ez71Aow8sMGujz/NK1h0LqlaRvpQre9UqpqnfEYy2k/kMpe96UFA2mU0th9vcyU
RQ6A7h5bOv0+u7WYs7UAVgpZH1BuiUGZ20WOhcCPVi5Xygh8lpfF6oEZhJqUvLN7cjwDgr96CjN1
uBwe1Ax2NNJ/Lm1cH7P3CATMtMSRu6Dj3dye9wNviP6v+oAWi50KKySj2BLyW1MqVUyExsCzR9MO
c4+wLIOwj25VRnK0sI8+Oaejw0eoTIPRgMWEixQJapxBuLWuZK2TsV+ptQZBmsovyX9SXskFX+rm
I4QlhfXufiYEMfwDjJvhLw3/3fSDiUhNGvlC5SZqhNXtAqfgBp9jPmTYa9jMGb+Z9yv4/MZkivM9
LsWsMRZz+8vTCBM8y8a3Isy16v4hz0oZPzYWIb+NEHsfCZaOKSjb5v+r9CZtyAc78GyUDLNek+0K
2c8cw+baavpkO3YcDYrNmHCohJ+cAhUSJ+TJAm+xqOIX3apq8n7fkL4DrTX9tQP3syT6cZ8orFpt
BVcZEqLii6DUpgBiRv07hl6J2nt2zH1HjvlfOwC+ZftY3LUtKBv1QVYfs1W6QxQM3/WNy0SLM0Rz
50lq+lN2ALRuYUCt7xhK4f1DW3a3nn2j3q8dxykvOcdJRJLNvuFQgUeBBXT3Tpk5I/YjIp09HtV3
McHzepsn1d1fFafLtlf2YnIZ0E7O/6b8M4HNKLsRBRZav6FEkAJZImagi6SyOUzRAfNOKpenq/jK
t3i4X+nw7x8ybr8vrGHZbCt2DG01xqQelECaO/bsUsSfQAuc7aVDkAOx8yV9tOLH7W6foQcdO4oK
EWfVdHwxkgY6kGEvImp/gSJvj0Eci8GcdlbSc9bjv+2USbLvzFEt6FomvZXtE3xLRR1GEgsQXTrU
NS2Md83zYDnAFENVrZVPLaeZREMapEBAOT+c7NzSp89JrwP6TVBe6S8wQtkrQVF6MGOZdPae4c4Q
PQ/MIV7ndaza0diZcg1FAU8FhejEov1YjwFOFvWqN6ORA2WyLzY605ej8U3rkVO8UxFsdJJLJ/9d
C/I8kHSQVoDr/PbBhuQzAvn7Hyy84VKwTwfe3ukLZtboyI5/RHLy9Wg9xH5SPtpH3QhaSs6RNTuE
8L9RZvi7/8NMmjsCZi5/C/JmlYIHRV3K98pnM+wGZy4mxRAjwVthcsgSCFGCcFqvZMM2unJgIffP
bn9oMtXXkoyVAYcuqug5emqrpdjnlwbaKEd3PAxwlD43f6D6nn6Ne2jm4CJ1Ztm53J6g8mA3mfye
S9MlAfILvToZIak05xCNKjsNuGn9CyYYnQUmMR+mTBBhwYtdo+bOUzPOSI/bqOqnO9opjQ3aIvrj
TgkUjOSgfyW8svE/bkMtsVA6XMAcXOf3xsV7uoB1i14ZoqbMeCYGNjQpB1na9a62wii6KIYTMxss
EXHLFWR3EvB6qKEUZhEj0NI1MGAtsr7m2Oc9dzt51fW6MMu2P/YZ8AqGXbPG1kx5sXeE1miK5VTZ
PBjwMYZnsL+Et+v2hSaE7F6BUbuLLsiOQaUZpLSRc0y5S6ozaQztaThyH9fdwpsYcBf0m4U2NiUD
ABGpzV/7i/lVWIJ9Atv49kQKXeACfQiygPYFFX4qHBhhWboV/C71ERw2MhIkErOa7RU39sAAW5+j
LMk4yyWO/Bnwno3MBR17Xn30iND+oriVf1DP6t+VP0qYB2/GE7mV7b7OjtTkYl5PypT2zpqEiPg4
w+gQ8cu3NudEf+MxmgHrk7WJPYLCg4SI8fNyQRY5R0yzYHYkgkWQEZiIHEUW5VZzpPdiKQ4ZImxe
gQ5A9YyzLcJlCGUFh5/MGej/N/GdGHL4xuz9MntIvNn58Wh7wG3YkqDZH4pmR6QNsVJmd66159f2
sY8vlHz3OsaOZ9PzgqAw659nYaGpf9g1NGmpENYW+1ezmW1onGyipyEIzxsh77GJDKo5BHZwR2WQ
ppTNMRF4RQazbyxCie4Pi41MMu2FqvP249u8b0wnKHTXfSoLM/lc8ZPWZ381cZR5UOKsFs/C6nkY
Quzrr8rjI7NSrM6EMO0Vt7PREL4N8sggGoMcwFl5CVdP7OVN2L2rgbtHDl4TDjTtwKoZEpsA0ouM
O/wcu6Och6YWFmo0ysAxID9wlZQldZWZMqFWgM72idCqLRXrsw0bLEuuKI+lRzy7pmHaMu3NDlv1
kG3R7KoScEWmPeWNO7U1zPzPxbU1L2z4w6dU+4CroB3vkp1JL02knHtHYe8SlQ0lVMSnnJIIu2Ku
9f2QXeDfB/u4KNhAkb2VfujCe9BxowaU3EHvJmIZYp+gmvv2XkwX/GQImA7TLrdEhpAT5N7Tp7+p
Og80EsxGDd15LYeXN/5O5cZd8dGdpBLH0cWFCeav201iLPmFArJzg3CFJSICFHmuoLyFofvBaRVJ
s7LfYLoaIBZzSccT+3J2Q4LatsnN88NkV3ZphzWLuosml+OJi+6SATLVfXDUcr2iDVch1vu6CCiT
oD4XRnkBdVrMnAshf7pVbrqtPD7DiwO9JNKJuuJIBlotlGuoIDypKDw7VcgOPuu6JIfBFQZ0JjrD
BLykAQU1HggNudaqgtgeVI6hoEiwX0DmJv6TfqFgdrg9ThVA4/XxdHr/43dXddjimm5tD/Y3aJjV
WEpFDunsmgpPY2o4gynTVwx+q51hfuoXnvmoczVtWNzK8OpJH1NQYlY9nCl4JMJArKnlwR2csRTE
Q+MYnlkKO5QIw58XCSMGTirw1TEvaS1UrDy80y21FmEx+Z7KKhrwIrRIhiCO3PJS6Wj/o/P6JeNX
3v202yDhUBPHZ8eCiNHIhk8AwI6M5ipnF/PP4cK/gUSzf3Pvt4aF6XOXmgFeaQ2HO/JIlHWm4V+k
EmLv2VfkrhRRGzefXS2QYDk+Co0yZqsxWoL3amu7+2BWXcV2b3MGlilcyWLf6Sd0ra6E8HYJvcDz
Yn8UuLSn4yB99NIWopuAUn0GscjYW4QUurATDrVcuX3IkXukg6jNdY8eVUP1UIyKngsg5Z0Qby7j
ua3GH7YfdVa6eAj5ehk/nYVFWyMhTVnwbfhSWr3w0OmciqHhd8rMj++JPsIqHB+51+gsd/qWdJv7
8bxyiTg2/GXZYjXUPD56KIM1oFA35bkjdaUBcS5Zrr+OYvU+UEzExSS3akcoe1qg2ry0srUTkxY5
mEqZxMyNpfpYaGlIHjpHAZUNi5Yah3fZw7fqOUGmJPNoKsnBGCQRBuTUIZ0ioN1cIrwXh2sqalRh
DJ4gOE9ML0cNMVY1LxojLmLJOAKppfd/QbyHP+cUuEhgg9cYOjPvs05svICI1WbNgla8959gbtJt
SdwHQEZcgfU4lnSXAP0SVTxcMvxKAMgBN9Do7PV1gYbJILUa/pAgCOKrclKJp91+ExXgi44YifKM
StUHjEn2I/gFB+J+aXLxSMXogRuMCwVSX6XZ6AAIA5RlQSy0EYR9+N21HhonGjkEOVw0jdaSwT5X
vDSKQcwjmmEma5LukiwZASJN/gGD5kx3aXPLMR3MIWcOYiTjEn+C6VuMHHyLdt0BloHXDRuHh/0W
4P1kkwthnDxwaVFMxwk+lW7wcZvqtKWz0c0Msrluzk1M1vFJgRMBGpwaymhtC+V26dAv3WME8meQ
gMcxDCVsY4bZn2aK0EnDL17M+uIkMmBTsl8c+aA4I2ap3fbb1163FyNwK5ppL+i5C2n0IiypCo7g
RsK7Pautby5Z4xLOE8xU5vL/OCBIYhhivbe/35cP6PlfhvhdNQMIbuj2ZZjmzJPYo7AT718S6JWd
+Qb6eTr7L++gYCfZgOJOr4rjUFHGV6VpQvmJlOo3ZJadBHDMFijysZ5OyR4pMmpLEVXFMmtYmJqQ
IqVD0VbGZzvQmEmnHXMHIHAohVOuNOtI0jCO89Ge4Djvx+ecwXkTqluEeIHIDeAAb6csp57xZ7xz
8rgwwWSwNW3KKSoUx5fcmBJel79YH95kiiQA0fyBSJsSrW+o+EoT07F02wRsKBb7G+VDACezYqQk
Yp3+v3A8o6l4QHPpY/O0KXtsg247A6Qrbo7q50+CiMDmvlP+D2H2sq8vRZp4KOQH/kiSHuM4DAg4
stFC6nyVQWJUEHqfr81TrSrsa9INMhPCEvbL0Vnm1/he0D9/n2/uV341WBvvJZvJ0PHyvQvBfAaA
/7mlgjtv8xpG/l04jr36KYwO98u5+W7EbivAhK4d747zusryzaYPpJ3fHM1lKgR8MHuhlGRueMkl
HVEzdFU7Ad0CRonEnduoQY9klAEM9LxrXtfeU0IJKa5M2HmrB6jCuAoN6z162LcZK+goU8MU5O/1
CIkkqQeQbiSl2tKZt9BhmmyJPfiujSa39rfJtamNnpMI5O85IWOm0dUexo7GuIbdxxxNHWOiFPUs
WMCpfsmYMjf09j6j5hKgJxZ0AjM8pt3BZc6btnveXbc9hEK1yrKDXD0HRJ1sYnpItbEnTamoLidU
SVsx3E7tEja+ldX5kc/4S40nLuXVY8SYtpNdBWFi1B7iZHa/8p13BY7zgruBx+9l9D8A96lLIeNW
fvBVe/xMUq4f3yd9fUAQDp2lnwHACvtf/aZWdluUvqquhUTSphSgONkQ57eQ+p0qg+jIdWqSSkR2
SRC8Xg/nJmeLRCQPOjJpDdhQttcInpvCpTiAIXZgC1ld9+PelUXPcTQ1Fh/BE4L++q5mTUHdiWYI
cOFhi7pYSKdKF9ndB18ETY1qVpdxkk+blUb0EeUfKPkUfsS/lhKzlwsKZ9Flq6r9sqbXNqaGAYdh
JkL45AnzK8tCmyEo/q7Kb6hqLdw8Yu8qIeA+D91WZPExdYxDItn6cz4dXtiXZZ/+RETFldprvN2C
yH/PQhnbhZcg8e/F8vCP4E3xxfhSnDM2YNgGnxqYwFOrFVqzojbR5IXHXRW6m4JjSHnnm4KXyI70
xyonyOLBPHzcpQt3SG8hBJRkoCeM07MymmeWQqNxc09kBsLKXeTIdNquF5PbGVZgNEtNnAAJu2pU
YTZcja61J9tdDk5Im61Jj3Ouhj0GvbkFRZNsf1MTbzOEityzT4wCm4pm/ruR6EL1q49uMSI69w2r
gXrbODJi5d9HQgJI09XRDd1lhxfFNH3H5kZGknOScWi66XYL8FS18zyS3N2k7rZKAz2XgoGPXFMJ
fX0pWD8BVXk60f1djCI8PYsrZhOmK7XGz5qBrRw0iobi9DTR97CjpLnQlaQeJEKIKu7dD4H+VFLf
dTdtMy9t4HVybUnRDWGKiWIstRIODyT/gmaLeEKavo5QQPlqkR1sipRnSuOJHnJO/TMAMKicGzFC
bugob+/IMpHLaFRtdTHu5rkFFIbeHAcxo1cX359fB2nygDE6Ek3kZDa89jJUrudUcoGUJih0c4Nm
EtfeLyGuiIZqkCTjiK6m/bO8lfsRcGncEvfc15gbOtr3ZTetaX4fFLQeL1Ji6qkbz8FC0nrRvpbS
kD81VuPnVMIDe7hoYKVF+qTJbSnqA/LBrGhSVOuuy3Cq+3ytI7qQsYze3JI8KDYzCjy2DEnQYYzL
+dNnQsY0XXyQZRIRhdoiyO6ZoimGz9RGonQMmF9KLO7sosP8c0DV5kqkhC7ACDX0Ag2DucUc9vXl
D99ybjtFnXbFGxhyUCsxib4gJ1mQUpKMkZR5oLmSPGLMZg+TJiOtRbcP33CFrRH++8M0lpEMH6py
D36FpwHU2PboqB/W/9AwPXS0Rocct6heyrSg/Fa4SFtt7U3H4bENixX0+c2eJjdQQQS7ZsLdFsp3
iqRPsuTinsxepvHz/nP95eBQMS6WKrQ9LOAMSIpHxKSbRwMRqb/krWXJKsTfVrYUC1iM1qW2eg6L
OBJsXv6ma0Afin8hDSih4yNNydzW8DMVCzS6ipJxDHW3iC1/iAy6QhPo8Ce/YpDGDbwwNdJJRH6D
mS7myXS7gIXU7MF6HtAxcXPpr/FRE7P3As0IfMF9fIhBoZQAMMmsqOK/eyp46h9hae53pDpgk52p
TU3LaerNYILMZH0UQPSemvM9pMtmmvaddhwaFAr3v8v6Ka5MIc203mmkDLI8R2RsBHsIRZ9uj4NU
MdW21E2B/M6B3//Y60S2bqI0xHLlqmVzQLroSt52S0Wrhfasl01aLTGVq2ZaFkYxl5wJpDC9UDsq
JafUHM19nRP7IJ+qWWM/eYX9lyeXzc1h1yk9X21JnEhm4V7at7e8JyjXVPR4jYTl3nOnnkBJX9q1
60gigVaYv2/d6TBPgAPGBXTdUWHoCJ5autgNp7l4qVJuF2rS2mdyYt8GBqDAJ9JgqXwEcrhZEusO
xeE1x2u+Cix6Yfn7ezqM4ifjfkY1WON/VOrLArh6JMdCcJTxm7fAZaMB5BUxZi8B9TE0uQ923SDe
Uz9jJiYAWr2zCqDgU+8M1pN1MBgawrCsZp84lv2FZ6LQYIuyeNuahaQ6oSCXzieBuRZ5HIzJLuJa
zAU4rIYMnKh2XVk8+yRUzoHHL+pvXDuW9Jk8G0C81/L+UKN4EGMwh1qZVGX9p5GtjE6dr8oH0/AX
hVuyoU9QtRbWyqfk1KqcvJ9W37mipC8NQcGm9hLzI2o1H5yUX1MLom4IAmP57WhrVD5Dxws1eSwS
2jigTLLzmyMlRkPC1f659O2dpWLCqkHJIvmpHd8mBJtQTMBsvZk/5wznkUYy28ATqV7tYc1pz7Ye
lmYk9D17SQloyCwSSL7ZiQYCjRF4wDCLr6tFdOvK2K3qCB9+tTCUrdZlfcSdFIdt6i1u0AK/1nkU
QedYT8KfVrpGyTfdGK3/d49ypIxF4QIGcGY6GVlQVGNKwoQSBrkIcgUcWqP/jAHwqkUY+D35JwUZ
PtmAaSEyGQN+ahUcQ0gpIkI1tOcCGhSw5eZyd7aXPMTvtdHB5Jk6PtNfMPsZSY96M9pJVWN6rshj
vHHfswgBqSakLPTIFoCm2SujqsKHb4wGESHJMpIm7k8VzQFhAJTiXVci1h/w+dK10crtMIcfEYL6
d0d/hWm7M/KzSR+dM4afTao9GFilq1S01Outanf+YcTt9GJwtfFHLflMJiDxOzQgsLc3piMwt2CL
7OashT4FRac8dGlIUXdld8Tb9Xn9lEFmtklrmDpZ9bE79VESgiqTxSGBm/Zti7r0aHeP+QhFPr+v
r3M5b9HqSGVCRVa4JgcCkrt9Egn6rfQ1NoK4iKVsrqlk42FUNZb6jaJqIXQhbNPDPdCaBHKYOtLQ
ANRa9hUBH9qwjuduaEq8huAbdSdoxManzLxryZKCt58iPZ3PCOJOzRDzdecbtSi8u3nYe9/DLZy0
/noRLW+ZUcWpFTsJEAayUjxoBHKbWh6yjIeafSAxcKXLRfF1/7tglH0jsw/9rDwVZdSlqp5JAjw7
8j7kjUHY4BQv6tIAE4ijeuz7p/uAgEd7FOodIr7vGQCBY3lTDMbcI3UOf1Mtbi6M00rjITo1BfxB
pMgKDpzH7X/Ws2GK0v3GHdiHWZAGBHW6Y9vIWkWyDa2s2rRYGOoCwf3uqOc04JP4yF+z97rgqLEv
J0kk7c32X4/ib6MJg+PGkPno/YhP0Vk+ZEU5A+9P6mOw7jnDSALJhMK5NGQJqbh6XS1UxkeGmAIO
2Pymz4V12l0CPHXPSWbh09Ob0kiDL/wDSq/KX3NFZllAMtk8gR2kFnOaUFCK1AiutsVJFP29s7o8
+U/SBrCJxxLkFo6yu8GPB5asYAWCnZgfxvVwF+yZjmfwlQKqo72pPF7d3CdjaEuvNVEbGEEJebEg
pjSi8d67Ck9wl0ZmeR8Jys2Anp9FhJ/uQpKTxq9QbEQqCSyPOUsDbPWPjxqSMC/wFzeILLGsbYRt
UuJz0kr10U0j4NUn2mtJFF/4YskyDIgq8VsHa1cRBaxY5n62s2FNN7XyxKdryEOmwQe403m/bj57
oiEtAdcTmKQzNTeNpmPpS4VncvvJZlFIoB1nZAqmR6GXyR5Kvcv89tB4etTPArUK1j9TqPomyC0k
YefzzeU6tk4mj2WI3BOFsXtBY/qianZ34B4bF5ipx65Om9dj/t/tfJ44yOXnGoT+UIT4CfwheVyL
K+AX3vVcCYF69PltiKT3//BMNaGmIYpPOBbT6jrZPDhq+iD9yKUJ+K9rnn/9ZKia2ntm6Fatd2lD
7sNYY9lij1qvN7lJ54wxwbjo30uut457Iq2nz/2WDOm3laMH8zbKVe1xBE8rKSq8sck/4HuDd1WB
bPmUFI29iAAAxa4PuZwfsiet2YGgfYVNkb+6VZrirxh0aB3G6Uqq7/TJz6gidOHdKaoTSui0jXrF
rviNZZ2ugh+xgy0sLx+rT586zVMnzzQWMJQgQvrqSCjQ/5VoPEq9NtJvLQ5HFvAvwZs+27lXrkvH
ljq6s4wFTYFjbBDVehghBCEaxZsjvu+PqH/aOuFOmw93TeXx39WaSpnbHB7ZKLyXOEI1mnbn3h9Z
jMJ7taWJhlVDGFB9CTHtQ4h6B9AxhRSbfULCZZoIpJ95O0fA14Y/TY4i7oiPp+yKbsuIA9VdhO5T
Yr0syGXjRCjAGLzWPlzcdtuwGb1wNu4EwZ+EfI16+B3u1vc25dAoQKUEqj+zzsH8leClcYgGQ6Ua
RwR5ayF6VGdVE5Te6+pWDn79pIM32PcExcXwe+t56um9UMDtVxie8eGyFnJGxh1Bt38kKelt6u9Q
79GBKXrWizRRLhFkDKatDcskXGqDlIbqNfJXio7V1m8poQ3fF/J0GhUP1DNZS5Qs8A/5ZQCe33Ve
4AcJ/RYhdJM7cNFqqhr0dDK1vMmxD7IiSVKcGBc5yTvT3fhbcZwFsoD5NZL4SPMIUvdO99rzMBZ9
wYEsKXBPP1R24mdsTr6hMcHSuHbzKPPxx27+BUyA6fM2fqZZpz04+q9TCD8ECOK+ZwJS/nT4kYjW
L9xrKoYS6pWAUSwPD6sM1aZqhpwGF1WqX+7UWrI9fv3/eimPyuymKA4rvAhji5J/gEWcTuj3rSSn
StRkHEdQa8lVvAEPyP798it91BAwKCEJvbVtg5tLUnPBZ6H0esQPLSYCAyz4o4vW8+uRb6CpqaNJ
lc+rDvzBoQ6yVKx6zTyxP62YEQjmywrx9i39v4WBptGAhuB8N0hYrnhbcFIpCFeAfRPbQSGl7nKS
UjQ6/ttRHIevdwnndvCVCIMVWQLgfBtxQTOiagkxOnuZKaASOagGF0MLODPybVm6PxhiVNWSe6au
ud1pXWUuoD5P+Y/zMf/m7ubHx10isjr+kZHyeKiTpkodLUw1J0Fstrd6jlQJ/i+hgt7lXwMXGdVR
iQvIkyzJ7wbKAL92y4U7hdo3ClwNLS57t41f7pWGApWcRNQp60ofhZzkLvEBYbwquU3y8snJKFlH
zFf61qeszBvVLL7liJRClY0hp/1vWXjxSaLRCZlK2GEJ5ImbCZ7c13PXKyD1LeXkzByg1OyBvjJP
rXpYlCRaYC5MhHVMDypy/AggBxrTINGhFwMZ0J82YhKFEE8AULx8gyYGYoU7/o0NRiofirpYzWp5
Bw7wDGP8dvD0Wlc0N/X+K/ELtNiOe4b4IDB92pJ/srOgOHISS8qBpQxfPa4VmeyPwJD1I1HCXlKc
gp9SsKKTs1jKX+O1Z1WEZWB9RAugCD7dj6QzHXfnsWsq+ABb1UVHO5ZRu1UOVhd4BXPZ2DNuCsHy
tfcViqbSbxiSYF5/uV/AU/EtLlQq/xkxYAQTWeWVz5yuC6azMZr/YaGoWUHhEtgcWpGtv4CubEe1
VfCMu8Ny1mL6adkZR/keDXDexzPypO+LbyzfrhE/h4/yKpThROUypb7/cBQKbUWKukRQBefP05PQ
2HSqVzathj31JjHxg7D8irCb9RaXD2gw3jddQt8u9isVr/qp1+h6avmkMT6uETbLOPFGEU1lzg0n
/i9RGMs9o5OjO7P0SuvP8PWS6JWPuY9y0uhs3WkyAOKMTdI5fBUm1ZJN2TE2I04cN10Y0ewrbpo0
SIZwJvaHnj7JKrNhpXr8owQoK5ZRu4A4XuxegboQl8wZFrO9mSaA7oxn3HjyFrZkkdgkHKdr1OAh
hNOGrKaTVAWbC4YZuuuep2nrkZtiq5tT+llzuPK0h3v4zczkzhqaq8Y2UG6Mj0ccVtE3uOV1e4CV
fefU9HBGfgAHrBLTso318y6vMfT9J1UksbSrH2nTzGm/YvmSFZiVJf80aHIuvNYCx3r6XEJtOK11
1LWy9v3QXNjn0/nZQQtB+qFsN3Fy1tkq3KeBWN+3AESsn49SkwaVOhCt/8MAEQq1X1twCT42+fII
Ju0ob53HRx1QVs7O5Bj3uiXe0Ur5rBgRU/qPaB0aSDnTSWhpe3PhZFb8dJkEZP9TV3U7wUl0qqb/
717v9jD8+1VT+Io8XqoeKeLSRIBbPDsJJf4VR6qWFGpNRRPjAVaywPNrrUm4wT5KuBNz9tOU0wdX
+fxdB73zbnTbOWxU0J+5P64hhCp+vrO4jqiLQzNMipHddNqRoG14sCmB3W2Q8ioRlXjeIF3dT4gD
uJGuo+htqKNNQ7KqT2Z50WIBy5REZ9P63/fcT5nJW3ytOC+gtWyHqohVQ+n3LSWJdMY2wQaFXjQW
dAy8UgUd7nHWmHPs4xghGNU/YxCb6KO9U/NCUl4I8iRg6nUhmTPZTv8h4gMle+nYKiPtDyzGIePx
LaKXAo/fhOloUrXni+aKuaofEFmfUOKS0Y0r1My50ddtY/PmnTqFl/q1QdcoCOyfibtRNrKR2BNI
Bfclooj1Bk7pU36LIt+y+ukFcQvg/w7V5wYFCqFx2d3UbOY3FlvsItsU3F0A27WhjrjXoafnhrCy
7qx6SCuVBg10up0U22UnoaXgbvJBxhSlLdqQEwd3MUltceyB5BsdiNtZGcBP4ZsFIAzl03+Ea3n/
lISY3aBB49TkwXnbAE2gJ+vJDRnbX8Zb8AW4QZwccwKHYDAXSqqq2ZQCNInF51A0z1J/pAtz/lcL
HGqCqL3C2eS6ZT2d2nueKlzodxPsYHORaFJTuTiXEoZXI9bDqtTzE2TRcbMgjqbIkgJK8NPZyE8e
OOmVqeQqetn7ew0RRftyT2kNiydVhUkBQu5xso4hbgqBY9djKFLewv4ssiOkUKpIQQXxaRVw32QJ
RjeXNUdUj23lEZYQ9KwQRR9AdLMyLwH7LrYG2z2A/HunDPVN85lgbDlc9rbatcxYN9v4EZbiDabN
y6EdbuLq7qlRwuqFsX8D/n/rUusIO1wOonC11JgkS531VroZwTOSSflzHvPFudbR5zIyVAekfQTD
sVANtX6m/3dnQEc1Fy6Stpo5xE7DqV6XoeJKQzwpAFBVyJm+Bs76YMMIgdiPemYtv3cuTAlqnKPw
HakXD1PT5KUEv8cCMwVFCGyhswJBT2Pr6RZsUMfVyTSTr+VF9kU8rIzsmZbpL63qfRVAxklOBUoi
migGJddwc4SWfb+CA7OZX7F4Onr7Pf6m2XcaW0J8Sd4YRRarxDSSLS3Mg9aL/erhfuKpOl7Cc1Ke
/BZsWOXFo4kc0vj2GBeqh/WYFC4kAvPak2A5uUXt1V/kYPzNKg81QshHZwx+DD9vlg+0ynR4XrV3
0OypxyDMjN0YA7LqdII0s6OaHQUoTST3e0VZVcnOmX9xhhql21H1E/9A35G+Hv0HCs4ItDxlzm9K
uOk3Ffk1/+6K6HvESt4e4orX4zXSdBAZh8Hs6utn+bmezDQBj/GuU0DvrGxn4P3tz86HXWYamxs4
IcDg8bMuClEe7BiixQZlI31byBlFCi+mPUYndoMt6K8SW9D5Tjg1i1Gh5fzUrNasPmj5bdZ3fZpj
GYliQtL8+ikpAzDOqWmYXTzhDhbyqmrNled33k2t1l5BIGhLTI0fh1DG1zawwMyuPUNIMLzuPA58
/w22+dlEPoZR6JEZbutQufJSC29txud77RWh1bEQNb5au+paco26DHcnCpHDVwRsOF71r2xmfpVO
4lPvwjQQXub/BB/Bvek1i4MNFt73cIQw4HrpyG6VY/s8bhonPWlhdOZ4riHMGIIcK+ip2DvDIAg5
+gLuwg7lhCUSEluiLxP5/PBiVcfS0PVvNIObNcQXZxqerOi184K2cHBk46jeL4HhPEUXaVvfY+78
pAUBXIIDV3E/ZOLHJyiZ70NUHbZHi9UJ/ZeGaXo1CyliewHth9S3mX0oEsgkk38JO8nt5tHXF1Pa
/ckbNRWHaoNVZbj1eOKnAcZ8N+RfUvBjMU64Q5tl4/zzLDs3N1trrdaEN1R2W+9usnRslUUeI/QK
X2zI0Wtpcwa9qbKdz2Brrpixye15aqj6dUpYAm8zoZT1NdIcIK7bTDl8Mjb7yAB2Z6sQ9GDyiaX3
pdQRfgr+ulN4S/wmbnOHgKjoTIHBG+BLagq4fBaOyD85Dvx0p4VKGVc0/6qv5Vre5g9HW9Kv36re
nIjnl0Dkuks/CPRsgYabnCS48di9nRvXbS40zlfOoj6qOfK9cXYlhx9HXUJiv1kSexCpASvYgcQs
JNoLZNvxKz5qzgO0lnsdGgHZF/8+2gZVvI3slAkj+aPDS/NvGKcUMSnjBoM3JhxaAamki0DVzwFO
5IBwJmh5NdMp0iMWHwLXP5tlWGDBGOeIAbasWveE5AfZLI2SnFIG/GPQHC9yRwYYqhnwmBZHx7W9
lqdQjhFBe3f+E6iPEXsn0MSdIXUnQu50pXBmYt0glXUsputDsZsQfeetrNcbzNSVUdI4wqQqNBZO
KDVHDsGjuSgDNwNnGmtdhQnzX5zvw7f8tq4FCHcsjxOTrGHvP6j6/kl3fW+HFsC7fNQn7gnmfeNB
E5LYY0Q+58oRnK1APfoFFRqP2tkExybdaQ69i4eYYIqMKdtxZcVdyhR3m8N6Ley2mltaQFql/+Yq
yKHZbcr8zf/SJ0vfXAPv8TWUsn3qfhH1m4hcthHdxpPPJeKj2ZiwAqXqyuLD0B1/Zbn8xOwjNzPo
tokmhO4dGmHYu4yAKu1wgSx6Md1kjLGJVP3gEikYTnKvrVJbiHKDWgUdkAgIHB/s7qSSpx9ANdjx
5xiZ/XJfYmAo3UBzOsBrJ+RlOm53WeHK4I0xEHIWxhqZcHXAFWC66VPBU7UbGf4icEzn2IfaTRHQ
tHiHZzcvyFaeISo4/ghX79rPEs1nmbuljkFAOEICNa/SLKEYzJxkbJCNTJ8ScxdmsSd1eYOY6WVL
V4n+8nwMxALS+LH8i+mVwNM/mtacu//nRWbLjMWbOBkvd/Z85Lg55HYas8IszYxtJFKmuYHm0s7h
pTT7Bw3Ye/+mqALYbobBk640csT8wDwu8MKKL+01y7ZvR8ikPE1Als0kD6c3Q/KBgAu9HuNhWWLn
GD/uD8Q5rMN4llzD+PnKMjtsA0JE4UMBuXWmyRwjcj5KqbTTOiQYa4QMUeorUc5JGv5tS4IrWJpR
SsgRbxQ4ZAaCER+FwgEaCG8yfqAErJJGcM5ocRrbBgreHqwsgOYd7bJWTXvkWyCR0r0uklLNFhH/
PLMViy5a6q6AnegUwDXpq7/blR+v2FVLRfwnqpksI6XEC4GGKGii+0xP043+LbkT5nLGtsJ57T+c
OgPcBh7qeMtd4LRingMx1t4dgrwYS9eRMmc27BgW1lOKuwV+Ym4dMvvzwshGda6g9ar92DT73JGZ
RQzH4CUrW4QnNJ5lPz1aN7BJYfVfzWgIzL6QneFOuC0rUpAW57BxMn8Mo4S1MLV7yaDcLvQDe1oK
OefwaUgSlJnD406l84mfI2wHAKXdst1aH2Rg+LPeZDdNK+mY3qbXdewVpCPhHPO5z/IuJZp1aIF5
2EzGplcvguISJ4tB1UCpTWflMrspqZ+5nySixOx38pBM6+HUQ/xwX89HIzsb35mx7NCvczTxaoEy
XpDNgSYuaC+90NvT5lI5axwB/qO1eY8KtT4bhUlIVlXXLZOFSol6l+geE0yMc/eT0NdypE/vm9xf
29AeLecCUjmt2Fl4LVXQFhyhaItNqvXn57GHZLbQnFX7kdbpvb+7DSu4hDeWN5wLv3GO/5hY6sKN
kb6YHZosWZVhMKMFZsrFM5cRtiNT3NPEZZu0nQdKgkyVabZkFHDAGDsnSaw6rmBABiOTJmIfknzh
WTEMMHS6KFsMK6a+rCIl/KrPHLT87E1cYrVNektBEk54WzKK/NwoJIOjaBEN2vu+8aQiKS2zXZmO
dAsCcbbqfxgNvVoLqvN0DSnunnSVNc6Y2kuMg15FbdLsb0cBLd5NuKqt/MqDjiPEQIrwsqYZqRgg
AqmY5wdzQjNN+UWyFWXsoR/FFoxyJsh6glLhGc2QhqXyi38L6pzbXObk0/R+F7dmv/cyi5tb+G8Y
B0vblnNt1w5fNP/4kaM002A8nRHLA6b/DbZxa1TbX4ObNk6Akpg1mRVi/jQjUf0jBQPuAshutdP3
XQg5v+lW45oBEti3xrm7IwC8pM2kY61yP+VOj9Rs3ROXdZ7JYBKkcwk+pqi87jK2ZIqHf6raGgXR
aH8+sqb9hG4sV4vHrH5TTzNyxbybCrB8Fx0uCHXbrA+Hcg8aScorsDZm+X6R+pxmKTJP8c2a3nSJ
e450PI3Jy/BboDtb0jIT9jQsRRNipzPkCDfaJgDMu7cuCdRVFi8K4DBGsENBqiYZGUz5J8WJ9yCK
Zep6aQU2k9OX2u2FhiVQc5evAJ19LC7CdzQMuH0udHYXvmHvY4e0ET80iwBpnusRXOx9utCLOeNX
hV0GNhyygQuMZl/MWn7ljAsfkUOp717HVqVmggIKywtUp3PPMXJu52Ezqq/19keh1BL6SbMeugBo
GSsM+9OPOCkGwBGA2Nyz9R9CD7714hBV46ituX8n/7VId5CiolI56tL+fDPjAAhW7FbSZsu/rRJD
dHJkZcVs1Gwgl8Pjgfb3EjpFUDIkk+8Dvp0BnFt9ViFsZ+7nP1WBGMf1QORZvS2rYpXdATAcm7/V
ZIwZoil23f53w/lDn0wRaPCChakf9MJDJku5UWlVmdsbTEyJ09snffioOmSOtRU+fhnFjKi8hAHZ
DqSPc9U4VnLs1iT8fV2KMLpmIk/3Qrod0mk8cnzT2Z9z+pgP1UyRKvQEiCNEdeRONC9BrdNfVQsW
dxatICA38XCSPeOBR/mmzz+Ku5TcZ8lc87BPJohw29KYjdMXAFvpYXMDPcGWnTji93U+qUjlwwOf
oiUJi7N5hf1ERCXmMu2YX/MYtZOsxaUpuvGA9Dlpmvcf+VU8Jynbgy54VW8dpcBXWnGrANp2dj3S
PisgTsegs7XXkniFrACCJOw7lkK8jaUBLKHKy2qZeCmDw3bVfqJlVj9DUS6xcBrDPtVxoah7UQV9
iPgyHtGjdFr8cVyV+CufsV2i0V5z8KEYaoNVXJysjsPmbp5XHry6Xhar7sBU2sZmrMaT+bU/OXQL
AQ6+C7r7ppfHS6RTdqWEj24P+wTLHqbehrmiGtA7GjWJiPD6u4/O+ZnpWdYla+ifiYJ4Zij2m7ej
WmY5ErOxFhlJqxbY9TuB1qlyMmSjmxzJH9efj80KJYHYEDFNuExbUjp0/db8yqm8jD734iG1Lw+i
j4jug7tAFPEPBKw8pdKkdXmuNdWJE1/j5oTcJQYpB8Bmu0iZGyc6/2U1G6blRzUpRSQIq79w7WIE
Erku1Y5TRAesxqqbw3UEKL07LGU8/uhqN7dTNiD1azrfWPbSkvzBMP9LjWjNcQEQ8t94Uop/4w79
85NBPTgkRfomR1w2ajU6pV57f76eUDaDmLAHt5lyoozoyOnF5pPVnr3ytkA6u6aaUzIQq99LarPl
3UrnAy4XKXMh/fd7a/G0Xdh0Gxi3Jc00YTxDdWjn8m5P9PigEeo8ZVeKYnYsXYwcv9z2ntS7tH/q
g1rkTGH1arlnnBO6kO9YII145j8N5GJUcOq1bs6LokIgtsAqV+/hLaii0ILW6Bxtp2zJxAYmX9fU
U4Td/00cREG4fsAlFsitY3xm8oGJ6XEwE698V5C8jJj1onBDtASMxs4yipG/Cm2T0t1Dctd3VuBN
JMs8rfPQv2YtbXQ4+FGDct9QXyBY/DNa4dqDHsVlYo1OOsfQS8kbQjbB/s21Tg1DWK7MNc1dEgds
VAHW/t1EXN/NqSKMjr6bjTOWmWLulFCyUpljEqssOrXphmpT/WTjHpWhleymHYMlyTuPmoE61qWC
BCxvlj1pVWQHuWi3vZOHvpzMJ15yapcR3O+F9XFIuJkmOMdY2CHQpZftOU1wiVwDs7rUHxC2Kbqw
q0upRsk4lwHPWCFOHne2rqrpxEt3aQHvpOxTVup0EEGBu49qghdqixElwu7AkGtRgrTND0ghhdq1
60GhA2HWlD68uERTxVaifvKHyM3MssFQBxNYs5VyYSyCSitXaMgXHdWpEb5J7IssvLfKtcCKeu6c
AcCOsI80tjXvJq/aFCBmmWUW+FCTzoWNLem5nJz1a4YtYAxVO9617kDiKFFnMl+9p+ddIt62zXe9
AjF6J93mQNMEBpwugkjY85Bccd+mPkwLlPuD42nw0oXe25Mr3KPn15kOZEu2WjqIrCCQBGuvXXm/
a4tEBYAXyxFHRfIt5jRkHw7oYMlzFOiHDrL985ZOYb24FLHxSeCp2JymCZRgMVtyN+7qVsCk9wwR
SaB81uJErP2CffEuWSbOmiKrv7KMxw1aPDhb31d30woiPqXFP+VsMmLXvcXfgmMBn9FJljOT3PaB
8d9fsE/Kfbhi9/yKJG6AEy4rpjudvA7m6xSq0i90m3/Q4IiclvLqJudzQR+y81ppPJlBUL7m+ng2
+LYLrKZhzMO+IQvZsL3kTNvT8wsqZvOzm2ccpsJUtJ7g0U74neyUMpFhPhRKtgSR8wU8ggMrJHaD
sF+h+aYl3ls07WTY5Ik4xQQnmuByFvYkpUu32EZVXJ0OyM0cgyniyoTo6B+U8typ7yH5TUOI9P+F
/d9RswUzkXJpZp/ki/YHy9yowmZ2fwobVdXeHbCK9z1dQs4EfYQcAuY9PbykAUaFnTdC7CR1ebjP
fx2Dmo6GJxxbt1fbEoJ3LZvUfoPkLekb2TlEKeDfvqHUjNhxjTvoj8oi5S/UgT1NlnWNIUEJvPRl
lawIjexeZ8iy8/+iQNF7TkYNlQum+Zy2yMaPFvMYoBa3yjk6aTqx0+wipveMSwumbllyOMw3NhNV
Ry2P+v1bMpaR3h9ekd8UENqkDpreQ3czeWngIuTvcIpSlDUY/wkSSAaz5TorL9rAFPQKKT6anfu7
zB6wlBW2YbiiwXBab0IQepTCxGoFc0WQCh/uZdgbPx80K3vuBvYob6fTR6Gtb8UM/GAtVTbzTaGp
cMK5+gNv+O25S3ylPA4Tidao9t6YUrM8KjQejfaYcVhAN1Kqj+WYwm1cLX4sBZuGWWLuMOjqFxSu
Tq/uTyT26Bm1P9/BXIFVGHYUz/B9qa3SsUZQ9TVKS6uIctGXm5vgbp4Z101PHBBn/AJ4zRhJxRXI
gMR86vx5cBbXeHQk1hfTERd0dadCSwTNx5d5rsFP/xezAa6Qp9dKOB2r7obRyazFTFP0fCVUESV+
ERqDF/jPAs0S1wXpukfE8rsw8THzxj6p3GsC5qTgNlnp/ntk3LxeV70Lu1b18BVPIjcAtZzJLuWM
CwpAG9yKO6KlIEa8ej177Y3DDJjV1ZG6bazda/NakdyfmPt5IwlsV2HPXMEUKJqDjGydNj1Vd0bt
PpAq8mBXO2mcsuwh4Y58yu9NT2DRhRJPVX79q1xNTDVCQeP6ubHv/TCxsE5AIlOh/cwEEds+LYcL
lSjKwKqypYn7+2JizYJMQ25yqfhRuaLfbWhYHu/eyE114/y9kYzut2n55IMu3enng6kRe2r9rUcP
5kL8ka6rqUNcaTVCa3KT+m/1xcUoJs6M9UhYfmXAiY+b4ayPbq5u+AeiOLWjt2KE5nd6y/1d0Sbd
xRpdeHGkZhSKlJHD36jc5GvxwbcER3e0H4dg3oLJGiEw609hxCzFmes8F49fSFqNXk1brJgPxZEq
DXL+mKh6fEpMKhMqbKgLsUDyjjv20Q269WLtK3AqDP8An+5OFSz/UUven9eAOXsKGmaFVE89sXx5
9Ehyi0kn1q/P2sFc4zZyNPUpDO3Dy6d/TCG+0GQsliOYRcJvcU7Sygf69lID0SIfph15hJq60rtU
DN0rzFFuI0C5+oKmFdEwic7BKA1dIp76kI8461/r6ovLgPTF5F2+svmU2HJsAoAJkQP6OQCqSqXt
NNWO1wIXRPM+eJbFamIVOd0cgBcMB1diym6KouRP1tsqeDB0ZsB9f/cQHcKCrbGMNBjpNJPsYtwQ
OboxJy64NO/QY+8Cbn/+8yc3M+BqYqLeCpo3sHlE4b1fzC4uB5M0mW3vFNJ7hRhDRqb2acdy6pXh
Zkvw1omIgDAcdTUx33MFY/L8+qw7+0wfXPDD7PQeo2CkNXek1nGm4U5Hx/b3FQrtXUP6IsAfMJ2w
jYcbk4YSiOYcyWik/g66513s0BJ2peGJLMRE2izuj+3TJODgZ2kt9tpcA9NdGBd3yLHZ79ZwDs3j
180NN8QmqkXJD+8uKijbTsblWBG09lPoot4yyvuzu3/xTLLJlRodkQng5uMDCDk30etOFodEw8F6
6c3qKAWpXtIcqZlFzrPNfyRclBVJB5duhjQRP0veju668G4YscIzNJ8j/r9I9/K1czYgR8HS9kg+
ypQ5fN7xMe8LruYa044vixcJ2lv+OmDiczy3sKy9eYpvV5ECei+D03DwhT55git0Vrxw5pXN4RPV
X27EOl1QpFlRPf4Eda1pQkVdPawhXBnvn3FaRwGKMgXxusLunz/NhFJLqE9f3lt2f4K6AMCxAX5i
mnH0/+a8J4rvXLIfBxc4tolQQdP7zv6kBV5S5wvJZOVhzNxSGIPEzYNSyqJgoQXVP//izCxTs3QS
lzYJ2GWl5C8tAosOWfCSObwmHl94MkyksjOJoL0XHxcVxWS3csSnwzu26Z3pDzaZSY5+kXh/TscH
83YtMCsJ3N9D/v8Ocf9R2Ax/crhsq3nth1b4NfWUC7xIjPHzdZCBSSRLG6306+JYNOzVfk30sq6a
aPYe2PlxRWS1cq4vWQ3SfB+5rVxYEHktM6d/lMFnTtbdY8fEpNQTaIE52XftmwYxvLo+uCpZz2oU
RYtJrSk9PLWezSFZkI6pDcwmWavcTsaKa8jKkXheS6Ut0tXiEDCcVjHqP0UYFy6ECSred6g7FWJ+
zpVK0FafK+qoi6FPEnRbI9REtvuWgusHjF6uDlwDFBFJrdHJHmw+9ysNM3nFPjDYPmANdV6nPD3S
0SWb91OMlkv9iKQ4GrUuLOi7ExJHZy6kuMhtVoWolC0xeYrTiBsHd56ZAB9g2ZnaJIrXIc7Bul+x
1dP0+W88xQBeRrM/1xuNaAybMw3uLzn3ZUlNkHYPL+t37VsplZf1cnai/v17DB64EYeTAdH7VlHQ
eIIbH3q0O0GLRAsoHFXWCqWOIJy40WvvqXEVAqZudqL1JTCV2t78ZkIf4LjhvDCKQn07yBjHlS7d
XUyKaPkjqm46gem5GRu1P5sY4qwVl+lb6EGBx2gbqA1uRkqlnx7278FXtmlQaUDuZQPQlsWbL5qX
T4HWLktzzN+BAJHHzmH4DlALTuLqaysBafMfsPc4bG3NvROYnyMjA0VakGmXULBow7a9Aj/gMEfq
eTa32kjef6P+MesM2j60j/BosVqbWVKnoFLGXisRwLO+e2nufo2Zwm8+8gwBdueCNJtzq9oqDwCN
Jsfc1parPTDuoyPhAw4PZKAJKu7cXXEWctxGQvdyTVMr5AxmaI8ECnZAboks6gIPEjyrs1Ugmiur
A1dsFy4k546hnV43eP1ph49vuDZB6EXYx5IbPI/QT3ltk/2KRAg/L3aYAzly0+2XVUe3iwmMxhdR
AZeeFpnbtrRUw1jU9KGS9BO+HAYjJ/aaLMr5aB6ck7ID7MX4hmQOIsGwS8/IyOcgmTdb94byfHFB
zjzJEIfa5M1aPF0ZQz8lqTnOFAG55G3hS5uVhvo+JcQbjU4O+8OQUQ7+Mvio6/PzgR6vnP+DHcA2
4agE6O3QS+rs/kgIaTHdHpOv/d6L1Dmpm37HRAG/DJflbe9D5lDSVlCgHVUHbfeh/OWPbqVAjHC4
ol/THhyzvttZ0fMuj/VRls2LRS8W1gGGI9KGI6wYs1cYvz8x4aXRNfXVK4qB/R//XsgVg9Zq2pgs
naxq/vbS7744+t/khMm52VojRA1Kh+1TK2i97iy+RRe/5d79ZwOmFuQSgl5po09bfhk7ROEwCyAv
Foelowc0nmNCTg3JAvK5U9AilvGWMmRVaO2q1sCJW2HSw13TvbRaluSHluelG8zi44Gmdkscpfr5
FTgHAoBT1sdXo0PCts6Hrq0Ugr6zhGhNtg/cNB5uzlk106hoUzuh73AKIoMPqlE8oVcY5+mKCit7
AzoxPxGoeQ4XrgGE8QZQWsGt+NyWGUT0bVM71DuExnjWFZvbQ3LEC1R7c3elujqoeghf8mDXNBrV
GZ15lEnR0U/0vUP3R1GfW/0SHsAxTTiEYQTQ7cYCjlaXpWaK9rg6zEmv3HmiCGFgDFWVt4mhgnhq
T4aat4OYb7TVhIKFitwoVukBtZDwjXJyuAiVO57AermL9i4oOMFUULFdVEkeZvTrRbTSbiQAhkUE
xVDuK5s8g1gm4HJ3lrsVqt2SVywqZBmwzoMoGnOGgQqC6K812OioRfMLjK3GExxZJx2yEuYUKySy
dP549ZM9OIyecxVH/rFe6q6tE1OazmuA4+tX8vQSEKJN/X1vdfNDqVWjOnjkhMydAKEoOcWz8DRi
c1/FE+x0uc3wT+kvzgGxwJ+vVDTZUboHK4CSx8r/gibjH2NNlmQ8g8xS+YTKWVf0Fm6EPeXBPVd3
hNp56Znhth4LY2TDRLSyJvL7DW9NzzTmEZqTU3UCA7vciHq0CGrImSAJuJI+cBxh5c9di/GhP/+o
HSSfE5ESQyWOx7iIZHJr15pNN1T0+peRfpHzFuSF7XYSSdJRN4JjhFLoS+psWo4nD25sEu2QuFQw
Gj8K4kZIkjNKHipIwci+ngirXuqYJ+M8OG1uzIB5LGh1nqOqVcHuKp9GxXRLul3F2zF7keuKwIo2
Bk3BYRXlkwVVo2o61Ruh8vCbUp4WDshBQTIzrnTKFOUGmNWPpwse60icU5GqMRGm5dRICK36chw0
B6yXmozqE3LVAnntq8CiYjy7qiYLhc38xB/F4Hd1FCd8kP7r3TyprbNWkdo6CZ6Uneyna4JTTBdc
IQmXODBdMNQ5hqm/o2UvmDCDKgRCWrlLHb8D6opUlOx1bElC6ee0VFitFlSBIJgs309EaSy6Tmj3
tThKSqOsm0ujJgWFg39RJuMB/3s0Np75YElVSpAGBS6hEZbDu3jkFu3BlMwFwOoRse52PFfnGYLs
LaJ7AVlF9xffGrGVL0jn+A/kf5Wh9wqmata+c5cvkoP5pVJ1KGG0MHwakVPiRy6DzPDNnbvnVwdY
r6bj57NgS0IKmJ2tEXFQi5AFOoB3qTiQQET9qOGR4g3XI50cNNvWE52qEE3lXZwONBBaOfykBAAu
Cv/Ohm2dzaXPw0jP/TEihO9Je9MBRKKGscUxwVN2CfXXZ7O/r6u6/RefTEY599H2F4p2zP2COnGS
miTBVX22/5o+IOm5kHkysncvekqfgZE36G+KIo/jxpEL9i7WDAaybVyiYKbhe46/ttCiJV4oL505
lzBbp9mtGpbqIAi5ohoJZVkpFtI3yLZR60TBp52X6BREQkvdma/I5l9khFb6SIlokrPqZlmwvOIc
27qvDXRCfzBf8lzqFwn6ZtohqLSA4LPEasSXW+kX/HuVp0PTA061tOhXb1aVonhYCkvzvfgWyZey
Aq48Pf6NBilFyIIX6n0EmDHa43XnTS5aIDiwDkYb0Muuf+eaH8MnDNmbzgGEjWQNhcPpi1LEnHvo
SqDZB4rxL2pafnU1s8GpVe6SKhsve6LDktGtST+z61CHEzbHYVVQ0F1uE7TxkpIx1h9otuv/Hlsg
z/Xup14snsDzDGf99vWKjyfzTkO+CIyhQqRYNyB7JaVaC/rqZ3bTG3UsF8gSskSDmBCZllc5tI9b
55oDy6dHkQ3rRsRJMJiwPqlmnvQSQcKwvF/ya7/1THUXwqaJroo57Yodq0iy9qLrzbSz63LXxgOn
fZU71Ebr0XucFA5xkO57ynfv4w1IXnG3tXMEka5HLFQlK+vauC3q/5gRhKQkESf42C+GeZ5DRBtS
3JUastiNUilH+J/dMVbZfYcLrLYwEUzSXrh+4R/C7ZcuuA+qBdRNBDm2Ve0ENCT0mLWKiBfV3gLj
8JUYUXBqFRYI70yrpSd39qEGcfTAorqk4rWV3p17zBb+d0u4vSkPfp5DPioujso+47QxMB+dtEWi
Y3ZkITzC76bZGSY+6QhLCG1Q8ThVP1QvvZPrKlZObCc7/rnopcP7yrPS0TLDRSgPAignZRsSB6ju
wztRh1iHcttHPGsNVwywxcd7rxvHPoyf3QbYsqsBRb5GUt+LzQur3lg08iMu4h1JNSq4O+aEbgsN
TYVxwbNMBXn4QBh4SbRyIfEVw9dDnCasJCkjEKcstwq/aJGfSZDescS7z7W0sDGJZxFrk0zmK7YR
Ug34dOcOq/1m5t9j0Uck/i/v2ARw3r688Ht67+o8/hc8r4EGhfU+TIdzTWdJEzdVArYym83rg+jY
9PYb/zj7LN6bUoMNRXwW1RoWywn+fjz7vaFc7wEEyz39P0ylVR6DT7yJp7FDElm8nczifGYbyYug
BHkyY/4vcxfstWPh3mZbU3QmYYKwwjZJWFZdNXUgH+PauBuFKBF17MRh2EHQmDGddB/kO6WrRsu3
xHKlDuVRJZqDvTF4/Qn2RP2gvXOzr6tvKHq54A+riaoqgxrlmO4HygR/cYSAU29TKe0QIv6ef+PX
ahjBfWc8IAvJ79aISdxFy2Cd7xpSbC+keR4HSwE+IaaKByvZ1usVnZEnPoeoukPcqrfq7OaZn54F
uEiH/mSVf9E38vwEtAphO71YTcJy3ym9g2LlfAd9Ou9BwUUGWb9qEEWvPPKjSAP/LnDErbpvYnj9
OOe2/ufhsxdgfmrGF+TPff9QOApIkTTw3fXcC88nbwH+2XZNyO3f+Us/laaRZZDUAIoNi1lGAWiV
hxGrOZ0VoO+SlNbnTmCpSeJwSXWLB2+TlZAcQgVgG6wTZVPqE5vIa9NJk1IHDzWOa4CJZIkNgrH4
mM4upsyaZEFVU7mN2SFJqDj01yc47JY9fqkS9KSOz3dygsakL704829AfCbyk4bq5FIEOq3kdawT
QlRUABZG8n0yDiM7fOaeDRY7AxdGTJ/kBaQfIBD7PUyKTQli0mPjhUeFTf/wfR9M7eTIfNtLx+Uw
lpxy5eX3GyzUVCbA+KMtAzwYTQ4Is3sDqU6oLRLWlYq5C3gkcbxGTArwTnHSISGXFfmkuXEe27mM
pYovdS/o1hbF+kDASsIlCYhtEjaTymvlH201l1PLYNq2Vz+u4eK7SX+Mms/l/6/VGUWcdtE8m31+
tRSlcMPIKCTOv3KTCcmeFJraSC8SwAqwa/6WzMcP862gep0+IzB1A/F7BushsES5KSnJvXuAG0uT
6r7g5MihhFGfQ7SC5BCJD/nCXZMxcgD97qNBdUJ9tqrHwH+GNXPEKL6HQzbTwJHND/xCPdblUYVx
A5WvR2Ey1oRpXSlo1uyM947Uj2EhE9gQZG+nlMOO8HhbaevpE4F4ZpyyzLOAR9Z1r5updduEjhsu
ZKroS9M7GxBhhmF6XysWYR1PgF+mKAV+R0RlIZLxB9UJyHJdzD1i+PS/SKtxkWtyLhk/yZWoC5+b
Wb6KcZkbG/xxJVLO8vnvqY6NmSQcwZdAXeXW5rvwMpw1ii5S7bwjUSiShUe4xvw9mMnzMfUM9Nnd
7JvOxmm+XJjI8KzGy1vyF0hgUuAdisQWXCWwThjkKqwDHL0jDtv37/YLlo1z7RguWtGxSBPIDBo3
W0QofJ1VYf08OP6XNyHDAqkdfbovL8YgeA/5O/l1Olbe85M/nnjPpQsk8oQZAfb/eCiIWzyq5TJx
RWl8kxtNKe+hyOP1y+XrMuAQ+DrnINOkJ+IIYMiYbOOrtlBlBYjk+pFzycGKhBikv42jWMMxkuXL
TjdpVAqO51huiD4UCMdFlMWbB37UC0ef7XbyaPPLQLHKZOQ280hQ10myHxJlVg8P3dcdnL5UxPkP
czvIhbtRDJsdWH3bbxSmi2ZzCijmPyZlxIKk52SB5Jav17iDN9SDFivn0E3nbWN3+1Vxvj68fNSB
HmQhFgXsr+512tjA+iShh35e2nqR3DNKN/gqaLDLz4lC8gLmA/9c6ko2LAWOb8dZQwqt6FjTp5SO
KBauvmVo0AGHcW9LvSu/HyT0s4UQmNqJp3cqUvFO36Werf0s8KpzUt1eeKMv6/69c/CYqB7q5UO+
+KXSfzLqUgyXFG4k0OisEFGw68oc+h2TH0+7ZvDiuJQbXHqVFximmb0IWOzN3Rm1CfK0DSA0S75a
IAWtTq4+6i2am4m5WBVjd+DC66c0aJEW3+cIR61wtVdfU/6YUYT2qUQZ4Bbi8a+LTSSyeGtvNehw
f2aA1FBBnp4HnxTl/PXvMdYDRq5/i3ZH7bKPvQLpxNB3MQGJmuVv4pC91oO5SqKoIS2/xP3UtlXC
i3cD0ID+Vxr10s0XvoNr5mJjG7BQTx9pjCG3WiAD5pwyno+rbnn1YI5SPBJX9CSCJkLftrop8kmp
v/jCyNUjZIqgxzJI82bn1dGUR5hdWgJx7y67FEfiSH2+7UsrkLwee23wd4xahKlR03Jw4VJT3t77
+r59Bdstwb9N+ly4JGmO8/01BB7OFJFDkZtdZB5/TvJFv60RS7Iqem+ldl6+VCA6f18pAh9yO/Cc
KhKkvePY7FwFIY9NY0fqfgv39qaj0AIY8zWewSAvbaOxX8fvhCnchhYD5DD4LQltUO+siz5q0Qi8
iog7brTOyyEIgaDwiZEinbkEyEdlFR2yl6H/v/jkgvEJay4zABbjjEWCCL81b/2S7Vf0yGaF6z0X
oq4J7uI5y27fCuHU+YkhXgZwvOIlo+XB0wmnROTBO42VUiWJLRFHbaVdEAWWf+sheYufjTqxalsj
Uxy9dvQqSak+n/ngvHb8gJJotech/9w6x+3rVzyvSK02V84NFJIeTD1lkx+M17qkB8WsDiYJuemb
eaHk+Ure/X9aBx6u96xzZ/PBwqZmCOKjNUnLAUeUsClQSgQsIBLcNxkszYHhpTiS6YOfd//542qi
And+yUN9/is478nTJwixGGR0ilOOS4dPOjhb+zO8eWnqjtkzLlqm7oMrNVURtq72DEe65BMM7SbA
ubmNVcdNdffbU7lmYABa1ZwIzMSsxCKG2gQ1bBxfcEaSlwJn+OG3tUVhICUG0wBmca6BN+0MXMwa
1QqjqzLCkZtQLl/Rj+MzvH2eckxefQYPv8cwVfJTNeqECrhuJAte6je+lTda4PX0WptUFSGCPfw0
QSGoxfTjAhmVLWDpt3RVNIW069XhHAeKZnsHQ5/OEcuRjyTfkEhLUeWfpQwzKFa6QOaodUs7dXU1
1WaThcLxlsoJuuw2SQ4qbhMh6nZK4AkmPRWrpByxL8K2KVXugKAzs4NBz3Y7Y/eagnFP4kM8lAOO
2Z9xJkOzCBb4W6wh7GWvOSGF3NZC4y48nU7aFYmwG0aDH49OaXKDqR3zj44So+GWKx+GsBBaaF9S
8PseABVhVE4nbqsj9yODHliScahfVsLXEALne2hD3deOiKXZa6AQK5stqZt2Ymt2BiK5shTydbMH
Q8o3RPNeaoPvH/xaBjPbP4hD+i6V6yLQU8JOqQ5dLrOjL/Mo0dgU0FcB0MD5ODyYOT9F3PJY2HJF
HCh3Ylu1syJA3tR8YRg8tjDSEeHj911aOEZ+6BopWSWM6KrBIhXtH4XBZgnLb/dAyRoexbBPleJz
YRgr1s2FwF84dRioqLeCxW7KBHArIO0IhJY/kQqiKggNdyNcltZUceqodKbhLCcbJlFv6QzY1NL1
CyT18yO57YFlKo2SBNYdxbLAL38p+P5kBlAOw0o89TWxXU/xnYw2UyfKDP1iBG2Q/VNNglD2VJG4
7mz6Xpk7TRpdENmOaLLm6sQQeI4r0Vh+YNBoI+qu8wLjt6EZAOPlYiRbP+dI2DTHeUNoeT5/vICE
m2EcVSA3yJRiNHAr2ZbLjbONOy0majUWrJ+bi74H+ELGFqUrKh9rchCUmpua1LM0tO83pJufZxzT
nu0qaqRXMMm6ubMkztTRDlUZgnpqVRCmGYvB9slCjgIMUjQxWVXURLUFCuKpwqJJZhcvHy25HKR8
zBN0/alXsf8sddnshDqCXXhJNJCv52/PWSL89hVafIiEx8IM+utmPMwwCsP8U4+DpLA22dlbTS0U
QBuT/BDnQifNDbFXycFOS5+tZqEaryrEueOlKTr3s+w1gAmJVCeQkJAxu33tLVMvHeGKW1Z4kVVs
QOlTFM5XKsq5WJoAcu0d/B7idtxlG1Pi1L+7cwvQQguhYzfTlZ31bx5L0oufFgAMjTYs9CGf0IzS
CvR6kKmyxrerkAVWaBjB7I3c8dVMlTYAqLMNguFTs1S2trWurDmRNzqqxLOekgLdMjx6PCbKrge6
ZVDPW1TQaDcTo4sK4qzEuEJNldOSBtnill+MyqiphqZj9Dwth/xtuLsON/sLxBRTmz+YwSrPksxR
OwWzPkzeZEJ8ZSszL9QMmeyWBK+lbCJzDnCzCVoKhKBPOy9sn892TzdcfY8DpFxJCWYFZxZWTSKu
A1m5MvEP6XnC6oa/baeE2GPQEO6SCRkQoXGk6qrWilbbU1o7v+9SbJOANTOpwZycsQswSkG24OlX
4z9Mw5neKFZKO6yoqyLjmIA7zq1R81sV9IyBTQi5SruZkmlRooG4p8sQM3T6trBTCQtGZMwwed5U
CAU4YJOaUNg1Ej2uoNnB5D7a0rjFlQe+UV8bMRNmDuNGIHpK1461r70KA/pYMyaUzIQ/frfM3dVW
DgtmZx07JRtcSXlMjxkKGydefDz8ZKBJPjBzmTK1p63lXFzYGGEWqFDQPa3Tw/nbH2m2/nLfFSaA
fTVtfYUvasfsGPcObaHMT2grnWHQbw+5rHVwR+2zNrT1jsWrWF+4SZ0y+5Pv5mh0vQqLg4tUWSF7
zjvDe6o1A6whyYHxrm3LSLmlVGTM+gh6ATzjjbTGVFuOxyFj6Tvch41ewLeei5muxLqdC+Ovjwdd
R/NXGS3/rRFF3PcVvIDnyuZC0hgKnCXr9aH87d+MrrYkk1RB19bduaLaaRftGfBMMBqTF0r8igCl
OC5hifqbcY7/0dhJNhamFCuIVtrv7OKqPeKRsgVcOkrKSPn58FJRCpoGz3XUzViQylFrGmKE81F4
yXwLy2pdudcTpN+VQV+8rbsgMf415aqdtyPk7LwDNIzNPzVkm4do71+11nXhD5ouMCmDVNKoSHW+
BoM82gBcpKz28CuPfWiOK/4Q2Fpphkd7vQcxx+Y5WpSrRpPQEPI2oBjmzU7+BZjHEL0qWch/Bewq
aPcGhAwaikouLsj4nQMDylhHN1UxNztUELiyIxwlTB4eS6DfMTKSW0/WHmwV/oYBG/jttCEqPupV
d8NTuqn7mnAIns/QYEg0JcQsv68Lb+/WsTF8UxfS6TBU8dAIJ+luPTz80T5WWSyZdwL4bMDFPeF+
8ujzYgW6zObFZWurpEd4HhN1j5q72hw8OAc0ZjWcIiwMnrvDwSasqlidDK9wzuGI/u2j4fN9xWuN
zLpP4pTzVc67dZGdXckNsLxc/oNaFvusuaVYhdDHZu04DnGlu5BxCverTYMCvz2mALFUloscJ7+n
YfVfufryqtjkeLX8rFfh/gRukfpXvwA27R/ec1+YhxvOaLxiJZbNz0OOReKVrdtRgAubRbUifL+y
+j5T5zN1KKB8R+3/7cA0KHKvZomG6q+Kl9BsV/ur8nY98irWktCR7UCGUoYQcRct+RaZfCTJi8SJ
f6/mCgJQeILb1LuinyR0vrsyUO1gNDh3sFj/pwnoUo//r3Qxrd/7A+atmHRjbNy2VS/SzWhWnXTQ
CjAo1UOWPSf5CuEiEEQsOjcqzYjPcGDaCcAOktqMkEQ3pknRYJJW6H3AXoeoN05gitZ6ldOULjaX
lceXmDo+p90NNdtItxvjjpJaQq6RwZ/dhnuf+SJ4E9fV6MVlBGebaBubj33DI5Cn/6+gGLbb835c
PTYGwa+rpdNnelBv4UvYzR7lnR9S+VAf1Nr2asAvEpZ79eEKROP5ng8m4sxqso9OZN+dIRo0lk5R
A+b3MUAsyBGpd9eeaYxserkNJ/hMSUwRWT41Wpkizp2v061RNY87A/lwV6Oxd8vptwOqNM4siDWO
TQp0Ie0LjfOagi8QqxfGRilDBtkboXYreG3Es47vQiJHPEbEdrGHhHiba/pgKP4Q5tnF0BAxiI8A
95RJY50fKpGvTMOC9Q66RsuEW/7w1rAJHam0ycURqBlakLxwFkUZreioe1V0gAC4OZq/ZeZlfKc+
r9vJDeVw14gKf+NfrUzWgcDZDw3ReRJrXWeIcjqyFNIg+Q4MMw40972Oh4qgXnvbVEd9IOG9yUyF
dd+RJfd0jOtZ36t1LwLyKQeNaddnOyF58O8URed/8Smkm6aKEsys7Fu2WaclSCy1VguM6vSXGoCI
xZXwzhxr1lXvpC57a9ErXVVMr5F6UCyLxIGLGqxJy8imAJ6daeqaZKdYSCKxIXZWgW1KIhpn4APK
M5FVLKYIg+jxV9dzKyhq9v2O+lDVmN/hF/iZmE0hVINXuD0SM1A0s+viptEbeCS/tTdU20LNN2Ey
firVZ6WPDR4syufKO6mgs8bWCVJbru+6bfaQywHs+gCPJaSOeOGACy9r5DN3uIhDq/NbkSGcIGY8
6ukMCiJ2JMokiNVMIm27jNwLkHbDXUiWA6Rjyjbu/zL341vVPbTIxEfg4PH/5rvjAJDWpjpYGRr9
1nLOJ36AG9eSTOETh48h/jLgIFWnJE4iGB6cqaIk95Q3vO/xKmfsftAKXwUNgWv6bg79SSx147yJ
W17FbPH5MybteHSrXhxbpl/aec7ogFSIzpPajGDKsudBnL1TBq9CVhIvAMfwMbS3isa5olC+NXtJ
CWlk7sOByS8yf5N5bVOBpJUaUgNVB/0E4Yvd3vvfPlrGCRMQoC5BlcluIHTe8J4zCJTEquoHJrzU
8tV7+nxlMFiKPIZJYRVPTp87Tf3ilXtcqw6zkU+eNo7i/iGrhHU2ogf+ntjm8QCEIynsvIlihSJO
H9KfvTRR+9Fi6fSLtlZXpDuvWT9QA4Zn35f1MUitShRY7PXgW9IsvU86DMSy6ZxHQs0EaSCIHgwB
JdDKIWre+GZcTrKSrDF6nuiChZC0FRAglXG/MWy9DNLFO+aDHOELCx3sxGx10hC+/0Wj9ZgwjWCj
SxHj6Y7DZm7aXIdqX243ETXkVgE9qRa/uzAsCoN3F8AB7dcDjYKHScctJB4mfbLMLBjFpxrnhGtv
GEw5/DWjA9K6NZ+rW9X+UqxRfjgKq4q2d23paBURqbrohsc+rjTaG6yaH6GNTKT0wSclScP3a2Wp
KmIe5mC6knltFmhKBuV0tii/9GskYHwP7gdo16WxW7ulIPWtwIQn8ksWVkFxhlHkbkJYjbGSxU0k
sUSXjiUZU3Z5pjcofoICXjziEPbpXiol0pc8UlYceOLD91JgahIe3ouICuM8aY4/Vev0j9beXaV5
JLmbWvtHOwk+8MVfi4LYKFnWgxqi1wiU1ZuEyalEdviaz5BDeDxgJdWBJqA57tEzGx66IncoKBKf
Uq8gxLoFL/NWvJGbEXM+cgCfCcz+/hiokZfyDVxlaA/w9ao1x4mRdow2IBGakghIvmpoe8XGbbYu
6li5MN473YF+n9aeyi5gsRS4joLh0OUjKkaBUy42uGhTyzLjSyb8UO8QaWFl8xRE73aCFh7VUtia
O16QuDCWC3EpU3NNLejYyHjBoFw28nim2CbTx90gOF0Fj1dD3z/f3KIPr4kIXVi68/3X5do4BQmO
v5KWs2x8TQRsZuZyQyvT+jUtXhE0Vm72rKRDNatDLfo56ED6TnNTJepKqiWv0oP2XWwjBP/qpomt
GceLkRek3K7S5eiJ8qiZjK9PqDx5KiLb9D3VD8bkuhnmYdaA/gDiJLWxXs1Slkm548vXzPlujXzc
PXFNQHg4eRzIxLGS1v501ZY/f4v2/43ntxfsz7mV6j8AHk7+2TVNFTxLxl8Np+qIYlRf+Si4WwzQ
0yuC+GPrCTTk/QjCqtqG0gTRzXoltFbqVXtexTgTQoUewFYFFeWHAo5CIvG+r/ZxMA9fLmpBZDoV
FX4F0zbrTnUbKff6Ouc8yQWkT9jym+hviT6u+8xLJO9SzvKbIcUnyhyJOebpUhT2VTDoxpoDnRqG
RMoj3ygTYpvgGdAF7LQxBpZzGnoBSsVzqasrp7pWzPWvK0gaIUNvJ+KN4cSowvyIw4gyQB6RgXof
mCfhwU2pgKR7DO8zieGvjgyasULZ3hmt+4KWyTmY75PU90TPQRYZN+Kxz94NgYxENyZ5V7WIt2gC
Js2zl2Bn+zAPhCnxWnnkQzQk18goqSFdzCH5K8wKtrCfP3XWHm04vxeAsQUIuPOR4YPNbGDTb/EE
q7eBIi+hG9H8LoGZ9jlvU0mVA0YQuWwyauwFTT8lJrJ1nHKVJwJLPrNNq9anvoQiJV/2Pb7y9lBx
h2AZEupIVT9xDl/o5DnEcfwK169wXJASmrCNKO5ZbAZ3BQuftn1N4vjWG8J/kFOG4pyfALqKKhiL
37QBcSNlcHZiTThqE1LTCzR3O6f1WSf9KnvzMGG/uzAdyeaYymHzQeMflwo9uvl/yhS56cbrcBs/
QAYmV9Vdd8MnO6JfhTOjM6CIj/vKLvd3sR21UXNJG5Xp/bAy8xofZVhf/p5vX/A8I6CMrCko8kcM
txBGeE3GzdIC2X77e1IOSgn4mK9useIbMT5N3LZWDxODTy3zLWRq491vCsXWXBoS570fd3wpFL/k
bpqGDIHeDN/YRJhekmRDtyhb0Cg9CMja6xKzXLLabKsYR7tl4gPO5m7fbINquj3NeX3o/9bNQK/z
UQTqjCcpFp8q6z1n2ftvgNYi1U/lIBeunCev9UWIg68MN2dnu49Oj4sxK3zpTi4uyEO+Uqj18tXk
2Wou++gKOzeXct9RcivVtfbyvRBHpHHAsuBJq22Bs9mAOGZmPSZhevD7r7BW1ZHkSNcq7yWPxMBz
x5+1sjsPkADfOpk8lm538visHae+xYilFrDBM/hx3lpasfVvteeOdU6280NEzNAWG1k5Ri+pg+Ai
9tGvpaZJtL6RkIUmQ9KaenDXj5BQgPoqygvlValrrjD437k0Y21c1Qmjy4S1VVKpWkq0C4CfO2tz
9Ghj1JMuOEV4d63CS68aj7IaCq0Gjl/f/v4N425EWYO39YWC6T+XmWiSud0Wboatk+KiKl596rQq
eF4l7UNS6Bvoz12eVewRX82bOlixQjh8b0m1kDvZfJDiv6Me8m2te6Tr8BrwuCM9uGJi+zDHr5yp
RtyPm/iCqyd4AeOH1KGcUkk74a7uVmLlt3jr+EPcYpFwaJzCCD+6lSvK2IlrR7Xv6bF4ObzqXw3m
OkRJ+t/fpNKL/CZo0uEJbIbGyAYCoeht7L1MJfzX0SMhEiQTodqNFjr8tR5M1lTTrgq/rQeVdF2Q
iUtL2NfNjGPfF5pvmDJdrjQLelg7U2pEasfQOKdBt9koJnkHbYL9VzP2AvCA3PtIPFJe9MnXE0RO
irkUzFqVKlAYArMCxjqdBDqZF18EMgfXMYY+fz1OTgnNcy3NdW465s9VQH+gUm/eWqn3XxVrAK7l
l2ZHyYVNjBKv4SF8MuwxD/rP0m8qWaCNBltuQ0XwWQStSIFvo8oPmk3v2GtSZ17vC8SxUmv00FJ+
lAHOj1odlsn2yXQHNo/gmsSq2U1xGgYtDnGcf5eVJTdLxDKjIu4LpXpU8qb30C/SIXDMR6MAP8Rk
y56wgvWjSFPbwJx38sW2Uw6l+TkojYBUiYSgS1V0VjLZcAPRdbitPMPw6/kTAgwfnf/bdhhBKHTE
E7OSD6EdQzN7ZfSPFfchfUh6GlJnuGKvVhS13Js0uF/GGOYW34N6mOSxRhfrRhXzzubwjVl9AdWE
rdnLB8yeH9V09Pu/gHgqvxHQtYn9bl4Imjlz5acN0g/6+wy1QENjqH4/lCxnbLFAWGaWOmY5zuUN
SIEX82MwFSWaHv7y1k7+Io5ujTdChk20DSUyrOfogxZsawVovapwpYk8xWSdLm+E7/nYGWJ8+x/0
BbsACjdeG12MKnCUZASzuaAIvQQil9QUQdCxCmMJm9AtkkNFQAjoL0rlCf9ez08q0fznV7qsQRGq
q/pkgcrCXm9QJJjlgsgfabg4OMmEokq0e8ijyYoHTyrqXKON1ZZtkWh0Wh4beyIoiLbogPVUWKpu
U8dMHoWrrS+Kqn+Nbv5Qd7GtXo6KgqZrnZz7ObbJG/rbdFLUMC5DSOgWH4pLn1GTHIKmthU9V1W0
QSiu3KXdFeSDQJawY96Itn92lBmzNIpnlTmR4KZMW/7rxwT5MFdFn6jN8T37lYk2eNT/QJTObBL0
47HZnTJ1PSkDeL2atriIAmGxaUTVop7Aufk3g3M46BjJ8Dq/LPKN6zX6DizFwAXVY/Zk8NSCUMzs
h+2KgHOgCWz33O9ze1KAStDTZDQgvDrYoIOqWRyI3S/SA5cMomQFhqI9BAGVtaDPtgjYu8TZ3+PS
lzQAxNDhlnHTjHJQgfzMHniOHCukL+Ntjm2Yy94UUMLZQLAVyxd1wFEF6qS8PdaXIzVz0ADfnIgL
mtvUbZat/2tNG9mkVgud065dwpN2uUM7kMx7nVmHQa14EjR3Ek5imT2dhCChLj8VTUpjCKUcSNBa
PueexS5Kr66ODACQ6eD946OkQqZslb0Px1Nv8Q4DJF/smvM+noWS9IJD1ubA02c8ZsgsiF+m5Wxv
EjvYNDLEHw6IRfoxUGpvUa2OHtwnDp87y1itgjGiBTuJgR4PQi50JRx02kuZUwjSPfOFgCRJqwF+
zesBDLyfJSkIvZz2UDVCGntvlNR3Ju1fELKPF4HOEFw4/iBgfPgOUGWlxMAJUYdlH65018G0DSxP
G+dV3+ARF20X2gYacnlZb0pluetpnAHQuuddsMsbV2tZaF80JQCQb0qeI1vHzkGeV5DzmaDLqL0K
vcUbUC3+ix6t1y6kv5YmbzCoYbb+/u7IQFHZFOe2SsyjOzGq8zIVNe1eRoz2HF6yoHl5SbHPZbdY
n20Yds634BrcKMo5rqxUdDZzoYXR2Vhio+9YdSfFMEg4eWn9Ztu36NoATbKBxqVPHrWndFvEalNr
UFVprgBi1bCZzNgIqzj6qSyoVjncqDkjlcUeYrtPSa+sDnYOtOUrNPa1epfwS2YJeuO2aY2J9OtG
HhXAxO+puHOnpmt8rTDYw8lqRp+ajrh7xJstW/RUArnvE5KfRB2Z4UZWO9qSfRyGiq+VEz+sB3sc
gN+jH4ZfT/U9IQ/LT3VdGUI54nP3BqugCtTdSXC0ngFVM0BArW6hyt6VHBpw+8eGnKICk/TX6oO4
HkVLzV54OvLxI1fkxKRBeqPGWl6iFI858hGZfQS8gacil3yCpIHdspy+iKchKHcut8N61+pk+lM7
uzrvMqGk66ZeLkZAS/yKxQB+tZWJStBNyaCjvSMxcKygs1k7BV4vOd4sGDOe5AusjI1+A5QSi0oK
rlblJAWu2gAVnYPxpRMtgokJA6Zn27vlKEnORpL/9U8+pUkdTA3CqTYr7mTuFZPim2G0/PlTn3jz
pDoaQVBQgJZrKQAKwV0c/QeBgz7Mrv5r14o2vmL5jUmo/dtagDcbIKS1UCEjiOUXRtoF8P79Z0+i
K6zCdIEMeot/MWTrBiqnpkdtm3PUdosufLC/MaG7hCOOqkkakJtSAJoVo3k1K5RLKq4zsYDKUHpl
ykLF33rV3qPJQrj//0lXbdKPGZntdOR4kqM12BKVT7uWJngNb1laKlgfwqg6d6DhbJrWUXQOOYAl
kpi2YNyX99+5ZI1cCL1mxeszTqX6B9mhLZqS97mtpXyy8rPa2xgrqiaqLtEPeTx8piYro+mf0yW8
91ZdEkWKhXLXfBOqR45fAp5+9sq6O2kIut/HotR4DhK2xvB5HazOm+GTJ83+xUqZ0pKwXGSRlaL7
915cigb00quKglpN0ktF9JVc2D4qLwxbWqoDKwATUvLxpEOKn3hjqSGfRzqvXqaIpglWMR3gsc7y
WHe4Ikc800ZIK5bymR8kTJglnGgfdi2/AbJOoq9WQaQqDBJyiklGzpQxS7HfDSA0VDxtjkigP7Jv
br4b5nfeznlVoDL6iX+BahJ/uUIUoVCNi3pDMixl1c2KLN70VPVPNGbFMkN5k3OWQ5doho5Un+rn
qQSWQztdNHwG7n3F8g3R5SgiiSORmsowRaqPbI11otauT/QSWkurQbQ9CtoZLnf74J0D50Q5drf0
5fxRZwdXA2NFFasRSMi7wBucBtwZY95D6Bszu+0V6NVRc8sbT8/959DptTycy1k8AqNtsa7eL7+5
suoGzoTkkKP7g/oEceZvhRTDN4G+QYZPfNXC7tRd3KoW67HbRZAzmK9cpJHD1sO/CkdwTWgqHIKQ
YedRmjtLbQ5CpTe7i2sY9uwP3yjWHd2nZRZqJuSfiDBTr+UESSViXQpucj/m0cY/7W0oEWWWNNVV
WxDf2ZqqmzicKMNL3tb+fiJmCCO5aSaKOxoRdCJ9ArjlYdbuvgJKJJfrJNN12rfCo+UuQcr6rGo9
s40/HPvsr+6anlp06sdeOmBNljL+N1FyEHriFG6Te2G7iDy15n6IKY5o4X9SLmQqHAZ5CN/QvFXv
nuGcuaCsanroPHODEBSiP5l/EgoxYK43LnvFGoMKKtUDgXzVguQJCS9vQuJjASRLO4PfIBggBB9b
3p0pgEctwTSW+f2PRoQb3KaiusepEHL3+5EbyS2nL8jtK8wACGBs+2jrPqzL8O7pnLBAaGAL7qkx
vBmJvkwPG32cV3SMW/dSq6Oi34cOnUjKteG9WdWKng4H0E73i4qerYQQqzmhh0Rv1oxSBw0NoLNr
jZzNIrIXoO9PFQ6EzlewesZ9btSbuwl1qY2cUpcM+wmc5HGlQnziRydDx8ECOFHOoADLqUCfw/iz
Ss/wKy4rUFOMqNMPjZ6SOzCNsI8IgxkVQjNCY6iV+7aKfKAGNTGNQ5aaNjkZjU4t8AKbPzTXmlEx
G4kQiRnSHJ1/yNx+eexTcoMQQsVWEP9d96Ai1Zn4yfABUdf7JqkTZqwkOgpWAjH4Nq6X262J7r1L
25C6kE+2lwZQgebdfNTccOkjn6s+JLnYcXATalQ/FaC1xU2h8ltBo8rlfzxviuSX6cCaGBnZ7QKm
6+EbpKVMYyD2KsWNJzjgig+ULprBZ+OzQNer04BwcQqp49XujV+aSwG2dXFmujdvAu5i7HXh9/9a
6aKBQS3GaNu1e6XcaQUqK5NXgP9ptlbhgW6szMT5qOgoqOMhIc4xIKcVq9LWZ6YAQjBK8zlk883n
iBFk5IIY25TlWuf7b0PoYUc63LgrjWdzv/0EMYAE8C07hAx+G8u4CvjKRwJu16gaBcQ7qt4IVjtf
tv8M941x7+5SxEI0lNAn4dJaupR+LbV+2wJIh55EiABRcTuO2Z9VaK9g7Ez2zcq70KAnlBVMBeiX
s0bGlXGEnQOOgcmYCSXVl+Icd2k7qRtuTNsjFToFzDCHyyRdHOFR/DpAD7l9zV7G6TvhUGIrTmg1
7MF5w4ADPZQtw6JXR3jNCbyeD681IjQ9xpT0VTVKG1KiEKYGJ6uqMbwaL5UjnekXvRPbHX/aDLDi
2a4IdQytDFEKxz+gNr+NTPHMvqs7V8vysU+RaSN6/B+huTR/gpQbH6dh81I3aMHC+xvYn6ExyLbI
JqgjKd81fgqPuUmmxii7BFeFbjpb0VFlqTQwTJTppPGpvJiDlvL1Hpnno5DXvcrphG2y4Sa6L0fp
Jx7Q+nvgTxMkXeA5hPgjz0RqbQ+eZ+j83Mmo1LlZgEo8RYU6TLg2MesstwlU1yrk8vJogM/VbqTt
OcE7lpcZlWmNMKNZx6dY5PliZROG+IbrxWPofJKz2Wt8AzlziKekYrTSiJ3Wyv7Mg51UIGfmPnde
W4IJeClKCYkdsuuFMuV59tgiQTq6NbXhYI5Yv+/VE2slMjSvU1Q38PaqwvmWYDZlK7PaAL8C7Mvk
AMJh2E6zHt9QPPsr5FjLZZvgxOQ3bslBC0FzLxODbKXPeKvMmYkI8VruaFvEyaQrQU3rJfO02EVU
CWCJzj/KspgMyNWY7I9pUMxl/XLwuvW2zM1Cnm9BYojFmYzPfdMblDJ/aS/sTjmP/U7/mwFzx1oL
TH88T0+yZyi+V5tuRLJmGdTp4gRNCnCS4nshaR0DhVSeBw2W1b/CNiNvu9YwRdvblkHgS1E/pPA6
FvPrzEvd3gQjrdR64eOFUFDTiqt6QSaLIdTaXVgXkQkaSGgP802eWAqySWj19HNfTVG5RQPTTisH
tXWg577JKrRi7ajb0HPooCqD43iyHqd9somiLtqXmLJETNiAodKZddZYySCHzaXNVzxP05mhoqhD
sIU30b6qV1OamZiVOG1oC4r//OQGFaO4qMlslLuEjKU3gsDx4TeqfM0oLYYAtSOKhgQQS7BaIgzQ
f8fKPLSYwxrh+NDCpOZoLd3hTP+IlxnHMY/xR8XqzWQ2sZMXKrSjZfZZeCdsEtL07psmKV769pb2
6FNQKi72hZUVvyiAN3QvbQlH/6I4JxcXmut2hBUfytOm+/ygzKGjNIuGTCB+brkyrpoZFjB/yL0A
A+xwQgTnV3Em/MN8BmOfEWisTtYgF+OzHpq+9y2RH2DdhGwOFWLICMQO+KYyTyhgHKcsIw5J01o9
4kGVXAd+7dFce8sixOxkk65yIuGMasAQNAOFVVJv3gi+v55obVdqxzveypuKSrj756NZoMmjs8wo
CgOodj2ov6zDG5vjwT9OoaEbNDSzeOJrRsjxk2DSsPVH4IFSREp5tBgAb4mjOmv/m/gPYO0vd/m4
d3RU57nqgkZF7HdNfXAY62002fhyPXGSVsDQi2klqpE55jIncjy1ZROnS9MLzVMYkR3Jkn8jX+kh
oXoaxlJt1NagFjoylXqBgX8LshzLCo73zejdr1SQu3Kr/EgSqlf6DHxz/VgfthIAjh+XIioNekLy
1MwtBFft7/yE2oZL+Ihz6949ljkrvy3eVeHYCrvGTv8lMJEt7vMiTBGoU1A0mFPG+D6CEdyoG817
nIP7RykzAopjCZrchwfS5D7jhpuvIf28O7JEqVBKJZBSvfTjSqf/pvrEv7x3UA0VeA++hzWW+895
nh8EfAF613qgp4ngLznRL76aJHOqocCQMmoOohE0jGGrUVgxdE6RPw/EeRzP9jbrNwp+MjvzqbK5
CsZbhWX6ewwaqylIhpRxsFIRRcwEGASNcLqDE8uPYBrT2gT5k17ighOwzTXJOCNN6JAjtovii2WX
Z63WmxoP+em/CFxnJpYP3QkPi1AUBUVGOSzjlrhdR7gu2LPC0M+RBCSrQqvFHQcURV+TIZcTTCve
gBQ0gLge1f96vjZtAmgAVoGX8M/Pquf5uthyym9UR2Ez0bro5u2JzznaQB63Z/cobGZN8YOik2ZG
9UHNVNmzUK43W5upr1/7iMiMe3YU5OSM0yucSV65hFrooNAPHcawpmnYxRgpOQ0M1FKmUK9s7Yos
NmcJ2ziglI6D2mpSdw2CufNYMIgX4O7XsC7Vjicb9fH1k7O7BBWxBmUT7oGW/ASAlk0HOYc+F1tq
O1APfL/pLu0+pqOs7EucHjEtygSR9RY+SMszcBXUsm7dzAfLUfiZfqXRsgMOMh2SB6J0WK1OUDl9
+V643lqG79R51W4PlXEGvCkS++xK4Pj65Be8D7Ezz0sdGhKg5ECC2eqWLwzqs9zpWhr7a1ipiGzI
YA9Qi2kHjICMU96r6P8o7+OHtd3om1TaBqahK9n53zy9I0sanz9MMSIqG+ZxaJzq2BGoShsIFwnH
nLvCAGK7i7z9k3ZTD8noWaKjSW+Jmbk+9UAOCLNiQNDKRNniHRyyadQlWcUgYVrSsjmB9Bzjv009
xv5fqDnBzUayn0IImvlf/1NBKrJMhWs9HJyvB92LxwnMcX3kQonmqzDxkVeGIhUwTaz8MsbEMAYc
gwp17zOP6TPGv8na5HYOpof7nOw3WizPJsMxptbkNWIng0Zh4lokEtio6JL0Raqv/oMdwRv+AjGW
NDSl3vWwsiTQupnbDOoo50RieoHjZJmHNG4/0NBh/MWSP7x110FqfPf2jWWDjCv2B2HUIl+vy1Cp
SYh+tK85T9fp66O7YdtMJg1fBAlX6ENxOfHLkpMGozvvOVcZNtqZgUyUnhuMLiFzmhpM5kP7ZjYr
VNOCOyduqOT6k+OvhTaWXZS/oiuOHSt28WMZooj9To3Bs3Il85fomPb1EbtXYIOLKASvx6DaefPA
zM9XVeSVGuB64B8y1Kt9s1fd+Ck3GPC/kQhgDSUafeuX9bNn0ysOyFFCpaViAtxTAFkX4OVkW3M2
pejfWM//xwSRq6n+4/zQND5ajFUhgdi214q1QTu1/4gc2qk0QazZSD3JZu6+5jVPu6GMfEqD7n1+
FY7aj5jELgWbFD7j5yLjIje4vJ42adECKTbjjOs8OsVRDJTIQnnjjJxWJ7t1XzfOjyeTSdc+XPum
kihB+E2h3+i76i7Q8qs2q0j9BnjK+MkAR9y4ZBiK7gmGVSa67YnNBFg17gW4e1tgt5SOd3St2p6b
Rmj3mJnhco0hnwJIlAf6VBLofuclxdQyAAp9SRIIoi9/i5d1aNsFXMKN8zJbEYIyeeufK5H7PpiN
9XShIXAH6Unwoc0f19kN4byTXwqBzw0+I2z+dqTbBUEjxPIRpznJSALPf3iAP4VENyVm4QQBkFyt
USVmIRgKwSHxzc3MA+pTzzQxm8T6B04Ax+LKbRbtvCFEbPRIiLKTrtxysx3578oTlGBWFZrmLbfE
uYrRQ51NxeOtpjEpZKqFz+TPfBpN3Ct2x10DIU4tjv6hkM3TPOD7E1Gf1rvcspU2AYvNWJVJam02
YNf3FooGYOodYsfIdXfGOacl3bldiyAegFqafxJlKIr+qXMX/BGye8zIxKk9hUYzqiQNS1ky14XJ
EtU/Vlqvzfj/YzoqRfvODT51T5GeoAgLmEaMETA8Cn+4SVC93sdDMJNSaRxv9exIyd0aovLnUc6p
9Oh+5G+NfQgmbMEVPORJEMitMkX1+cHV2Be7x/dLbR/e+KAeaJXO+ylVz5Ffw9JfleEX5I1W0v0+
wxT4V02atgw7qp4M6V2TAfbpu/XfArqfbArhjKBmzk2Qgsrhzc7YvkgjwpzBdQM9V0VZ1S7JQSfu
/CAIE0CbGZUd5jzaVE8VwcQpeCnToeAFH6qeFnM9cAIM3+bW1hK47/C+0c7vHs3xgHyKLqdhvcwG
vJzxxSpEFxfBCeiwrGNQrJSqy403UYpcxFP32xx6loUORcrdDrP6y5YeWpHZrJx1mIphcVoH+Qvc
HPsLP0zuxmQLYnIDaa0JqIbXzNx/4C+dm2ufoiWJXNdWcMYnUyGS1tXupMVDAnduVZ5SwpMMKiVB
rJnMEueMvWFE3oMuYoqz1PQ9DNKVdF0oSPYakU43+Qd/uMGdV+F9PhVi7Qud57ZytHi0d4q6Qvmw
NFzx8k5ktw63g+RJicc0bLmKFjma7HEJnZQAIQpmfvhl39ER9/+3RplYgYSdzySbEMGq/3IrNZ5D
T8EyUNtdDyI/iq8j3WQ4H/vDNTvuA4U3lyEr59TxumH7OeUOSAj5WU2y6kQUghSX1kkmTM/X/474
11xDgBR6K6nnsqk/JEgcG7yhICabprSmXtjS0JpsGwCA3KJ8MM+h+CzFwdk5zVELFMhgqIKyoVg3
xFMo8N2pINQ8t5+W5R/5tzwVxe8kZpldTImIQMsDEDp6tEeJsnn5DHs7k7YN4KnPzBrWOUJcggRg
oLFC39E1Oz2/Cdcr6rFRkDs6pkb6bf9Qr2dMA4K4f69QY+vXiZI7z5KnqSYxUPECkKbFq9O7gUQm
9KYbvQoDZJw/oR/B3R+QJBB1YtmGAjci64T+Qus9nJeYcWNRbKNe4S5Fab6sjEZ6MDapA9hCXyBT
awp3Yql0B7zv+x0bM0aayunohAqaeyPuIWKzr4o++0NsLYcHAqKOKkM5w4c54VrOFwNghycY6tti
g6kuh5H1Mg2bTuunSXk3C45h/JV265zq1Wa3P14CUnPrx6SPzyZe+h3NovBffpqJ9EobsiUV9ZM4
LlTQWsLqljiA7Somba89J6hD3Ysrj+6EkwP4ipAOu0y+FQ3uoR0RnVESZ+WLNuYexpOTwnssByV5
bYWWt5nLy05Bwt9o+JdIzhNE++VUhvX5ht2H/jU3uxIOFHIHU4NRnjcZ8xBhxbDnMOlCRM78g11v
GydnbuWd0MkqklNRlZu5UopgbpilrWi2/zmCQrvq+Jmo3tmxA+Ar+mja257Ui+qxE4mQEUaBPO4T
7ooR0teq+OqSc12hM1avIROup8aEBpqMkOknu8eaoqwjYYOX73vWa+jMcDsFbbKNP3rKXwYCZiEd
4ilkBbp81Hh/UkuQH5VKxTxsnN6vwZm3q3BiqoyJZms7zcFFFLzftBsDl1JOTCyr6/VSUB08GJ0h
jEeUWAPCx5IA8MJ4f7WScIk/qvcGG/MYGsPrf1xA6p/dHDDAGhJgM5fYSyc6BELV9jhaoea0b/hK
j16KlmcTUQoq8BtbUYbvgvDE8xlrCIZ987RYAGFUZkHYCYUKongWF+doHuuEREgcw2hgKZvoVFjw
C3CfbTfdFX3Z8C8DOC3xoKkMJGrxyb0qsYBBlPweL6jrj18+yv++QZQ6HaxrIEFtXUWbV1Akm+HT
0xf2Y1Hf9ihjd3LV5KeQgajAKbvS9lDUjKpM2KauKapuuQYDZqHZrqaisNHMHPj+uD7n9rByCbwT
RvHaeVxhXYX22CPjl11mbA7xwCU5ep9IJ5UP8UUqY8CT1H4nGjjVZYGJdqbDJxiP544n6385q+YC
DPP8LHAVFOSzsK+9k0J6irRIzJt2YCZjk3OmrVkK/FoYSBHaQuPnxI0gcCwk6U0RBrZi2GV9F1SV
22FAGWcVPiaFNEICqfnRRJtJPQhVb2n9Cyflc6AsLoQoGrHXQpo4Se3aY/KxEovJFaR2zaN6VpAg
aN722YsNOFRMztzWpVPvxff2LUjYYtBfulgXELBr6I00m169D3/wca7cVtEidX+0kYs50KjVe3+f
2GRHCWYydEI54pb00XEnB34nYZYEfmKLaajKkXYM98sp82BPao42bAdJEbERy8Qbieb2WWBKukZw
hbj8zUociXpAwmRZkVI696iwTPw+2pDVwk/lArefKsVR3ajtOD9eY4A1pcqWHkVycb7oPUkAmsbI
5d8uDrcnOGLZRjjALF/rJk9994UX2iwXaZgnOTXdmJLwu/FX07pDmo5ISvsmojqyuBIwajlebCg6
2560E4HN/WDnMeU0gs5MZq5gB5w0X8tc63Ry09ogjcA+PlxaCzCXTSd1IUomR88ctOtaWDTAB1jz
We7u/YJlp8Q5hp7TNSf2gI08B1/MShU1ZNmCEUf+q6+5KUc38ozFR0YEPDAjBBhyKzZOezl1Aoz8
K8OmGynoA3e2hmHLmlse5YFFigXEGqKEmmQR2I5y3zfOraQBHl2bbawjYcmR5e3rXhgGOIfkKVSK
r0XGt6Mx13Ar3fKEdsUNcnm5B/LYNrWVJ39ezEGAUh0Y0UJxFRdaq5eySUJ96XYYCTFB1q5OWvmK
sPYr46zA550OZO0rhu2vTJMhwxiUbaaycnEUc6J7G9R7PptHc6sae9bHAm4Oi8qCtpLW73kbaOf5
Cq5fd61vmGlupWA6NSoJgX/p/VBoMHzWeR/NbjajxvjfHsIZYfrnbKX9OMGIp7jb/laAzdDk7IAu
KkDNsbo3OH6wZdF1OC9FaT83hqqfQTn960jgJCFC3BP6THJSYVohOh1AjrTaPV1qIj0/3lJmCJ0V
2tQDe1VAlEieeJwPw8cZitFVLqW0gn/AYov1NUW2MEjIOnapK6E6embB3mDqLT0qxjb6jpyNlafr
gsJiwB63aIfSdR1ZCQl56Al9W/uqLV5Sgxw0qB0yTJJbvs6e6e51M7G3PNXEJuw/gf6qaat+Vka/
AdaeqYApOyYYpmJ1ugDmVO67IUJp5bj9m0yjs8am73Z6RZByUNnAn40bzjb5R32rSWgIIegeMjiD
LprTSU29hnvHPUQEE/a/3PPdwej1GkH+95/bP1tubGdf9UJvwiTLGv7u9Oe1LUyL2Gz+1U/+hxnY
SPs57xVfErR6pmTV5cjfj9jNccDVtTHyjMQXD7hGJGh3IJn0KP296716XGbx4gBx/PmjLajytsPz
UCwU8GxZBjBVpQr54ffuJThvG7P3Rkd/ejByXbbhtQdk2kSew6/C2sUePT201zXECjV//OduqDks
x+ShuCbttJONVgGaQErxkgYyEZo3MsHtKdJsQCKud+rfK1gIEOSyFS7HtKTIT86hjWxSvT5DCtvq
Her3GWTPrBuj7PR6RJwpTOwlIEqhDJNN3VfPvmCsWPgPdL2yDXFSHo20+Th9vhaIRYsQdt1w8PgF
Ei26tWwWc9xe0fTJXAihjhmSBUf0bekznjjfWMO7ZKXxKBVNDDfvOnSxTHpjaDlSDvEn04fslQcP
nFXsNW2HPegpUY3VoDd0FwlNwkV4jhDZ6xhVPJ7HL8o0i1rsm8oH9KGPyvmPZP0Z485qyaQg3Rjf
cRNRj1sr94h6JbAXLXj87RcI21mFQOjNv4OeWeWUbQ1NJTry8KPuqYCwNo9HwM6P+0zHdpXfGLSy
OEOXPyujaaWYQdt18J7XzA7vaTZA2t6q8U9sXHX/0lPJgbmov5s5VsMN950K331kVa5LD/uYDkdt
ODAYYEfBTRY3CR5LXuZX6I2UP9+eLifrDUPXgLn9MyokLpFC77TtJD7SnKEuUe4nQrTm7vX6GT3w
ZfClg5HBWfkqx7s27eCujYppGJn/5Prbsvpu7vUrlhafBAZulHvFHVIV+/VDueAQUteiRIu/i8+p
/vImpI5PxKo/vkz8qsWKt3x7G8etWSNi8pm+hOfD2N0Og9WBXGnnrWlHcNdU6ELvhhYAV6+0WOMP
qdtWWqnrVODstY5DuTHfRPJ0hiKS4ozzGzPX8HMBl3MMFo7KoZ6j+groSzIi1KYaWM5mFwn2EyVk
jdNocmhPGsgdSXC8Oxqw8KaPGua48bJ52cf2sejbL+BKMQOG/ZoZncW/S8lNYi4DO1mmjNneZB1t
ithHTO4/fr1ADlCYu4IjW0VHRvhQQvqkYvOruBdUbA5iTNNT4s+VH9et0vO2D+NP46Z9dCC41A9E
vuQuJ5OK7cHY2z1UcLuhkiR1uWwdvli5MBAKTAPJZbpJE28Th6gouJSkKMbNtWLDijyHtBVZytkQ
89Y5OWe1a2+1iSPHdFUbfTBvgVYuqR57irdWX6HChyXIft5dBeg2DSQtH/42rZqpPBUdLK8j4Ejg
VhOnQnNpKXts58gCTEIhGE5I3Jz9L1ahLYUYMLOGK5if9FcEIIBPINpeIvM/UaNcocfi2QJ1QICG
h5jyWmFnrwa/LW3iQjiwzYYOuaoLtGPGbhpqp4H7JWGN0VD7NzqtLQt8A/BCHUSG73HzjW4qWF6B
M13xB1Nfg0Lcb0CooBpznrgyZ5zhSz5LOeTfehs1AEKOYhA/CFyu5oXueTEaZf9ZPTs4xRWL9dws
GH4gvqgBoKrRkXjwJ9HfYWWPhlQdU84QwRBHafCyvCs0cNDABCOl3HCD5LBhwxwtnWPMLBGOLzxa
XqFcDoa4GmfQz1cit3znZR1AcGOy3iRZQgW4EIek+M0FhNuVbP8grwVKo1SOB+U3Ha+L0b9Hidl1
msN/Rje9cbwogfM9v/6Kp2quuGClFLZzShiKni7hPAtDPBNVkLqliUGOPX9UDKi40+mR/isoNkPh
EjW5svJCkL82+UvJE0jd8O061GDuT3kpmHPxm5chItMQaXzTZk8DW9vy+Y/N6QW4HwZruyQotDZv
WEDzfULdCwz0SCEO6aD1gSKpBwU42tJXttVu84W90F6cFHSKiYQYdVvYIRq+PoJJXObXbItXK5Fn
SBHs4RSGfLyjpoNcTNjWGUs4MTwrj2qm2aj0mjTMGcwie8mmxJs7kFDkom5nqkBfXWcDLcaAwx26
JF4m7RDXGS9r1vOM4ydviVYBrzpfnEFHw34JdYu23600+WsjZIu/X4Ogr1qYVtXMCnfhdtkauLc3
UKVaXVyo8lHP77YEAyZA1HoFVF3ZYMYFJ6wUPWW7KYk24iYmD09MLLmEPsBa9BK7Mbi4Oz21kftA
UwYTXr6surdQgrLzd+8SIPgoJ4ItaBqGtLdTBEVj6Lg+9gd6mvLoaiO4N+fyOGe6yYnLaKihxnAS
e+08I5pcp7clVkDQjh2R4TvpaIelXz4AeJYK8bvO8bGFJQyPcfApKel1qEBuFMyyy7YOuDEkCt9T
mp99PUXlLQmz7qoxpKpJfhnYbahcq8ISXpWFHPholJi5wb9lJLN6s7hfVxll0UJVlCf1GKXXgci9
VxB2P4OsFCHEYr2Og8VTGRjh4JTcYDUAx6ALrTJg1A7f2upVBAfgNcZ6iUtQ8IT9N0Fy4wd0cD4U
jMT3O60JDOPhjdsq0vhq+5cc61B1yNcd0rL1KtgMFwItKysSl2jC9m3Kcpxo1Nov6E3qDMg/lCBb
oWJB/8J66G/9ld9ACiikDUuNxiBdb8wA1SE71WVpOvVPpHEcpC3QyBNFe+Hef9aEBh32t7TloekF
abwAt0e/f8H4z6n4Y1Wdc6SNfjdQzruyVjWZv1T/n88R/X0itM/Q6SDAgu+BBdLD/x7ysWcUVu2L
6w/A74kMEiRosZPbcRm1VoReoGyL8HTCum4+S2qaBfXItISe7AB1xhN7vm/pcG/z8jbnl164cSW6
C75ZV1pP2x8c8RNDgrp0vuq+f+xt77Gx6hU2KIxiuutUZXsBey4lBc/copa5uJtT3netIpT1a4fL
flxFi07rRU8akXX/ncxsKEvUHPZb9nKs/SwbQXRuW5t2Y18fbONo0lhz20vLt2m2Qc1pdfivVoxf
1X2TQDrLFMRr/z9JqTs34NAAYkYNv3eBWX/rNpfjdgJbhUVrAOXe5u3wyAS87HIumqZWgEWejdi1
M4xYmuWhIVcP+S47PUNzZqths4HdTcRaeUnjdRrcrrNAPH8oTkKlfe/WACx2iAJ4YOqpap7n1LU+
UWTPJZMINYRgUj+AudG6SrPU7/k4xXGouM5rtQsjiMZhP8cLmXHbu+MeGOq8w9YbFfH1kywn+/cm
cchqbJoJ988UV1D/ljXrf43H7zwddBcqpfjjk6rsopCrDrPrbW8eZlH1VoqVmsJL/dCEPbDm0GHS
xSEMAWxVY6QB9vNnadimP58Am1hDOqQqgL+HJBhTChrLuFC5hQ+/FHI5cQ8Qs+G3Y+zx3G3llKPn
EXYKF2wmo+cCUC/1Rxo4uf1eUExzfABhSYl0vWjlAAPcim/gg1yzRxAOil7Sh98/TQM9UuIReJ7Q
Pj/iotcefWYAtFvrnANA1OdJM77se8r4DfwYNkF0eJ8hqEZBSEiYGLutQPJiMEljuNbwLnaq/S39
5T4lQAhXw16j9fwCazJZhzQZaz4SsXk9p2XGK1MjUjT+1oqCiUeB4gHQJMHiIfdanbrK3vppYoc/
I1yaLm7ghOBMGjhioPMBguplgAFmIXCMqww8hO0V3PqGZMDLURL7n7X115aPKgI6Wx24/skZbowj
mKdniWn65YV9aRe5igBtNJN6i4pBjjEPqiXqVSile9qzEMw6rl0mBT6kamhu/ZUmKyhwX6v+wgY8
lch0GZPMZBSru/DneJauqyZROP9Ie1e4ktPiHND89QaOXmw9CBjPj/DGvZuqxEXq/dYJAIz0SVM9
BFCdgVt5EYHN6aRIvmD43nFN5jezU+deix/HC+/oPFOW/2IGGMUKuDK26vJpW2eoT84FBECNp39t
AdIGOhRI2U3v2SleKrvRUZJ+D27Pl8a5xSc97DGaRR8sEHyMv6SWehY7il66TH+n7jbJgXZNI8wt
ppesGK7xPm8+J3yNYV7h9Pv9miZNYzjhrRHlSkkwhfx90+bxUBvA7GjpYylvmV3xWp54y0ymObbU
827/8mV24zM7H+dGjxHhbPq/YijOQCwPyZiYwzhDOZrYbR6Xc226BLBCeO4UPnrv06qHMuri5ygC
Xa8XEa0Z0hHwZnJomMs/a/3jAC6R/4Qb2B/MCUb9XhCwmGSo75A6tDLCHPcEt/uddg3LNTOhNVVQ
7mF+0L8zm8Zy8mJJgFMcw+tjfUsfGcoLWyrO0E8/bHdkrgCcxGdnNl1LCjOohZoPzaQhipSrrutw
U1i6qaUua9MDvpj3T07l3vGjHH+I9ocAK05SVydD4Xr+hc7vZ4awEwC+T6Y7UTL73mRtjFOA4Y4J
Wqv2kOR4PMl155Uz2CtJupvK66DxAGqIdqOGLiLMu0hhltSse/k6GFWngnqyzv9Hm1C0rI5y8FIR
66Enfz+h7NxA3gjDmp9zvQttLWJxNvW71M2w9GqBh4KoZFJnJWpiyTMeGJY2b4vCuz5K0g9cLK/0
0I2FNWWNyOap2Qm4qFg6T3ZEAeF670fEjiEMUZYIE92NBVecfmat4014XurLAZp0RISc/3pwW2yL
YlXxhS/CWPh15WfWgF3zYkg0rDoSZ4Iy6POs5Ie6R1uLCiIKvZ8a2A8rVo1vWaVHLTnDy30lg5PQ
p5yygttrTHGFVSd8mqVDUC1A0kLjfDyKIHAGW/bTa+/VA+ZxQ+4MyJIV4eeUpyw4+jpTepQVuVYv
9xgBfBq2rbG37Zoz4AwBouCV2yKpT72WorBC/oRx1HYsMkaSe9NaRN7ESohOxrexNz6/xVaZrBU5
nDAGqu6yNEh5ThlAki4oW3kLF+u1pNHy7MQGcUxa281bfHvgpU6SCgAMz/cKDOFv1MHLC2v5A2WA
Edk2NlgmwwtjA0rm7vgsrg/Z8ImgmpDh+vjMXGHwc/U0FMrJJ+JOSglT/9Yrh2W3Ms6HqTOkgwEu
Hz0zGseL2Leh0ZGgZmqhxl/Oh8vEOs2iLk3gvdecC+0WSZAG9sjrEKlxIh+HBHVX1NDjtwkH76ui
/rhFvls0mE/S3dQF/O021woCBFd29ytvBpy551bTA34iF4uIQBfySt8jrauanhBHKVjBspLTR4If
GRH/gpBYrQYBXQ8OIPfVIxOAWw9S3f+micIWhrC14nf+/44ERCR+eoOzSPuCcJXPNbGNcYXDPQAu
BM82/IaO89RxmMATAocspGBTlc/GEJ0z9gtrHQolgzIZg3/tuiphbDm3rt5kX3INgb/sq37+O0/m
nvITc7IVgrJdb/2aXdvP5H2KcbMQqX/BV4HTfi9Z8sH6TM62p7Q8+zm5amkEDFnrxksXEGu+UXd2
rLYv++s1X4CXL4h1B9Zo6OmWHiSZ40R5NmLrYbbxov9RHHVYa9dW/KWPkY8vufQmi3s9sMtJk3uq
E41rxkdCqjRcwOowWVXi4txi0KnhDkmeY+bqI6VLgb62v+AmyE+WmaBtP6EwpCZt9WX/MK1Gxm4r
alLPSMpv4baB/8GUzM62/fUikg7MvWXek0/sqGEkGRP68hVDua3SljPKxmCM9I4Lr/HXkYk76mit
Ce1B0QFfWWIWBSNhzGqcvUt40oDosAzHip2rkmn6HUcXndUxpj0DvUVxsmnlEx3V6lZcCwlU8QUe
k2oq5+smq4/Hkk8Zr/DZ58Ld93P9x+3dLywN561WKzybQOxLBMYEaCZujvEL4uQh4TXo3rlXrtiQ
kakN3c8XMo/M/okroxPHF4ebYS0WQWtglLd2BKj9qYjp0dnBOV1HYHeJ3TxnCf4ykun8Q8EzHfC5
g0uSjJ3zQyx59C6efINSGgLTwlxLxq9z8siIOORENMHxIlkfLQft0D6l5R5xjpXdpf3Oaf9VySm7
IBetImmQGYzP6LKQoLENUvremnfP/dcauI/q3+0ejBCRltgBwG3r79RXzHQzHXcTxjXMwRiNyZTn
Ysp3gGs/B+X6HeI++SDcAjQybgtb4IBikq4GH4cBT6xO8CX73rY2N2EbCODC5sUDoy/O2DZQDj+I
T5RGyaSNfGJHdSfKr5tDznN14sNXIwvSrUFXTr/hf6wAtA4xZF5g90F5i17Le8HMzKVl7Um9+mjh
yYXQy1ixrsyAPz9hj1RtYVejz5yaytab4U7h92IbXIhOSBa7jCI1SGq8izRqL/fAbGN3XlHqM/c7
EjdUFdeoyxcszxDDCS7v/m5EvEGUu6grukFG5jKfaWBkrgq+7zpZ/O8yUR0dUyZgJ5hU6sq9KR3c
AnTvzXmdIepOOWKjV03HKF6e4o6gFIiqsGpjfaoCUOhWxGCuZAdqLp/eOzB1eHShrhbyj65vzgBh
qBZZDPxl75ISMFKNo219mLZMRUhy28+znfzUqFiVqju+p1c8e6r+140+LOOvmH9GbXOIRGuljrPo
MIxdN0MKGlRvDvUBcqa9QUgvPOoy6ofbMzblLM6s5M/AjbRNuoHnql138NjrjaiLBGgcJ4MKZj/C
zmre6hp+uAH9Xv4F/rmQ78oWdVfZ3QZuNfiBIDs+m+ZKL2MwVQB9I9MBarNB/dOtp3vF9eTaBTVu
a8KVvxfK1YzakzfDWX3DVtitqrRxbE+GGFZXdaho1W+NhWeziIlL5H+zfcuAgP6fqN4IRY9UBHSu
Ny2AQtIDzIDRDvBLowc8ZZXFcGwDvCURxB/5qdd4Hlm1aOHP+4Rep/bL7GdqrAgDFEp+kQhgXME1
0IbxRLjG6WCI56Aj5bvbIBnv5ITd5IHnQHOFbjpRlzLDNLVi+30JMXcSUs42cHa82o2tdwWSSMoy
Bn3kN1Fez9vqae3YKr68DjElsAfLhBtWBWfJtRpMCJjSo8tSNg1YdReCky1gitdzhDVJa5y7HQIe
2g7Pz0Ms8JQr/Mwd5K+1jsVDX2NyswmsmkIuvIlNiy4U4IzOrfjj6zDHs52hVfciMp2E3oWPeAbT
fYkJrwonfhw5c67BLsmvv99CV0HxKRtU2HmG+Id7MAzvF6uD8FAnI5LRAiq0cpe7BimsCKck1Zn/
mtAOzs/St7IkivJwvjpMgjPP7dLg2ghksQlhQj2+5SVoR283VH9zxhxqbLtl03cjZrRRB1Zi1Axe
ooSdnadETfESvgN7DJGynbipJqNL/OpJQUVQRUeD5Zio5+h7TBpUZFptrhrR9uEDkUyx9naK3u2M
Urftz7WJHFcD5PTG9mJ5I6B3LBPO2PY8PWZN0FZSuWY3dz68Bo6zAbb6lm9rdynR1beCXoMEc/kH
yLexanI/UZUGQnUn3Ff1XskM0YD0XHPN2Z3Iv5kPqe768D9lCQ6rRKs9z+NvLeioeHwBm0kft3PJ
gB+UwcOnJQipEytVTkgSRQez/mZtzOtKjciFJQrNlsI3FtJHu73Hrb+jWFYRqhQIklg6dcZi5QgU
icQL4AbGZl5gTTRyThrwrHnIicwb3W7rL9wnaxol1YnxizN7us9FHUbFXk2d45//y1DfSDnY4Nt3
5l3K6FHO/7oYQS1m0XFaWBEcnSVo96EcHNxXPIkfuyZd5TXfnuGb9k5PKUsMUBNRpCdGZ2Q90b9e
6aoGIBS720oXXNAZVIGfOBZB1s2xHo0Z38xAYu+FtiRrHcrho4cFny/ZJmy+TuJWvE9406pc55VR
wpAxbtzS1aukYEU12FiMsj9BMbY4bmLV3kEyKiGoxPcNz60frShxqyg34C9MN4Of5kYM8iQoKEXI
VG7keQXNt722knyjdGfpA7MGP0rQjP/ben/pC1g8TtkAG9DZS6QEq+TjQj35SjsV9D0QeSImf6jF
14BI02vPwLPqdBIy6Abd3yFDhu/rqqpZFbc0Et1xVfWnrb8pqy2NbPgMW40pPpatn+Y4Oh74uu5+
90xL1XH/bjXpSfvnFBlvvFQq8h89v8M/jnKH5Gx+PmHB2f4ot2o/QtViCVIcCpERFJTGpTM7ZLZQ
ts+8sNJ0sZYMWyGtV2dva48vY03IY78c08NPYD7r0Qmlvpqt7aEHcKBFG10hNsNDDqpP4Uos6IA5
EoouHUm8Lk6i7A7QdFlDMJTGjJ4FY4+2kZa/p91EvjnEAh/rtSGS/0ZZcyEuxE1o5urAeRrJstbr
wrXQyhN5nkTJnXsqSuduNSYZHsnXHnGgkUqKBBarNgfVL9n10rgKpdapHwxpwjrstVI5WqIDaDrE
u4Oq4Lrmj85sE+OGDlbxQqh28EUvX5iDGAEczjzlKk6tezkIYf6BQJhdyYWaKCaHCd0jIIHFUTM5
By+kWDxkpsOJ5/58BRCIQdyu0hNGPxG1fe4K3Xfm0nWA/S7L7tFRmXQxBpdflIg/DgOwsPxZBVcY
aZIV092eGc0Af4Y2VMs7HDu/ftKg40fSCbXMDAyi868nWXdr3Dhlm3VueyDbsZrKXmAt4gIQWB5T
ZK9Y1+YH28SB9oTLpRhKDX5Ciw8ZHZDPS2iwBnXSPAE+6zN9QPai/eFhqMyoRyagzwthI1zYJ6jA
OZFV4J2xEOOc/eniY0KkZFGFr7psi7Qe2jhkeK3qHbqm4/p1b9uogHFZSviPc4ATPMFxOH57+2WV
8OpINPRm6b29VQFonjafHHIj5oM48GYNQ3oSO/WHClsh2k1sPBl++HJwCtRAIcVssgCpBnxEwUCS
lYPD3aFmOXAm+Ly8TyCKLJ5khLvoPznAz32Bomq9eECWbm47Mbn3tqEEVOBUqPj44NREk3APb6S9
NSCDl47bt/T5rn31amGFEo4WQZe18KiU+iRe5pn2DoXTuErpEt/ztlIbLKrHAROCpmaWSujnkZvf
6TPLucX9MC+n6VY9YhN47FxQ9ybDn4b2Gxg2F+KCXWQTTCJHD8w98x4Dg55uMZ7f0OZimsGf/U80
xzZZGRgHy1glKpfpnstes2lN7pjCWvx8uncRmYXwJxjj8GXwQzLa2nfSc8BocFywDbwnhnYuQ7IF
SGvbY1m2gKxZSJqrdZi2AOaMnzCTeakf5QhpzH7M+aF3wqWbD4gU1zLkIGXCpay+HP0KQxcDBPYe
3JoeSLiari+lINjK3fQx2HNwcPHjGvY6G2aKi0ic74yWF8gg/kh2EjMISDo7gDERQPxH/xCv4MEs
g0ieIXD9agoYSVF9iZuS43ik/gVhVfWa/YMf+p4ia67yHF20YGPnzCnCsn+sULafQ3Ch8D175TfZ
3eaC0p0YWj+c9WP7TIFF3HHQsYNUzEPu5vqfd4ee/23ifE6BCDxKnSf55bUI7fZlshiTZTCYM8iW
iS3MxZKJvUkrj+eYsvQ4Kc2p+9MOW2JkiWROeJ+GbbFtrXYb4QSJIVDFRuoPLovZK6NECmOFKdSY
1ylFIrD+Xb8Yl3ewn6YibxoimTDbzxRYwFgeKxkJg5jl5Qv+piBYB0IITvHOsPJDm/UkA8mdMmjC
ubkcw1yfIm6jwn4ityXhs+3K5s95poJbzVLVudJH93X+ahKzCl+pIGR6vuz2Dug7TMOzE8SpptVS
DZhhEbG8elFAvukDzN/cOME7tX2piufipbSXdc1kdLJDB/mgz6mBt8HTF+Z5y5D82Z+mVUtWEgt7
qfQqn8vCdZb1jpwZAWZO7A38Lm187sR/Faeo/LV1dW8QCe6RGtQuPhuj8rEmVEL3DVZXd+b/OYf6
JaYPWJ7GAmoDrGAS+MGZfxIEUtjM/cgT8+IpGeNcDi4hixvgJJesFfqJR9pBIj2aqjU+/th3zQ3K
LfKdSOR8bVeGi3tLo1K+VAbDe6PUsHZ43Wm4qCNP7zAmIxb+jIQgKHYYq5Sb6DMgLRIdM3dVuPJo
ruFg01fNqjl/zhqp4T/lOdf2HAENfuqcYUGSIqCXsHIVOmldkoc9VFFXNWZJtBZoFHQ7/KsnK6rC
N3uXPokfZgDjveQz1FsLYz2BlOdvkNhLsJsCK8qfSZXedyJyjDdtfKwUpjtX3RHomiCUzk2OSzyS
lBaN4o4n4EuEiwOluzzFkX/c9zBjxV1XP9hY6W0VxUp524pjQPkxDM6zYaBi13YnoVpEG5/Rp6UC
E00E775NZNx8uU/IoXgL0AaOR4bNPngUhmNntckKGtjRaFLfHjqzH83ldIfBvD9V0kQh20jZW0R7
ZJE2MJLwOgfH3wOynzvKhQuhzTieNH0LnjNhcb1s6t3WaP5ua/MtOEgbrxWyftlqDjBhefe4Pabp
9KE7g3Cuc9LrskRCB47J/i8yBSflYPgPYheLMX3n2ddD///xjT+umjTaGSk49WV/Yoa0se9Mr3Pe
Fs6mkuMwzq6mJsAGlF8CLaG5B11MQi3PICBjV9B6jYChAwlKJMS3fmUu3LPonYNCOW/AJ0fzUpsO
0ZXYIWxQqwA2Dry13f8FQEl8xH2OHe2iIvjaLaH7KxQaSD9WDeIpotUNSropqtj6Uz0gkoShCz+W
60aVgNsGVMSx3lbOjC4dco2FNX2wg8ePY3F4of2oOCPu4BSGKbLGMprZrPhbpKV3vHhx7Vn5h5I6
N9fgHcX0jQtoYJkzrjzmcV6XDAg8j5RtVJFR0QoAXoR6/lswJkmXd06NP1i5X4n1w3FGEzg0PcoL
Vm0ykbwvXNL78JOAGX0TGOo5ZNDQGDkbtt7wc2bDz+7LWxPmKZXwgYimTeE48CdJk6RBUltEn6ep
XTFFbY53o52/1MGPzqS1FqND40PcgkZQloT0S4lNp3vb3MEEsYEdz9/lEgPW5/1sI4a8OmokMV+9
+yDmOOQ1z/eaD0olBC4HRqvnj1PlBFFuCyDnSOHZpewvcVwbGRxL6tIzrYQmbmAtKf4GRcLgRJYQ
ipoHhDZRonYo5NhDWCmVWtUsuP+266fexR62EFY8CPQby0WpjgoCoiRrLZEpyWEqUCdTDAbdPR/B
RBvS4ZxvOGDz81Haqye4sBHwERmLDIGbaVU0b5ennIB1Qf0iinA8uRJKobRaQrFwmbdOCL9liqD3
ZywSU6EJN77NyNbHg9zYTCSxAymJ0l1iTpHdbpg34bFClg8FVrQrAExJyNM0K2TXCqfaEBK0OAGZ
sYEZpu26aK3d/L8qQDUH164TjHisIkr2IMUbmZZtFyjEMdQuvXvpq4Ed6mcwcl/kGoaMjSOQLpah
opg6aDB+OJO+dSoiVnSccfT+UcXddVQswDuC9WVL/tBItw5eKZc+uqRnBJqfh+JeDsq4KwzDjeF5
MD5Uq06OXK5uwkJCBduzWNtvdLi+KT3Qcssr82pAf8dBD9cfWKzNI0TirE8DXIbSpJgCasnaiekD
erD9GdzQIz7tnaByhXqg1Pnm/SX+51DfP925Z6CI6k2w3tqbDrUyGvx8BXedpK2aIa32UNf+J40g
q6mEpQy8yZaURV5LZkgtwe+AGZfM8lNkZkdwEIN39VD87SSB3GCRgM/ui4ajtKFvRrjlDpLrwjtv
KPnzJ/dfRrkAtb9g7FtKWgeLhSnhXt8Iln9H9L2V0POh4rBzn31mjx4JkPLPMrWf8SpCnoYYMK3Z
FSsRVTICoSp+cLjx45mMRErFyKbQUkZyFBNSn/aKhAnVnml8tpDpRSAWi5C2IoYlG+6RmmOxAauz
WYPOSipagfJbP/ZgBWjaJ2Bd2oxIF8HMzlND1TXdmu0Fq3gPDG3H9kgDVYClNUTTOCMfkwP7Qn+b
aIOfFp5oE5Ki/tB9CK9MAzw7YTZZYjqnGbmqrYeD2QJNvH/ML+UT71uE2s+NzGLiQnNVeFmFmfP/
ptXShjTyqu8Ng2y48KDBTtWA183FlmFPn/SEVtjcBJiY3M9g96ByVnguvzS9xMgt1we52FEqJed+
g10wMlzbySPO39YjozcQh51XfzZdBIZKBPpXaCyW+yM1GWG7pTlHk1Tv701gw1MmPKF8cFoqD/5B
ECxP0fbtAyw/L09KA/3XS3UZMN3GtUROSpHrFJhJVvT+07PNnsZxj72byCAIU1Qfm6Xg+FE/Ke8J
dFpibZu4NO/p1y+FbTZCqTFoFXQLXiw/pBrBlVpL88NM6mFbxggw9/J/duguo/51IFPl/JyyPw9a
IUFXUXLDbw1enrEPJev77hXwSYfT7MAvnx3orY/px92m6L97vooKNYzG0lbrLKUNQiEDDDjuUNBi
MTSzUxFGzQjxXuq6pqB6kkja0dUBibRHnXzSYjg4bA/d3CMXt3fAjeNcSCW1oXyYJeibJLcWfhie
yxk/y0MqZXdxwcBrItkBITF8CPecm+k8dr0wLX0CIXWQ55qNy/0n9r5F9kIXFIUqaXPFC2SuFQN6
ODfZRRC5HesFjgy/H8rbvH1bYjGhEx19PZr1BOZYh86FbV9xcWFDJkU/6ofQ4EaPxbax5ybeioUD
yIpZPAcZLOLIIZxc34TGdFy1jzu3F0P2hIJpcbuREjZ7EJd1Tvz4dwnYEG31LlNTffIOEP52oklJ
EcxFG+qlJbRSKrBUxdWjwuJWjabXgBN6183wY0LZuVRsgivuLX0aDw8rNWfBVAYgIQ5iufOmYbLS
XnCRH6zd9mqFPKbhmTk5kWjzri4VJAU016nUlOchTCsgHgGc0nWvJkmPyqwD8v+lYwmGS4GtoCXo
wJCUusUBtp2xFHTLLiYKRieLH4YN4gUhkQ4FDJCuVf1rVw8Saw5+LEcMufOZ0mobd5Hv3eSHeAPQ
uAK4XWy659AwKGKJUFSVVypniH6pxLzmc+76eD2ijH1rvuyMxKkrTY6dK1aDBLLPWxuMh6COfuwm
aQ8q6LP/3qYCrvrMnGrl56gDNo8eeji3xsQnnFf/5ltb+g0vpRSCUTt0cgzNH86O8UKI5L2PcYLF
FcBWETh/IXidLviyjpkc2HEexAvmBbIfZ5Vi7/294Chylat+IkrJdj3rD2kPzMOHYlkgZOZbfF5i
fjkQ/RZiDUahd1jLwsOF4WWI+cnWB+UZJUuiHzzfd2+RpURlHam9tJsXGQkJXb07OJznGNEArsRT
miiH6tcTuBZDPPn984S7KfTzaMbTreeiDv9WAuDQ0uNYP8aQrgt/DtTdW7jBsS8R7fAv4yHzAGy0
hx1sq45jqoI5/WoqMqHpRg8+x23Q3XuclM7Nge49NiPIjScXJAhG3Hq51cfb5hMYDYGelm36/Ux3
HRebgljE+6FD0Hs1t0u446dDxHW+RWlNnFqU/zyMqsDD3MIzgBH5/7VMA7lh6mkHIuhvOHcsl4bw
9U3IZ76ZYrLiBNG+46vvkpohG81zx9tAlMAdqaSBtpuEEZBur76wuT7WJYMYMPN+lg+hDG42ls2i
ipIgz8G+Cemaui8nfR5C8LQbHVIIPnPl4hE9HAU0bCCLcHEWLP7MKNk1ZRqakx9ixe1/u6dsP+w3
oTtbvu+rqheaJuXb4CaFGK0TRtE56yRG/1feUB3Y6CTiK9xCnH+UQvU4rH6BG/SmhcBNLT+Pf01M
ITTUYh/MK1hMj8D2tjgRh2Ndtu45YIskwJhdOhvkK/tSH46DY3wDHU9EB/q9hm6fLRoyn20+X7Mk
POcs96SohxL3J5Rh+nQJTRrdvwYoQV2Fd6WbMVLlL3/V+Plr/XEzUenkurkYSJ2Vf4Omkty7v2Hb
E/UfCRrtSKrGAwncSls3vnK1uDU0gnUeCGXXa9w1Trw2HXDyRCQd0bT9pPKJxcutzuFqQVNa1WC7
c3Lnare4DtCscQpwpXmkqrhzqwNjUJnNQs3kcwvuhrvKBSmPz6RAailzG1lvl9G382luFKMy0eUy
YkaVku2YgULsPdcwbOEnvpFWClA9gzAPmvM5PMuKPYfXyFi/uoYjy5/ITFckNjt53gEEjKsQtuLA
19MfLIrPRKYSPV9+Ic5GXTZOcW0is5RE87p6fk2M9od7B3s/csKenhB0RwGX56sJfjeNVkbbAlqF
cejYXI/QXyATO5zgwp0LOy+8quzx8lf57PSv4aGvU2NTaypAfbLh2XwCrECTKs8Ka6cWGGPZxh3q
LXigHoTkgbPBl9r66t2tR5LwG489DiI4/wp7bgR2zEGc+ofesPihNozSz01Ll8RmmEJmFfryOdQo
HNvwTgDJalGAUUpD9OdFoHqTZq5rCaLc45qNrq0OwGbk10ytOiRaDGPy0lJ7nj/0PfuJud/CW/7J
hM4egBRIx04u6pmQGIUwftuELExi1tnfevR0/653C5dvLFlWRT+KXc8Ohm0feS6Ojq2wPtaeBbqq
CxMCaD4tUIVdoVKJn/s0lWAGFkqt/V+zvK+mgohc5YGPgXUUgRk6+ytRmXhNNsWc1dlyGm/KHlAp
2gPyk/2/FBL8v9kmc5ovn7howaP4kISuGo8gdeOXclx2LuGSbcZ2C3JJf04CF5C9hTPK3yc2G1O3
+LsPcsf+Vadku9vLxzpXCTRHc5QKtBB2Xdno2AZqw1NinjQybPI8eKJU86w4EMEvHMyk9E1svCQQ
tpjxHFmuzqAFQPXrp0rJfLZlfbkKgXNUAgmxWWTpaRkyUivf9qEJKI7Oh9D8ySHMFX1jl3SR67z7
+6KrgVO0B6+FcJ2gOOMz3RT1c+AdG1x5jom+SElvKYYZ9PkL1pTji1Q+ZAWQvOeNNsliiyGBdUhH
zaW91Iu1+3uq7hnZqG00SrjUZcaxDZN0nMpNgCR1cylXgsU3ewzrvlxnUHeVy2IUcaLllDIWeZEY
OtPUpx19p9J4D3egshVwD9wECe5DcspbDtQPbqGrncE6zZzxKNr3irZN5WKgdzLoaJBn/7qUrEeX
thxnf/X37d/U/D0w25xmNfA2L8jg6vLNAqtSvQSgboJIMfUsfjJIkbe9PvdkgegKnZK3igeneBIQ
jytbpFDjiICvs8ATAMipq2p8WQTWWK4f0UOGcVbyxBKMnovwAkHsSQlls7uzRhIKmL6Y3mfVzW7s
9TykxNK9QmwhIOctCH8Isj73TjLBnRQCJZ5+z81JEfmnd4ac4jcq31v0w24IpZ382tE9EiDKjIR3
F4nRyvvyBdeNDB4oP0vloy7ro75ZS1VUmg8nR4XcLLrr/ZFWKH+MOfvwwMXgYD9moAZFJYo+kR1c
UAobx934pVnr1G1fgE7au4c1RupZ2HTqdQukX/ENMTxTeH7zBhWkPmUZYLq6JOgLTcTueOVEe12+
Bu7mODRJVM05HsGdnN3SJ8oyOdkbgRc/oAo0db183yhz0q3oaF2caOPAp6A3Wm+8r87rpiQJEYx0
mK41a1BiBV2xUptwjry8VCkHmVGQdAT8JC+RTiY2MqVsUR1xu12GME4fOLU+O5bPfIkvnmVcq7Hm
PC6jE425jyj5g2YnCXf8yaoBLkpgi+U7eZzX7jhf4AjCx3B3qpyNlXHnK/Y31F1FcIem1TVlQ8/V
MdUQTiEDOl+xts48z8cwPTanhZZnnAtHPqVQ0KzojnMbM/MiRgBoS6liHNuPQkUo+xxce2797p9O
9td5rW44MCLPJOnLQssZR9mFZevxMdVkfMD8RlCjBYVKtD76pvZkwoPHgroohymzvs/+cCWj0S8H
IlNxUPJeaC6H1yyWP+fpbFQGcDIEi70MoC2tOEqP7WJZni6I2WNQ1PGhueo8peBqLK0mxoXNpJcf
TFEjabo9VHbXmEWrsDM7Mi761TX2FihTwj2Ly6liMk4dkFcBZmdjb+oOmU9TurR4ksbqVZuxSlKa
lefhtwd/AjUjFFY0cRm5NrLxQnoigjgtnlFQ7UwpDEO8ITkD8kmEJf/sAU8YenuKZlXzb9lBu+HL
ydpWTGoHm37ahb8ocm3+fv3CBWEVCuYLv1PdMMw6GiUOrfuhWekn9GYtqGgsep2yqqKrF0avxGBQ
jup/2lFp1Du6K3D1sq6xTXMF2lYZlU4mTHqtOyWwP9H644ITgINq6WPJ7QDy8alZcAhFdn9+8CLe
Sk2+fWB25HQxvIB0eC28hcTRk87z+YwIwZE/xPGlPIVA8ArQkZc/n2yjvUTVSr+FR8m1bElsqlYM
rGzj79fzX6Q/yJGxQjbjJskXEl5H74A+rz3HU5Hvlul+C2g3Vwyk1Qd1PwwxcrbOmIevutm/+zJ0
YulDWZwhn9L6/b/deWHLlMvEmHy6ETlQjbDOAj27YrmaFpJp6l2Hmjc9NQ4+CagNIGM2PDdsvvdd
shiCwiIA36b8AT8yuYDd9flE4Av7d/HqyKxaB/X7yh4j8OKUPkgOaajcbLCtIx93N+Xy3edQa+v3
MuziFq2rK9wsIppfmKsTSidkXC5QRqybk8AHBAlZWxxQ/nWqkYm6b53LdRgxsH6DZsK7v7ruq0vu
//3huP9IsCL/y8xDa3j0iE04Wep6Y3mukMe00wB1lodUAcuKyLFzOMfQNFaHBdo0We0MYWLCJL1t
LV8wmpyTQXKOLJO7fG4H9jsKvYYFamKrfeXuZZH/blbdN+lG9cfPmrdQL+ZF2/CACl6mXbom9SG0
xjO1nhbquJsLQmCxzASoblsBlUNeilg7DxCv5aQ3ejcq3pKk9fBb47eE/+rEvrENGguTHjE1fX6m
93ss5QWPZxCOYN0LgWbMWZq2pJS0+PJ2K2K5j18xmylnSICQxHdeyO8Psdm+w57crGGtbw2mLouo
cHmqv5NP8lbKhx2CBPA6IVePucQk3DOvxogImQRViB5dqGG/h2LWaBTeNs3ARbrrtGcMfscaKYuw
t5mq0MFjBIg1Em0c83XBFDaOxbVIGz4DM0JesIlM7wZfg+f5vtoii6foLhqriub5iUBnyIjhgtKK
uDROCrLCVaFESMuU/w0NBtFxj7J548xxmYJS+gfC4R5dZpACgijOhozqdMKb12OAOfnUYODkcHcL
Q43x77kL9mCUlSnjojt1ep2sicQFU8Dr8eRaZJMJYn7BrIWp2trs9hd0jQjejP8g0luxXefFLf6Q
J+5vh1lFh4fLxjsuEgXsFXW4dxRF/bCvKTrTpMQj1+VYDvQi6rqPAyBk9c25XGgaeuUCJh+F6A+/
pWtZ+rzel7BVQTfZcIlackeiR41UtpQ80SK5xAPnH5W5ZkmXmVQanw6WCB43cFEfH/1PrpNijSJk
LVJiHN85reTXxvb/heSPjL2sKHdd7wWN8Zsuq98BMTe/jeF8QgIyuUlys8bCk/lYKc03iPXrJQuj
/mn8xokaWyQ1QaKyv4QSVD8/8ccudofWNCDZWUJ6P8QL20GPFzXmf7c9Eea+DeZd7JYB74iBLgSi
wmCA6be9cN1ibOjV3nhkbgoXUY3flUnPthTC0f2QpBcjo9gOoyDIdW7unON+vazm7RuCY8rBgYKG
neU5xih1ioX6edc6BQqr+hUV4uP4DuMid0odVQL9unJaPPSng8syXKJ07soXGfpuWfzkO2aDBGVb
lBNedOJoBKmMUtDxl3IBa3OSpMtoCNxoHRerJowdieW9xJJ1dFsBa0pgLw8DscTwUjt9hwzzCpu2
jzKfbOBdR7Ajh8j3bUyWMVbN12qF7QOJ1GCZ4vCH9brQwwAnGCUL4SWxJQ6Uo2mIkew9d6yIgVLW
svJxecJ3c8sN+mNi2BB0Zx8K7/JSIqymoePntR7Ux01gJCvY+x6tTWWwd1I8c3ts4tDyTfxY48Tu
YF/9RcJMwzzFORB0djyGSz1UE2pTkP3R3fP6SAizr7KKixwuHX4D1csLzM4BHbHQSVpE0+zIaMPw
wSrm1WdOTr0J/4bgbkUkYuyRvGOQPWDULVvVmOWCHL0okHWYFziOqt6P4YQwYfRcXnzGnSGJ8ahl
Kki0JJ/kE1qlvn4Xo7gCvYEvWSUeuyLkDE9AlPZy7kXwhUzzN/9UkC0ZTnHz69hWkk5IhvkWquVv
4ri3dLj/HdUXrb3RuVzT4oeaaWC+p545QozBCfkcNcmoHJ2t6Jh82expBmjvyUK9rLD6LC1s04l5
waxtBdfJX+rQtPqda9VPgHLRyFkI/PdbYP0LsElbnaNhKbXpMdBAtVmpoVIg5UWmmyv+P0Xz1kMH
H4BRXsQ2jq6k6r3ivFc8nAZ+gB+5rfFg2oqa9TcV6jLlx1wdg5tuX3nQl4xzJgrKimoPJYpP3WWt
hIpKJBEn41UlGb0Z1yKSxcE/QZOi3oi1akM9ei1USiR3WG+pGTJPweYneU2D+qRdx473OeTsMaeX
4J6x5ktJTzQJBrtOHmvd1ieBoGYi8OzTNN+R90Or0RHTmqWrjn3G4Shrt0+7PlkO2/U5yqHsqI0T
BFyssG7rXr9OiskBd5MUCpB0U2RYuEJMtfOQNOUGoFd9kK52Oy9dLDvRQVnH/ai08XtN2j5R7tup
83/BsjPNgOZhsEHYxyvTJGw+HYs/dZ9ey/shsTGb7h9B178OACU8GkUFJSsdvG4NmW0TyiAgkF/4
utzkzs2vannEAcGUByqxtp+DYgSWplpr4dBizSRYw/qOOk2v8mH/rtCk4GObtZuZD3dNrUYwh+43
WimPfCLFZS7sMvlyGCjh+dcV/VAb91FwnDhRWRkOzuqE6zRassZxQZZOaImW0CEsbga+8Urn2w9a
/JPz+wod7qajx9/mEYMe/GMLrmBwIuYDvs2XLTpHB8OSjokI33m3HXerFGB2+ToTxXL9na6peAhQ
d3kemPeOXNhzJsjvp8y/ogkp8Ch9+bzEqQZ5rHJOslvV7rY7FFDLGsV8ljTW1KIU5AnVDIeWdzAW
zeizW4mIfLSOKdKqSnHoQiAyY/WWiR3/jJV5YuvJfISts0vm4r8EyCUm/krHnUCfOFYAj7uA15/u
lOKhWZfgfpCmGbThHFDhm35e54YUknk/k2zyLACq0hGfYXAwogvg5o3oaAQ72GbLMLc+ecepwOVg
Sp1b+JMUWMhGbPBTAyVJEjT6TQojlBc5oUYW1jxbzlOfZdkX9zds9vK9wdVleOy+tSgF0QE2e4NB
3ZNfxAx8iWmVVVQca115FGtplBvWQehbrRNNdkaUAXRasGauCQ9+0Gyiblksh4K/RPu/HnPUM8Uf
ZfKj9LyAWV8zA8Prt2N+tvJFMD+3N5ZmVYAz2ZMGEjVB2lZy9h8LxudvPjiXAP5Ysuve0WvpM0rC
ZxcOmv50/D2TD+g904znZg8PCsFRDONvKw5p9mS8Zt7YSbjP5c/sLEegAgLLJiRxh3oGowAUYBsI
6AJfIaOM1DbSgAUK/fX6IQNnlVm3totb4Lzb/caE2xXfUZJGkD8/WhCm0ot2mG/82HqL/vgbNWR0
gOh3zzDrqTlybXgjcNnXliwYD1ILKND2fGllTS1D65uQ/FV2Q5BgwoRxq2Uhlw02hsdj0US4wnka
MrBe+tiwNUtIYmFOGReCLHiKkiuXEx0FJItlcuxOgAu/Xatmw9HK7VP8YYk9Q/HnGxxY3xRvu54J
43tsjLofTKuVG5SdSyLCM2V6cJccLD4IyDUXVBUbV7DlNjDyqNAq7zOxp0qXCtfAwXJpzptWrajK
h4iGIveUhfD/4JqYZ7RwlLCOONE5uMCqBxBoMWN4Papf1vr533d0J0T550AHHbwd+rlP8OBdcY7W
TLK8jRqS32PcUOdZB6OZLaRd3X3yN3LTWmXupdBVJdfWSBAe9p766VjABfIAe/8NjSZDEK5JopQ2
ikXcNzNIhnfWe1JbdZQLysnGsmu2jhuR4fmnAsjilKexT9A73zRDLBhVNc3kc42hhYmzMDGBYbJY
ixTIklMIKEmlssIt218nz2asOAgSQ6e/aOEQHSe5w8k/8D8a39TxzYiBnVnUHVOZuBQIfpJbgJPx
Qym1mMjbetcGimNvFSfR0MmWKYY2bL9M3yKVSYMNMbw9XVjQvwpBDSJNYpXiq5Sm48rfyDCKAPso
hTRZXkr5syndfHTMRo3UWqlr92xaJ4J70wCPaCVrvUexRF+RTjThpYAR22XTmG7Y97FrZoAX5BQR
MFhWO2pFT6s4r7xaMPpPfv4SnkdLsT4WNq8pDqtHDGTr5UmgaKvvvPBstPvBW+CjdTsoHSsF2BbZ
o2LyB0mMSp0BijfJSF2mf7h0qM1k1zm+sItpPIAYCOaX6Fjhh6D0aMyldfbYIMIOxkVktxATAHgn
somKiQhN0hgnLFOs+6dUUwi6ymoWGFEMcNLJkh4WZiKB++CMBeC1cNJ3/Fgm63Qu1C087z/YKW3X
ittO7KEG5sgmDy3HZf3hFsUWUFHP9hd0XsVmM70MuC474cdDrOfZNQCNsOGyGlPXF9n4xRI9zUDi
ojgWDtqqp1jai9z7XWC2HvOYvKLoqliQSsLGi/9KIdXvd5wAd66d39sWzegntur6522On5l0l+Ni
R+E/Lk8BB7SLCp5EAv+Ze6CebMte96gFxgksEOOeprs10pnhM+LTxrEW/y6GRhUfFthBkdFvkqBq
HPqsD/C0QlmzSa49QnEyBV1TTjorOWpugRsH+Nd/CWcdvii5s/3R4PcQ+e7yQllyeeuJ7J83HOVS
BQaRxL1jq6+fH0B6hVz6GKCouWS6TF+kNOetXsULsUZrx4ORtIu1O2w4KYVlrybbZD3Idhct1ljM
Kydbl0u995KmjB3vTGCCrkxVNwC9WmklSakAg+H3KX97UzKO8mVBHRTJ/gZWs3ENR9mK7DnAFEkX
U9QaWF3VG3usAP7LJn3N4UgH2kZZkZ8UOdyD5sYowuf8tjqCCTwqG9T6YZqSvhouHMkeniZP47TR
vYo9Ao3KVS+30VVbKDLfJ8vlpOYycA2uYbIgY5FNWwruCG9ixtsk3br+AGG5s50EplSRgQVFgFWk
opprtkGtsAV6tYAPnYO2vvfFqJPp/btLyH8omE0b8PMAowrLeD+Znipn5MPa7dfEBBGPFDf8NKLJ
a6qMcPjDrZ82D6gz9FtnQ6RYQJ10BcSy0pY9TP4J04sgVGcVb8+2BUwWs/XXu+w53c0drENOZ1uq
l5QnBEXL1soAH9Cw05eFARDc6h3/zTJahkMRQCpTF9D9A9rBWx6wao87v25ULFx8kgel9TIfeolg
u96Q9R05U9uMRbVJxh0TltKbljRmwmjKOm9VzFakXubEAAIOZPHTIWVtyTYQGi1Vm1KG7UUrX8TR
EKCc6AulsIGbwbmRquIuDeYv4m7L7v2BE1cpCe5XUfh0XzF705Qs40aK3ana04HHc9VUizzzvR1b
2DUz1VfgjnY0jXGaYCtSCT6AIg3f0FGiPW3R2kNF2YZsrtW2XgcKTGpCNxMnCXGY++Vc8fqibPeY
zU+d5JBpITPTWL+dQ6rLR5WpYaAM/Y8UWAjX6fe7awPYbO1I+yCnn/eOoHJTv43VrrO3xPKQYo+k
+kpZfqZP3BB61OYaBRolYo65buKS1lIKK++BCSxX3mJpZRG7r4GTwZp76s96v9XTouOI7Z20sUpw
g5s2PaB9uOinzfEJPe8y1Mgs3nu6A1zhH2D2jxy+6L0RCPHxdTwQ31aM3zRNW/58mgFIlnzEGaT3
FfMzYJx49YPKPXsXY9Q0dILxRrioBFYssy78DMBazG02qgLb3jEM9BUP85+X5MdMnl89Xc2VyASa
GNIv6rvdEwfkXHolVSAHkBtsD5uXMZzgFDYepPYDd1fQc3Ee9eiyI+HpsR8S9r1GSqEaWSNq2VPp
WuDNbaeePIN3pxKyOTwkG99P0Lbs/H9J/hJmqxmYNDJsUVeqDeT//SO84RMQnw3s7hB+4gSlCWtd
Dg0Y1TIiQtUd9443sNQs8VuekDN3QNMDRqTGagrFV+OLGZXD95eNTZ5XFHiHCOAAFoXLQ9kpQ/Qj
gzvdCD7IpQ71GJvInSsGTvLYfzgMvkVe7h1KaJa0mZnYbI8ldFJm0jF3oJzu041HtqffYAwM86Ir
jd1+4+jvIxWSrzUkRNee3wd/4hvZDkHqomevle2m9BwruCDbTGREui4ztD5rbnv0WXI6hMueJrL3
qO8A0Jf9A/B7zm5Guv/0ZGIH0if3eDSzTP1vkoZHK1vhZ50KJjAeO1Q4rz8WBgl+4m/eVkiLpnMd
6laRUYAdkb/Nv6kMVwz8CQP7wxt14czxl03uMsGJvDTKAcaj9XT4bYr8z71E1M5/ww0Z8KcLIYUJ
3KHDc/J1IY7/ILufldYE03schJGn42oInV6mlt0VMnEa7QYzCPfqk5iAUWkAfaKBvQ/FfTWB9ye0
06EB+aTYWdxg9fNm53kss8H3N+pByn903SQVYsf4Tz418toWKYT/p7RwA0PbKvnWkf9dW5NA8NzF
Oprhznfn0b9+Vw1yDVPwyrvwAq/oWzlaAVqnhQTao5g4R6uXYfxzOHr8OVi3JJcAGDh+PM2dF+Gh
pkc4lMxoG9HgwaStlx8GEqAssFnHQyoL7j9pWkLgSM4QqEZKT+jF6IgbeUiym36LvZBxKkMFvmpS
jo3SUBydkPiucKkG4cAVp1oFhvtwyrOOnRbQU06i8mfvLaptsNAhd3Onsb/Cu3Cqal3jg2qZm0GN
MzIyxWDxK3iQvq6mrmpkN0dPTuDqrYUDWQZfZtaxWlY1ZW+kStubcOEv1eYl8kNvqTEZDCoRMGc/
aZaw8lN3HoHGjWCqQ5Yb69APrDKl30o4mlp19m8ds2blZ3u+IGeyDmOonRtEUWpW6Mer/0u68MzX
f+Rm97BZWXCjER/SPqmnCcSD15UIzkYuMTh6t9YMqZPUT7pNQZtwuEmQPXNDkRQ0yEteJc9EEptk
I8dURZNNUgRUD5HJt22CwLNdbjEtSlRlgb1W1yCCIm7wREIktr1Et2ntmjDJoHDV34lRHk4Xv4dW
niabcrO4OrZjX4ieai5pbFrp836zc+3IiRgDsOIW8L7BiWsWMAfub3fheZSsEmGoMXUV00UcZJhf
IMysYn9fL6E9gBYuglHe4MDX+QkY2X0CXRlVeu3DTEx04q7aeRsXW9B2EdQrMSLmZMZywcKasIOy
8sNrY16XEVVrjPDCnSbnXP54cDXh7xQpvyapwYJnKVP78MLqPzegcCXr2wdT/oMgVX6zgwRW+kpL
uaOVOfw3vFdusFpbK6FJ+EsSNdgWChNFdE0zEav374ssHYVmXEBU3WGd3USaw2valSPI/l33fARI
6E1TZxMc1YDR0iPtKfOX8hvqOPFlySqQoi9J2ZHRHwT+67xLXkKTZ+XV4D2l3YI4rS4p2S+UvArI
ZMAsJ0C2YNkjyuNCsiO/6sk/68C4ctdbbGObgvSiDRbLcEIn8CprAFbTrt/8Jjn2IPK8iw9fKv9g
7Vbxvz65kUA2s5PfBmEStIns1+Trph+382tTAsjxCwvwzA1p/znJvqdy/2jXSUnwfrofbast8Fph
rV1/83L/FK01BJ7dWe3WQ0H9VSxNblGY2scECefhTCIPFKbz7iS3PFZmIrwZA6PADAT3cXbmW25e
6vUi/2VMQ0MvzXEqfsGmfpXeNVSfhVjGoZbAaqelfG5eF0IrhLlo3ue/CV6aptjHNVUXU1n1zXqj
5LsLl5E64uh9Di507tGQmAU9oZsDvjZOcVrnTqGYGmP0xuPeWgey5eQBnYAmPPS6ubBsMmdaAc//
rPdi4HUuHDReBpY0/iFWMNUdW3BkOo5aqbWETEmMUHtvFVAPnFR49FStVJmqPxWcC80+G+Y1lqaX
KiLQhx84/R3SHVM5zRA2cY6MkUYRP4MZ1VA5/4tKYEzlb2j7fMOxeSL7wWrCZhhS5inujNnPOIHA
puUSUOKJDSAmrH0zw9mTulyURl2PZKEYaWTLk2v9pJ72NLmqSMjiAJPHoyl0eTskLGT9ZmVeL/cM
GtJulenMS15fkK6YGJyKBxxlXbNJgsOr8swKJeJ6sbIcCxeM+8PTdNPdaUE/7+bRutU2E65+Hf00
wB5xTk/wsVNcU6tSQH0ciHU86LYSV7gOiYl55BwlsFAEcokRPcnf6NtyKKX+1pnzQdgipBhSjzry
baFmp37EkckpYgXtN7cTL4ysEWSzBkqvBantIv9x5h7EAw1GS+NY438dfI2SQiF2f6WVOLHQEHoN
6DkElxADBsbiGwDjOsIB93wUC50f649l2gR/JjagWJwRJz1J7AeGs1Ux5TfiJB4AJ/BfLnJ/Iw1q
OUe7n4PbjjshpvPTBkp+jVOGNWKpasZKM98dsnkwWN+zv8ecN1Dz7rrXdprsiO1oEy34pZ6nVVt4
5iYm95nNXDzLtGE81TFfu7xJR4wAvYnHplJLMbJGCVE0gBZ6LflPP6o2jgh6MZRizRoziZUDbihX
v8o/SGZQgvxiXzjxM3Bvxn3y8lyS9YDDgwvJ/VLNeTz1YqGYrmYUKLsWCZ6/pI6NwKE0MVVHJUBx
y4sccpXq5kOT/znYUlxBJwg75Y3cDNx/SjZfDyFclIvrP+r+H01NygBWAHD8bVf0D4mWLyAbyAxP
Sb68fpIhhTImed1p9OcQAVOCsIX16XmffKe1FaUmLnOpJ7sm/TVURla8P2JIhWDBS7HuvFMJOmBw
VSazIspIwsls/Ko0dBwQdUbE/xvGM11HsgHP/pZnAZX/fw75Pg6Gh9TxsVyDAFraPkj1a9mGtHrF
IYvmf2PG4ONyXKyDqJX9BDzSYqb6KiiPLdP3Rlv2Wuna2kGod30YBbMYv7le0s/DdaJwnXfgpd6E
gCFtq3yugiJDVRNnHGxGxxUo003ieas5qWGUWhhRgubFTGQcS15HZxx4SSdIbS9Mw1nXJGZncJSJ
I9NmHO1wJtC2rE8VRR9SnAy43PcTAv28RDVyDAhm462BHPxc9V11KDuE0XOoD6CHI0XAIKvj3tRN
an0IruiwCzblh3V5ThBor6NFSoIV+PnZZp2IEI19qaSnBMajXAoowMwunYkWgM64gI04GupIe77P
Dygu7gdNm6gSBOR6LkGMKR82pwFNiX4kcR8oAHv7KmrbeZkNAZ5ga80KsG4UIFM4pLYLbfA4G1ho
jzpQ3yEGl90DizHZXlN5gxvdeqa02qdOpnqKz7a9TQhc59awAB3fHxAfyzeYDOn+IofAja1/suIg
S9u52P932q1P9qegsyNGefbEPUltln9sXPWXApBb4ZlVgW54DMFEoyZ6HI8u+vVe2OfUAicqLED6
HF9BSfPm3ZBJ/CdWxJVZ2RnzSuxD16iC5desWIacynvHH8v0GsAFoixM3qQNqwXCBe3BTPfIiI9I
64rj5EUiuZoWxzcjku9yvMnDfMc4kQJhO+bJK5rRg59thQbwui9OzYGTwu/4DCl7itFYRIZYNPqH
rL82NNOOTNX7jWaHD7Rjgmwuy9WM8oBZRqBZLWJeK2tGwpdwTprbjHphQbNcnw9zqV0bUf/6dl42
y5nD9y/FBrJgq37A8y+QRLB68rijkaR4Jdjv0tOISU0PU7IZda55N/uGGvcg2brCYifu7qz9Ud7I
Hnrsw9wTNJG6SlGz+COAVV1BiqCwfioUb18+lWIuwL3+PjZQ+GbLeYVZQIuEzM9TpDIZTTqcJHaq
SaS+sK3ufiU6ccJJ+Ke6pbazUinyL1TfyCLfnxBpb47BS6SatGf6y1t00m1e1F5G/6dmse8v7hiy
EVKTHa7h+hfTY5uHaYM8sVGytpVirGnvs480j4ZXNo6XsS65N1VZMqPBHXpfVSyngnweCfG+k8Su
MM8Pb2Ix+y9DhAA5hyqsGSyosLfK5SJ2zlyknU5lsHkiKa5ggT4k1xYOHzk4dHTooWNRr6nx26S7
ufcekjknv6X43mcT84rXfHrgu8a2mQ+Gl/Vsj4NRHn3BsSOqTYrP2qi8sN2WKoaQyCWq3z1sQYtc
rUYrkg/WwBk8BHgi2q7Y2sbk7LG+1oKi1zvt1zTL7qvkizDVGL0LlQsHqvjfMrXn4bLg4DCdvEOQ
Q2vcoMFQw4LvxAyamvhP7TSjlDftkOitcYGibJL9aYptyjFs7d9ZsG037nA1ndNkcz3kU9BMHg37
AhSXjsN8B0G5Kvw0EjTrBEDgGKBRQmpy2Tfxgc4iJmR3Akls+skSl4R65ScoKjg8ALY9ZCzdGdZn
4EMshWgxTeYABHFAAol4vS77TjykN6F/EFitgnymiJvW+iKxRwqsVsipXn1XJqGmwvwP81pk7w+I
4FFDyoMDHPHSAfmayBaQixzsCuwh2Rf7g/mLWfAQewFxyJ7/FxDGsNFhm2SuJ4yjYaJdnZo84me5
nxcOQP7oXMeabV4nC0it4WTDrtWh5mXxE0z1CQMGWRHMTRKwjQipPXQ1zAkgPNsHnGINIsRZga92
6TQgXl9ksQuqEb6UoHg3+/yQqyrh+Tq0y6hLt1aZ1aW4xz/WBfFO6xtNQNpfssI1A3O8SGDmPG6C
lk6vvLoY+puICbr9cegUPuz3ayEqHg59IlH3YTdMTQN83wNF+GfU31RaB/nyTu3ZbD9GjrVa5taN
9gEm1hOPZWDT6DEOzykYRVVcxBEwk240aBv4dwVQLqD7qVtOY+uoUGSlvFTolz3xP0ZjD6hqQ8bn
sgbqv+bzDZQfZiMJHhGUTr/YHqwQbOMUFF2Gvsnz6ihrYfgz+1RiekuwwlBA8diaNwqlcwYkUxNS
MkYOZjflvkWMy+ZIqyOyP9d2y3lKphgDju50SY+B6eOeGXlZOBRrY49TTofvZ75b0Fm41Z9VlvyR
S6FT/fqlX44+huJwXbXR8BAIEczBlVdFcZoMjSAjOKJn7mfsnWRp9u1BC+cLRZ8c/4ThFaK46TT0
iGG0eQKZqe1cxSv3XUVJ99PLXOEncB9ACyta0y/bzvlqRxvojWFz1c4PcTmwhPjMw9b3ohTjkHM6
2GjanVYd+3GRCM3WuNRJFFzxp8p1iUwjej7B88i+7oXkhy7rOqBpGxV/fJti4BmZk/1kUjBShvoA
am0llnRjs53s3jh9OdwOZEHYqpdYoPma0fcPMplpsBTciiN9WtTdQrWBKcxU8jNv9xsVM0YE5XOx
V21pk6CQ/dbGbdzVbpfhpY9t8tDiOy17dDFu2m4WierURplpfNU/o/+1Ho3PmB9YfHt/fwfx0txx
7DPF7DSOv0mq5IqXz1QzQrxbNsPIAB7FaAvS4bLqdSFvv9MO5evUmhe3N6oca7UIhZsG6hhwyrbs
uiC16upfIyvnRd28IQLokbxwrloB/YWsKa8x3HjFxYosWsVawqthjVAbwOjF2ZbG3+Ll85EIgNvd
wY0XBhZhPbhlZ4oL2H7tUvJ9CukOnd2y3oaWzbbEUDTAi7aNtYk2ietr8lA2O+R4zgpjX750+Ong
wRem7hBdJtwogD9CrVQrHw40UR6pN+JymPNnVmXF3cXz41lFRe/77AG/OtOdaUVDIZmtgt4XJeHr
1JqR4+/eqoXcrG5v83TRZ04vJrXavrJRdMY2Kh7s16Xly7e+BK7qS2VZM3qtBoMXr3ZhXSPm2YM0
2xfralN9IN5dGKtq20TFjePyYNhypmFzJXFF6lqKCeerQZHBIiWcw1vd4GTDhpE5VWwk9UWeqfEZ
ysy/acxuMksCIrTNjh6HUghKvw0JnsFJQSqrplvhP7TKdI5DXduJFoGQ63aSE9yP/KFipTSG2cti
0ie9Jhxtq/NS76PGqfTv2gizikHdnEe40qSyYVGYk585YHqPeJu266Exj5x+efh/CZhNHd9UMg65
FY+ElXK3E8ljivDG84BwrWz4kCI9ztpRQUIhymvdBf6IhQS0i9kbUjg1LKwqKbh8rQyxV1WsHe03
BZ2L94AbP3nJB9hZf+1NZKpNvqRNt4EFyvO06XFZ4x1N7/DAYpwn/pf/ZPIMGd9KUy6Wif6YwEoD
qJuvyHbqllhbVLziPa+VoHzP7RR+KN2CZd1cNbWuDw5Lbs9F3JLzS/pXdPMSDAc3YdgGV98vA5U1
RJy3HiK6eoIybmlj7IgPr1GbtD/SNHRdwqwKjt0m4kK5QZQbNMxd2i0L+V8nA7lGNaLEtXu2jVnO
ZEJRCfUsRpDZOoDa3ZBzNAyffbJdba1RrnvBanjC1TUY1A7GzBIhJPotRCE2g3y/t6b1GwxwIiHt
dLBNKHrV/2H9cukJRJY8JTcpalMfEGQYKttBUufNIIy0ceGAxPYVjCq6Yl2sMY7rvuHOZ33bwsUU
WkXJuLP5I4j8O9cDE1CxJ5jctaZEQrZF2SkGWb7Sk3kzNxYXAwHtamv11kyoVFz3foKDzTOBFVwW
ZmY8xaFArJs2j6eVs60BLURjYbnx0t6CQ8DI6af7kDyuQqkb/+7w0XM9vj4UOb9aRoqEnBgKCI+W
Jp9pp7eilitR0xQfHttR32yT+2pRWNurgO+eUkXhnhrZ0bNC9nK4CeZwMnIKLLRqg3mofs1oyK+1
BZQztFUJOlFazstES0liskwvlfrpyxHHfu8YT7P8oOOVk5ds0qYr3epE747iJC5CgbNyphRNGS7a
bYl1IU1rzwFjj6Ge0EtAnNvfzAMiKzFmrxtZoBPFm9Xy17tUs9KUHLQ6815MEAaLSTDeUa9a8RkI
usZQxfvNW+RmirPkgOzF81rswZE1aXY6Sum6yIiVpgAYIavgieAK34zr2lDoLEzu6kC+MBx6Ly7h
weArNdQsUiIvgllvganl0lI82hod0JZ7oMzCiJNbFal2JQ7rtW6o2EjSrKq4VW4DSa5914vOSC2S
2P5zZEmku8MZIt+3XyxuJBVoUqRJ2DPg0SAve5HMfoBIcmBvtFLKpNBU+mnidyanM3+E+elJlmBl
cBnIUy7brsSUIJxpIz/BTEWFEkAPmZZh9NKTyrrwMvdXrp1BV1CX9G7u728Qi6Ao7OV4n6nASaKW
Lx6bOxslJONUjyLZ994+D/zK9SwSIX6ouau/yDb/+/xNoPg3qhVTL4Mh1Cq87vaC9USGhZWCqaTJ
toAaGUSkOqFeWTA2lTp8X31SxgqjYsijOXhlPqEypBy7sCoSwMlzK/C5jn9kZNIjNXv0XbA/ERnK
pcV8+t3op3ERMdweKXojRTbTu2NVFrVaNDjsw0sdgCqdYQIe+CMyjlMyJddCKadmJGC4Ty2GXNVV
NtIpUyoOJxrGfoWfmBPUlUzdNoIBG/v4EKCoXXXWofDZwZWcaRvaFQAtp4ph2KbJhzSBHR+i6Z5T
R6zVQ4gO4egMFcgeqw1vaXZbeMdSmA0AlZRMJCJy/X+WFGUyClHbba8Fy+vZFGHqT8Ua4YVqZbd6
3XeyUGbJytwImk4yJZ6shGNMkm97YIyvUzyR+5KcFztAKe5cdFJo1Oc6ypYhRw82ERk+u4GrjnS9
BQ6gb8JsNqQW2rKTPEeVbln7sR1fLuNADDD1XfPuLHEHi6dpobQTaP+cCh1Fw+fvTxNa701IR4c/
osgQ5/ijpqPaHUH1zEIUOZXj1aeENkluxfRcn/7WwefKXbUzZrfugsQ2n72CJUZqa36+vgs/8iiz
pBHNTlmh3kSvmmV6YQNiyW6aaZyiQR5hYK9EuLEqBqtiPeU5oHseHZsmXZPRNdmv7CJjCQ471nUv
47NJvKj1/ZfkJxeBg+HpWPEgz979EqtgeZQkiPQcvL1KyX1hxvSjALkdr0u9PB17BwFK+iRW9Ja5
I3qkb1/d6W4Y642KgiZ1swN73UH+NhtBXWvnvRHa9rLMWSh7mOvjErZXT+5M97Jki233/Uyjssc9
y9Sc7Axf92HwOmfduKnMSgkF0eJlClhKhaSVQghptZL+vvM0yFk2vrVx3YfKnKPTT8XexGGkMvkb
mT93PXKs2r+TjMQT5rSOv76PDWwvR9rXMxE7mskdV4R5n+hJOY/FoiR1RJP8SgTHJKz7mAp8ClwI
wpvMNSVfEmxGJLnYO+7RXtoeqEy4h8tuKUWy6vrmlyjW9h1zXEnp2BBFAuYt27QHoF1EVYx5MLtb
LocRHX98OiMzCmon6B718xby6cGlvPezmU/zjrEWWM4dJ0Pj6vWOYMH3T7XaQ9w0Ogr82apDX4+J
qwaXnNkjWHz+SWIHU+L/Q0XzmCbJH4J1+yXxZeIPJyQz+MqSeGnlx0mo65A4HTkSKQFx/sTayISI
vMXImXeGmcyvlWMue2Gn3kKvvPBI+9xiR4kha9meHSseu7ehOwKTzjGZ0NK2AQx5LlEEQbOR0FWn
TBKpSWlS+bod5se+4Iu+r77mNB83iR8q+0Zb7+bkv2ZlACl/f2m3NSMQkqOzg+h4GvSJ+71KaL/7
InuuHK3O+aaD3NaYs7OKnlqlN+S7cXyqTMLOWj5lktPYzS0LpFHqCjwO5A0kwo68XMcowXaa2JDU
xjLdtXMmasu3JOjqywp+28XmOmAycQ4PAokbPMAUMmg3I43T2JXEFkHtgzq+ewZmsH4dDBl88LAE
qy+R11jvFHoqME1f0Ynj/z8gCnq3s4vEOZhuqI95S/ePpKjtjjAXGURZtsc2bofKrPRixTmh5EFu
1aoa3Ee6Q+oll0AsLsrTznRePBtQRTqTXIgILySAD+Ndfw3OnCEZMSATLKP7Re+N6rUARJhk476w
5Ev9dHLS/pXdUyHVM8qmpA0suTaD0pldu5QPj/b0FVmIFQz/6o2VOIWiutglUoFvMynlqz0gINPJ
QotdbHEalbTluuZN5LWrWZl5hKZOrc5ijKPFQ4FDHTOBOQBf7M0F8okXw3yqlbgLeqyodmeq4Cbn
Hc60zTGnOitK8HEFOBQpvoOsj+6bGfj2waFTt9K32Hpzf1bZkaqgCFD0TwqQQ+Ie/MPBhs4WPKSa
pyFSxTLDnfaOKkAX6+g6VhtBY/TZNECHXwbJfMFK7iXr+RNbRpLrpW9Xp4VBt/CCQECWgtb4lM2r
ZONYpiZeAxj65ka19S55IxUS3nV0NvzbXXo4vucZxdah+rvUdK49YBzbQxety5mbr6N0YycGxQ0I
xzFrdskxh2JreMuMDU0zGfsXc6ThQS8N/FMt1xVJ/7U8B5ur/tewL6TUumT0I1hMrYTDK79Ta1/f
EKyB8vQqP0JJpdmXDCUgT6MfkpY3Uipbk5MJZ9vTrO8oNGd/TtXJGixYm2CCZV5hVRkJfEhsGpO8
MIAVlqqVGsCqAr6mKgIMvPAERJCVi2tBJJwcgblOFFfzcyHiTpO6h8K2Fcxc9Wra02cfD0K2qH2N
uLp3iYRR3KPfwYc/IF43sAk5qzDdIrVerBQMdZTKqpUEJuIYZEQXIdIIFhLR4fpgP8tlaaEuk7Gh
hdnxw7Aq7bKoCIjcXe7kXGb4oLkDHluDFoJ7n35iofmImQcvL4lh9lLP+T5rgFQ5Jp/OOJYQglOq
3fo2rvhiMCwrUrbK+nGG3MW3cNW/vtSMdExkeZVUby1nPqkt2ZXmo2pHKnMK35q72pYuShOnopeN
F64sk+XJxBRkTYhES3Ij7/7+Kke0Na0IhOu4yu2n/bdaXTi70gpYc0FEsypO3u2k69CyB0e8lY4l
hRQZSbNFjwB/78ZZsCqkGxI/FMfP7UncmQb/mdaVH0dhJXSNwYWitSWaRhn6oUXZcA/nNxsFkoH+
Frl0+WsSEsp6p74I6Wfvl1xa/xuqMRf1EPoXKSbLexinQjsdYCYzG/uWAGTc33YKjCe7dBSxTTjs
TNt9X3oX8eueaBvzEKdmAni8v9+BskzOOXhGV0AyBlNJF2Q+wBPPISiYB/mEUP34SqqMQGnHPPkh
ucvUMQsu1qAd56QTq1aWabpptpK1G2J753jNd/BxuTXCH/TJY0DsroEgESQnwIPTdfuSYbOMtoLP
yLiqdsIwSsBbsLrV1Q5GvGSqIeamfbU1+0G/njXzg5HGuyP2rcok7KL5sMxZnl6CQFUVxU9bECHt
NleiywkGrjcv4Vd4JjMjM7OB0yt61d+n3va0lRac0ZLaM/TDfbo20mmlCt7gFbWePOQoh1jTvBeQ
GyuWx0NimOUBCqgQwyiskGfTJaObRIxt+KFzwhVGpeYGF8Wlveu4PHPfTcOGwNBLl1Q5xG2t9pVp
FFkqVIGGar0ysV4/eIFDhqUjPkgsQbIDDFqDExLwd9jKsbKKCyB7hUROBzPuUri6fTK61zdEplG5
6rRdcyzVF5bSmcmNJwBX3H7T+sy1EWmnFtQW1hfbZMlQmwr2xFVJo1LPYAyDuKgrh3Y2hIUAJt4H
XcaDz4LFJLOZKWNYbf/k7W+VwncJEJLNoNgtdOq9OyIz/DyIJ1mJhv7AATz9MynfkJjB5vcSW7cb
eH8h7ErULM8aCkQco/wHZWZXIyQbkB1nhuGGfmaCQl5CYiDftgO7aP02+b4KPRIwkBALnDTE/16F
QrVr8okP4PppSewuswi3RC+jX8bd3iDQL3GP2VV9vJIjcdL/+vJkgS/jgWSHMJjdNXp67240Ob+C
xCiQ8rsfVnqVrQRbKrdy8aD/Bq/xYF21othWO0+1tUR9M+s3TjFlTFJ3nQH5KvYQEx3hQrstIvIT
H8oru0KFD9Do8gozAoxCGA2Q0qGApbT3APCClaRh13cCepAXxfv/wSBFGjX/cDE/ZetKIwGNIBkq
/lCth6NBkL6pZ/gBs5j60kB6P1Cef/DfZMeNSbhVORmtW4/AZOviy735q5FL8nSiL4qzGa77glSv
g6SuJ+vs3RnyLRjD2+Ew/ha04APM/i0JyQo6/HIziiQiwvSqf6z3dypR41X9ztICG9UdMrdNCFR4
Gxlr+ZKtHxGx4uquFyvV+ewIIOUdbVHvoZC5s/scBU0zFPlPRltDKy9w1chNaXT1zJ9LHmJttsia
t2qM65X1sAq4dMuUUN73ueOSVs5QrO6Y4p9E3xHk0a+hhRsi+O2PfWfietrl4V5B85U2lOvDwo/m
ec7InSKKIrH97my7P6qUujREMrdqiSJfXr6Dttf/osYYozLbFDKkMd0VxuwCANO3IHOLN4uJmhk4
SY06df8JuCSMrGdCsi2EJ+qVLCznc8cvqt+NGnmx6VmwIQicMxzkjrpM93T51/xHTuB/+qU0O7hP
b7DlmwVTlsnQ2Bg8PzzrMuB+06fKysQOK+y1/1ChYx6zmG0MafxmIwB2OoeH418B466S2sGHD6xI
WTKvU3KCU+XLZ6L8KtcuDSgLKmZWj0QexfzJdpZQK1nnwGHD9epGxUXLKEjVPBwoOkjmJhO3i3zT
djFLsHiVTzKZAlgTlXOyhrbSpBByL7z2In7Pa0MHrSBbwvKgyXjdsXq1koVrnGzh7iQlmkbklHjW
c4wqqGVWPjJi2++HqcwY+M0SXEP5AK3At/xGqV2DP4Lc9I3T3+oK9FJgwD4RA05otCpfXrbDC5z0
GAkoYjcIDcwSjd5xw/zXbDHqtpIb8vW/1wJjKwUhSmPcl3LpcoVu4tbaxEEQGFL9N57qN4jVYusp
nfpByz1TAkg1EE0tDMilaePyolU4XT+CTtgWDqKvMuDYWHwafftNGtLujyTO1kVepom6+9osT73l
eOmO+pX7NvlASFPX/zke72VvbkGMhEliDHl43aCjEMoiy8k6QlixwDvcUYkQk0RDEKeAUwfoKaYD
z8EKsYxLI7S6qK9wt864EMo5mEdiZUdO4PSe/sLg8m7dgFlVvPZUmLGfi0mYV88jhYz0vuBGlB2z
H4jbNx108Y5HMXxDDVZGiPQT5+99GycPv1SHPR+PYRlndjv4Rn57kdi7MZx86rASX81NLDic0B52
fd8pvSXblySPVeXf835mZ7JHrRAptjXNadjrquyO1yV9lqFSVUJ/M3o8q9WYB1WoyMNwFKlGCvuS
Mk2CwVrTqRB9b4f8MOalSlRZObqnr/GDcdfPtAZth6XzQM9VcEqEEBjF8MtO2bhCfw+ZWqPuCoBI
LgUjqINPuWMydrj+Fof+wJMrITjXBcDe+ydXFICKMM5Ms3F73wpotgX3vZd829/on5zCtjzb1Y/D
C7zZ5UYv9AzPydZbaxRDWTb8hv7OCiZ+dkGSBXCJ78TA+vFKPosmjOW9NcMz1O7sAV96xfR/pUnI
fHOO3TzVZ99vaY2R3lUd/jEZs4Lhs9YgN3SH3sefH1GurSEcMaFGIc1CeDQ2Efxaam+6XglbJa6h
MeRHBmEkZiPBa69nmDaglxmjEpXBMznZpxMRmnGT3D7C+hG4Lq4Y/x3AqmiMRRbQP0hqPkvTgyuj
Jxswl4IyZhmZqdnNfKCnpa+rVKzZ+gONgLBOQA+V03l5lOeKM4d3cm5dIl1GnF3br5t/O4DNBrep
P6FO5udtWKnddZOc2i80CKmJFpFly9hcpAoN9ZDRj5rgK0N3bpT9+Uans1fqmiIYXg12hrqTtS9T
IYByOAb9KK1wlBQY6PQY647YgLQ7du877ClbmR6ClxeGQn7yEZF6kw1Z900V0E4lhA9+cyGDXaBG
Ysa3R25yIH1scYKq92JtnqwIe2+x2IWI5JFN1G7TyW53iHDXo6lP59iY6lzWS12Zy5kvn3Ji8Cjq
dsYFXBkFq0y4pG72O5OIFYTHQIKKqo4z97nGr3o4OCUyPBZt0izIGuq80g8/LBaLh6I87sltf1Dl
J5I1CZ08dZARNJvZH1sLO8XkI1ITCnMD2lcpyTs9WO0jm+qBKSwvfDG4AwgxYk2wvMjSabPY1q20
W3ZLOxxzc4lIp2XjBx4FtO6785xFLxz2Ae+FELecLHpuP8vfKfBUpT7nFLi8QptjAZD5fckmRZ/2
FjtsA9UkQC6w1csWcqpJAVn96tzpru9iix24lKmbyaiNMTiZFsfw44K1l4PcE+PE38tJfmprBBoV
6wEBO+iH2HX42n0zFBlzIUzKErNsQQINro3v8QkT3PGQ9IL+psAWKNKtA7qu5HHjD0gNH2Ptu8Og
lLFTCoc6MtgC1uk3ptzzWlNuSkJNtaWX+o9FGHHNUYxHqLwOj6lTThCnJ+jcBlx9m+UfyyVlYBHK
jz62c1Lfuq3xOPQwJPM798HkLbo5A8m5sx1GkwWLAVSaxemB+YQ5cHqoJpx/wOQ4HCGbmKySSJB3
E+RMeM/hFwbLLZB621NtuNR1FlSjyH/4DrBRd2VwlRZ7sLljTK6MxrKCM2sSnl+afCfGWht4Ewdc
OPET4HtYSaGdyL5+OtPXq0A8ntchW2zocFvWLR9Zj3Ss75fsfDFNNAHG5kT9lv3T1lSp5QtPnfpr
mQUneLG1R8rL+Gb/6WNcO4HHagEKHt1fKs/DB98K0vTiHi6HvWDTyj+sumn3bCnBTl200iHf5PMM
aaYFujmEbgOxPjMLyN014mv3R23mk/Pj3Ow+2epbPIEMo20yQIbsREaetpJNi78Xh+uJt42+fuxa
iwwSk1YsevWv1alqK2WtHJhLj4YOk0lG4wGc+5vHCjDnjKH0hqvtPtb+CO5u9Oy1bX9dUFoMEoR3
ZAtM+0TEqO2d1OXsCwBLf2WJF/riDQSM9VCBhUI3SRZ2LEYwyhjFJk39j7mtu1sZ5dBWKRxf0MgK
/v8cUqeQLKCCPSRAPOqS0kbF/L6/aqwHpprJGRGhevvXtT1gsmhobMgJHmOfV0QRPxNwLINwIB5D
MGuB9kCyj2K96DugYUSZ0b5sb+A4+4SQKF4Dx3BYzHsFc7PiONLcVQUIZrZx4R/2K7BGC8Iovo76
8aqOPZMaDNR2HguPZzMvvB4r0+QXs7k73cC+VLT3otZ09CmsK2Fz92eyWv/3u+5POrB5Uxml9O5s
3/jjjDaqKrlDt5akbslBfcVoSQVDHAXdC1n7beVc1At7OMiW5OAYSLHVFAtYZrK348EpTFGuCOM/
PC+/Q5jDD4Tv7mTtHWrx5+KOdOIVLSXQCgSbb3ujogs0iyY4JAZr6AAyFhc6QBS5COtxaPBwnTW2
TgFcpOOUD/hkRicGnGTcFms2Fx6yfivEDFtYm8/4myrcwRj25guwSWTDYvLXEIXMjL6RncKc2PUJ
G3NEZBheHQuRkmXqWRaPeXC265u+qQg9tYE1L06Eo5u1ZjPnm5DiwDpLEfalTR0SxfIvztaCFqFF
GNWj9wKAJEwUbHGZq4Fxuj/qL8gOXnUJ+O7tJ1SKRtXK4N+n4dQgf+32XxW7e7jBVdzHdGb4k7qa
VF9NHUHrRl8kQ8aZCttM4WAINVGt/9oj0Zns3e4Hn1PpOvicXLazlAC4JX9Pum9tSCuhr+SfUtih
XI8HPetVJ224ZozIZUOMdejKPJz8HLob39GQvusGBHtC2JF11l4a8/4XJ5LfDvKt36Er1ggz0cD0
E5A/8XPKO89qZNwizhkxLe+BeVY4GTWVAkd+TcMZxmUNG/5RnJiCDYS7pB4gScz5V/BU/ILcG8bp
0+DRSY72Jguhv3ZLkJOBtDTXWcsGs9i0mWV7pc//yoQ/W1fVuv5rwZWmcYtkSWOFSDm8QTQlq9Id
u4mdufMVHvAb5/2L35V65DmA7WkZX0gzBH637cxfc9e3YqpInJR609yL2o05K2EbjWvrsEd5pe95
IM2izhBWIi9NKmDa+CBhZpmFV0zC1B1EE6kz/nISEHniSRnVMMYqn06O3q63vpC4SUo0b9eDFQvZ
4t3RfsIehY1ikCnRezmZ3iUXsOPa/Vfkh6ueCpccSk6GjJpOrVNg0kFQ/XPbARk5OJ/S0SHKskBj
hYRbmlrxppmPOYRjNLYWRAQOn4L+zNywvmHZA/Tp/MGmRSvIu6rJkopvkDbyn61SX65i6miZnfkn
mVBZ4TC9WJkl87Xo8CIgLM9xNq0YVfjysvXy9awc821BkPtE/NzXwEI51mUZEkUbnZzXWgslSExW
jMQB+vRq0sC3/OoiZzDeTddTYL0bFiQh0Kct9BHq86yy9EVQM5ZGC7fboHhqRaJak950fKn6TtuP
70BgH9HD8Rl2zRft2qYzwmGKwom7a5MWFjku1G3135H6S1W1Q4YtRwxWVJjzc8Eh8Z3JKf0U4i9A
lr1XYG6hLHaxYjtKUMSfn7ZG31oaZv7Pm0wReW8KCw7KffVTTQy+EPOrd/cbUhHfusDp5Cxn4jwv
i35D9g3m/73i1DlYTY2XIhBr41sxfi2nDd1zzaY+G0H9wC80aiaT4mzb2v9lP2rhMFHffELYb2G/
A9x+xmgpmGOAEK0UYPY+sQBYC/Z/92HLanz2YKdXgaJjTSdWt5iSnf6QI3NoAtrs68GPdYSbFc+l
dTVKavzw91IeQtYU2IyJbckG/ilE/pWK+2QGqqy/ggM813aMl1lB7qRupcw1KC2droNKP4/YbdPT
wlcX+nRJZjugviJcfScCW890ZVQD7VmaPvKdjDqb8zTqks9NXb/dY0yf892WXTf5hN87gYzBMeSw
S1rsvpqSp2p3+opnuz6GQ2RVHH+a7KkzL1Q5+lKz0YxBO6BRFdLYk1Q1HdUxTDsPmjYNTEbjcEpG
yjE8Th4WSR1YuFbkcpChJSZCaAblTlYwskJKFB5fl6oGiytQ5QD0k8X1tt3f6pCJ+N2Tsur5yUtl
QnCL6VolRFnfFy7GQQpouXlQee73/jyB6Q7wKp4kDuzto9tcTTSSl3prEZ0ax5gtgDjYieej5IcI
ET+hyQXuXre43/Z+9Tzy928T3xiKtK50l+sSG8BwZtDD2VSp4jXqk7VXozvc8TxTcjFau0z2m0iW
fL5KaIgrBJShfNgMr1ll3CfzWNBaj/vaGQd7JJpFtKSKfaw4v50Np218WzRwxlg7QpahPR4NGlMf
JWywhen/2uIe7q8uFlRlV1MjOQs2E57SmT6Nd1u8Uw+y6vif7/DCaPq2FIQ7fvlrZvhIRJYx/Utr
89uQrhugkkAEx3ePzImaVg52TxpGzLeMVGmQQfJQ/rAcDuFt5/6LRUSW9YRXyNJ1YRuZfceTScPY
odX08SArVYYmf2Zf1URCyy6wi5ChDAGS6D9xWBv1ULkcBaQpXr8F6fObywBhBEDQ38zzf6gHO9g+
grp02VA2Iq+KJd6maTWPOCzKW4vqv3Grit3HRzbbHAKTQftLrEiIPQhcDK9nsBgyfOpW6kOrOcUO
ItQwhz/KSzOq1FAMByeSegpS7ixh8DymMrNMWjO/lZjd5p6tf/RJ2WjZulNvBfhTWtkTITFjWohe
Zw9V8hKr5GFZX6lVkzjWhKmlqIaMwHJjIyOhYts2CSA25IO7EaGoxZsIH5M8DOh7N9QY2vC1b0yb
tqH+wE0N+YQtxmSTtINrRhqyX8hQxvsLifklmfXWavybCcqY4urWT1sLfzpImyfjzfn8MwW91oao
ucETQku4s+BizHqfswwKV5V7CaAfG5Wg6C2BM/AasPAnFq1GeyzkVAh6Ps1u+iP3hgmmw9jXO6tF
9sn/M97nCkf2N1RC5Eu6jFZo3sJekYS+4+7c1U1kp5mMpBcW78nR12HMMToVakHVaIbVyDPsTcET
XJGJiFpDrBmjMT04vjJL821I+WYn0255Lc7otJC7hEFZtN+9UfeItvZJojJM44gV6ZE0Vu8I/u95
waseoUfzUl7+k1dRkHCYq7PpZSzXbejILEyd/TXqd7MOWtAGGv7YNd1Mivnits9aa8GtuUzNS4Mm
OGIjMIhGaLIr//x7H38HPUqJ4T1bkdSJy6K0cVsHyGFxPXDVqeWJ9nYLGR9piB6mDpSx6CuJGIMu
FmN190RWNeNdZ5y33Yy7f3ZMDjvps1iyQqFkZFcOKT9zzVQ/PQuScO5s9wnsLw5rZt+5/n32e/+i
P7R4MRCB8uXaBT5NSshwR5mU6tBDBF6MjObGGFckNAADmepbVbwLJhZS2sYSit1lcKKaiUFoSUtu
S9n2j7C154B/B2a20qwOROfgHNNuKsQAxi2+QSYsGz7xzrGPtnOaHcNmQLTGAbs3h9sZGvuqcZuM
+uw2MZUkKGDAHR/Ig9p1fOhKTTfXp2nUPHzyNtcSuhjuMgGh0on3lpZpBpHovkqKnnAnch+pKx8q
VWDemMIuEz3mMvRPoWCpg38M5ZVetDNiEGlI+CPV813lz/HS0HsPOStdLFnDGZDrpFKoTs7Nimw2
zE7tgTZVbjbme4SO7UQYL5mtufuj/AaXrMATkPTeOIzUIuvfugia7K8jfwTHXs9NHiqa2kpETEgP
4t/Yp1PPFKXkgYvSe2rbN4bORhb+2x7iyFDnlLiYXc4b6bbGbrpob/vbJNNNBLht1U1A+dkCvY9c
aTssVj34MCnss9kFsIM5fJqyp2TnlwMJT6WEsXjMVErif2cNZKEsjbgkPbwQTuxamBc0fMIRo3Ii
ihqwISPjOfiPGjFxejz45BZl0nYVBacN/RBSmvPFtW+Fq54D3rjyZryC16Be2EUjHJYTdDhk2Ozl
p5Rt1bb+lycIQyOUuR/ySo7OZNZlYo5YJAybXFJpnVA97s7i8IqzgaIzqLrm1DG0rbA4pUZlCCtC
pe9U1Q/yu90RVNTf14UogMAioHIJ4yRND7As7VztQ9fPrrD0xBRBH6PzXajBDQw+JTgRCCrlGqpz
k8w8SMtewNcNWRa0R/dIikvtBX5a72NnCPAxYB5meDqaH5swIq9oB7HVNYkgTJQHCgtV61Gt/frm
qidz5dpI1tbXTzCHotexkhMSOVig2YL436daQZY3KWkm/mZLVvVi7WEXlWfc1UwR+1VKsvCIPoX4
GljHYF8Ko5+Y9D4nYowExBUZcTFeMw5G8nDXERoDy0mhzDJcZXO96eIwtT7cLyaPGwWEw6F7SSPL
h4L6YpOzCl7eGIby8odaf4wLTE9JCRxat3nlYzNHKU5E6VfyiqXKthzZ/LvfwZ099MHtjRtZEWdx
dnyfZnHNwLvOhswINZnyNNbzo/BiSQ2E0x/o8QypbLucUrcggngfaLigZU1NBIKuBJc+NmC7n1Tt
8w61gMqERY1rhZVk9mBQNxAvVGrpTmi7+reTSg4y5QaUeBxnbTJGxxpxT8f5WJyW84WjniHsm6xT
GAocvZqZwVoSF1ivfP9/g8R1pJEKlw1pvxpZbNM8a0SQ0MyvgrHBb9PWMRdJRbk5HkNvp9DB+Tuw
6PHxo+sxSmFqleuMLlQLpV6sFYZYnrTpK+Sb7+u04XGZXImh5A/4pH3lvFQPHnBpsdLF+zGdgrNM
MfrJ7Rlw4YWLFnwCrJtf3vDjSAq8fL2dJ5hjcjGLaljwVcCpCAWTKpr4Bf6vqFZZRWVkjFv/O9S3
l7ybpEhzNH+ve9e3oNIMMxV2+73Ch+aTqHWebyreunpTLZ9lATrum2ZmCMMYqNedRpfwA4T9FDlE
Xk/MckEB9Jff3gtjSwA8l6WZowj+5OS6KkADV+nUZDpIFLt3itS0chDtsP4c6+biCCeghWTuFBIJ
QQ/9SxgIeDoOLS0RVttiEC6IhNgKxJOXqE/4uLHNOxI33iuMj7idBrX1Pcyu7xnsA4XX8su8EeUo
1DNyBRMl1HFldyyRFJsatx1A+RB5/W7UBM7j+JG4jCS0hXMvjEJe96hQWI0P8cgL68uXrJQqOy6I
m7zlplsYhPGgLchQ+iSQgegLDW0BsAAlZeOqNGvEUEKmVc/OdplvKzwdii98r0pWTEKD0dfxrBUN
RU3vqKVXMI77pQyJapz23hRBhp+I117HJ0S6aAamlpoaJ/vaAapRc1Ll4vpiIJsDjWsEcq7Q7cZQ
ggVJJ5agwxzU1RW+SJhl3dEnEGfz8cYdnRIciquzpq41DxEMOdJKd6i6le6AqClDdkClXSldHtBg
RtZvXj+yNCo41KFjKYqBaySkZ8imRC9y62NrqupaWY+k4bJCEnIBxWiJEnuOfx4aNDuPDu2na7Hs
e3l2JMyU18AXVRUrEpZQcsfu8sLVoxV9GLWoDj0jqNDIEmej2iVk3d/fjUgKsEsl1l/gqCENHV5v
xyCL9UUlRMMVqCw3mJ/Xevv5jLFPLpbARw9N4x4PQ3zo4ZF1OeFGUDI9FBXMzus/adIHsALdf5hF
mg4g7ggT4//DkcmacjStkhDkvNSt/5F6DJLr7m6a0fsaDQeoa5Of9qdOy/uxVMllXgnQHK5pfdX9
cdlzbm5XPkjEGTDaijdUalnCQDI4cgj7Pm3Rqx+2eckgN1LeNh3TkgBYSpXabCR9NV4AX+h9qxwy
EgAG5fcBq//qqvVfTKQ+fjH9Gjc4yeIOGf9Vr94fIsdlvBvdj1FtLXbpYchFQMk+mgIFyRi7Oywi
BFBhQytUvwoVfOVkrc7VK6KcBxOPwsoEwIfErfozYo54kQvIs1mfIngmvSxPfBypsXPRUQE64b3P
TVmDHCC+SyZHJQRBrzSK1HDoet71vEPwcDUwdJB1KsK6nM4wtijaAFo81q1My6GnUnCHaGH5R34l
jbkl55FIpnQrfum8HHfvLT9eKyUmP64l9qqU17AAVQ3o+jyicedMxPSLCac5OQkJAFW0iOexTz7N
BXGwW+6FGZ70RPjq8DW7hHVfgjuYAFXHkO0YPujScXOcEwfIfih+1laLZJVRIBkAec8XzJHclhsl
4BiIt7YO2DB1YbgBIF1OGYYhmqVZZ1MI+gadRlNI8Y8GB0vq7qRCt+wW2NTMuvVnMk6LiQRHeqk7
GTFuy2X6lM7iqUcgY+ZJidzoW5bBXMP/HqYXxjvgadjgmA0aiNwr5bUwkh024E0CBdAOohFTk6oE
E1B/Gc+FtW4qBacSIDqntIlKJK6b2EAEitL8zRL8cTTKK2S/pvI78dq+9OMlRLz59OTGeJK/swoB
GmbDLhAAikuNVC/K+zvcb9FEScMXUo7nzDzruF2K60hZaCXAhFdDi815trizSB9m2xB8FIVKW/s8
fLHHjA8POhGnYLo/WLRCtTKdaawSQbqZpE18/udtee4td/AwTV2M4Ius3jq0ae5xBK24jdTypr/P
gsOxARMMBCFOd+IqsMoSGZg5IJEKMljwp3OBlTjZW2Dsf+pGH1NgIgXa78Fkwa6TYYNpck89Kntr
cZ2oC0fPYaNqT0kE+qGKJd0Q2Tcwh7uTST/tq2NmEUUqjnh75l7X55Vik0L6FcsIVcFgZbyukc66
b2XgwxQvNfnBnlAC2p5gswGEC0RJU67mW2Ia3GrUtQ6HytiZZRJuwf1iT8V7+13u5G2D/YKUdWON
OzccRCSl5zFJ6zIj+6qhw51q8dSo9FYZVqPDqcw9EDI6afadB3zkK0V5wK0g/snREZYurkOmiat7
7CaQH3BcD5DcY8nLMQXSp7qAZ+LpolzEwwFaC4Nhi2lTuutyLzBWj06O7HY0jm3BNbj5SGNiQIEB
bR+C1KYvu49BIvlwlJukTloBqZKtFV1pxjmCdlE564TnIOB6IJCs4zHV1crftyOKOaJlsXyUTWan
ugiiTTPRhJUIsu0w0a5TuyqQwQsM3EIfLndHHISOS57UWJit7ZtmpeXwK7/iazK9WPXgJcpSJh+o
3rDwwOb+e2Q9IT7Oat6cj+X76f8XuutWzn1Vrrq3gmqgy7UBfnYIH7g6G+MO/lPFvM/HZiMHF/D1
hXi3i7KjYdPLS2g1fPvVx4vAjJfQ5EGEYGt9yjRrvsWL4a53t1pbtx+nhZigRvZI2K10ZhLpx4Wu
J/Ck+HaU6x65+utHW1I8DHKMrIea7c2N04AWcg2jVU779nZXomQ9qyrZVK/Dfps6mb/5SN4rxpTn
Z+ABzrQV5DLItag8uBhg2aJNctqclk03Y6a45pqTgKczB54LuxRgX7jtRAo2Pb2wJdXfKFzlwrpy
Knaaq1HrAIQgyUeXXcv4OZpcxTsJvb7WpW982VSyFN8JwoBPAmeeexVi6nDT3bJah0nbwParcsb5
AFy3Pom+rMHeWYVuGO7X4LHStJsC8iJbZxfvwnSCHKbnD1x1vhylOYcIPJ70IXWVXrbA2QxFaRnv
VjYWlzR/b6/uvHIf702DWXk2aMV9OrA9MZqLV4JSei+VPIgRdPERQf5rAP+aFdzo9XpqDiUHgDuG
ISMZewFKMhHC4TA2dFWsugoTFvakmWdzOOqw0rIshHC91DwHYEB9cB88BT47jYm7vQRvyqgHO3n/
eHmpiXQkzglNg/98G0onN4g0Yu1pJb4jc1eX+MUI8Y49L0RY3GiGMVMKzzBIWm01SD43EnZL9Gsr
Ql/5fqPpBD3p9GDG+5YTxuATJvJlaErCqhb+LjB4y0C3XEbmCqpzgqDwofkWPvIqjERVWxWbHeRC
u2iBW7ax9My2R9vtm3imwY+9v+TLnsTaTaLGgzTWI+L9BpcXrnwnLM2k0b7eRxKWKPoQcDvOwrkQ
sjFHJ2K6nT2IgprO84l9CZ7Hs4b7nrIpEhgRFYKSQWml+6luRfOLDtdVWagFz0Zw9cEXJ4/yijTG
sPU+UFsGaZpsNriedOPnXXaHPVIrYGrqsd6HC4yT6wTxCWy7xpxyIJpdf9JzVnnBtlxIPUdCPY6v
BRcIzzRyRrrXmDOYivZTHTbr2zRnfLRBT9SbZTq7WMOxNsQh9A+F6QVFDM5hxQjaQH1tSehe31dQ
6Z0OehmdB6l+8YI5xSedz8md1g1uMWc+wdsSSvCPgfGEcvpsYb3youBSn4YKzcRmfpXml6oN9t+h
95vzmZP7f9+KFF1g1wDGVd5LEI8xYbQfVp/lU+TA4nps/tSDihVSTxBMvotwqNNsTldnlykvpSgV
z/4tj3/ffG+520ruIOovrKd8HV5eueZ4lqT6B0mip2CEc6ZFmWfcsr1o0xYw2iFSEejDrDU78Vkf
xv8X4IcfvN4IMXTRQZ6viiwaDmRzBpkq3u67zHJJrP4Uwrc4bPicTpxPtpcUifeZpvKZskH+16Jg
SmGK73pBQdZeVmT+y+ROzcuuFN+qdoa1eW7CPKbzRBQ5bN63V6TB1U6QAWh3lFbc2Zo5BJDoyn6e
9zIuo+cY7XmMXLKVmte3l9smOJ6CoKtvVHUEUg/f8vybb+W8wuoBYbsH7fBFpwX97/OcKekZ2qf+
O2yVR5YVJO1ap+mW/bcbMM4cI0dtPc5G8Sq9xjKroNXApt9tQIMUI311luEpv7aI09oANdDGYOfJ
wlNwm+02VOzCwfEPV54gpsuL66cpLtGr8vBnqK5O39ONtXizaJ4N/SZCkwmY6Mrv0jOk3OxQlJ/k
Ta8NYn5p8GQPtk2gHUgsjGsinLJpOG6n0o6VDovDAXmXvjMupWaaEZ3e2TcAjN0HzsAaCi58qRo3
590cBil9kcNWDGcE2rFCNWOqqYtq1EN+Yw76d1RBqSqHmFP5appgR9Vf6VK/1G2Oqeaea9BtSlFr
Iw3ePSf6YIwVVwJ6n84C1ZWpMvvWN9yvxghPUIpOBOTBCdprRrqr7XgasB7yWxZXmcinAmDpH1CA
fYWJqO6wOoI2ukWsq1eFq6FbKiQTi7wvYWloqw2K9EMkMJsNPE4Mx4kFc+AHcAQgX8nb7AV24z2H
F2jn9gxS4Hpt/6msVV50pvmNTzq8i6Ab49GjSIkNXlZrR5Fq9m/2l8BiZbS9raonZx4FvMBx16rf
XYtpA+U6LF3/Jce1l8sZ38zKsnDujJw/d3LcWSwMCSiEzjLUenHrIhA2oIwWbtyAhd6m73Tqs1ql
34/2y3mzGOURnq2kzl1M2B6b7e80dSoj+4n09Qctf+1u58TaG4W4NRlk2KXrZTUVpngDPfeOw/tx
NYdsxNH/WT7AN3lfoRSLAk2GVu0VHVxr3a8A9lQ4hTgOR4p0bXLz1s/CM6fMmZO4bE4jCxpNP22J
P3o+KuFpFbgXWwmm7x02tgBx9nZ5zrkKNpuXVAyyO540EzPsrsSVjzOlN4WvfwW6GGpI1p0WPoar
xi5SpKOC5k85QPDVr8+iuNwLu+INWoTkke7QsqJQ+RrEppizvfujGgMVmNWbrtrzit3nm7EGqOll
KF6ZCjtjt0784A7FSt5xAc6+QWiP6nSxXD6o8njgiGWjNb0LsIVyvTBw4PAE9b4GC86MvcGB7I21
EWSRUXjOMfDgP9o2iNR9BRjbI7it0EMB7xbRCwUif19Dp/hMo9TUkNM4XjOe8ksczXaETexJeX3S
ZBDwq1iB6P/jVHysGDDarcAeSRyVmOp6Uvu5aHvI1AsCdtVdohKbWvIpIYRuODc1F6rhEOy08arP
mPbRZqPBHgx661xyB44Za37pwBTNeC54MUaXwOb3glgdZmyYXAv/ENXwTdZExCUjXu8YCdW1cvy4
1Sa8s3kLbY2OEFBj8yOzPKDAul6QjEcNl6c98ohnSPHBCBUok2LcyQx0yetxd0cmY5nUnABlqwcY
OGDhHtjIwLtVT/7lMzM+iV8S48L+waPwkRTI7sAByHp8KM06OrkoOQ/APw0CLY47LajVDhQ61FhZ
8kY8dkVSBX4XR0YNyjN+Ob8QPQ/VQLbIiExJU1tLJB/VBCeUY1wWlo6rQYMgX25qIpjxvJWoWGmm
oS9xxIegz8Rap8oU4jfj/raUQdHlAKVFKNDwyD76i8uO295HR3hVW8GrGz1lkbAc+T13qt2hN1Is
y0PsDQVoL75pD2EA48Dz11Mnj2CZSmYc9WoWP2ercF9IHTgcWrxZ7XzXB9A4zkf5O40HzYZzo+NA
J1wdyThMto4lN4JMdOLpquJcA1fCeYv3l+U2B+TzCmcHIXK91oN/tY8lYO//mlmXqe+mJq0VCeFi
q8aECJu8hGjMvc3xvDpb7NiPqw1zIwQJoqHg8kd4iiPxz0we6kutE+eN4JiFNshZUjZfScjZd4Mg
rGa/C05Az+wRSKPtsokfgi3Fz6/8BPOun5GR12PB5APSJ1QkDDGACJZyPe5Pl2JympKQ2JYylfRP
vvnwqwYK8AsSV93s0rs6wtxt9+TW/M8Br3nHXlEtnC1/XD2Aw70QLt5YhqVi7zn7DBjRHr4VZgAp
Z9nahCf88FjNH1fslHn//AiLLMehBL2hA/ESPu0pzLq1UCH3O9aTXFb2eV6bPNiC12YdK5sIlglf
k7p3Js5/tGGOfjwXQOxxs6LzUNlfbnf9LW/oUaqTNLFVK262QdzlEzSEtd0r9XmOxsPSnuacusKg
i9OZyjWRASfhopF7IpwmNZRHnYPfrwwvaGCumQpr/E+MGS3yMKj8WPcN8N9TdAaA3iGNYCKH1nkZ
HGhMgTPBDJnK2kaBZ39+rkgsFJoU68FJdt0lzpNXzWkg5Fbav63iiSdce/+xdVlRvsxhr+jZ/Kvb
jIJrsID/AwT5HO+NxZqH6nGJPpZOmb0bgFu7QNd/LdC/6OG9lblzZ4AudRTpeqa+YkUgTAF2Q5Q1
P8NmaM3aLkvpRlnQufKHY7rsYU4bM14yca1fTn2KIW6J4CJicdsBUdxixqfQKzLeQpGKcgEzYs0m
mSWnas7uVcg2iii9WxMuvw1VrSaq7G9IQG5E5Xbhaj5O9Dzr0bFvhgaow8u3SN/6PoMbIgvTVcH4
tg4ExtX0SLfMdV2ZWvebb8PYBGm7JqdROyWDFsiF17Q69pueVD6ubtaAbLIBBemNwT2VJ9U5pMES
dtaFvorJLrYQ0R90f8O/yUQuTeTN0JMqDh0cPSirYbceTxodPZ+Ant2Jdq7aULrhDZIabsuFB/PW
qUgKuQrnJBBO+quUS3Saj8+KyJYixbeqUyCPKKLZwH9gJ3Ng8dtRV/rr9I2Q9ujt7mT+6g8YbFex
YvlR4HT3DOAAS08fXEiTvxC5pnoDxSl3EdqWD4f3H515K5+/2ybSkveQZ1lkl/B71GZ7eEeUSB/Q
HEuJ2otKF8mcSzfx59ASD90Z/2p0gLJ41d3U02MgndmJANSNHD0N13gM2Gcg6dfvxa8k4IT8L/JH
K+Fjny3PRKfspiNCBa+7sfNzfKLE4xevfeY0D4uYkA04veoRh1XMqEuICdeNo3B3hrHamzpD8EXV
tVuXXkfrPhhzXNhAwX5zju6IMseITPEgXXgDGuCfPqZnXdy4QYpeH1ztCMO1Ll8+o2J5KPR4VoWn
CjNpVMgQ6YyABGGjrg+y83dRGFvKO4t9oegBK5ONZ6pseOLpJkHlUfxA+k+a4Y2BN7c3NXWhc5WP
h675MUn5OhjkVD6pjEIH/My4QXYXBWeMP3R+uh7BwJ9Cp9na9okizuLfi4pH62Fm7l2GmY0blMRr
5lCySGIwlFcv+tUapIB3LK4P3rGd9O9LyIZKLlkZM/yW7Df2oNTm72xjZ6+Nd/S2C7L+LW5DTu1l
4fml74jHYvKFpDM3QiZDgpBJEuyzjOLir76vkyLpcydAbZzRdKKtvMDzZ1becfv/qmwjNWz6FiAY
gkGPs0n9L1aWL87KANzdXrMEvqgh3H2WCyfZ3+n9zZsYhE1+rDGZPKBFczSmXLwQyBPcCJk6cRb1
EqcYuwCQ+xuKdGCp/KmuTYkggT+l/OHX5wEQgx2GVR4mtZpHbjy7koYomF1FWcjlO7xF0KNuGpEj
hvmcs2R6O5R/21IjCGWw5K0vyj86HCRGOI/cnQV7i9HUTgKwp55n96Y0YYzeccJKI4/xuGPM8eWV
/m6HMOHvS0gN6i6ZNVKcQPXh5ilcTFOQoA/x2HItFBublS4LGKwYSWTztr2qUusdNoA+U3woEPpf
y+e/j6uAoLiXJqERBnUY2zGvpc+h1hMNmCmaH8Ql9VkwFl9mLyquoO+W8XJzVppOEI+0n57rt0I6
TagEvdulZdJTEDMH5aTu9JtpbCoJYlGJE7X59LdpGBAB5v3ke03QfmL1xwHKr/Nic5fA9Fmv10aH
WEHRaN37Otq80A58Wb2uzJmsmimFbGO4gnvIAuxZl9y4EI/0OHXV5tfWWuXki68Ki9YOdj3b8b1G
kaPaxNDbICI7TVYrAOnhrFzzAKOC6GR1q+r9XvKJHTtQqYHWjs6YWUDrEm9xCrJXWJEsre8M9CbO
mmupoXdSVDJaRcGQKaq6o6OratYGCuGO0r48eZvncNo8yp259icSLmbqaaMyEtn7bMk+KAoOKETO
cyYSnDGUMHeE0gTp25ikIq9WbPy8envbdNHWleArnyv3vmHwJAUOc18zP7G/Y4vC3/At1oez1KeA
+BYT15lGUE6QOl/vbZmgB6qHZMzJimLYAECdAEotGNzXaDhQyXrM79kLmAUOEhXMQhhnwGFfJfwY
jb9TtHrQOO3ZR6NkJHOX97WqjnLPjEJcxv0GHpnZgCOmysj4LSDE8gswUkZlS1MNgoHM8w5lXoEk
tyjits8GtAYdDD9OK+jP3g/xKok1wEYbkh8eV9b2F5n+Tn4YqTBVFKPDDTHG+T6dRa6F9pQ/vOwe
Ao/ypOta228mt4IkAbjGuYJd8GpMbNk06MAFSSZd3InHV7cBR2v6ue7J7nEJVTp7QmZ3J0qpmznq
+EvmhY5zttBErFplDjX/ukNXXQ3VUziCoXEhRAwDfLqGHpRMFwZL/7an4QORcLYLShXBk4BrHgWF
qK4N868rv2iEmyBKeoBhkssvxEL5vujjd4/5hY5NbOXSTuohXqOBTDL+EoGuT/LSrYCW6It5p2gW
4VlYl1LeaIV5JfyNR2hTBSIiV6WUNZAwjt+9L5KeXuVy/4Kwtxc/HTrFcjxfKrOP+LUi0vlseDuW
szL5MUTXKqhOFAFZGgJchvkPnfRezdbAFT1H6elRGZrvKgvb12xVY9xYakK1aOUybGlWYz5iV8+J
l8mdf/MZSFbhzc8yKq7zOvdLG4Iockzugt8cvqxV5D4e9BFeLakht2M1K8AU6OLkoG5NhkNlsLYs
/LHALDZPx/qAVBW9HdveMgji6kWPlfZ4lp7nUDGdwkuV/yzlQCjKJ6vE9rmN1zhke5fna/uOCMQl
IYTdhfzpSRuQ7mM2ymRYuRomhGxbmuZvSMpYhn8rw+Tgd3OksRc9ErdJG7q2X5k3x6AjL0VOD8tk
N+vBNV6hjJnYnqRQSrhHntNhOh6I7mNb60rrHQzweN7B3FKD2aDlSapzBFW+aNdTuHX2Syih/6sC
hMUdy6nsXYX1Ayycrp8NZla1zSdjzU+oSTZvrPA+XIbIUW8FKaRKRBFyWcJz2jsKVjHxitUiXzD/
kqLbaA7NrmK3IHLgDVHZYRDt8+gOdbXvOj4j6jJ9y/GZeRcuOtU6k0Z/RtZzzf/Zlc2zZJTY3wc1
78V9UgRAwSFE6V2u2A6I+1cBITf6hNbioLG7G1iAl1T8Cb7cjZEQRt+mCNjcN26U47IH1PlPFJs8
42COHoxT6RWXqEPkXqteXkVi12U5NBwzxHJypLz9qKwuxYPcX5BMvb/r2M5SBPknVEburVmHmolZ
OZ6JBW2DhzL6VHPHjoGSBVg4s/8TdsYHvOwPigXp00e1zSPZ3AV6LV3N6EN0y0gEPdGXaEs271nx
2fN/7p06FC6xctx8nWQITAdaKGyiu2PdwvK+bQQLtBcr1cci3FCZiKjvMk1YrBlTJ5BWg+EtnPb0
q1RohiwdQr6yjMgYaYacd543/C2grueA5ir526m5BaG2tOQJ2jCcX+M3d70phPoGu2GpIUBsSy3T
7FCrQIzbCVsKmXlRRyrTS/43wZsciRWz0w/5wXOGzmCPtiZePpyqi+pxHFVF7Ch2QnGckiEh8XfS
aB5Nazge4oOWzpZfHL51PFjShAcQuU5zBysadrh9hDo51Cbty2W3u2xkOh7rEdkGSlXzq0AW8dlB
qzUjqMfPTTRrg/2+oMtKhDy9UwDQQ9sJU9Jewgxp+1D3i1Tbbn22dFjkLSmBRsw6ssnAu1zSjxK4
CCs30ox6CZ9EPtj8BPe4V6Do6Oxt6xJAtm7AjZK9xqQFAt34VIAIemKyTlLLD7jvY9nD6odWf7h3
yJoxjBUngMPfOdId1Y+qjnbR6no2NPz3CYpBh5XUikrIeharqVv65/HwXUu9rT2Mq4Ze/ELQIeth
jNCGss6Gk5i4eBO4mw7VkWFCMVngTgJS7Y2F/UTPlfMIxn6mIJwPINYNmibgwNuBkNjFpcz/ppaV
qLIRQQ2KGmjkgx4qQOK2vXv59Xq/QXYgKfm2ahhT8VS4GqbmhMOSPePsBvWITIW/SVMMQly+0+p5
vPk8/gjMvYXKU921BStPT0qS//kBVihIkp0vXVueda0aOLxGSEFko25X7ueHFg65nwvR/FSoeTC9
oPknEv5vPiCGhl/b7wbrd5lRyBSgHV/tKMwXp5n5iHRW+zuaiMZCJ9nju9UtnRoZWYcjmZPk50bJ
GWuCjwkrXYo0y4xjHvfeVJ09Saa0U3LFpMN6cqXMxl4U9/5C+58wgvggybwv2OOV41zfkP/qeD1d
ptyr5eA9KpfbcRh9VRkj94A2rQaGavOfk6nMPqax9MVUynnn2I/mVT98DkeWkuSqyJuh2rqP2yFd
QJ/bPNUa3+dxp8HFy/+nqoo7k/FV/jWTAGHsztVPntqvzTsBYvIt/9awnI+pfyAGLBbhFa859n4Z
xt6V9Nv7HI799dyn5XcYrbAt/5KDCiKSdYytahtK9gHgyaOKdj96szeAuBfGG1Xl+Lg0BEE6zHtf
S3/AY45lSv22a9EzXQWhxMCtCI2uyo4CI7K33r76frln3wcflm+qhdCciEJyCQCbHTD387aq+LY7
x2KfJfp9i/7wiykAa9AHNfVah+7IM5CKRvhKRU3KInvly9bgmfNoYSbS+uBMwD2+f0bg1ka4xGvh
LPDtyT+D6YssbGIbBs5n/emD+cvt2H+b9EeBBgCE4MjnMNsCqmF2hBDQZZM5wyaOcXB5xHkhKUZO
1ienoEPYmRKqQlCPrRHm/gupA/hGbfYyhtVUCoIEMAm1RBAk4S1N2AgSSC+e+vQ0OefM+igDACfm
Ye7nRoX9UW9LCdHvsr6ZnSxsK+sMP7v0RQzMUflzxVfqLvKq0sdsAhz+S+crVWOdbLSb1DZ04cKk
HOrCBJHEKvA54bkKu50q9OWTYK35noKYz0KAL1sxgXw0e392Xt4xsBw1cjNxVhWjwMsYhESii/JP
igBFoUDMLTdWEG8CeNYdQo06CX98G5vucfhLqAxFQGvqAawrvZOmGMg2/1x5zGCk5XjxBoV/LExp
4fILnnuH/mbMrwufBaPE0b1IId4+BoNBIISlAdF+fNs0MB9Q/Aq1BCagkAkRe6PhoIEihRr95/Yj
lFGXFZFYBBlkN06WUlpQmqo25nSnwcylu32ju0LiKeyhwWQQ3hGNDOSrmbqZkAk0cKKZb6VmhWjM
TkH6sDH3coJtCJPDm6u+ojfAw7arteBF+hLerYTNL8jTUfv6V4tfqrtnaXF0P/NAp0cLkoXgDXo1
afsTWgdfNyD6cLcgiFPlLcKGBz/uHR3DcY1f4ibraOnovDSz3pYfLJyBnug0fNn4jNEg1lgpvd4j
vAp85NzDeow45MHCEuIM4oGhvfvC/g01EQZVQ9l0PotY0lZlC+Z7ELj7UFdMvTwwauXu50e/sZUi
J9rxcrnr879TBFYEcYvfvNcOz6BPB+TP629kREVm3gVms83OthFFEmwQ75bOHoPVtCZqQWMYMe9j
LeujhAuXAEkqWshklrZEHNc2L8g0Mhm1JXh9WZW8NLJs4+fPOvZ5OwoCGi3oay/pdDctfKIr5U6g
imya4UunjqIxGr27nDxEcCbsxZBYphfhHeon7fWG3qEqgmMXogIhg7xQEhtBAyizrwhCOmM7Yexs
qIBEUJRgCNeRdafHz+8KGC8ITOILKBW8i7akUpgMXFa35aiz8t4DzD1VV4FR2OF+W1ZBovJnwbsu
tUTqU0po5Rs5Wbau3VaNMnzrLfEN7CvYYQM3eA2OiT2/DnLo8JhPe6P+TnRzPzOmKsWPtGdY+bsm
SnXEeOXdEat1vw+T7UFjeg8sNrWk4IBSkkc+YyBCgNuAALuOTlefKkVS15K6TceryDLRltvQmxn9
MCcFb/to8pzDnWKZ7JSt33sG3LE3GQg8KbKZ3vAqf4YCx0T1vRV3hpEKG9OBV8HsoSuZQoXhrHVt
q5VAuY9bJqDm/YN/8fEq0HwqZMz+IpiE7oFRdYNYiDKbYLz5Vy0gwZeS+LQgmsvq+Aj87slNoavx
SLq/Jjp0dJoMu3k4tbuMTzAfTrAl9r+8BhYvkmjxq+OvhPX7FIkAeXXg32dPwk6wNxbLDG8gQAzt
x3UgkkkXjUAMR9bpmw52UqKicDrW5+4Vn1xlaWQJC+pHfQOQG3iQJHe0UNEL1tVcURQTgFjHq5Gg
s4DV781DgN5HPgRO1Dx4zw3Y1nuEB1JCN5fTflqt7/I+0igXPJFvO/l4wf/taJeLTTpFKT8wHxKk
xFaNs9lzmnGlBW0F5GT3heWHlVtc6o9xpjm4sixB0MMLOKeNRAiNU7ER5nbDjwbyFqdGtuLMWGtQ
DqsJ3Py3fQ/6So+WdJikHdbxKmSKth5J9mH9aRFDkT/+53RSU41HuQjrlp7PP52YPh2UmZrgZJTb
KlCTrX5auB4heUYp82STYrNXZ8LCDQttDG0Ievm4hxCYYN7WcgkomQ5xES/2WZytwTnWQc992D3B
vEIq4UmWJ3nS+QJGJScEda8/LSTSIs308L74pR1JojHzAlHyajgK0VH/OoDM84INWOUr6gWejQyV
BIJ4xuza6a8Hye45RqE0gMlvE4hamak5SUZtm0M7NbJ/sKQS5nxIj+K8jYpUc6dnNO1GKyAWMp86
qUd4prPehLPWbcXmafTHW0lXKcY5Pl3Rc+l2SiDvEbtivl0RufA2U9qPYxvosodLrf38qh1adG6F
WoFmQoMn7qui9gSv7edB9TSqkzvOQ2wg3afAPpWtL16H53IBJKnW8Y8TgnJeFL/xxw5Cq6Cb1ki7
8LeU2t9o85PpiGZX8TpaWpDnx+n2OJnTznyxW0AV0X81rf8lPHtO5c3Wk9dOxly1WXSTONQWtlMf
pVqexFmxJRHAtASuX/UWFZ8YEnYxuhB6LjWgwA7a1OrbH0F44alrimlMATw9/YQ9a0GZy2IcRqd0
XgidjSGLkNA+mF/zF9NBcN4kUl0qq3cqhdXjZgtb++SQcFGMXObFsBFlSgE2Gs2XFFAwfCZ9ciAD
yUk6WRpuz75MVDx42KYpxE8TMbr71R/2Clqg2fzRqudBrkvOaUF/rd+zyTXU64rQKDsKnVztW8GY
UsrWTZTzBAjc+AUHY+tS6vWA1E5fFyjyOX0FGaZzob+bG2i2q2xJHlqabEZI/mSBOBjxJa0CRJsx
YCvo4r4GViNaEXWHtx8N6/POi0UWwOQBxdNMuEcN/kVqecenjvjzXKXwH55dRDyB8MW/A/2pyVU6
Xd7bElt1sqS6rQ+Re8xBymltfovwuRT0mSyxvukHh8ZA4EhOkEd3AabZrhVn8yO3V91z6uYro0gX
P9dpZFhbQZ7qSl0KzW7h9Wl8AK5kRQcRxYKWoxJOteAtAz8hW+XPumSkhTozWTKL/JAYMilBTPGw
+d+1sOpXJZXLBSXZ/FNXksyj850P0fG3NNFPZYeeJWjbWS9tOauWCpibJ7B2GaZ8h4BPxBaqAZKn
8K2vV6JoTiG795JYp5sD+gngy4pd5HVqoX8QQgmeURBn1TSJ0PZSXTStvd7J1PRp/RPR1P/zLVhT
s/QmN3gd34I9+Ynp9yogbgpF3Xr+WmSk6up/C/AAZ0baTxaaDeWjE84M7BVqieYC3jx6JOqXHACC
bq1lP+psD8bjvrz04ruQoftJiBe63rXyYmdFSguVk98RKJhaozVgjWt+23p14HUopAhKO51tybYO
KiVsAZR3Tx4zn1XAk3ZsiEF7N/Wbsq8lvH8yYfZmiq07vOSju2Yei8QnXTyUms0BFjdQCSLZO9Qh
XA++mYYUtl0KQ/emCoQjwPmcM6a/02/c09D1yRojhoujPh7PBf++KK2CIXslNu0012sSaxKq5W/I
Vdwje6QrDk21sSO8uZ9pJhfJM4j60WbcJHHqPBWP6nxgWD7A9uXTkLupqCnGHneXtiME+wZRfwOT
zDOeqszInNlhunA9JRFhADiaJGGNZK3p/w4FIGNmD7CHgoBa6NwGHE90/LU6GJDhdfGfHJEnyz0f
yDXB9IXi7WK3AlOh/MFArLpLZiplFl+1ecboVPK7e+8awWOuKTPUJ1wp110B1YcstZjqzz185H7J
QSpOuASOLCT8R1f9SvYfhR9yPMI13OqgCJdWUd3u4vd/guDtGtz7IrVqzRtIBC4sUdARdXnC5R4s
e/YHaA4vq/31n4RcLJShM0FDzOBpmigHA1T9aTEblSfELtwu6hg30gnE0bHpqvGu6EFponKYXwsi
wgvOx1AJJv9ik8WC7NYS1mTTN4MKRiAKVacfxosvlCte5CH1Cxmk01NFmRrFV6l/dnj+IVIjN33M
5GA89wscsQZUgTAKOumFbLEZcWgQ0OvX9w6CL10SgMJEz5vuFujY5tdJ1uNOfc8WyjkIPb2HLiv6
vFepoHEaSGFXtuKwgO0lKO+8uSZ00hb1+2spkqWq8b8sZPZMIdWS2c4Fg/a4wrQkIthHPqrj4q2o
0d8imG03NhRxBbi3VAMlMxUF+NaFfIK8NHGZ/u5S66NtkM8B4P3ZCjpOlYBSRq/byhcZ7YXih/my
6ULLEYe3eTTSszehth2NlffFouEUVega+XV9P49yVXXJDj7urNjDmduXkM8JpsgT2Win/DcMYw3K
IctUsLVdNYpFmYpiudT/Sc5ItM0T1P34zsjPlIW9g5OThbOhfx9SdAgRGGKpV97lr02niyjY+lun
qrMfh5xVYCnKgj+97Erd+w9Es4hCL5N8o2LMclq5jiXoIaAYcqqChcNjtfmmFRSYIAAcZO1287SX
Xw2hQfE0UsvHXoCJxhO0su0Hwu7sg5msbHnWDiZJ5YXAdp1VsIVh4Z+DFp+gssC+SA1YiDZcQCmd
dHOU02UVQlVBXYkgvCqSnIgTJQ5SvOg1pkcYEVTy1nmUjBWYNm/cFtGVS79hX4hin+WPf7qwCMID
5S9WnFApSXSma4aXSxXmFvqJJQjFSfCFYwOhyLW2B70V+mKCpfSnxX5yv9zghVjV3M6ti8WDuHV5
eJ2lmGToxB6K+XT4SOGEFsBxI0aaLwXEN2acZTNMchPb24XXjTYGEtCbBXc0QnLCM7uyMGqGxfnL
Ry33+UvcgjlAIWUnhHyevCDd9UA53vdwb2fKFZHHleghIUpz9YGXjnRrs4hEIDP7kADxwy6kSt2P
bB9WWRuWynmBnvJ4fxa5AkN2I+dhOF/bfydKKyk8VOgr1Y9iRN0JPA26XAPWsH1bP6oZTtzlV+ha
IxngyfyfckdCtgQ0x+XQ2izOcK1y3a29PJKBZ4BO9ccqKNu1x1v7sIAtoENrFZnVaLj5vj65cjOA
m4uVA9JeybDIN8LY9P7tY6IsJXTARCgmtAY/Py4kiSYfrF2+y5yox+OrffNhqOoiy/SRQCa8iUeX
dlZp57cfnZ9Q2D9xU0EdCMMfB18SJGQXxwN+KfD6WGyozQo7yJFaBOFj7F03l4itJXu2PSKprFzp
ZDfoDBLPW6c1IbR0ASL7jktzf1pXhnpKXx96+r+VYXq/y0YwjhW5Nq0+QPXXpp650jOn8EwnvFzR
EleaPTKwPHx0iLHJbZSL9LaPZTdJ7xAWDl7P94jvKDCpJWyqZ1MZgIrJGJmRv4wNRC/leDj9MwtV
AXSshDAqlul+sKLrwoPFtLLujo+6AZpavNDyIvQ3YYW5qWp8JsOqGBqUIAP3DXs5xeexYtWvpT8g
akmlf23Qw3Di7raFMX4W1LpFilQ4nh+mzhB1HFOA4/ZjUQfAZ2C2udUIcRKv/haQSQ3lEi1YIYVZ
dyhOuXhxNyNcD0knMjuP7aMtSlRJGYYHnP3qX3Gh/dBF9l5Cww+5N+xlZ4YZnFUoc+qYdBgorupC
eNrfr5yoqwwB1DN0mjL9JL0Jyef6I7UyLq+yt+/UNdtgB9AXoxUy9Kcjd3XlsXhaxOUlK3oerG93
5qkUPxxoaJN+WV+93X/feRJtbqiwjcANZv3diBbSdxOyDYj1PoLY4TBPjKy6SlULZSdW49d8ELZG
lXGa7TKS1DhH+wCXio/qAKCMyKmTlU0MxAYPRITUqYHvyVJaIcUBLWxfHVZ7t0K6OJG01WuKiNHq
neddc6DFZ3xUp0L7tz8yuJAUwgmGly6MNso/au2ORP1WUxSO2C8m2sOolstVHfB7TJxaZufi8z7P
NnAOoiFn4UHyT1dyF5EDs4P9M83JKEVFa+FctV0j3oKki4mOYf2qfgPAQ+ozAKpAxxLoiN3Dz/j9
4YhdJuHsmTBJEG2yOk5ATPfEFg+21flmq6eZClbDJtkitobsquqhPOmsMd/20c6D6FKeI58fm589
6lFC8MaFuptu5Rp0eaTosHaaS4U3uhqb+7tYrxWu9MOXp5VJQnoftjhNp/xHL6Hp2+5JuKjwJiw5
oouaXFgQ+mYYhs+F/qdEYJtduXGu0PZbPbn1cyY0ZQh7g7F7/8gyMR2lq0bc6YLalxNgyO24ZpEm
F4SvuKr/C06jRUsIdNFdhLXKbzidczOREsY5/2du4NFMTPi8Zct/xocmPBxzYFI8g5+Gb3ClKVMw
pT/G9by00SC+rtztZViTVsJfoVQWfKRR4x9eylfmhdPQQSwBVlQFmjA6A/SNdy5pmqx1KfR68ocC
PlTngSK/hZpP7zkEOY0pdyBMvYAGCzz6qSxoTmOfLDLidgD6IhYfUYcdLtUpnxCZul1HdwUxAffH
338RA9/bYZ3b/vWPUwcoNF486mKj7viqJBd/mSh8C8zJIB7qKxudXYroJuPqL97brchxCqrl/dlg
E33CIL/rdedFJbGjE4bcJ7Bmbne1SnzAvgkPAT22AVA/oCZXFqLY44+FQS8w1yDEFpwTvyngSqUG
SVk7VZEMKxUYbGcbfGbKswYYH/6Rh4DDFLO/y5WCSUK/KqbPzdLQgDD1JOfQxPJRWXIMuBi6vvRd
Lqs9sxLPAMHjnw0wbfpjJzZAOrCsCaGT7n+IXzy7E7rqnLopa4rWW2gznOVWqREZYA8cqV+HE5gb
FRsGJu2JzWxqQ7btAxbRpiz7jPd52ETmtyZVpjYqaDoTzYwQ/uZR05e6JDtaomRzX7xWXvx6Z79u
CEyB04ZYeMAVvfKP0qIMIkH7e4qN0MmRv1aNkS7kg3uLf6XTuYkOHTIEXNf0+yETq4ZB7cMe9ypa
60FH9cQG43Lk/QjloduozZPLxfBo+yB4/HMNB4ZsufcflXqM5t1a2Ta2bxvfp6bTbMIlStlyBs4F
9NmjFvfTFjQYWfd8kNItxwPyyHHnAKAJJzDPzGyYmzlo/j8z6JHuRw5ZbtExSO5d29irimPHno/K
75mTey4GPrSZTW8Uhr8LT30up9R5ANh/ThBpPQQ+YL6g4hFSUthJ7yPwxd31upmH8hcMTmvaOcQu
xd6A1Maaqn9khGAk3U/m9hMRXOIDvfDWLW8xTpFDyLnz0ZwzycQQ+0ya7/blF6etPag2s/WozR2Y
YxSr6L6mMFTw+Uhv6sTjWpWEJF8IpW1naqLD5JKpZl4YLCzeH4GCmy9Lgn+jZ4c/xL1sQYTBQM+4
D3tUHM8ERKBq5K9+w5vk0KfGwgak/d+ETZozRY0nifDMnVQqthH2rARepEqXQxZUhd5RpgCUvj13
orShM8/bdc0OVepixDWC/GXMHZBqwiQ9QhUjo34e3ZrIyekNd1jXVJufiP0leP+6KRqf0Lodm/XN
/s3m9jc31LAwF/tDYeTIORYZZq2BMHHZRR+IMcYAHDsreMcknJ8BC2dvRed+FFoFmMTXyxlWvRHi
SmCSsGufgj5l4wBawL3/Jq9Tb01TDvrKHIhVISmRh9Ahj6jrIlybxvQAYDSc6xN5Mx6QofTxRXGD
8Feves/E4+1R6+8Xnod92wUIVj7hm+NI1Ysgw2PKhr8w7qijETZks1DXG6ov0Is2uowgjRtv5LCS
IQG2iNy8NNX5T3TzAToYDvHnUxrW/4DHPNvJJ68q3HnJa+Jj1SQyyeXCLC+nvE1fNFpS0Fg76mNj
HROirIUiqmMF95QHp7FIOwd4N8Sg+RNU7089ZPR/mo0ekgwBYMKkjKZMi51GKkM4HpdEfBZpPeOw
6E96jA6fi86ZcBfCezZ0lNcb5nx+n7VI1kmQLk+NMWAQAjTJy0Eg64xpfLp81gK7TRUK0uAgKulh
76qJlIUTo2J1fKz4/7KITa8FRnpfIHm3Wl9hvZBvJ++Wo/Ee+DVJYjhVbYVZUMsgf0/Frx/yVdvb
/hZHIeUlkFDAkP1fnivIhYUFFMPBimP0Ug2Fm5DzpTbv8sWDbG/coaLZYSiZEsn9RyJjBpAwFh/p
CZ3YKeulPhjbQVh+dSb3Fp5KwQe5nssmkpAsBdOvI/wQBvfudVTjZ5FxBGjm4k7fELcrjgXVtb54
wNstv7ELk9dlG4Ct4fTx/tJW76R/3WS5aqG5lZQ65r4M2VMSQ85QSNNmsoIk8CNBpOvzbQ4WNncd
3ZQp9cgRd0m0iiCgJC5T6yrJkzf79YRQQuiLFMarmoJfdLk4QICHVSsuqRFivjLap+2tb6ryGSRG
5alblQPBAoW31gnTdJxlXCwIxs9VjV6KFRjFTMZF+WqTIcoYl12eDtodwWEWXGe8E9DI8ZCf9jCk
MdPF3PAqrOGmuyGptJoCnVqkhzGV8ppqVFh4MfsjbltRZuMmjErYTiGiVOBZMimNyaz//MEJHE/G
on8du+3UBG5FXWfbJZYexaMUP+/IjzXT9+1brMypKNC4B8loajVXFCFxxseTNbpRiYqpHUoDZup7
qSGID0QhC8OahM0BZIz20yrXfUZOwj9v14VyhFX5dcMx5zFljY22TK3CMFt1sBo81mdQ6AZnq1CA
yrsr9ZQQ5MtqjJb++SdTP2syOSrPKGlf22PiUF+pKrWksHVMgzZi6Ry1BDkO4ssWHZNwq4DHJZBZ
OAegYeXsYyzfU/8W9Hweg1zsc5ZwGricq+AuheZGIHOu53It0VvrSxPeuO2vrlrYJWiIGWRrabKd
6+yjAaG2HDK8yaB7gYxQRxksme8C6YVT7ZYx1zSXtou4OtssBu2M4/GyBbd7665dL+Q7gbihjc3I
qaaTeTmRVQ34sFx/t0Gku5DBq9nTXB+JJ4Toy5NnbGImuCsIiSUDBlV+LWTQJfK+Y7i8zukqovPy
nsMR5Nw+OGxEGlMzAP9eYKH/Fic5fHZhf07f00oIUeh63kwuCCf4YNDE6czuXpjnyYPrqNlxLa1N
l0FCRPB9lpcWvl+s1GJxBq1nGe05+fOI2oWIl9VTxKDyUoTB5aTM6naAw5NjOYs4bNEftLRVQtML
sHCX71OBYAw9iQ7GkdCk/qpJSXhNs7IFT2NAYUBcr3YO5MaQG9e1dIzowUpdluZsY/HcTMYmucxb
BiJOiwVwR9Ka9Qua2k1b1X7dNdfEya9XyJDfKHL61gbNaOBOwH9GvpVJ3fkq4QQ6DQEWmXkBCTPj
SEO1TklRxgwqxHRiQGVjOc3Xp0TnR0azGc1RqX0xesA80w1JWG7uJUqzS9eE1DyiPuKJbcpDSojH
JNGz7c0uESgiRbqOn1IHtzyVUW5VaA0e4pd+wZlKfJXFkqAYp6ATYAZSMsdh0kzNp9M6tyQgjMq9
ykhmNKu4fDE0zwY6zzRuAelYLT83smPBb69TWbAQ8oRwCZsNg3Lxs47Hzv+pTuFAb8X0VcmaD4jy
kLpr9wwvKAzEnbvWXK3o4o9kLjWK/ZPw5gkpl+0ruXz7xnfsNBrAZyBzuhXm6LxOFg5hes7dOiwa
eOgZDJd4Q4ki3F7OiCF1AXrJppIyhrnC48nfDSbvf5NoVVlHr29KPEZykt9Lske/owWqLWrFNNRA
TG/Z4bQSW7xkOV+zIvgbQreCco21EEu996ccKPXb0z3gNiyXfTXTNnQgcPiLfPpf4quMFkjV3fqO
GLwRrb/eECWGPlPUZldeIoSYzMIag6OQp6LpVgXXfycMle2klsdsY8JEAd7rCrshvvpYlY4e9DP0
yGzF5jiffDtYnng1ArqNrelGprSxQW5o/czyKdr6Zi0dz/0ic3yQu7ynAHgc2eI4VZEll168uGQO
CvFRW2O77JU+PXL0utaVxOfOsQqgXJBZq1yS6kiMIH1xZPhzFp0/sG3ZRoOQ1d0f3+RHMkCJMU1x
DjUsFianaE7OTJj4+CueAGhrZuzXKs8tKbfC86pA201S9B1p3kBsVN4a93kSHEFfZSWIxqd2SYiy
CKcWlsVdN9sIXKq+Inu8BvJ2yi6RN9bSIVA533XBJpEpPbGp6Cs7Fy+redeaSDf6aQ9/J+zSGWdm
eO9P3txwxCDJGwDmf2wDJz1vO08QQ8TlNdph5Z/Jv1wvsjak4Cjb3ums+T16MRAxozk08d8prIAT
tPWX6wSHGfgCQSi/LJplHKOYH4sG7a4Wjo8VcPRhFhC4xDxQfXBrxDfoUgksHgi6f7hClIuEOcov
8drNOE0IlqIguodwYms5FHbZVq53+J5at/NyThyBLIBNd3+Icbes9HFgCqzoYuhhDocE37GTpTTm
aBS5X7ZNUGO9ygLFd4tozE8eRePVbJ6QY380Optp7HJTPWcyOntTUIgcLQHSTPl3AV6Exz2rIEm7
JQZl8+fqm4sfrIMWz7XkSlbkv0Jtv/pYduXcr4lrsj7upAUq2UyUaCb2UINvP7M8UEGudrH3hLPg
+O17QrAArNw3+RadVqagjQd/pWX9OnTulOp7fJP/sWErWniS2qfCVDgZ3pjEHZ3BuP3iWO4U+cky
dKr93iqFxXJulGMmqPuOgCMfNY5yAoVWgHYcajNzm8iOie0bZr/zdjsm7pyH2buKQXwgVrDHkdbY
IMZ99C2hnk36meVcqi/eZ938WzJJz1+odN23amCTt983Bd7cQKy9zJ+4YHBAq245GRwFPhqvocJu
N7xrjaFmJu0lQwfj74JfddX842ZWGwk0q2Nh8CzkaPl5NvkcWb325nqdUDItpl7o6tu+Lpey+xeH
fNfZ6tKNjXx1sijM6ZEZd7IF6NT5D8yCn/yEgTnXBA+0GS/vUIDXerxCiLkHPtU6O5YJs4adTOln
pqDdHanAuaPj2hpHqsYZQT4sGCThmha+dLHL56+YYFy3s2+3DBTSixCPUNgb8U0AZA0K6RQq47Kn
58qZwD+kQxnP94hWBh5Jze2KNBiNJDyRYzYD9zwP3b4FIL22OVAtfmmobV/wdY9J/RRbQoRqiIeu
bWNG15SvKdV1++ZLhtRf2HmRlP/AFAJEwivI49Ui4bLlBCskoBqOk+Iraq5fK6psWg3hBzn7kyym
S7Qm9adHKRY2zs7SAi5sOIwbAfBXK34aaKSSLR+SpeeN4sPXJLraK3GL3LluQ5HCNaIkUN5z1KM4
WZIVh/VH6hVtWa/D+0MRKugGESzm5yMTV1iQmBKdkeZUkRwrd7hd1gwwLlgqSsQXWKsbL74wdvCZ
ZmHk/7bmWbzRjSd+WF2qLgx+7SX6vGIhTjeBFQLbBRaYa9OsFLGd/ng8tmjV8gQvwhVBlTCf0Pky
j6ZCcual2iVxMN1JtKP0kLt6osU18b1/t/kQRsXkJsJmwJqsFg3wdBn+XkDkKFgDIYWMZSqsSoal
OwVTO+aO5p6QllElWwXkIGyL8zt+UWVZnJ/DsO54Ap2sqycguVIo99MFVZcoTpzbcRh2Q+U3ffr6
mplaQcesEAGgVnFke0NZTEDi3sWpRZa+AAbjJYQ+TX8+5GcQhaO/mcIUPNx0ZDdLiXHiTGJuP4/X
aN/WVSlulE2+4Nsy7cWxLkgCBLwwtmVUfxZkvPwneIRZjJWaEQ6ZRnzMqKzRbN0R1WvkncKmkE6p
xIYqrrryzFlmgvHf1/CR2+rLsgeRve44IbaNH6rhMxJz1KOS9JxEfVVQ8BCMnoU25qpM7fBAU9Wb
8pSojskzWhkekc/hSjObLU4YjXHCrhALwSwtKeJ5Fk05tEiXQSO81B6LMMJIV0z7FhiZNdASbSWj
Z+VJHNWmInB6dNuvd1QfBH5yJ/pywTt/JYxOMNGw0NJoWQkXXt8WkxHyT5/YXkjRf0JJEPwZLF4/
gY19KVz6n6pZuZy1PpfKz4oIVTfKiPoyXSMZoYZmPcPbuHamWwpDe5cRfK+7fUGFwL6o+ZL1YJNV
MQd3rsAcIcHMyp4BnfkYSYu+PLZDFpF6uW+jCO3lLw6zFvHCu4A/vx0Tjrh4i5ElcfoguvW4/QTA
/gqyGjsvxOTFhBzPCpFZjGsOo9bSC96wTDhwflvAioi8Z8b8u2+OXMkjXjPUI/f8L/JGBJMvs8Ht
B5qSBo2CX3TGyRhGrNqjA+KDPVR8WtB+/jKckpRlPzKgUIKhs/FUYE00WjnWtxGb0k7napqNfLes
Tf0T7z94744Jmb03TJH9S/XVDHb/5bJVDv6YCaL+tazkeOYYEUpZ15U8v6LS5VDVHZh3ifiGSV2L
X19tgmNyTrJJSb9Jq5zmGL+5CZaYyTbIAxpVce5wjkFng9YXBXdtfPjOQ2HD5Jwk91j/Lqm0LIpy
VLgymzdgA+Ayz9sJMmF4gwv9uZT2XdllRi/Az65dQMybtAl2RTAa6FwL9PftK/7nkV/t34B7UxcZ
ctUCAAn/hzsfy9IPvAFyRarSzUZGl9hqPLC8WIingQdGsm03EUNlWfjZWTQ6x+o0jugD7d9bnrM/
0OL/5xLmxvoUYn0kBrL7/ruYXTQNFWrEKi0UhlK/G/eL0q3Ehut7qSwt6v6Z/l1uqusOu5qQU0Qu
86F5mXKH72WcwAr8+WSP/rvnXeC/NBRXz/SN/Y+e9/3kOUUmikkaC/XTPlnqT6uIKGCSO0/VKK4v
0kyMlQUq1PB0cmZZ0Etf6SXA7GUEHMAjE/CPbaea2iUFwShAOnL3V8z7dVn4OQO/x9iMCHzWwiv/
K1MStqmZ22wdXHe7rrMWYQv3gr0ydUZsBdKjb9hSfmz4cDuDAoQXtakLl3dGFRFD9kBx0mTe4bTZ
74vYc54gMeYWJiq16MRetZ0JvvGgvvWVYYneG/AEkOVJ765ZDBOXJURTHl68vD+MDmniVzdtnhof
Q8xZ7M1XJS+aINmSte/JIKGtgjmXV9LTfAcTazvhGeMp/xZfTl8U5cYLHmlJJJSobuH6JPsNgbdi
5puIXaR1FBZChAvP7yEvxeosr6+C+PG/vXXpq7XbhOysyPKlddQ0Z4fXbvw5R7YVvZjHqQxz0nQ9
7rVnlo2uLkHqsNydhxAAYIXDSdoZVFB85NsuV/vVqefYXvo7WkHT0rN4W5R63abUgpzJvtXot0US
PNWm2vbNa6vT4xsnilnUW6tj8nS7H5Bjnayr7rzt7tK4aB0Eo4uBkO74DC+7EqFMrlROyBOtx/lT
uqEe3KgqbYqW5vZr/IDLUlI9+6a8BXWDUR+haUYbDibogrGsLeT2HNVR0jr0/WKQ1ZdenaKDsTgA
fB7Ua/pDzSnwIeivXW08fjqv3ofpaTuwlzri02MTAB8auBc1ZOIAok200QuUfyjW9ysjp8E1Xabm
9yiJrOHy04FBWoxQLWXQ6moaEU67ejMiEJoExl6Y/7K40psFWdD0tEl4OYdYJ+hDv/QOZdGMc6dk
Osp6RTIjSxdQgw+dXW+q+mCTl2oPGnfR+3NaGi6M150PV5GNsMQh3fSv9kRjiqcVOwYwJ1fDsYx7
+8tSn0KDs/N3Z/eX/VGw6iq631CsVgOUyBG5uFfDo+GmllNCVqIeUE6CBVUimUriHOh6XvJpiVSZ
3V209DZdcHEpDCfytkwgnf4rTreSC2RVPBBgb3+qYVJjgHHEjS2b/pVD9jGgWTs/i0zm//R7rA5X
NAT4WKNMrs+sLoibJUWcULbU5Mvke6Yr5HFdb5YL/OUC0h2t43749AVbGJVOO5o4ly1qsFK6sxrh
1G1jMnwxclILaCJa8NXTvlIiAWnr1sMJctE4P0Nvh3AYG9lNCxK8j4mW9gya/9w3QlfIRn6lwTed
tNClCrprNkUxrhHWBS8zzcCb4hzSleEQafd73jteCS1dVOcsPQvYn4Bl4qwTL7j7BxxtV7uU8qyd
7Bc3VQheOTK6ih0BgIAR3wlTUXY4JaLMdHAeW3JwLDNhUtXeYxR3lKDapHymt3UUHFS4+VSV4ytG
tPAW7MmZ/EbzJBxF7/KUt7XtPBayAuPWwFAUz+IkUVE27iOs5XBgFTJu2UpUn76HovHN/18gjp/V
zjuC9rWStnBzhUT6hzvteFYDo324EPtolaOcjXxXkHIygq+gamtWmSVCZnNfH27QDJ9DE0JYsxMr
WBjLMn6PIlKCcs/CeoRRd68aQy476Pqe0ePIksaibQHw+b5K6Fx32OMSSjfLU86tFRIt8Mlde6Ri
KNYCSO5Byog18TKV/nhNHIkR/Us/+8MgBtdGXnkV6vkKANGytxmMoglL3n65iXGuPhIUbjBs1KQl
jATb4i9N7lif5ADHr/NBhaj8LXmKKAhNQhd1Mdpldi75FJjhub3smV7nLEiezv02ZK0Hm6CYCndo
Vw89PQPr3fYWQhGAmQc8lWJ+zAZAAV6eG1tzABC4m1ssy6C8zS3hVgz/7PrPftJtIws6VBBgXOLl
9/eAzcEpCnc+QVrev1VKeUGWksBdbKT7cjdZq8O88myPYsHf4+BZmg2rRZj++3LMYletcA9l9ppf
Ij8VwrldjN+p/jNrJHgjmdWsUkG5+nsyAdOTwxdRywVHkG9eES+NaDZK0W1Vglb/Z4+sc+h+BFks
9WPnIfjW/H//+HUdEZfNySICKTkSgtJAFTXpq3C0XRVerMAksW8VT/SXzZ68rQTk3TMIAcMh7Kg/
KBtDGg/NSX1te8xzndk8DkTSufBq0rUM0mEr0efyqLZRlPSZJk3TsdsDP46hwPscMqregjtzWMLh
vR3Y52P3RTLiy6N6JYMMcgPz9X+XnRkBmJ7beUmalbst6dK50MyVkjQxKcwdRG/R+EYStDn3MDUp
6ijtXWZdGnFJQ7qEaqMK0p8rjbSiUpt1eYw3Z2ZDEvOzJAC9YsyRCGUh/YfumMb/BX7zEs4jfNvz
uONfAG5sDqmgtUxNq0BWoZLYVeEmsJ10aMoum9CXUlgYfzLhiqAgLZdeKgP0BSBEX0BXyeDt5r5E
9NcmDGNO+ZOZJRd8Y5zhAw80e5YnryjBFFCHiYO/K5I2ktb9P+WVAk1W7cGHj5EGgRjkbnx/6+td
tdIqzJA+DtkXnlELOTLbJdiWhX0i21YaVQ1ZrUIwZJGI/AY6Vfqg5b+rJ0DRBbe8SW6/dUhdP4gn
8K6mhey96JzOzsRzT8kywHhIUBI54TyU/LkxJ3xPafRGzNIVlIervf4Ro0cXck1cKJCih+8T5O90
JEJAtFHf7NpD/uFL6xU4GlJV8Rf9PAMZU1lTP6q2r5Mj8K7vKNx8NZEkd5V1+HiUW8NwK9BHt2cS
2qo1MxhHdZMp2C8elHCHGAWW9cd8c9VbFdf90b/FIrX8rRsLD5VxSf/pbISTEienZLOM5LAv3Q2z
oJRrUSfMFZSMvGGhQhDkncbPJ5NFEw18IOQZTX2TGiPvrnK58L7Ah+RoHuSdkC/iG3mIRaT4bnwq
DoBGYWsylbY9IsfL1et4S6zlextaKnLagUyjVjV5BLw9CHlaj7fmE8NQ52qbu4ZHrkj5cvcBocAW
hLYEt5iXg4YMlAWthyHs4vQbryWq0EwQgdwMMJ8xKUJEXf9dgmd2DEiNC3O91ZelhfcNQ21+Lnmp
59HQK7csx5zh206nkFx1vgSaFZTZNNMKyXCMx5kXlBDjjRBKzNbFkgRyfWfPm0Uo3xBo2p2IVton
rJ7UbWQ/zYY61/kyFFSEG+G7+WkjGlMUR7xp8cL010vDizHiFdtLRwDP18CH9WuQj4ahSfVmZGDv
iPEK9Zb5jkhEr+upZCOAKLiAa7HzDzOj4T19sUOHmKOP7OxZ7Hmd/X3JH9Ugmkk6uomAfth27XSU
KIxzbxOSHodIJG2bIk/PHOsNep1wkVJs6gCBtUiHUiGIux68YKbkGpif7ihpgwOBUV0sjb28IYVu
46BCDwaVYaAF3R7poczd4QggNPMTXztjGBdmqfWFlDoCfkx8C11BjhGuO614xfj0umssUFo7xGsF
r5nlgJ98AkLyBR0pL/vUWpdAn/BF7Jv9IeaIiIGyYMHHoa5URT7T02xW2MOGCq9kot53VWpLeJrY
ol6pmc/fGKSquZsXkUE7FDNWuePkeQyAow9BzlySQ7bhNTfEOaXFKp3GqBdJ5ShGUoain9ZVInBq
VSEFFrNrjxDfYxAiqD/QA5F98sGegZKV+RYw4pCFqOPppAmxpvbDvvriAI2Pw6uq59ifY9xx2+jX
7+PSxoUhAd0ocyBoyy3N2r9Oel5YGof4fjuW0Q21rAFeVakIkMWRrsnIPujofgzHN0AyFbnu5GYZ
FlqHpD6NY5QaCMux2tKFv6rukegNa5eLKo6PDP42BjC4cMNYqZe6YX2uQmtMz7YVtvWM8iwIk1yo
GrrzVXqMCapjhiEtCve7JIn1TaABVLlN2J55klvW7TlYsdA8Z3RC4L0cVWdd/jtkqEsGBK5xTyxg
rGl0Z9UpOoEpiiFTLw1DbsiFSaJFkrTPS577sk/tCMro9mXUiXTRfQylCyg3Gpf2hekgS75GYtxa
/1lv7kroeeXwozHHvkeHLk0pEr2kSGpJEWHwgXSLB1SThlWcmMmhrjqjdFrTyPPN+TbIQj66LOEc
WIAQJLUcOUEm6AgrnMYu38vR7b6BrfjFXNocM26jQjOAJjJweUxsujMI994H5QImoZSfUjOYzRCG
8U4AncwOIDQH7XYLnKVsU/jrbU/UhJkmvV1K7GyjgXjjmQ3brvLXOLGIs4vk/TI6IHiNnwdk3SV3
4AB+OwX/GeBEa18Qn0mcgh1Zn3a+jVIbioJgYETCY52Dm2Z1Abm8urBlLFjcavLH9GbVu4Hws9eT
N9dT8252RmNhzpAYZrmHX+mtelaTaIsSyC5Tb4DccCvPRIGityLLPEmWSyapjieEJUl9Mf9arWe2
1RAJ5dULyZfnzaeKilSVBTUCmW/1ZiuAjUQZjmbPd9FhjJSdA4LiHPBHNb2DaonJBtD714SfoQlz
UDtPc8Ov8mw6EM/sjzfdopN2gXBUNNMsdWvZTcXYQWSVgBFeBxjem70a+YDRkybk0U8xB2XH3Ytw
8tOR0+COKFVi9xxVSNPE+yExg04v8dhEu9bR36NZr9d4lmOnkpq3pDRwQVGWXmKgvgXXJpCKorU2
f+oeFnelQeiIG1xLlNOORBzfpRuUlNRrn4TqEG/DlNEfb7w4SYEdTTJkXJ24+9tiO8UrKFxvVYUh
4JL1NtYVCApzEkX0ZEUFzF4duSIiTqSggc3aES2A8KhKOYerihqvg/8imr18Rc8BnorplYIZTHNx
L4P+HbQcfRwQDmQKt58Zr3FfntF05+VTykzGJ6gxDmrEjXmVdpMH8RRyTtYspSbwjcn4hJ4jgyg3
AdCCwMZFA+7IT/2BxCiw32XuQzr23gfLQbystRPjdCkBp4MA4keOZRE66se4F/kDgqeU90sz5j1m
k7Bh7PjrfGohiToNbML4SuiQnFbY2u0dQ+509exJG2sEUYQTMqYPeOyoTBcFMm+bkkzYF3s9v2mu
jzc8WJn8/Bp2SN7Sis2DeGfiVEy5JmwgmDaKHE5IK0vgplK55K33AWV70grjLU4eS7gQ9h11hPvz
gOzV48MdVEiTQlG7Djwiv5O97qyRpuRRqiSdJuZVaKg2BhKNWXManUQvDpvX1xjrC5TIb+NKGUce
HY5lTyiQIaeJKYO1Mrffxh095XxOd0YdnJVYibbFp00sub6/7bq46aZO8p+mOGPgwWW0KBx8RuXC
WvdU7+oQH6Lur9DDJr+QkNDPvkz9t8ODGkrHRI7UPdmWVbdXBJeQtRv680ymFh4ICc77Tp/DoaDX
+lLvwFqpQXAWTYHaw43hZdefQFb33amUdx6I8Plc081QOBXCblr/LixZH7MN8pk+1MHr9+gCFQ0j
8qSVTNgQgYFntbgY2prG3a1XquuG+Yt8UIT+7bzcK7u5jJLcEayK5iv27XYMAWn0aXSvxULR0dUt
9eLkYcLzYpM3bP9cN3rfazZ+w/32TZjgt+f5O9/HjKQ0t/OXIdfNA1hgBnmPA9RJtZdGGtBu3qjq
FIIeQYgXaqSetSzyzZmjbVaMTZOgrg7wKSRzEzOYW4kAsff6JZNwoRHtXkn8kVuCzpgTWLlcEaf8
eE2JhUQRE62JDLX3x5MdoAhl/xmc4r9cd8FxdvLwzzS3SvamxQn+HcmjWjhLD/bgPr/jHkgeZqyE
WUFDCkumNZt4L/wZop/ZeRYHj4FMIszd5b+DPx1Ty3q9If/mKW7CXgdshwt386X1d5RbwNZa754p
nn9M8vBPOoYZL77er3ixBm6tyWbX5WyDAsWM3C21WZaq2oQwdoTTKbJpOO8pUDxGikvkgi6A+duR
oaWDOjxrio71QV67vRr6qzYIIlNwHXXj/yzvUnm9RaP+DrfjEIpddFOj6Ld/nyCGxRUGRg2zwSPu
RdU5Bt9xzLng1hRhBqJph00Z3juNgbN53bqS2oq9WdcR+FOPjvYvA9m+dSLqaTExR1kt+4rTih00
SETrkx+bYKznfxBxuEgQ69sRnVoqi/4v9BlwQcx0AjFAqD9KmK78efWjuPSgIjA/ZjXGQjVIAB0c
KO2ltQEwBwfSc6RsVn27WacoaN+uZObKRTqA7Ul/1WBk9ftR5tQGBpPVJgJAimcL4Hn8GTi7ypQR
PEOj/+wrMz3e7C8nOJfGu7usEAS9J7qONSilN3hbbO/B2vG+4rmsdrS9HGP+fabuR+ZL1WVdfBil
269JGkGRGcE/qtEfdNZcFR+eSjYTd9wTDn8V85d6BVCLwK1ECSuCwpk7yqpfmqP7cdqXRnAGuVm4
YGRQVoY0OYZqkL2Pee4YBVicoBVDk0PH0uQhVpktlNY3eo8bLAtNyPRgwaWzRzMC0E1j1GYRsZ+n
ESN4KFmpO/Nh7w7+vBX4xU//fovoskI6FkB+ouOwJXYrZCvOpKs1Ve2l/QUt5PHkvMxvo7e1/oF4
4qE39RUp5ni39KS18TtpLTnnHYV+NFt0q0QbhwvLRWKmFhaWnrUK7kxWzjimLvt36Jx3mzCan/eY
WIQmRpdLtRfQctye8ymJrOf3pZ8D1owi4OBZh66+yxGopbFrbiom3SWpWoVdh80+l13QjLMssW2L
X4DhrxYCMY+IxREWdtblHnGwY/rOrkD+GeAA7FXq/WQBupM72sE+H6GC11anNNGP/ODYR8d+xX8y
1J+U85fJ0URpIA0f20Y3ZuZS9dWd4tZUlHORqX7ptkEsHerOtuvRi5FpMk1S8h5klqLLcFnk2Zfx
KxyTRR/L/gLuUU6SLsewMxIMSiosiLTXYMQlo4VNraymEXd7Xvh8ZSy5HyyPBtrzHq+iKmfhEvF9
2pA6GPYGh8OPVpCoaYRc7kKw/7JTYinAeJRlBaguB1SW8pmawSxGKSKEGU7uLaibLZmPtgVn9iPj
32cDwhDhVQ34azU2TBFzO21AY/d5+nQBR83FKw0e3ePTraKdoJwpGI7DH35BGUcTM8C6CoSF8KAd
aJ1GNG1sLluIoHPlyatEcgN4JXMIXUWLYs6LjgyohDryiBqnsrg74AbylGkXwPIDjmy9w7jMONTq
0FcC1N3aWAa1AsYyZVb3q1Okr+UTkIUW4bWsaZi7jD3jo5j9DSyr1FlcCIcnreRkEZRbtzjAsaNd
bUqG9xpyzUl0HyIrirAPDce1ulqSHq41fBFtwI3XANc2V9hMNfUQsPGTFVJixDEJftJdWTXzgTP0
z//tlfMdbY9LYPpDW1IdC6gCwotaGporh9plGu8lWgNlsqd3YBXDJz4qabjXZGbdhbn72vLm+ecI
lo903aOejLY9EDYfwqqUmG3Dki3sjy7evBo7wO6DlX6Hms/1Oiq1xqBizE5npETZ1xfWBU97K1Bo
qO4za8E4OeYBTig8JMW64TrpB9yVcq/EN0o++kqZytPg7cF+Ap9cT2gCAWpqOfqpMAl4RlPJgbCP
nWaCSvroNEyQGxuR3FRLm4RwTqCxVonfs7FSoROA/+/KnH57gpQ1oka7PLTkOVoDqPKZoS5+jOns
hmm4oK2kLFOi0Tg5Lr2c6cnsyFORMYs/HUwQMmbsV+PoXAlipJB43DCaihkd63RSXbron6Uvtiqd
pCLjgQSW+UswMGxYTEVqtkUaj/FuAMtBMemvZAreskFXag9VzFDH2wNKpgCdWq6WR3mZTmegva6X
mmhgV9oRWTmgN9+iTsoUNklZN6FEBfxpYtRK6Fd0R7Be4axM9yZHoNnfZU6e78u4Jtqs/7lSq/iw
H1H5/1jTTyE7sa/RFehOdU8AGu6JbhBohfsBjRLwy6OlwtbL6hrCJxXMBC+77EkCeRWMOs9NBe0o
W8G3on8Bq48bBkRhoftZS/n2023XlZ2L9a1NGYcuPBhDAcvhJICK4UoH/SH/A1Kfo50OrFIeo86X
MMb3wXR/ndorOyRoBSLax2QfRvXg8PIdTeUV87mMvwZN1t1Cy1BfqsBuRRtfstq2GtIYlHJntFu0
h9JLu7xHMs2fjnUalise6hmGCIKXrEG8CCC5NYLpxlR1kVWWPAOFRxTAaL0pjuc6Hk0wd2BWZe8e
CwiToXDQumnZ8a71tcQG/rvrm77VnSo6GCXiFyVuZFGJyTVU6xTnB48lYBpF4ttbNCQlTxZJkPWX
1iAiZNGriZb1+ZsPKzTpHHw/UJgF2K0D0Eg7NL7U0pfGz3eJvT9eF022dqDyewHHE8Bpk8AsJlQM
xh+tP1Nk8FqQtvoOaD811f1/5ioEXtMLDMCo74XEnlNmPC0Bg77C55SH6KVkeDniPHPQkxqVYfC/
4JGP1kiKmS1ebHa9i60v/AVvLWIYQ6hsZD0bwVTFn7I/AWbl6zW7QP1ln1SswkCNWb/D+0KAF4LG
S0nUwh4/kzLKFgP/JgkRd/TETivcwu28UfKIRJ+yfhJQDmyOdLxnPcGNZXc3ljPojlkkPSXPkeiw
B6tsgFucXX7UT+1xGZ489BZ3EVizz3+JUUJm+eOe9Fe+zzPKMyg5ly3AnkuX50/p1AN/6ghnbNd0
xOQ2E06O0LotDvIAHNyd1cvE+zv2cYc2Lq0ydgF9byl2apPofFjji74/sJrO9uvpZNuj8OwgNFni
RmNpIVKH+IPP13TC2vsBWtaRQR6Rgb/AQbkjmARVeYmzQRBlxXgXjMRu3srEgqUmz2OYR87iHUbd
pg9fd9LA5IsFtdbrRU2MxChdE1mH6QKYZjrZaHERm0YwhR6cEKi5xfxhN+7xtCsCiv+yyMT6MP0G
86bmbLvXewtO0zKEPPSKzJT0YdpjljysmBuIGXOcwQK6isvHvSZugXfeWpfYRnuBtoLZFPRMjhtD
31qb/ZgL6/ddknAHq0sbGVXMxKjpsfyVNrkopb4cXsfE+chepO40HR3dFIhS8fibY+G4rCxW8kLO
iLW3v0oCHHG2iGFI1JKRmYE+bOAmeZpo9qlRj+ZfMZ0PxL+BQgXd9wZz9YqdsR5TL3Hbqw96NeFk
WibRkoJRnfRKoMSFpeQp+1j4Gsl/LBNuZ4nhqF9IeUsHyEEfQo/XlgrRPUhPvgOWiaLi9lXxtqVz
nORyzLVaQrhEUsiuqKov3UFyv78cxf5rTnEFpZMdmSzdi20qYxCsac/w6aYqPF/nNG4aVdGa7lWW
O4CvlI6a5CiRN8kpe/AEWzHZQ/ZWOIIg9BPFMroCq9WoU5y2TyJ52c5ZXzdNRJigzk0kkgA/AGRB
EC8Q8ipdIogkN9q7osaZV6sTRUuqcu0mcZP/YTLnGa2I9/fCwFF5EX9trPCFPVktn+MygacQvmLN
2SUg1efQljPKpcDOz3QziDd/ufGlo5pUq9LBtLNxkuGLSDAwLEGD6xEnBgHSoOsJM/lpGr6/9L1A
NPcb4BIwuz4SYk0KHxjQjRuaTFJkVVceoTv96yf+UjqmkXp7rZ6Ly3ZFyjmnnoa4xzxriyQOyyCl
fBKxvRDXwNBK3Y6szj+4gKsyeipPfeIUxW9fLAiLJD5SFm7w3Ou+EuHeYK92ZAMuuz1Q6wlJnTqF
8PW5JkvtNxpTP7OIIs58UnIsH+prpuzgpFxWkMCUH2a3ndk8Dnogbv5t12Q8jB9UIL8KcvrySOX1
MlcAQY036EQKq3I6IcvvZ6OaMb9Tj++410vFppQu4WFT13NVnwc/D6QiICdcVOj3yK6OZ3wCv+1H
PeijkL5GNpftOD9uQVv1+U6ohRcVgduZ0c4ty9YyOhernAKgf2tHiJKird6+Cf7qvLKUhu+ZTm6c
s23lUks7J86fnycruygW79FuLAYUgn9FAceUdPr8ygCnTSiEoY+aHFBWIaQ79QYrPruEUNvNEgPR
ssU1zIgUxejJLP7iZABmYUM1ypYkJi5NzBADIASgKSHvDoPv7hf0RAl4Qb5K7dWBt+wNorXRiSzF
k7S0gxTDkqSy34PH0+JXb2rk7EBg6u+G05acELvWRuQ1psaCxfXxlX1qR728ro2IkkYQOHxtjJ44
vPrl6Ugb25SS9Z066WCo7VMOsyJ4JzwNbG1W4Nh9qKNfjfYyFzd/CUec9le8P3ap+w2XjNw9lMNc
1p42EBW3Jxn8IN/WwsA9Tg1lcJV59hBKC2yuneQViAbAIw4+SYdFcE7wrYcIal9m1+yvwHcW6d7O
j01z6uK3c+JUvYTf7np8s2pzapPHZE8FJ3T5MHeg62jWOE87PrvPZ5L7t6uVlGMhkzWc0SIGviTc
1LQyG2dGXDymFgPgYyEtgXGUF8oPe7A+GXesDd7Z/XkXitWvLBNNaRBOfPgir61xRAJXJmF0IDPK
HXsCPgPzWZ1tPUsOgkKBfoueaf3KL0mSbpcElc+3IF2YKK5MxCEwqnYBu7Lol5+I/U2YiS0INdQ3
yS7ZGLB8eL8/zrWOzL50scXnVewyL4fn09pEmkfrme8mRQDZQAIDr/I3sbQ489kAZTFBQm5/KJin
y4j7R9lx/WUg29j1Todwf1MbLh4IgEnZQNwTRNgCZhv/qsYIcZ0NvNK2zeBWlmBpzwRmh2rZZ8J7
GDwB2xv7OmhxtVRp5eegJ1WlUv+XkVN3EeQC7WegkKKWlAFTtyt4B97r1sWF2jPzcbDzr8oSTd/S
m4MvaaZsG570ffptOuexPKiETb2mCLvevY6e8kF4Y5LD4EhbKSmLGL4s6/HSwTVL0qgU3YW7yNEG
yYiUUMSVHV3MLcWCNsfdQrWH1RkVC2tHNRfxYIaXu6rBJgPfjdmCIzarS67PhsuNfybdS8avCk5d
7wTwj0sLRn+UR8L0/z5NDJLwPAzh/dV3RbevVAvE2L3I+cMMw6R2VtdhUpaCVcrUEgIxcNQyoFDo
CR9g0iecxyI4OuP8r3mly4sMO8wIc9q+nY9Lg+KJeFtQxWJ2bju7eQ2mzzHkhLmugOXndIHoEe+M
qp+KXA9kWaeeaRRGldQLNiFVjvhSPoJSbA5jayFEvt7jZWVADh2NQa7NuFSJBXfLcn6eeKvChO42
l8VLDzMMnE06/BQ4IIPhgPybLzLbygk+FNfjGWgtNYuPLZOthWmq11zV5NNH+6HAjpbZq74kj5YN
3vPmfRObI/1U9ljPzRe9B+OmNBum1s+g77Hb7RQ98YMJFXH/Yv9YrQGSroICezeutNbpenrAkTTs
xYZWvLa4k2WRM63YO81nU2l3jc3jaHDOgRKOpEpyDi9staDu2W7LaWmOU3QJ6sd2otx/mq+zar5u
QkJkVXjC98G6u4LltneG/rSnU9KBcHhVZibchYgKXA7oYavM3zHdR8ZDILboM+Kmit+v+G5Q1Zl0
F/DJVj2oJd1LSW5Rfks+CFcURH2q0fufMrwRLVJtYmiOVxK6oq5AENcgKjqJUTRzQiiFJ3E9lB/+
1vjqMUW8rHxKUgwYjPBhtqSv1RWMnZRnqLC0L7PjlMm4i/9Je/jkEHz4varGC93GPxsTK7Sp9HOi
luEzaytJ9vUV5sGjDR1YNet8vTXlzXh8R3iHjRYL4s+3fHEZmqk4DmxouXl5rzKSbWNsnAPep4jJ
YcvAyAdRddhM8Iptd2bGnHoTIEHfMxiRMzGWoFI6UAfBGHYnCTA+5r3ktbbEyCCAVl8yDHncnoYd
JPIB71GwgRW4FFGJIT7jhl8p64VWW0TEWSNAija6ipuaqD3IhguOr9CEoKuZipKld28fPsYljrF+
/HiME7gdwYevXnA1TUvpfTYPJM9TtOP6fDNpkneDhdgzRCDLPpxHkAuRBezfJ8C+wz6IKGVjU+JI
k7pu46uvsRM56jpt/aetk27ocSzKL2R6QXPqwHePGdSLRFkwfXel4XkhSSH0wKnnDRGsJc/81CAa
GqllVYkU2ajeJ+9ciYQ7usXXyxoAxZYrKtnWHBmXcgQwz7PH2QBpRAhQ4V5P9Czl/hxBSf2tatK7
Pcylf0RM/JaTiizJxgp5p/71bfAWQZllq2sBCA0GsiEgbjwUNsJ7o/2CICnQyGPYkdeKE90M4CVT
3XP9urh9fKZTWqfkTy4lNnXxY8nN8XnOScmdG5xzmHfPXk5Gdd8EHA7WayRs8rNyf9inaklHP0nC
0yFoLUU3MUn7aihmnKGqJ+wIEj3PniZwLIWp39LssfzxgBYdN4s3APGqBWbHj1gd7KaHmKyPNxQw
Icn79w/bmZe8o9L5RL4cN646WK1rg09r95bi+GE9OQjypm5LEgX1H8rSYRwg859xYfCRLqMLjOg2
4u4nx4vUPx9uch4tSX0nbMUswZnowF5CgmbJJ+VjdzdZJq6ZKBo0lrNBvEOaZLb5F0uPDsN0EoI1
LeIO7pOkiWX2IBkAQE3BskH8ym3z4BWGsY8eg83gsxdGXE7Y6tLLgCsFphVMk8C4QyYSAMQLz7wL
XIqau8eFH0M3yhru4CpYANaHOYS2N71Au/rzAPi3XhbiVrOY15ODIqBcasl/u0EI/CDLkAcGJtm0
lS9KSXemSQyLTjca6cT0mY8Hmv3vkQZYgkL+PoZTFtbLmWgnBKG0FmAQ7+MJDUfGwV+kBZ+iR32C
M5k5SaH/58wvNKtrlTvQi8eE/+zXavYD+puSoT8QNx77dBk4oHWX7CYWKkXlhxhsXyxPxsz6K3ly
8R7IXi9JpexOyJg0DIsONBnRgLT7tOjn5Jg0H5L86xm17uEOES5z3jFdk8ilTJzFsBMPTXkeMbqw
ergEHMKZwE5qYwrpfnSE9JuGkweF+ApZc/CHLdSDtKoLtkvn5PpzchU54nxRxtwuob4yQgN5XRmU
E5uTrd7Z+dquNIhtuiU4EvumO57pJZIDbqTgouphao6Pc14MvLd17Xp7Tm0hEjGzdLg9ifWow1at
0yYywyH2b2SuL3m58KP7qy/XVwK6dO8ALt6O8/O1FuBiE36h6f+FMMu4l+6/q/eI7Gh2nfS8FYBl
gadnb6X0PLT//XlV5VozpYJxwrCQKeRwQEXH7av0P0B6/HEPomIDJx9Hi75DhDjHmlsT+IHS1zXQ
I11pX196+3zeVqP7boxqxjwjRCS75zuxk0t7c2E7l+vHUxiqmppcpsW5Z4gBbjxUM0aP+yVkk3dk
HoLOaOm810IyVQFgdWhgf2rqKMqlNQcCKUA1MScXidMqnrflTWRv1Y34ZuqN753kUzXa9Vg8oHPi
1F5k2blvR19CTG1bCxAgT41770IAyQJKUc6IifRUpsqWb2PvAQAHXMaDDzWH94jrjQLg2NQ7KLpU
0S328ggLMJuFcbQiz4eXpnm8dP+ocqo/1hFUpUwDuZkzXr47brOAcJvsF5ja3gyF+/3I49uen2NY
Dzsmktcy8JR6acr8jOVdGfYPasbUSbW2F99tW41uxgGcT+jSMzHuzyaAiJEUWcHKfkMDdRehd3p2
RhQtB3/jhSEHteL9X57PGLg9n5q7PblJwXyesUTEDLWI6BuMUTOEyLE70gYg2Sf1k2OXENtaiqBm
YWlaAV5xy9dWG2PFUJ9d/0c0FENiNyqLM3XG3TaeGrD7c/LjL0pWGYhxWm94m0TU5gHBlA6k+XIU
sx03h9z1yrl+8YQ3SD6fE+pqx4ffiCa3KXzYwB/UADIaR0kaWgiYXvZs362neCyPPqTNAzjFf9pN
OO1KuP3uZhOU/YZ4GFJzlKvyuDGAkyNtQsH2xlwkoRERkbynv6auo5XIQ+ztluYWA+hQ8FXTwJg/
foIE5hrtZ4EXrfAxTmdHysc2oKlWTfLGoyTEIg9eDZRHNgMUh5ExnzhbvwbGVufnqD78KQ9gCsUC
GvrKKIEC3dVesLsG9Lhkx6h2VDQeEIBohHami7hCpB7XA1aa8MeFf6iYm4eJq/driuvz11nC1OQe
GmUtONde63993VSzbnoGjFColS3pigYQrGsyzkNZmLtlNmtpKN7FrECv+Y5atTzJ1btmzYKNS9NP
K01Y9BhqhqzzTguj4Lh5H1lgrtFApcd8HXBIOSUDwWiAwjP4SLkf95GQsHjHO3W9awUsUQQ5O7sf
rD+7fO0CQaT6PDv8OrsC21Zpu4/pTUx6MlU6xaPvapBNz6owF73yjVbLmabxNcXiPuL0JLWq+0kd
rf+qmdeTOD85FtHxd5+nw8ua33kICGj6eUl8YJvOcT1UanCpJLeesTZmZvdxSiMwal+hlHRmxZG8
nc7Old3D4b8cVVFhTMP4FEBCf5e9nnjFmlVPGxPJ+xwFKsALFk4tp+aTR+TIiUi7jRhwG5DId058
Yy1rxl3yZOpjnv0wraTtOkjsS13HRxacl5PDKQnk+TQ/4E1HTpaE/tjtXnrK8jTP+K/qSzJkFBoN
wwtqTBPIBMn/e7sHOktWzaj7Sr4d6dKsWHmXTrJxDlKKqjZKdbJJqrl0Xqo68RSXGKXMvXwS9pUc
cnYoLwDhBVZC/HZUXG1DyuvhVVa3A3C7IIDyA1kIhnbwEdj1vAx5+yw3SilXToYYWnN1+gbCP3ad
nxqsM+hcjddChFii1dcJarSOdjqyjhmD6LhQB6/4SdesfJp6mQAdYNVIIez4TZ4K4eN4BZlZi0eL
ixOyb7SeZ4u194cL2wiWCKYwTetTKvPoD8pcXP9zzE/mu49bSmneTA7niC0FOpZxrXF2mmbtQYbG
bYF66JoFoO5uWa5UkEADg2aR3gl2CkaL3HNtKpgZ82sjWi01E87gQPFsg5v8Con9MhHMQ2B/WBX0
CJL39U0exIcFd/6FPgmJMXbgopmRFZzd2qdZNDJZJwCZBD084a+ubepVbZnUkxKuGrmHD9QYA8E/
4+eDcri0MBU8aYxL1tTN6V0ZnA5rBbUDfVCgKlurcAYC2Y92V/NC79bw33VSCDeefGqc/bRxcPeN
ZrSurILFj3ZKvxljNSU7mMkZbia4GhQ212PzF/Kfm1rZt5VgomOfjCWCNnHhf2n8pG6c5M66eiwC
tMQOIJ6ioj1hhhmr+2BbopTSShsK6TdZjGIMIdrqCschbylzMYgNfIE7bhfwZztjld5LNLOI269i
uOZT82zEzJFGXZRWmzeKn6BBCCfeWUzGwfXDdboErHc/J17bNRohOuWYXbm7DlL6v3P0wJbS/Ak7
3xRsPZYYJ2KEuKjndyAepjUA6fQ10zSu1X6yYXwRlQMDEz3E59iwX0iyiDQfv7LTTlyOIu1Y+GJs
TZfqSn/EBPL2SUfsBbOvaR4PAtFsR0navTAWqHHrIvwEECvH/Fkr8gkj8d2y4gFO3O+rlIrvF2ii
CXSa2azu92rJFIy+ADqjMytI3PCnLGypDX8mUWegMrZB7IsQ0VZg3oR10KHe32/LhXC9lWjBh1xc
IlF6qHwymjkbhO1DOmrgaZkl6n2I3waq5GFWAW4oZrpxfIhRbE9W4pbEWmBfhYDGaaQKAs9MfPpY
yITLaa7UCQJiKgL0EZSVNRFkKidrNKBVNkTsl11W1Jxcox6c5kpfeK4rW58s9EDtVF7o1MA2/lHE
ysm6M8B40bR/wtFoV0V3caO6C+C9RzVAb6AFjCLgutMZCsMn5YqR6HbkpeQ4roKstZw3KUXyvqqi
A81s7G2xAVJ/LiKnl1Mc7ub4IO5exqJKJICD9Pf6v0rDDu1fTHf8d7fwQvxcJhkPcKhKqEjLd1cm
CnzYapgUyJ5W+KavvGO74OQ2HJPmBfbuDK67cLda6ullEvcdrdCI7hEz4ljIbC42WwYS6kwViOwA
nfLQqivgSUR+RLzMlkUjTZ81+tYONf6Y/UyNiXt2avnQavJwLeMk/2h0HG4kjEhuHfj4DA2XGyUk
uHlTZ366aDsGR4dwAvDVhyg+/UP5r6pn9dV32w3JBEu84jCRSODmoKVKfvpXYAy4YY17pzEuMh0e
9Yf1mOnPPKocjiv768i7VbK8C52CjAvNV0lmulOUTGPjfNx+0jmo9MchEmx1tHyUbd347e/+Kim6
43Kde3in20kOskvCRWH/YT3ubfovx/WKaiKNaDy+iNnYpZS+vFj6+CcDOfqvx0rzTY7mQdzmPzw3
qWZwISwEUud9BEDWrin+j92AUrzzXUxw+rgnf0KWO49Z/hQP9uPOSzcBpx8G8ZAKH+31QCOpbO7W
0L8UsX+EXILsPZPdtYeyhjS0Rk30efAkTe/YGhq3lZHiB/+YfWKRo58P44aN4pM5EmysB1rLnkKJ
QBzPXq7gfnSS28EfJ7tBrDfn03cIzpPoDRULSz/OmYrivzRKUVUrwIfAKgalkanj+bHIeNkS3NM0
mcAI5ch+LFiJM0QDjQaoubzXVqQvUlR+sC4v5/drZ9AJ1LS/KNZ16wdYeKsP8w6e243AaoU7E/Yh
RxpY1drwk62z0bXWsJebQbPNuV5U1ue/gocyKLTAOAdtYvwKone5AeUY+73ge89CnKmGADiSiWeA
imDxkrmgslxJkFSXgoB1zFgF4sNazhKuUcw9McomCeDZAL/ZvZkUtAh9A3xgiOMwKpjK/sxZcwil
A+tNJmYFbkCGUmdxQqSm5cPmdQ7dzd8kra6X7TNyZsVvvQvpSGsrk414ecotiHD8Y+sNoNZ13BG6
gnQJaAXODHsj2cy/yfR8w7QgdED7yRVkOfPf+kzelkX6w22jWVNGt8Ikwsw6SIqgDBQGYXF0Udqv
Qrk8HgcL4SrluQSadLbzQXyPfN4KxhN67dEawAdJq2WKkVZhsAnlk2PGVOAIdtDaDKmr/F/r3D3P
M+PUO30PxyloP/zPBGzErKUykd3RScTBwmI0BB3to1FLr+mWEWtbNG1z3e0oBBdN1aVOPGTIMjTV
oUsN/i9eco8ZgBtAmAiuQC1diAFQEit1SwP++NkF4awDxwTyABItw41VaiQUQ6wUX0rwKkhFGFwn
vpH4jWf6EmHXk44RLfiiSaDu2FCdO4Xl8pz8dQgGr5zol2Z1fI629aYTpvnFVRkfK430qx/TC87w
omlF6BFiUo+1X9GRR8zY42ieZFhz8UadMvzWzphM9PQdi0glHrWxcd6aA9UoNu1gAQTVG18i/YFo
BXGJI4hudtENgArLZg2Y/nSlMhraSOrFheIWUVTSho4LTrcZQXyDgGb093NhTzfgw2nJY+GrtItV
8pk3RGtpOi1T7Y1xsDDHyzgVtEspNo1yIexxfcjettTepR7H36rgJVZKvIrD81EMMleLAWZE5PCb
3KgWj+DrzeWbsDpNZmj39jY5s9vVVgfJUbxelMmfN//DmY6psk72bOTRFmgEMS5gba4p6MoIdYpy
590DgHXsGIg28wXBe8fIotTmsQkAMx3u+3+K90KvZXeiknaQ0I3L/2wWgUxyxs+o5CIyEZLJfUUU
wXY5SNBucKjIuZcHtB/nV4tCCx3p+9MNj1rxmCR5R5EFnALUm82UImtJN04yCoN89irvmXJ1lUsl
+931RG+WwW4Y9lL9pGhzIfc/SV6305nezEwkd62xSJ5WWhCSwYOcZREPsx9VMJLNZQeI4yjBlEFv
t746e4EbA0j6n3RoDm1zh6BR3Anf/FcDWum7tTgdpYxxpowdWkRBlpFdw8fnKm+uwux9IM29d0tj
3XkzeA5Y5H8aJmMjUut92IIbiplubJ5XYSZzxFUIlWCpOMuWItTcySj83LXwvExFrwkc9JdfyQ5+
rU/7d01W4mlMhfkW6Nry8Ac9JmAPx02F/vByHhJOrXBb3Qj5o1TRPqG4gaOFbsSvUw8z3pXsV1Dm
hbzvd4jfuQ7O2s8kZDTSrnQ/XM0BkJ7pEXo0LdehGOYaO05BmDfk0TI8bu2LoK/Y0PT4fyIoIlEb
xkek+qnme95nLkqeFPZiHFjJrbhY2guWrYFnuotXsgyWk/Gn1ex/YwFPHW0nU9OS9ObbsL3yULkQ
hAU/nnTPDG62QPIy3wNIEmsEIbT9iksUrEZFEQ4RzK4QoSWyEXZILJEMHTY/lm3aOG/bn3oGMiiH
jH1Z5w2VqFjWl8sBD9+zvmcbR8JZCDMQK6H0ROnXq2aScFI0XSQY9iWhdOVQfTIy8EJI2loPbEmx
i9FidVX6EJJ4Yk3yG8x60le7UWQWpnpeAiTEzsEMkZ6op9wdF6ElCfp5TfAp6y59tMIaouF5FhCh
gHLdrD85bYy5XRX1XTiJhFw7MISwFBpE7UiewWkyvARSwtVwIcxCQFYpvgxfQDSCdkAA4wjoRd8o
J44YNgFVooxuOu2u4ogUAkSCNhzgPJN869wL4Nz5BpXqFfxjeHuQvommgArKZlCEnAWj5YakYDFD
nfRAQ6OGiLGIhkalVgvO8xGOAm6zQePTp9mpzw4B8UK/jUp45q8DXLE7vjoNsIj6Ds59ryS0YF3c
8ymEYwIwoig6hqlq+uKanlmw3pwil9Q3T+oByHzqUFlkSTIiCUNWjFYvZ4tcz7ffXGVHnF6lfk6l
nbpx0/6zxbHkPXurQjUMPcJygYubJK5so27tPeCtmqk23yDhXqqpFxlU4N2jeCTRkzjuxCuieate
GmbxjlqlCtZUntqlBpvAtRT5Terd8i6swWQAVGu57MF9vPfb6tTs65REo0q/lXJjknKc2z+BePXr
2IGGLLUYb2REFqF+89IyLaqhTGaViPQ3zaGnJqm9FDHzd4TpR/A81k1NeM8boXmzzHkqzCjIAzhl
OnmT/Hog6lfWo56F91isvTD0nUm3FemeTftHKN91NNnBALKtJhaD6DZPrUEc1vriou1WT0LGKPJo
74ION+kXo6RlX7WD1s6DzEKElJXjWXrGpew1UwpCTm7HaxRwdQmSyYRmpl6PiIneoMpypNB91uSM
bcNfXFqhvwz1lPSiG42bUkiZAZS43ZXL9oKuFUESshSaPneY0H9JGF+oNjpq4hTAeejuhaoob0nc
xu/l5TQOrTabyyKQrwXucm1ifAPsm77oTJ2nSBJeU0jl7MUChnC5WJ1ZKfl+K4qLqu0rj79ohE0V
Wq6f8KajABoyQYWEXnJ7eW3q99759tk5EkHLrejfW2ZdsVdVHdbltxi8Dg+sI5g+Zmh/CtH8YGpv
HQCMv3ms3Yp0xhy6kZFcK0uIe/rcpadsyijiO8bamN9SbXCcLWxJXS/M+oihDbjtwUaz8Ogm3pFm
Q4xDEpgQqsiAhzWn4Z36OuFyAwHii6wpezdsHYyrBOXRhr4rEONPE7g8eRuE+CCAm6K18mJvlqIH
H0mcj/mEcvIy2wjJdNmiZYSxx1bu5Pn+UvllCegvoCMutmnfhERCtPqCb/2Y7Ostqo+ixsUIb247
oPaRPaqxnuYjmEu6/a2eFGkn+CZsyNX/VCIEiuQgIXUW6S9Q2n3EwOKOhjIjn5qOupH8C0M3glMg
GvcFaUKWTc1b1s7W5Hqf5N5/SiJN0GUE9xWLSoQrfVQPUsA66bZqRP1i9Eymf8iQg7Ovq4j5yHph
QRBdVZDhhXR9K76XwWYQd/NsDmSXAnV8F/REmFDwlf7tRlzpCiVnwjxX1ECA4EU4fih2UDQbrvsv
EtPGWJwAHZsVflWpNi7M/U9751aEyAyNCIhbOTUBLY2r9vYddkrpd0KWEKIZQpwtKUeFGUCBKAni
nPu+ofsjWVnI7RVHabxS8xsM3+LPwVPgAajok8tOQMeuoUCtIF11m1Tzf99nr2eklbi2/5R+fGP7
aQl96ZGRvfmuGuvGeqcHBERvCDQH7iykG9K8ob4/WSsAe225CF13nFF+7Du+pEk3/sVWmQsziFGo
LUbpKqugE7itvOxpqHq06auWjQs0GTiDXoxBStbBjYABfKg42bPot97vc67KL4UXHuxm+WvZDsyA
XIhRsq6lhtljKQPwvGJ0Fm8yOQEy6/v1PDMz0LP77LRX5HvLOqK9LpECU64TQ643WRgl6OOdcsPA
huY34UKtD4MHAkeYLKabAtWpMszUGWWPwlaQ+BQyN3mkTbXhfpfPGKU7FlQvN2lp9Y/6jFyy4Da2
KlCQtaUmpL/QDInZBbFQwa0XTCUMgLIOnPqaElz1SXDwbbuMwhKFyF60TxegCGRRwldLPbmwYWru
tlk95qPtoUNd9ibuW5dRBr2wtImSqZX2xMZIQzB7yMoNqrnk3qf77/Z10jeVIg4VZDyaN7KIbRSu
XvS+ivf10AdyuEXmKpDv7PKJe+RfUyaPO0rjqS+EJwgTKXWZaJW0Z4dDTZveVlI6LRVyCKP8ONrv
j+i1JZv/4V1//Jwa2MkcXwnFcer0kNwdwnc3ROu8JJ9V9EjieHC9wZ36y+7LpQX2wwIIP9Rt0xuD
+6p+7d3cj64K5b35Ewa55FJVtIIt//H9YUtB+vP+xRcgvsaIjgEcOsx4vgb9bBXnx9jc3rD0A4Mf
V+wTwK+1veEDEKkdWPzJuPRq4MU8y7Hwrh+Qy/gVxDIyrHDCdVvEwps59XdEL+QXRSlwI2+O5Dzv
OUp7gb3tGUqcwcdsgntkJi/iz8aCTjdzY33m4xOA1gwKxKYqrVhxWp4ssI9GekGIrUDpIiJwDMi3
990zrczGv3sdxb7AAVGm8/8aTsUAZD2kpqoUlp5TMlslnSJiwNkVklii2ZKPziEkzzwqwVO5Glfk
m5iV2dU0SqkSdP0Kd7VWQikCZZtePfUDOEW8VbyQ+54p9oB5OPiRwuM1dv3ebUYuBLQUrP8uhANG
ykGeGvWIGTAgSKyPt8mTcaXhu6SmBjzkmRKCfwr0ghVqVuCcZHMrLhgm1E47rjRgfK6o44Y0bAMV
JIBsyWBcSWqcO1puWR2/f3D/5CGpnpmlEMMoFJHsDLHrxMlGjueYbsGGGZVyZLGjuXgMQN5mcVtk
9F4N1eiMFFXgnkd+7ZB3LDbqnndMP3/Gl0ajDCjUYEppZG9iW4cCnh/16RyXLTVvPxyphxi8xfb4
7CuQPyg+bGB4ROOpmPEHmDMVy8FWfIKU4SGAtPb9zjMrdK/lGqLrQipn3pAqhvDJGvAF032Ny8tZ
IIkYXzzKoP9ezB5Q4LB8ux0syx4BGB3Mqa2dIy1Lkjd+b4NaIMOefHBe6EKSYdjl1w2K8ewo7yrI
/h7pV0V9HfDFsSKwB4enLTujRwzLS1KGng2NQRuD2Z6fJp6mgsfFGDpYJKkfem8Ai3GHiY/96RCT
U2frRhsNslvvUGCvy5uKvjL35e+i9l0fHRuVbw9m7R3GIiYIcXrfB0KmNJJIlg0n6GwlN1hgBqES
AACPWz8JuEiUSrmvtTXLC98TWebqPnVn4Osjo+GJaiTnF/FcMJU9zipAf8mlaJgbkPEAk5aOn8Mt
0PunkK8gg79kM+5LQ7npVm44esoCgvqRSixGf7WqfmGm4Jl7d5wDGbIhO5gJConyFFolAZEa74Py
CGtnJo8YKmB74jO4icb+Ldz3kEgi2O5SQ6P/NhU4fGmRwwnafYdaUiRkMoccgJfj2Gyha5N/Jbhs
0uNg4LnWd0OVw1cfFPSpBqP0B1k9SBHkGjW/x0WaRzTCnbTA71nqMayBIoj2V0ygCatXE3s7MGCI
NROd1CathOMLI3nmx5lH7gEX9CZbH00KnGXg63p7fCqPevYOU2uk5VW8/0W60YBeb33SPA9AJstF
qL7WcEsP+mp+zelJVuq28UTRdoCYgHXnrnes7G7/SfuXmQIcZiEmE6NeF9M7gPpewwS9WL9q8CP7
ENHtbHnhdP3K8zdDrT2Ktx57Y1X+aAB3jXONGSdfFSFHUMY0J8XgSHPCW4tAkgpuAnPVigHgNTv7
SF5rSIvQ8/NDxLo7cHYA2E8ZSpDlC6lDaP+aBm/WplvKtqxwMJKe8c53KGSifG8PtfHgyUNhezfT
Q0ZLELfTwnBKJ1vw1LwjPm5gbMlYNPFBZRuFmUz2ajhJm5w4WtM0bQdp7yPW1lN8GWETY5wDr/ji
NsIxqSbJzHjoI19w6pK+aq2AVixI6YT5P3vT96G1o/b+Rt1QoCGTQLWdkOTuz+xY6i65PrCQ8pDN
RiRR6JZDWbM1XSXZSMva98jOcDYGjbD1IQyUKIxVhHdt7Zvo/rAomnKddP5LKJP1CQ3TtjbzKflf
Lwj2qLFFVhnHrUzUrYp6msA2yTfJd7VbhOr2twU92oLFIzgcPufIL2X6uxjhhItTg43Zx4LwrDfy
SgLmHZlD0m4MkpfvLP4u8hQLmhX+vvW/b0tsEXBv3VGU5zqJ2BUwCFtetqYdcYUgCCoDjCBSwi1F
5tmw68qLUah2k+iJqxmt3xPTgZIr1SsHejMVzAFcbXsxmRzr2vxGoI3dV8nbrNZ7EZrcKgBsoM7L
iFL4ZbOapozGAbpfdDe682siN1iKxbgfcOGW5y/cUGtOWA45Tm9B7QbKsgHBFKje7NhYs+52El9W
Jgatdz8Y15CwRgAYvGrWdoB1ed4Eo1KdDzfdVyC74cAFTyfItyb/AmaRBogKrrAQy0mARqJO5hiU
1d0vj8PgDKnic/gDvHx0yOZI/VPtoRvuU7mV6RHrkhY5HMcRWj/ylx2HCFLV5zWHrbj17aUO1BBJ
aKB1EQv4lCSmddbXiP5KgemlknxgAPDD1VWXLpfyj+Y/QdVGbQ24x9X+fxiHw/hUEy8gedAdae4d
QACawrrG1DgpomvCUSjGPa+rx3gxWIlw/udhQj1XrS7wJmiBh54i+GnCtA06OATXZ7MTU0H6T7dI
rYWizLohSLXaVMIPpr5ir12gTZc3NNhLTsgHb7pk0enxQEx1BiHQ3eEOBQw+nFTuLV6a50hCLfUx
B10j8yrFNV8xg0Xn+0mwFSFPWulS9gIFcL78Y68xt5KHZ/ymC05xKOfnOOhcxE97XX202ugOi6nX
fJRPuvomDE5ZB8OcMlqHRSMxFXutUNAv7gyoaFrVJPOQ1IU2eWpnX+soMfKWrJHSHWGyonJ00F5z
Recb8rjUmpjgbZ/O8+PIt5q5xsb+Wiki6eqFEBZ7FvbiVkPvqcBQLn4h2f+peGX7CyDbc7oXBvQN
3nwqrivkBwcYCW0mVZVHt9JWv9D9J/Y/P7+HNp4lwPOoSWh+hUbSUrDBWrgHPcRMrDF5RpXLPba5
vn97vFwouz2HzplqDeyzxUnpF9AuE5xGCxihb9WJfj1220inNxKwdxH7SikQ+hGzKyM/l7fQ2rwn
+2D+sL12IZpzPFIXb8Qu9wJPTt0gIq88nsJvbLmZbcqlgkEF43+lWvlBJj/T0iMQfuF7l/EbouLk
qeGmp2ga5d58LI0EaO56ELM2nBr0l46IDsCwsR7Hi4zCkze32JpelCBALEVFBmlUPf80AcVYKWsG
k66HJXdSUyzi+m4nMPUKfq7A5f5VPlgF+fIh3NONc4x7ohSZ5BYLr45TOhfV6GfCwh0YMsvCVZOh
bIU+eE7cqw/lZEJeKFIIf7jFFtnOJSXBCjDKm3RxoG16S2bWf9Igg6vG0DoZKnLNIOhPLQ7I6Vdl
V6Qn/KvVGgx31LDBwcK85YedisIxYknG8uXX+lHf9jRO//q94ED8zzs4lgiYc33wYGIDX1Y3foAA
mEWVis8ACIoX48VDdOE9zhewhyfC+inyiV7oLqAXuzN9mavG9ohb0FdTTFTWKztaGF74KWcFlVz9
7wYch2P7iCpy98cjXt8oGIRG9VMGR2Ed/JL+KLc+DgGIdd+1kDahw9zVCvCBe7CZIZWVSV9IXc65
nzJUV2K9O0FQnBa8P5XH+y8q5zwCkxQLa6IvV2DBaT7yj+Flnsg3nDyTi1/JTW8/TpprevsfDoKJ
kJdjBIvwCrroztgN7qaRm+HmjWrCU5U599tmhS4LpGzVfMIh6pwJAy7ODmLybQ7FBOlt+vzbyVm3
fqK7ozdoeP97xYMVD94vdfIKm/48mywAQrAYNQH02DmEnNs8H2YjxYfdLHdICqxmUdnZEqPofjre
fnFpBrWqxHihrg3dnvS8d6juLbNsW7Eg24SabK0BknLkw93ERKzUIoBBGPkVtruDMPuyhp4hsn4I
sxEZ1oQ/k3kxGWJcY/4L9HZpk4AlR3JC6Ufhfx2eJAxi9JpE2x8mYF36Ab/Ei/uKRocsA0FfrulS
m1e0C51e/6r7VMBwYQ/IeXvqPBIVQqXWIDyNu1XKeiUREjw8ggLO/W5C+60UeSxXvNBn0O5TLBr9
dFivd+KDs7DJJIF0GPRPNbncr6JJ9Uwsx645muphxWHivgQIyUHEmh27COOYqREqx28XHA69cxEg
P3jGzazUe2PJfp7+23WSnQ+J5fn3IS6rm/5+8CLiPdbWJ2nBoP6Q9AOTlxQf2snEVEHrE74PuFJ1
zF6PeRGaSjq+h8U3GEZ3dBefdDnGfCb8KvtVGa2lTTGvnRx+hmDeLfu/UQeBTGBptzVjnXNxoIGE
U2IFSxUqQaKZSglmOJDkw+OndnWDW67HV6N/sLXo/ljGXTieMB8AV3t1XzmDYHANBAh3bq9SzMK4
iOKrkrWfXudvj4Dut83lggPCe7z/5lLqegDy7hFIwfYY0yv70ddgmLgOJbB1jowxmXgrovIqyDec
8fl4nxMwikp6Li/zKWQrVHIOptAC0jcNy5O3PO3hTrJXmGi1g1VdAaAqeYriRcmEJS9lTHwGPu1o
9NLO8ZnIMKeSHH2fuL79qWL+1UQGs1acaS+jCssiN7HHCWeDNJhkGXgkIhWBYlW2xlpwHpvfW06T
ZpEx0+71wHwIXkRiqqj6EU0oWYpZwOd5gn9mD/96YZ3M+DfN07BstcyT24NOlk9E28CIAMBDahhM
6WrpwTy0vt2GMXlFym9pu0DdI5NYfgInCjS9hwWcZJIWqXtCSVZ5W+sCVJZnsI85HhjxGA4hSQv+
icGsFskjQ8Nrs8bL9xQLuRe43UavIOk2ms7RuF8c/YMi64BVEz7gFc0xjsiAccejIPRlNTK0FhsK
S3kqeDNXeh0vYNsTrslTpukRNNH1zAJwCEB1q2Xgt3K2vZ9+hg16uGAxpQpSRoFBI4XnKkxzrg6N
XbYMA0B9Sfzg7TUT44XjIpRQ4v8bZM+2Eo/i7JjWmoySNgv6vUeMx6eFJ3OEOLUVjUUDUd03BV8m
00ie0ZFq4QnR0SeG7PI1EKaoWw1CdvGsq2CzjVM63TZaviiDt//5hLsF85GMy09Mr51SdaI3Xdz+
+98R6zDmO2hsija5sMoW64ppmr+2yB4e2U6PW7kvyt0A7cKyIEl9okTan1qL0jIezN8+BA5vGSPj
cetfwkfdDzm20bZ0QPahyWFiaUf7mQsIKijDOXTTq5zdHC74HUO5BExn/rUoPV4jnyPBzbpc5zjI
kcomabppNs6tpaWZBLR/mc0wLgjAoICgGj6vn6ScxtngEaUr3/F+8FyQ8o0l/lA9VofJcsE6wMCE
TV27HFqSscRDlkbTMXGdba1vkL0nryzC8sgttz3xWrVYy975DfaojxkdlECHJypwX9DqNpUrfONt
CHba5sxQKuvgEHS50cCXJPuDNhrIP/PMLkZXa8N7Ch1WXlOnpM+E/WzFuHLfl1XmtjT8k6CfrBqM
joOBBh+742g3v21dLf546ida/KQS2Ylndb2MHu7FNdQXC0p/cVc+z1M9bE2mKwD/klJZpWvnCEGc
nrUh7BUhf/yfbawZ+tqu6cgA7w/7MqeSEVsm4cF+oLdCuFvKuPwecOumAm3f/9zKV3BPQtZbLbyh
nIfNzsTz4uMc5Pz3NC48CV6YNxF1ySRB7qIzi8eKvrR2XJQ3Rtbpz0Z7iC3pTN9+phRu/SrTs8+F
3SrkJOU3kiAypyGL1vM56HNRHLuTrlSZ+Cmq83tLHfyHZdg1scqEgt3N592kR7dBvnFCPguyb76B
vKoCt76SPPuicvViKhpboFteKTxqFlpUiDwZV6Qj6Edpive0hWC6D/bsGvqmGeARA/am7jT0aaQn
nLB8sMbxnYUnzX0LT0EShLbVpqKFR0ZX5kRxJSESExQhacr5RxGH+1Lc3XJuquE8cK7NCGRoQkaq
RCTQQzYrYsJ3uRivYp0DKusSKKGrDKDH+QApiN9z0vJuYdPU+snnBnNewmVpZ7Se2rIb7Jo+fu91
TOsOS82nxJPe5ZxAFaS8oHCS76Bdsgd3DQLqKa99r42r05gpKzRcc/XEEQiV9wgChyjFfAtY00u1
Y2AwxUUgXX8lCnnrSPDR5lRVgUv2MqvsAexva2GNfVjjc+imd/8d/NRrjk0Yh653f5odCCHnFpH2
R3yF3YHpEMn2LP7XaJuLyDTbcyuADYkiV2tPecWJ1KcVYnnmXhF0pU3pIys4QFGJtKUlvbn6KT1D
o20m4nZsAOhc5aAl5vjffBkuV1Z5ECL7oKnwYi0oX5XpV55IA0Lbkgdl0KJHMoa3lK2jqjML4DkU
jlT1jwr3DWsnkc5prwcfNdCT7JK8ObytO7dyHJZr7aXZlhzF29UXitZEI76l19ExM1CEnLLVMakJ
uLroLFFQQy6gRKIFIbXW+FI7hBoUuEmm3uzsaNwSWuC7C+Gw7AeR2JME+GgVCLlCJOlmdlr1XURU
Jfh8PQy6t3OmW0SjItF6gbu6oaxIzk9zAVRvI22OygKrsF4nM9Mgo8ret3idYjl8P+uf9KkIU+Hg
t7D1hp5zjakHzoH0PByo7ZtlCa6M1vv1RrsVCD/KDZIamxdWIiekHn0zCnSBtdYAJyOBl901sKlG
CzrrUHSAcysdSIfsEr62thJsH2oRwxHDyQcuxfDVfqrY0TDqZyNuRHZHfC6JsCZM+XdUBFtdGMT/
k0ds5crkp3gN6EY2pZ64Qd3W+JfIh9wwPj7NZ6KShtHt+qUpVhDpfggOYwrDYDf8BZ9mqquNvUdd
l0P3fulf69SrPWmxzhmFBtnd4Q14Kq3YkP3FPXl790I6L0gjgJ7G7SEXH4ggmZqVsyEQ0dkUEG3L
ZPtquJKutmruqi2v88xg+KjAtfXcNojPI1KTC2O9JXRGWjYkL0F2RFWUezbDNN+CrOQkG0IYtGCB
PJfEXFNOxxMMmuASSmIsiFWYSKxVIdVfIBlpdgU3PAKG+Nq9Etwy8aJ80lE6HMZ4xX2Y7AzkDmSI
e1SCsuCrlRlDjehmasGE6zeEByK4dy+YP4N989kcGFDphtCYPkRDHwWLj4DJ0WiT3pBOKK3l3Spu
FbhuOQrOwIZOF0EfHp5edeSLrCAKJqoBDhzBPQqXqtUq4ZQQ4YfO00XLw0L0AcPtxOvI3Kug0hhk
W9pEtCYvFyUD1XNcbFZy+rEsL98evsmqPF1FWk+v8qIDET04RDiEqJOsS1H9A1k8Hd7WFX61ndsK
GsY/xFg0dd+YLqfkb4OkhAqfh7bpxs9rjxowEnrMgfwdxRTWROD3Wa+Q5C5fGbw0EXWKTduMjPJd
fhmXOMHPjfB1Conhnt1inu6Qh5bkRKCcr2cHAxPqnGQ30mzWGK0R9iCHq31jutWQvrIM9nuJrt5R
3wCldfhu0mRY1L6Q624dfUDQ2TLZPdQZkP28ViV6IL74JkJDYTEsdeUXhA/6d/nBLhd8kwtkUIr9
DHzmSpSQN1itM+nN9is/kkkNskoUcdnFxwDR/tWBoLLyoTMRgOZBLoyEUk1nvj1O9548YE2MNtAl
a9J1HLv/nh2X5+x4YVxxVQgq/JEvBScCeYkRYHe4Renb1QkvIkjzr0Q1ELthKFkpKWDJHXft4t8+
V0YnP6dI8hd8dSnvExwnqEh0XHgXUnw1ukxIdQDrw3nIDtWLs44L0pMqcG3Wl6ng44UwSdrWuZEn
V8SXu3gimJb2EaTDoOJRJS1uCa96+6N9qIzfoDGhAcdR5jrEU+uzEgB7ntPvPTlr62IYHRlFcUdf
6eEFVudNaqNR/BydpwrkGWCaK9wBuu3u4+HTCjLFRNSXxxFKDc3+dgCPcphVswgG06z/TBV2KP9B
enX1X+Cu344ZCxerOqGYmuDVBGzExF2zYoDdV2quw39oJ72iDLfDJZhl7z2dbzr1/zB8vRv26d67
0S3Pdur8Sh0f2YhDHkDYgllnhtZtzudfzGKYaOqzDyJ9CaXB5ogX+kjgWieG3Yg87a2XqDXkAJNi
ab2d7QzO8tvDruPodJGPccnCQbp8r+AxF1oRFYa8f14YgjUWJlboiYIH6qzuJG/8MmMGRMZAxy66
hQE2OQ1Zq6v019mhfSGQlDCFP+ZWIuWHirEkvCOJUI0g14Lk4QVynuZ9CmgaShbsfpDyAZUDfyba
i44O+xFr31mcyYdepLJ6a9JiUSxuLTcKFXH9dAeCgjEN6RY+TXbncUFDDw1e5sZ1d41w7tP3iowS
rjsOKbhHB38WHp2s2GDvyBUSi49PMGNfgbsXfD8p+cr0CvsZFgXLfQHToWl5pxy9UxyTtTaIB69b
Dqd4ECH+JeqjkdOncs4powuDTH/QmZIMMY7jB2gEDbfJ1xDq+jGEw0CxBWkgvnGbOA3ycKFXpNHY
843C17juKm8Kf+HmlT6hb0OfAVnKXgm0Ww9DKEqMNyDjHEIDuYd+VX//OBHy+VC9NUQg6E0yivpg
BHU8ozmwhnKMl9zvm0sivv8qwW72Tn2aIK6Bd2qWZu10ghBf7omB5C16LRs3IZFAyUwPKFINUtIP
V9gPti5D/b8C0vk7DIHH7HBe2oNQEn7Flh0Drm9htMrmOaLh52Xbuy8TMx8c/kDr48Wa/J3aOoBr
VXA8w8Ct9drFywr1U9XVG07FMnh0Vu4nsICIUM0ZwazLbRyvo2n+fOZ5yGrB9s+t5K9UOvrC6Ure
NE0ZCe2gWLr/me6C8jY3qgVF4I6r2TWq43lr1mHovNc1uepJiRA87r63RnT6gT400a5a5VZ6Ik+T
dLdprSBWPqdFiGohUyrK1uUF8e96zth2FOXZPS9g1EWwfHH3rn+SgK7IjwbB9HJjrAYeuDohjZ4P
wbaL6zvCLhQZivM/TORSSD0dEfAZiiqm+hKPnckiLn2X7Fuy5mTxgcczDVTzhmm1ZmOnQ+gXJAoh
y+u1akTcgKFsKpWYFCNGXrMrr8sxqVTXLq0W/4tAkjaJPhs4jiooo5uJV2ckzACxDe/0Fm15H5NF
40B5ml9cCEWz6QinO7/NruAfxlJnZ7AryhaIMA+ca+tNTDapW+6sP5ZVYjFWarmGxYmMenI5HbPA
lJVc9cvzVRfmZ+6GraK5zjk/LQnN5Zwp9+vXRjFQdDD9mKOuXRVMRHixsmF2PXBa4f9d1YDCilja
kHkFmgFj6Vn9hBrss+iqCZA/31d6G9qJyPgkkMEHjCPW2DsFzvM618+Klmn2wXzU+vLwCuz+sPyR
T6JO1lObBFxeL7yF2PUWLjJS+JnRm7IVBYEOa3NbVq7Q6DQzGhbjKeuO8XK7Fg+/RskPOWohN4kV
BaohakONhRYHjinYrs5GEn4DBMWgAbT2QInkALSyg3kBoKxv8LDtOPDaysFsWKbjVh0uKxKNVeYW
QSZYoBsAZXuNuGkR8Lgcx8Ws6b5bXc3B97D3JZT0ySPEpt62bU6/eFDTwic8R92zIRtX7hxshxQf
HewMD9G2zR+nSZXQ36K/Llf1QjYPX4VG0q5i7HG6MLD3k7kxvjWaaW7MC+Xorx7OCKOCEHS/xdhh
p/4l98bcN8a3vBIQe2mCCIVkKY/XpIMYfCN4j4oB0bzjSz8Dpue061eBp4aw9YahFr/AsI4cjCpA
clzPyIj1jH5i4BNhadV54mSPnjLNdpzOh+0gOH1QRJs0uLzxJGmD7gKIYlZqImzQavbNhY2hSA8P
wzIQlmto//nulltkgrRFQ67TeDEpzixxuFipuj4YvU2qfFFUQCEaQjvKPb6zRINbD8aRUAF0mQPD
XzOSju/af8tKrS6VYl6KfI7ItjkdVo8uIh44sYAVGGhQTNAC61CYLq10BP19xKKnVTX8WvSGZRAU
DuzY/tedSi92FClxRi3LwhHV+Z0gGACb51GNADcawczyr1FXgg6486EA/W1XylY9tnk8+cD8UadH
nF4xXxakX/OTFoH6F58bb+PbzO2NnLkPAXuEXUK3Pe7VCEJtVyEnaXOtxL2Xl7G7a1SL6bD2UUT7
F1Dpw7n+RQh42/BcgdsvnNAFN+xTUT+R36reaiHnOkjtQ0aayUh0w4trrBYKQdUrZIfhQuDWx5FB
xxefQQP2lxve/rHxgVv3myXxNLpBeNc8fxTH1/sed+o5fqJZD0+dIykiqBtTvRGTHdvCmFIMgfjm
egyLeiRsLilp3sT0XiSe+9w/LePiOfuXMh/HWa7exJZHoYbiMAm4B86oxXpb36W6wsyMH4dLmP/t
vRbAwIPRwOydilRGtnUNPpSvOYr5o5lMbI0lZnmHmgnDuM+Ibqtw3HbDM3iIziVutYxaW9IqWvtR
Tf0L8cPOrba1cPQnEh9SCHPIIyP9w+pamorU4y6lxDrTfh4et6mmkccoUwagkIm89EWbU8s7JDCR
iDOrXAAFbtcmVwPr1pI+XCrKt+K1Bx9rvHScNnp7li/gtdwdsxaiwpy4ur88ZuZs/9G5tnYqmLxc
qvNvMZYxiP0kJNujDu4Vuha8UtEp/LgRwHdCPss8ZM+sWtR5Fij6XxGNYtVAFKe5yDQZIFJFUu3v
yL6p/eQZKDQ6arjatlLOYn2BJz/gvh805R1JWZebXb4f67FDOCsgPzy67jOMgq1+gBXFaMtfCJym
lTcwf3Yo7TOwM74K7piLkneYptRkrw6AoKrZ1UXqZIAxKRqow7grWNPvN1iJoAxHyVctuUCSoQXh
WWi9RO5AO1is/MbopvVvRpU38yc8s+ihDwEQg4W/IJQ2ISRmcu+eSPjioxp7Runz/QD6euvE7XC9
iquGqNN1V47CbLjKNRCv+EMKAMzi0cloi9kwwNEBpK61Cy3uVANbOWY1WYRpkzGTZisC+wnMDmiX
AF9XwCQcDInMd8NdfEpVn/iWtBNQ8GEEsz6WIweQJquPGzhhjEfUfGTSBB8MkWxwLJ9dGnv9YAdr
A7QEx4WPaKKFhCjmI5YSZqwfGTE5llolOcO+fVMZfJHw+hONbN1APWhXOLRT/p8FLFHyP2G3f0Z0
e4lhMbl/5mLwrKUBnlMQSiWQxiIR3LjGb1OL88tf4nKqUV1ATlAaw/1Ub2Neiq39EVz6vRC9tXUo
kle2n8EDy8RbNL9QiMPTmy5+Ow3PH/Y+FMULIsHQKkmSKanFLWBSARdO7vpcwSjwDOCV/TjdZCxO
BnDhmWzRarUchK59h69t1Wdlc49CKjO0bMyOwEPSbnxKG5kVg2PISaCkqcynvDJO/QUGHdUcO2nz
L3SnTct1gS/cD9WGcfNiWa0qkOtEwAZzV++wGQbZony/26D4B1fvUOSlZZ3WgbjRDXqyAvatxZq8
rtDl2n7hhTrqdAIW7dCMXDLhpMR4662OyXWPcLEKdCc89e95Xqi9dwKX/pfZQ52dam3dBRezPgUd
9hO2ejlQYylfD9OGOy70us3+4qFZy8waQLa8xfb5pJfOLafsjZMZ5Vus+94c3vzmCaj1G9x8C8A+
L7ZHYrV257ZFBVIm0FunUKKY5kYaXikX9y3yggnSPrczRfvRGg5IUU7KXG4zhVsYHyMG98amMtyJ
Ouns7WuK1lbYmwmbIcToxgz5pm0JwbvJlHGSOkpPC5HIqcAybU1RynEnGSULflKyIg1pLBwjl37F
AeqZZOJb/v7Xn2/otaeUbKxrjarhJ65HL/ysOQxdf4V63MtuDoA9sCaCtz05c3ulsKDAnpMN3gH2
Hn/WRJav/ksZDU+Wmyqxhmn9y2H9YX3u2kxcAUECIT2F2wOOBpnbrLdHtWEbIlavLaEMaVtsJ/Rk
B8vY3hkceU0EwGnKjmCLk4/hYWsQ//3SLAP+ir1sgo7kbs4U6DC8tVu7xzgzp4dv+Bg0bnIDNRPc
mLfqBeWyaS06cT3JrQ2j7J9HgTi9fvzB69qHoPW96Og+eSkVuImhpDw8EeLKJYXFs4YsbNT0FdAS
1jd/7DyDOGJaID5Lx+8EosiUHF8sm9gkXGSXPoIP4qNQ5b9cJdOXFemiCMz6YmKc47qenEgcRKbJ
xOhKrIxyDNJVw8LpqzGEzySCglAEumaDa8Ayh/WxC6+jnMwEweGmj81axRtDzXI39A89mpjYa9n5
ZMVx7Oi0qI3XHPfSbbiM5mllX840Mf5Dg67UtW/qdPy2BPvHuqNqjFgXuVs2e5ig9BSOzzWUXu3K
u4PG3fsU6hCrhd/jorUNnmo/6hYShtuJUl4Er2biRy+ly7nbh+UeNKiOLBm9K3n1q8Zd1DJEbSHJ
aYctkLUgrwzoTrOxsuNk9K3X/vOe0hSwPVqJQpmAXo4kzRPp6ZJmFm6gZJxIIzOrzABpGAbFgFEx
38lzHa12ev3fbyblf33odIV6FeLrWqMGo5DSkSNz28LktqbkM9TB3dvfBzGVaDI7vIzoAyDAjzZB
gMVtAXafRZq+xw/fvSgrgb0z9FRX0X4L/is3yAvUVk3ceFNkXQnlT/H5BtiS0yi1RPVdjkzDVKhk
f6bPz4RwuHA/Xp1XPx9UY/Xw/7TouVM1g1WvwIhjp8CL0Wrkqgzfbw/3EHgCJj+yXsDAHl7qcV+F
tASiTTALQ/XjV3l0FMbfsju7ikP77w/tXzihveDrTyTCPK/u/XoLOxyBIZMVEuJsrCTYhh9zsYcb
ozTxVhoBFBlMe7A3w/6iPqIlq57RG7Chpc06/V+stlXviEdp/VgZpTcdx32R1L/WlqY7TnrD/Uim
h4PuiHdR1mLW4DAdxTEBMy2HtIFPLAWhEwcgWKtdvJLhiR4TRQijUidYJvtYio0VQecPtOPjJYqt
qW6hgQT+N3EX5jdlRreTu6QPiqDqeUuZqQeHQLYInMhy+6S1DibHShA3NZEOmXE4bt+1iAAMC/kH
f9LpVP8g495rbHlEZ4tl8K3KjHZLSPO16qXDUJsMYvaPcRGuPLy3o/YCaYnV/xHmObxPy3kVI5X1
H0UHWN99HCa6Sn/xsrUQqwFDgPTZNWrBxD5bJfVGvz8eWsTElM/bliD7sz5BU2W9YPZxkzM9/w5v
cI+HxJq/+DiHjcTfMpVb7MwsjD6vYrYQudhkKqMMKE2XgYVP9J5FkWUQvBlvtrE1GB22wrC/BUgP
1SDlSk+YvUwCkBN2q0onnbrHlqjXRw7qeFJDm2rGuoLuKaH5dazDIYWKGkT9LeYNwdC44vpY8GEo
bIk+fir6ho5OvGJ7gAAMIK0WodoFCpms7tUJV624MTPgOX7Ws/2Kt+LgkQK2voGW0mVJhLLp+3+K
mXHIvCGfHi9Y2cKj+ZpDXO/owiDChqgl/97VghJr5MCKQfWBOJIcuN9+AyxIBqe+kuIC7VkKY4dz
/MEzrmlwYYmVdFNjJAk44+Jj+3VgJoffH7q3svUWBr60J3Qb4drRIzRAongqW6irf7Z+PHE/ms72
fcEWuWHnypiSfN13JaqIZ2zIoEpCchZj4EVWZtX2tbIhVEU1brCwHTUJwQ4TeABsQur2zXLngi8Y
zWiNQscQhR+qeVKgQSf3+hBYoJXRAK/J35QB4xrP4fv2mYSPzPCI3twVVMlfcOxUY2LeIcoxySNH
PL5Oi7qinoRmyBShDmCUa0zB0FxJjXoo8sLHGOCTyIG1yRG3rqW4r3cgxAkNiTAMlp4su1G6ZIGb
AaNrevW9uU5jKfFuxKNZgtIS84ufqAibmKymgxwnpGDCgh+CQn2p+mSpLu2M1a3aGO5MRXyOmTIY
NO7ocRHAtQiyYw25Gg5Bqk0T4TNh40SIbi3Rp2pgd5objWCgeqPOJNhc2F4AdRDEEuezeLkpwubU
XrEkpSJtOBGwe65G36LFYl3/VKJhWLg6yRsVTO4CVKvenPXX5RsG1Umcyi9v2bThLYIYb22hUUbm
mzFv6TYEWSNx5rNnBkNvWJPGpozR94ma75+sDOXXOlDtTvjBEzGkQg/ym6TMEKeDN1WMftEO0kzY
hpNajFknT4tA1mLOCUHlD3j4pCB4ez4z6K2BJNyYx4h+fVrpRvQLy1pRax16jTzMoyR3tepPaQ89
Qhsg/H5WEAl6gb40ui2Ch9OXAHYWxkXcpLAM4mckMr2L71ywy6jIADFeIjKdOe0NpFZmmOOcqsop
PG/cZJLd+se5CrZRm5bbMGK2uojt0e3Bmn+OVNphwPEqQkVTY27BGqFjo9n11KIHI3xsOUVuT5jy
DJE6afbljFif+mnAFOKdfAU/jp/M/WwV0LgJ+xgvZmpyvzYCRKHprlh29sbkQhGl/HHJyL5mxoMS
RwEgKp0bS+ZUKwe8mKA9ukILsh6AbNmGJEC7Tdrl/EqHZJmES1MTLlLlJM2aE7Aiw8YfI/InJ8ml
nKY1PVu34vLQ9uL71i/px5cxMBD1tCo5xgxeYOh338G85yOUp2P6EAozunR1NEEEF5k+tSOAiIbU
cGoxKpWRaK7cUxfWW+pNhJBvZrfM+VESTiuM47yfTuflcx7z6cRI5C2uQ24IbH0ebA7KjJtWU7Zn
2vkiRRDRC+ME+Evq5p95KTofYdqaiVjK/Pvc9hYme6Ft1L6koPatwRs35AsWZO9d7e5Ngfmaektn
68pApbaXI9u80xJ57tGG22hHx/gxiwZvsU8RZmf2pj3oTB+yA6oM5vlxmBGg8lheJj5fLb7KDmbV
itejXYIvtn4o/rv5HQyTG6qwruqNPsAR2cE8LVJIE/nxRvK5h25xNxlryyXR0FefGXoaLcE/1eGG
1rbheZFIPgzTDvxXekkd8yTalFpbrYPtAEayEjJhfSrFsAgzxRVvFxfhjNyflZhM08waXNQfEVph
+XQ4wNX5JNXxkdshnEdFeDOjf6nQQeT/tcqJKvM6zqpglwfrphC6ksO2Bh087NxvsRFmbj8iT3VG
+hKcN/jljphaec2rRqHLPwFAvSSwyARXwVncsDwnKZdaSds93ApYYzskT+mkuJc1Fnngxx5s+RT/
Fkg+rDPd2buWknT0G4aUfR79x8wlTWSWinaiYk5huR6tPpVim/8mceauPt2d8Sj6F5VVq7PDIvKw
aQjGyS+Sc2somfdKsejNDhGhWbDrdGrXqo70u2lAslMDxuwnNYTm/Wy5auw9c2+OzBpK1JV896BD
1XuMSEtVc5H+vsFSVBvbf7Ts5ql/bC5cNAYWjysX+4EK8EiysbfK/H855M6lkiq5ojDvKh8Ngv3d
ZmEXlkHnTlXQrfo1fIQtM/sNGjgxYpkH+a8elflCF10hsZtnUsGtbt6ewPI/P9c1muc05umgTMKd
TC28gc6I0AcgjTeb8Fgi9juGudN+L/bhwK08IxS+pWRAXDTc2eD94gFQWfZgoislLKLDsHBupOui
2kUkdQSf3vE6NaZ6YXs9mIVk47UyHnStzaigm0CkOhfZW7OPfKfH22mXSh46qhFELbSr5/p9dOGb
uNHD+N/qnnI8jwXH1nN9PxMxQwKEJFihOGkW2S1MPwInsEvuwrsOeBKLhSc/O5hOR40V1I6rZDmL
hcbZLMOQT8F/gaefbbSLsN9S8byr1MFYukzjxIj5rGUYTZiqheDKDS0+8XzxpxXn94H/jZVPW1AD
6accB3ODbAjKmXV/BcXf1aHlclVWKBbZVGDxqmUCB68/Hii5zKCrzdMZGD0p89iaEUi4tCKPGStA
uFbtN/cNWC8P2dJQN7xBIoCMYSsg/bWj407jTSOIdzRNFuulcFuACuxwG7b1wstqFCMSBCicHJzP
nZfLBj0knPAthnTUAnDrXXt7Y2b8mfGK3IIJM3VEHYlRaB5J/dCPyzPczPMNJxKzwhf9yXMSd1UK
DXX5i/es7oXOSsPeUNBC6yPsaHIsWdWDKjTsdoXr0dZnfq33qUHpBNIyY4WBVx8VlN/fUQNCR6T3
HL4XLz8S7Zx1Oxlq2XjAvAQcOnE3rSxQr0Hd8P0hF/UChqo3eFkLuDSOcCH8nVEC3MWfFROGcUDn
uBzwBssei6UENBNKj8vFpdNkM8BYLNwINM7DZzdsESmqLAn90NWX4VzL79lPb0lZI5eQiSHVx/fe
1M5gb9r4Edf2D3TpJLFJmmfZzoECQROEI0vtYFi4PCTHOGN+BsxlWVJTeVn803YiKCa5KlOxMTc5
x2wrYWKSpSzXyf7m8bmh6Y3S76lbUWIZ4sai6JvU/tA9a6zU9gkG7HMpBXhV6rgXICrCuc//P2Xb
DLA442K8GhFAMte6nYfuSJTIshlNt4yLVHCk2wyEgnlZRuei/u0+dUbpjx0CetoYNiVl5Pvp3tTj
AV3Khu0oLK5ZEK03nktlZmrtIIm1q+vnjydsO3UTcYkzNDpZ6+bbz5ER2DjbyCBcCd1PKMO7MmxK
N4ydmTwSsxFH8AeQKGBIqP63G6yn0rX9JmSMYoLbEfA+ELRSnN/ACqwdZIprbIxq4l8qQbPF0G92
ASa4BI0qTzfz6+uY9qt4J3lRcH5L1vQsDAdvQAYuUfusODR5YMhDZky4FpAJkbQUZCddlXUc6aSb
jv1YKEyJXVT/Ixgpgrinqo0ayDe0Y9ZHjezqljKSR95Vsl17SfhR4cV0BIOvn+QnyT0wLQWXmE+j
CMg6e/geY0LrA2+GRNT0sIPCd7npxZASGoHbM36kBZ7ksuCOszZbL6ECqCiPGarm69wZLP/0NBsd
HpZU4WpgI8vnKP0LOXeK6B1CMrQy8KAmC6eM2aPuQEOnT22QmVSLXgdvD341vzsZNZ3Kl4BwQy+3
tDmyVRI6YyN0xzrscNFkO4j+pVNJuZIA9UYZ8SliXf47U6DZG2EPPlB+1kc1iv0wdbGMnBkKEo9e
++rnoPxqXw1Z9Ty0R2rsDwbZGvhT0z92abs8379dZI+BxrH1h5sfdyDMdk83tCyLGC06VR38wMuI
235AQQFivKOu0z+iI/7U3mfBPwaN+M9A7RmaOQ2e7kRxAwx+IhgkkIYn8MbnRHdrVslcAN1lfkWA
kcwBZ6YyXQrvVpxr4cEgkfXdOCJuIciN5fI3x7WcN7HIzEnOk7Ea2UUSZXHUWucLXvElshVab0sV
5aMPTV2f7/lzYtLu7WalHkXZNfExI/FwCFuq/iWJZWkVC4su+LcCcDu+9IfsR8hGJkKZ2heJzKgb
szXVJNLD1lw4B5nFbz+GzwDsZjU+G8EbBOYY/2j8KcEgPygY2QDQN8agbNxLe5rMWlWhhuajGBRg
L2d+xgbOcEPu9VFRZy8xTYUBbG5wR24rQDjSyOEYd2k9sOgB/z/Ur+Y1ctIn5drV9mtB3rZCUNKT
IkwaZUfDMgTkFzxpM7y+DOKNPLG0kIS2G7RSgUEFBf96eVlfxDGtlHqiiHQISH4Pzib1UetbZ805
js2SBjySetobA4YSdBiauTUVsK5pRHxmtLTHxLiMrVtU72HtnPsa8c3EgJS3HG8EAvzJUDyjFjER
dm5b5bEr4Eex7v1EK8EwfU7B9Qppp5Z+KYo4D2i2oiSIjf4qmHzsdi90ccxWpTYYH4Rvhiq1jno9
KF0bLvfy875/dgSW9kpR/ZZ+ADYvEzppuUt2R1HN7vPenQKGcYPtyQSNK9JkAd9BEi8JSLWZVfvk
YE5AilL7lUgtzPsrhjp0xXki3go+4sxRolxeMoTDqXJJchey9WEV2l3WkK/kGJ1v9T02Zczf6muD
wWv4/ALM5aP5pLukX9jLS2o0DjKa/VCM3ntnoQnvoEQ0pj/3mKXZcoFoVIxDk/gbFxJ5uJV4uECT
E2Js27g6g31mTcjqnbu1SKNLk5xC+HyIa0MFF2wGboTviDu7h8wlAJYW5HtxbtxxxiFwqKg6rjM6
ZStqsj3opPQvMZRtipWjmKOetGSCbPJS7oYiiylOXQVRbOOR4V9z/KvQM0Y9MmzadceTxVZsuTcY
CLXpiCGsLpZjkdQ+enEEdvaxFz4st1kmtC8kSZuwYGL0c9nFieU9Uy402pCt3Aloed4xU/jAX67p
EFWEforicz4ahwUMmyDnuHBvQYRjLT8cHzHZv3iczFBTu5k/osvrSNj8Vx6iu6I6EPT1XKCrU45f
YKv0n1kpxnnDZw2m5Gi8FFLeRMgkLmV5ILq0sp212iOzNlnD4Ca4DDRAr3isSsl1st6JFqmKhcfN
oqsJSUIeFWCR3nF9nRm47BamE+mqCBculzZwhOt3HnK9OWHiLa83PZrBhKpXpbit4JUyNvDl942J
ODb1ypgjfOY5nd12MZczOg+mpibGRKxF6pv09KvVvcH5WnhZ2F8YzjJohn+vgXzgAYbtyaALi8JN
ai4wLwnqimxbvPmqMNyiu4c6J3xlV/cryuXGQXwjSMGPehQ3Reksz4wcLAuJCxhbiH2tXVaytkXu
sF+xU3dDPhF7WIcGosQBtb40+/E3muB9sPJKYs0l9kErzEKq9VvUP3Qr33xsEYzCBSJfIBl40F8O
mX+5jeixAnh71p5MctmTZhc63KnARTgGRiBq1GjxmNjZCWb4OCNoscr9V1kucpyBgm10V/ZejJRH
Vr/g1wLr4E7Vovi5ym/F+XsrKCgl5+sicjoFoWyy98DP+jdU9pwZRNmZ6EFAr8AsLZT8RYOH/2Yv
zRKX+XZ76Rsk8ivdB/659//xRX8/icMRCOmgXccOUGbP8fxRB1Z/Gbi9esWPawiueE13X0JbNotK
3MfsotJjUSw0UDecz5ccwOGKafbTSC8z9cjMdok4/gaK73D1/84unYKMsVay5eEhhVzDtn6Lo7rS
jcKpgKmTNavc22WRlPa2TkBmG8Yd4cEmpMzC2bhMm6LDdyypQxudrD6LERYjvAnMKTN/2d9X4USi
sKO1GzEhAQU6EY/QfckZ49vgKXGTlCdYd54gQrfnnR6h14zMkL66z/ZCX+gG3vGNCy14LMImpSWm
+CDZ6WfAK3Yx6iPAnZ41EJSaDmJ4XqdOwAcQoEU7oUFLmxG4htOHyWDAczmjMvycDoEcT2Fi7W3X
4SzeZ3I+kfnVig8yQD1lQtIMLq8I/gogkcwQtqEL3/tkYVG0XX59fbE/ozucYUk+eTBKq1++v6Hf
gN6bqFVqlx8ru9Wp+OW1KwHQSpZGs/1VqkS/gujS+oR4+mXViNR1kdJ+6IPtB5EbJLzbLlm/1+Sa
o79FKTQ+ucTyZEdWe/oAQ5dxxQdlh+xBhogiBqgto49uKkMH0uSNqqyKqGpp3mHNW+X2NFGWCMjz
6mTY7g0yBxz3d2QqBuB7kQ3mNpw4fz7jUCZjoatpRPFMwfnEZBTl+fwZl4t5PNs/bHy9+Zq9X7Nz
+DhpwoF8tB5fZmkTNihzyuJVe3fDd5nLOGpyTmV43DNxsB4t1m6I8Gs6qIkQ0QPJ70XoUbAH5hPj
4P3KsfTQ6KubqNPELbC+NGm8xT08H5eeSBUEy77QvwvF8zP6X5sD+0JzRNUs5uGBm4X/5sRZmjJ6
kYBwF9k12MmyFWEtqjv87rpmqfhszPOxQYk5iO6ctQ8qnTfbnwWiprXVyMoWymzKOyUkSbvP4Oro
cflRpcclZWajMZdllBMKiJWPHpk7l7Mg57Tb9ZfRvau3VU3uioPulQRPxSo0R+bofxypdSwq3vgM
XjTiFNgAQYud9n0t/O9OQZmn6B0ZDTQMaHoFLBrq2LcOzYqRwMMkoJpYsFqXjrlctR0e+xHv4SsL
N5P7CAQlXxvuXEwUGbeEm6+RA2/3aq/5VnUfnxWQubVwMtTKlb2U1VHKPL1uZMWzYxgUS8PRVUSp
8rtT1xDiYEeUSc5OXx+UpQRJ+eX52oKYgGhO2C3KKEzdvipDtvmBbrIRC1lYmPzJjwSVwoMmEs0b
rZGxk+6oFSIZPr5CklrrzI/Pgh7NSnBU2YajRDeFvMrhl9ZkuiUFpUbRuYFWCPVDE/RtqHy6r/iI
Gv/P6GVPnyETq7xZgmOU95/yrTbe4HtB5KclgHCJztgiFik5c0PBN6xNJsvB2KUa6bQnEjiIhqB5
bAz1c2mOdPt2OmY7LeB5lyQwq/xZFhIzLncX4ZdnW/nghilBMfP/rQo+i9LH3G9BNDTNn4TlC4BK
FGuU1nqVdhM02ZzTsjcYMEz3BsTShXPX/h50VHlRR5ql9FC9j6kTtjQqVItCGBMn7fsGCnT7dTVo
PGxcBdD1uE6POSozFza3NTDGRHfvYKTIfZJyxqPDtZ/2TiGtRuuTHNqfaRkrQ6DA72Y8CPSkVhA7
STyoA/kVgU828bLN9H/YOmyX/077BakncrnImF7hPPdPRPkgrNfvm8/0V8RD3aPskggWnj1/ZfiT
5hKlvdrO1mZHLUNNRcm4zXj5GKv3ht+zHjFKshunMeEveRns65POo8OEBWUvQgJ+U5vAUZhL57xz
PTqAE+pGQ/dYHB3mx89NxX+xgg5UYw9nUFMChWBMHZDBQt+lvHFOs1yyJkI2CRv+93YW3KZqIZpb
wmJRE4GyuAAn/hOLjI0h+u9Fi+4U39orza5rqsz98T1qdIktVN9sWhjl/4/Ts23VTi1N0J20iteN
5Nx82ENZEnRxEw99uti30FlOb0h3hsp9XuvD3igt5OdzlKMQYztOzoEXK/dM9a/GD309GD3/4+/H
mSAN31QGCMnZh/e/LsFP1OaILeE2CPxwEoZ1WBupt+wKBHkTtNuIDePvPfM/v6JChxRNRAWlRB5e
GKHz5OH1ZPM+hyP4vqjzQinY7EvPkwjydbzYpPgsXUE0fzEWLmmIr+wDGta/Rehi6HrraxZCMn7z
3Id2queWMvVVzw1G/YnS2tp/i+rYLclfn+0r2OLiwLhZAQRT3N4sycdOiMmUd4DEOKVcr8foG9kp
Dkgm0pvKtDJwlSTOKiw7xZYqUDEWJOfg+TJzVyBtOpggdE+0nFlEwdy36KrDxXVlhisguQFk6c2S
b6LYYAq/GwutHyNZRAq2yL6l4FN6/Tk9wX/MESArNCYTPzhf4XCKXzPlR9+DUPl2xtsG1PKBFm2k
/s4tDJJoyl5ZSia74+lHcBOdFRdfcpVKJx+IhU3+CWGw4/OrFDxhLTEyN13pYzGmLGWB9N4TA/1Q
jPFzCuWqWgYa7J/OP+OesP3aeOeCp5R5VUkfLap2uV/0bep+nhyXuOhHiBFoyNoXdQ6LpSlT5bw7
S6xIqs+dURmsyuRuY/B2yCLQWKJAHTCzHemto/LFq3YxNIhWK18UmVRPnolsTkHu0t3s/VIZ3Aay
w491uRNNg5lO3X+F+JxFVJDOLIcGqys/OVIs7OG9r8Rh7FsCrJsKcvJy0YHRBlvOuJHkDSUfp8En
SBE9D9hUOMkt7Q+zKQz8TMVLJVzFpEysUDPdqoxd842/ygxFlYcT1NGgAaIp2yoVi1VdGmnAS4S9
jwExZi6KBJ6q+2JIsLMh9wtdMHAHDnQ2TKpaWTptn65guGiO3OcpKTQ8U9kNZPDJUcOZcMmjOG1o
yxODonpkun5d4zXFXqWGMgsF7nd+nVDha2CDaiu5aK2wK3cablFxBHn3sVKRcXT3Q3q+9adknSXA
eGzjKAn5r3M9sKCEuaRF2E4xiYAIoIAYmdb8kMm87pPS01KAieX7usAhqhULkPuJbkjpv/BppG3D
vbA/zaczfUmClIMcaH+OoHrTLlZrJdCT6g2b7uJlsQ51nV10QnY00xenRJ00Lj9+rRj996gWd0Zx
84fVrYXlvKbue6lFznXyq3/wK9FAe3HI/a+aqACcAAr0hIHn+IkcG1OWMGkDXdskXT+BnHOrHCiv
XcAtP/SyYCLKnJP7iMCutvUbZluoo+S1XRVwTg8GH6GZhgG8YzwB/MTxzeMAGGCnu8S8rsrLkNvT
CtxTL9VE+4G9Ie2/PU8vdBraT+KsJukuVoBbiyQkblPwxdtB1DCKQ4qyuOBiYKBlKbib0M7GtPj4
iVa2oUyou572jPzxY9ABy8LLJodLQtTaXsV3sDQKJPhEuJ0U5/bhFXF0HlGVO0NzYQXcsAu29Ttf
Mp2l9vdFl+ZjYm3wMRW2ibFaKbGULXb3VTlbuEFl7GSIaskiM89F209QLv7vP+xXeOT4hSHdla6J
54CKmPeDZUc/cwRN4SL10tGNdr2ocOujuqGpldQSJAhyNEm7kvUVFgZFv1GYmGcVVHfC080lla9i
j2DvJwfmC4o6WYwbY6v1EMT6NUBQgXWsPaPHLaTgqslnl9VtxUaxhWuxjx8qiOs0IvGYyYzlDHkj
SBRWJXRDIztz+SYAI/aOEBvel0zApu3wOUb7OeZl4sUb/jxtNw63nooyvjkYVO4Zr6LmJ8CyeUZQ
eL2OWQWbFyChIoihNFaEClJ2cyVMvMmBDpm6ktMxT+qMRs1zszTXYBqTFuiDSdlqcFPSj7WcEM/K
2B3lDAIV8g/QlsSkPHSLJySFJaKmwXaAXvkGpy3HrwCdYrhheVdqUue9nnc6CCQ/FLDzUAPnDLF9
G8qogkda+swMvld7TkxE5QAs27ZneiJodNeyMvwxDR+ZbbpvgsSUaoNKCnCB11TxJbRCUf03bTv1
yZh+68qM1b7eTaKriKI/2PdDxMdJmQgnThlU7RxtDKRX+3LOejt90ETBNCkMSK4BYq25OmhUOCIn
ra8J3fLpvlkb6u+KNYrMfbkTD1GOIF06gS97UrHPFNTmKTzpjnuNb0xq3xWK6M+dt1arVPNmBHOp
JmrKkloM5RXvQuISDupKBJ2PHpc9HgLs00Uwe0F1Dt8mlaxI+S/oawBQvW3uz6An0WauBD/FxtBT
5leZ0hAd+IrhgN7AWL8WRvER2INRN2ULKPTiBGk2c96ZGkmgieZkF1GfFp1rqk1c24zYNeuGYZn6
OGSfgputX9bnxzG8EFnnk5DmNPnzwC2vF8I7TPM60EXtBB4/U1nO7W/NqxT33yhxjNrtzlqI04vB
stUiLuyW2He6QxXyO2OuO0Wfk0+abbCibtSCsGCAL5ktQpuBDiJ9qlylXWm+Lrq4Q1NsICVQM1VF
IOpxiDhQo+yWOYTSMU/hqwcQ0xsMVSOhq2tuwxdFbXDi7D6s0gfIK1oaXZhNPR9mr7AJq42bd73c
qIuMaBRctuTo4TSQHFYEVSCvJ3oLeXn0G3X8tK0kcbYiYqOLk/65tophv3086gxnlG2VDAuvFMuA
+yUFyOPfxoJrL37wG/sohRHWQiurxjHV3juAIDTY73E9cNT7P+OGpN29Db2V10iuNQjBEi2Aizpw
XVfrZVUQcOzym1rKlaDfkDhKktzZu7SlsyXcs00d8q/AJi53R8T4Uh0okiO0FSjFLMoPGTDhZO9E
OdL8Cqpsv6tGm3IYD9Jkp7zJTlKEKu/sgGIG3sbg6YV1/RH0IS+C/pIJSD0OnlMKp1g8MyJT6O+z
YFExcvrp8JEluZOfMHQXoGPkrgXQI57ZiTINpHiC6QcuK2OA5mrmb3GKg4aSo8E/bdlQeGekEqXV
fmQQLVIcLEazmGxsG9/ZZP8cdbVky7fk6g0tmgh7Urj/XfzhR5gFBBB7MTsE2JdeqAi7Z2K2+mAR
GOH8c3lGJYtNVJe0e0MZfxOQud9Y5Aq/F1JCotly5Tw25iVGSHF44gP/dhmDYB9I73equMZvrsqF
1gqTnG6dpdyQJGyr0QiKDcxf2r/E8qN7AnU83/s4FIQTFhONNeA4pz+dnuEWlDJ9dI33+qzAnYLp
DQwzdYv6WC8cjx5VbFk5EFkVD4dl2o6MejEmVQpOw+5Tzi8g0CBRKwPk3gc3iy0TLJOCMQjvqZZm
ugju6x32amU3g4J36UX52jHu7V0fIIsgfe5lgSz6epnlR2fJz+8FHcFTEYkZG63pCv0YPgHSKpTB
mnAoVWbkpUDh49UYquyat8+rTGRmNcWecJ2Lti8uBnJezTpOWMVNNkm5xETTBZJFSQBOiAYagbsa
Mo9wVoZsSLDY8yELLldCJSmkUlL39QXEJH3oWMfI6XJmweZBCd1NAILX/c/kNARuBRoz5yGA5JcU
2qo9PaXDv9mKA8zF2Yl4nHqObwcqDnPWTGU/QprfoW570Nls3dqjzlBpijTChspHXQsD7bzphwny
F/0TpQBLWkHgysmifki8y1fJYKVCEfR75JJBTwWAaIZApoScoBFSznjIpyMIi5LfpHmtsMktHMBw
t/ay1QmhwXRiZAE0yda9E9ysd+GJi6SFjud6DXACKRNr5B9i0tUcKz0OsGlsRkchAydJZ8iw6MYy
3PaSI/1x84JmXG0skpvTDTMh8RLS//GavSjR0p1DADwejyv7UoFuUjVkUoZJatIXMav4rInl+jPU
QMGzIGqgvZFaLGgNlQSuVLxqK++YmUF0Iuui0nUkFF5jSoHzc/MDIGhgFIu0uaD17m1GAyfvnibS
GoHmAN1R7H15EEtNmB+pmH1YTJ1xU4Gs4IUMteynC7qFt7Z34NraHSF+FFz5PIlvtjz9LklX53F8
1sf/zg1lAvI0ia0Y2gWpGYL24ojDwGVXUQBA3V94vCXzIH0yWJQXAEe28oePjxN8UwsTHrtwo6Hh
8EXt6y7duQOOppGEFC5/uOpjasYYEfGehv4Osxab3X/QzhPfCs9Sj5Ilr9pX98ulRrCV2twh4JCP
dBanMRuAZslpwVyq32xtl7A2Fsaow2ZhrKx6UaxbILGrqexY6pNHn5HR+we6MlkuTgYkb/p+z4+Q
m2C10qf87QKsoCzSUt4g3a4OvWtCAAS1P9jJC/T8hmluzQuRmBsbq4UpWnUGW4nKo3nHI0adWfQ9
lQtM4bp+oW/IVqcWl38M2rV2vKE+Zk55Ez42HIotNwBEH4IYxAYIPbGbLLTopKaE2Ek+YAeWSBve
fWbBOd7tcI92WikfIrltGlT4SBEsjKaOB8tIAj5vEj2DjgzGViSQR8xHOECI17WXVq7MqyrcFuGS
JvJsNFOcC1wHBtdoS51+y3tUyExiVMu18NNVuLxbxGQ6W1wiKzpmfgy998TosQ6vVa0tFiFlJC45
yrVVT037pKsONXCFNcm6hbSr6XsSl8dt/nN2nni+WQc72cb6gIvHS9D9J1LhnyPm6Hp7cF+JIzF/
Cv195vF1gEVmk2a8GqTCs6Cwhvd4sskSOpSRlDC5XBCvttM/5l/hc9V9n+8a0SNsAF7DgUayF6PD
Bq6aTWGpjCwDyNubgo6YTdKcnUgKD98yZEK+n488BNZJ/v9g+bAt5bV3bzR0HTbN6HxqKtVzVGVR
slMflpVRl/hIcLFTiIoXSHcuRd1q6Fk2BPInMTgqyt+PFsjWB5NSiXSaZZgix3Ni0+5ZQrBSMPFf
4hoTQw0NtyV8P9Iateh1+jlTE5ZTikJQjAyCqKR55K3Z+rhtMShST7j5TkpBt5fqcUn3A/YIJAQs
neMOCvPJqvwZfRTgpeTjdGrZqeDRVy/qL8q+io+OinIlPax28SgAchvYqHkTGROmYTJPWw5yvQNx
ihSelbP5+7JsQWNiAaCTHedkl8e8Rpy6H15CCcVNWuWm3Bf9Q3CJeu/ar//r2jDNZYD0P/NTkklF
aC7jdMyrEthzEHd92nbjaKgE55vQN7C/1aE2HM18dfNRvMuJHVCZshGaGWOC0Mwi6V6KsHbL/PDT
ek9ayiCnmfRzj4CM3ohh+XAUsgkg48il+7dcN8DV18K6I1Sw74WyKEEQgtvCQrpdEpMQWyMQal/p
SaDWQa3i9Hnly/CAtBhGHMo7DcYnf2ZV9lUBYz1MQStdSYfYPCEAxt3HmI8nLlXbJa0xXjzT/oC/
LRGxMiviAk/9ZQC7+qPDuGCSNxbWr+/eYUGS81I8scGYshBpAhSQbm30F47VHXbFSWwp4Y03AZdB
obYpaBNB/zvxmlsthhJCj2pzRNuzq+L8H8jjZx/h/ZRGolWkDJrrf9NDI/odX1rwU0SHztfHtWn7
RDQABT1VHVFBRq7UAJYVxolScUbKn2vwyIiWLpLJZyVTQ7AtcY5L+rB1PYfPkShmJiBHM7wYwunW
OnmCfqEYO9bUctjBd1jvKfvhrA7sGY7tILIoYztVpIPe+JCry/lhbkbVhPtldlT6H4QR7h5aiXIZ
ul41ZZmH4kXi6/dHNkQrhAoyazn3tMot4WYb0Vz7phPuhitX2lxs8DAuaw+9VT5pOzudZNc3fGpn
qgaAsb3sPx2h4UmuaOg/ZZruktk0XrOWQOJufM25BFdcCOPlKMFU6SLK56+r4m8eShs4/Zfr5SPm
1P6GNFUyLPBhTp1x50W/UihlmfbXch7tB66hyh760TYbZqlrJYhwxLE0s+uwHxT0WN1vmwHOOB2O
ALj4I3Z9yWPLbR3IA+j48YFH/Q0u7PQvWZossVT9QS20skeIaW58Wi+scJ7yzLTqJK7DK6zhBPp+
Al8mAcICuPyWWIQDniHGPS6uSHJYTD5crVY72ALM8kXg2ZG+vK+qyJbIilIT7nJdeV9138sYMvr0
0W3Jx2ZuTiMABhtRCrpl8yYkdlqNqP9mDzIfHpYaxHc0yrTzK8bqZi+q5WWlvYZoMXYRty/6M/w7
KoUM/6f3L9IYpoxkLRyouqhWnulRMJ8BAjGtmMu5yhe3AbXe7j8uIo+isqtb24HURPMdck5ym36A
yRaUeCbkyjiCPI9G14kDk72pQQJy0hM5M1ynwyCg1OK4C3gaGarH48+ekIge9c4HrkNehWLlgzdI
ierjruuP7gfVr1eSv0+Q00aECkiKQBqU6Z3ooTyYOhghDCDoFEQRWvp1WPzg/qP9pJ29HZJifV1a
Pkj19YT2lK9aXseHkSTnlQxcmrSV09uXC25nU/JPXNhc82wE+5WpwKIOAZBAS+ZUucitv/7RsQUw
OKseKAJbq10LlydImA3FhjDukVAIeNbkHPIsm1InYJ+Ml2dI7Vta7vG+Hv6VppDmPrInILdGTkyQ
2ga9xjZerhLlO7SAA4nRhgAuR9hhNTyXUprjKYw2TznLmeIxrWtkf9YVggiHLUgvNIu0zAkx4+Gh
NU6KxZZirQ0C3lVIq/zAjdcTN4oohUvs0L6DrQge4R2HpTGfXdQstYtU5FxPvK9xbLwRcBfHC4Gk
AHykTcjOQK7Gjj9dq6jOfskm4XA0JnSjeZYb28ifxqtAaB+sKyWGuPQsDN2xwTqdZFX5En6F8KfC
sqYeHiexNdgeqCvSB/WdhBTZob2yBYR0I/+Hsi23XDzSSr1cvYv/OymykrFx500qhW3TqAXuyZ5m
QFRkHKS3Iv7mbTAfXlJk1piMDm43VnQA8iBITn08P68VXx7Xf+MYDdpd17c0B84rY1w9Rtn3ALxo
TskivtAbEfM+xpqAvEcx8Ro5QMJNG6lLKDgj3FQE6LGP4SB3UN4K06cUvv4Qj7PaQ1pVXxB+1WQ9
Lg8OoZ3bAdw4e7HtLjIk1uAMM4rzinvP5XlKsh8WKH3oE31gd1vAWshWY4ViCP5AU2wAzZoFLnzN
wdFuJ0ewqfN6HcSUKPKkKnlBPnZWe2vTSo5R1zmblqxm9btMpqr1tH9UsiEe3KswlMKBSmgKCgrm
6rXlgodRp0HBObfa3Urg84bPdMBiAlgjc8883TgLMG8f79lbN9aVUNwq3Jb2lFrwt1WtG+g5eB0F
KbSNo1afxwIF38lcronIkwo3PXcmcwLRS/oNsEgBviE/JJVirRUhQdqk2v447C1bVK7y5POL8Gna
YCKzfchEuYAvfe7B2RRrHiag5G0hKaP2SQ1+DBTThBF2osEfh7T7EwA6dyDtSUaAwT3GI7uonhqr
6RR2VRkCrDGTBpufl1SbbRJIczcnnBLtMaD3mF0BxCHFILKSbNjIhaF/jXouLqxa+opfHKGjJdzc
h6iXd84zN8RFHvfTug4TuCnzqRXFdXE3wb1Re3O6wAV2coqDt+EMs0pAYsyaTLKeaTYNJPyNvkLA
e8tN9FwNaq3j5zPUM2FxujulqijM1QEZPljxiqoeS6dDLEbCm7ZVMxvFS3CTkgYcYRp9Hky6GQrF
3/bZTZm8k3APnzK0WSYfLYgcyYLAIeQ9m2G+ynFZtLG2WTb3mUJBY3K/wDIz0VoOnw/OpA09e5Qp
HgQ6g6K0HTP4z0Dq+Udv6CJ7KewQbnSAF8aLVVkVYybKAHS7g5nC6LC+nAVOGZFh29XAm4RRMu/m
ye95GMhE4nwS1qBWEauqG9F9DQ1at7kGd0B8/qlRx369AjgW+ljj5nRNhD00Mj9uP8/v3izEqTb/
lL0lRbEGS2t8v70l+wR+Je9oEKdyn1ivNXcqbFD5meKzXweM6m4ARHvn5acjJ1g0xMoMyx6OM0qk
PNC2UWqO6BblOzBZ1+waMc0l4zHZZP9zLRnh1Uqi+jEirW9kkktLookcHAeDFXePuHP+rWvrUcwi
0oCVxtEvM8NdE2CELeEHIxDgucufOEAQ0RGlpQY4ncI4TwbISZR/UZXdV3vOULrkW7YXjb8DXd2A
L84ytbu1Hv9cYT2WIKTv7QNtrw0KLGLWq8U/qK1QQgAphtq3u5+1WUDynHry932w6feRVNzOk13J
U5KJvM4eZzYg8dlsf9jpfCy6x16raMknNZ+mE3xtSEGCMy99Q71Ld3j2bnZq/I72kRe/5Kcvirpo
FNv4GE/DxyKTvLO8lZU2ETKdfsWdo+w9jCUOScAFq6+rGcCloGWTkE5/lv25eZPC5H4AliZ1iaX0
s1Zh8gYg9IaKhkH3kJ+tkdCO3N51/oLVYC0SOAVfxfdn+lZd5lHaSbXUq3EAvWsxDtIwt0PiMbYK
S0oZWvnqnDjc6LV9fW2yoIHf1qaBAlRhtXMPcKzdfqmbxyr+xpkXa3haKCm+oeG2/UOPKBSlH5YX
VQAdlj+ESYoHz+Pn48fKW925eOqIdZVhxPfCGJaNmo5AKpwXa30Y5OJjUIjkCTXKOMTXZUuGsFhb
0si9mM2mvgeZVNSt6IxiLjtTaabtkY0Es2Z0hP8cgBtzEVZ3r3zBiFTHpoYa4o4Fptfr7+f/2w+N
YQ+fHI26dfptfLZpik7tVvrrLEi/qPpO08f6wuylT1WSVZyiM1A5hqyrJQ+xG70f9r3yWq44NVak
E+VN8sL5C9x6vBtUWw3QnmzyalEhB1u1yIoKkd/Rlck5rTzXx9PMLYlgMt987W395JAR1WvDe0m5
TUtr+lnvaB8lAb0c5F5quMSG1/AiJogKzlS3f0+3nCM/PYHU6/3ux4nhzNhnnSQ02crKV0UKaQhu
cJ9j2dmz1CM81/urI9z8HOF9vNTK257hL3dU98s8sJ2iZCX3oXgHwNft+mMvfUbhqT3XZSGwmCxh
B1ZepPKcbfoC4FU2PWkan66nxskdUKs0KCEllMQkid7+jD7dxyqkPapgzOjZL1QjssiC5Dx1iIdB
OpjNQZUMDifiGhSKvnttdR2Zq0xCn3MWkzUg1waHvJ9Zt0oijHeoLsV0bb7wIHoyHQEzB2B3F4wY
juHs10TZwhMKJ8s3ZjhhEbexVEQd5oUXQ7RzeywPrbXbhVQTeE+FblDhEq3KMxVQrTbOEf8jF4Ax
nhskwMRq132BdmmvDRqUHQC2xZ7/jJ/5G02izJf/fnGZzc/lIn8y+kKS25JdwV+FpWEN6/Ei6Y7m
CNP/+l4iY39O3183ERqpXHOYMJW9GYVTTrYbG6dNvWAiOW2EA/oehAybVUZH/ISMk7KLZ58RrSw6
DI/AYkSw07BN00RcvNIKdyDZ5jDfbhz+DV2UON+62pu85EBbbpVxO0fP/7a7zPsDSVZSYyqzHEiR
TT7zp8J+X/ExveZv694MvEteScGO/74mtgbgH3KoOwJc/y8RR3NnqXBd2mdqjQDsEY8tCnO7Z/Od
NWkfoaCFa03xv8n/Icqee+LV085v65XvAhuQNBBVbWxug0+ellyCl8kj1DQlnAO9Lxbd1ehLK9YK
2cD34OomXuQir0yl1qyYl/oFES7Wv0LoXCoWedWSNRGqwgnenb9mF0hKKGhcnZ+Zx+pKYWIRVbjh
KqeiBxRS+EHtOl0TIbobHz4mOm2dorOG/7SZD8s1RJPUNx2CZKIE4EYvaFMbTUsv7XXNwItXZ7lt
qYvKuk72OD79BU27ois+hHIJN+8Yh7KPlcZo8ECA5fGEmmQy0U2VHe4Z9v1b94ojSz6qbknH3dJ3
eQZ3Ohfkn0KD4n5yBtcjF50SIe7ro5yT6cuPcoaIgd5RAF3CX272tp461u+g4IOPXyivNaR8MNpK
I81sjbIhDiVDJYtshEGot8B825enSH5zmT/7MWfqtXb3E7jN+JLAUnRvHRXVCQi0zEBveDHPfBf+
A1SUN+9YH9jr9n6gYD78aupXSCoXK/T2NkG3DLMM7gHrm+lQ2Cjt7Zl9dWtUJc7F0BETezIHT+A5
vjxbZqhv94sx8KUGm3vqMC7/lFwT61Z17hu8zUJqFI7gmbbsN2LIBrpaL0Yu4WknoW7b4mXXoG3s
I6TM2fc94L1dqC1guNAWUb/hpuhP+MmAzmApksP+7M8Kp5ogTjT+ofXzePpgMDux7QAmgqjfcTuV
rYPqyLzk13j80RC+uxQRxS5wqT+mpu/ZIeEVt9a2jL3qSD9EuD1eE7QGedBGf5VsoaknT38rerMc
yvYhAiWxqMycSL4EtMtG2/ovg9il03mzkB/sf2vTSO6fQUSzsH0XOocJ/x2dJM+vw+odLLWLJRZF
+q3L31bwHs+jhdovxPXLGbTPx6tcqAM+hRLdlOV0GTaycqaazUbkRgxH0vkGCvP02GFzrrX2tBUE
+r9ZbdgGihhtN1hN7nF3P3WQ1KqKOX9R4Qk0mOnrFXt5ZAlQ753i0MsmdORNk5xUkwUQiUHa8Bh1
OSorLTXgQFjSO5Ub8CD4nW6+vykIws6NQWUfVZDDhsS/oO5HVElwrkOfe7chViAsMbf+63uTE1Ft
VBr4mJgN5XKiiajUQEKmeF0XehBjMsoWT7+G3QoKpWkGRinD/LU8uAEaLys9ownSGiFZJ4oyDX3P
mSYGg4zNc6lCmotYrfYm9k7cQ9ekDs9Nq2VRmo4Zf8Vs/O8oClDANCCSSEm1W6qsIfC6TXxM18S5
OG1HD2jlzr9nuV/YEuNS+/y0e6LWdBBcWGr6AX5/UAN1ymD1RVG9R+aT12pjySaIWLyeyKVeNe5C
0gCBJ1wD6Q7PYqGrZdthjHFo/NvfJ7uQ51FM8Kc0XS4P6F2aJm4poOU1591xVA25QkMES+DNmLFD
KLXXazyKeabbTim4BcNb86xNcrYzdg4aOSysvB+SH7JIsW881JEPUfCOuaCy4rpd4/YwzkRF9M82
sRwuTZIsjqcnKcx3NWEkRaGdH+BpY3EPuTy3fm88zNyIMDh810qxZLtBQWpWuyMA23gd0QPwk9Be
R/CBUKKjVt4tilJanFzdI13arNWBG6Ad96FfcRpcDkNdbVZ3EcFMHjHtZ3XLmhsbTQLA1SC3UmBY
B+8S1Vi8dtDpLkr4BXQbvgCEWosvixzRICdXrfYRkPsdkHUaKZtBrzzDB9hL6CSBd+04LTwNy3H3
k3juur9iKWb3g1IeFE/EpXYwkJCgQ12bFVOTM7vI0i9QQLShplR+8kcWHBA/euhg1Z+/y+sLLWlc
0pg7PHronSOFtQZSic8pS3nVxUs0jorZLKzhAr+Bzr4lxnNpmHh9tH2ijMQl/ponveJ/6UFBAt3J
w0OjXvTQo3KRE5a0PWBL+k1x0apKDaZDpgxIADgL9G34zQZA5ImkCGlQNgBbI9X3LVzOVL9TQpNa
0pzv7xgCsdgyDQ1QjdtHzITg6Kf0IBYM5AQygIzUw78bgCAmBRLGIp0c+pRHe9V/MBz0Hq7ZsQcc
9INXMGtnTDCNSTFvtHtjs6jEj7MRVI6pBbx6uQQw1uHtlfbDlrBSv0HotKFikVqUDNRVlRJqKmxn
NEXZrt6KSkWRZi0UAZF0uEIej4ClMtobuB+65Ww2HTbzPnC11+tYw7wmvC9ZgAEtzLTPznWA6KdQ
d08A56l7nl2VIfD9YswxwBfabHdL+I2/Deo70SZjXrqTg9/LyM9VSYzjawk2bEh10rwSEqukNAvB
39e0fvnuyKjFa1Xtqb4pUmeW+TavevDzk6rJHS6StUSD00QpcMWHZ4lbFmteg+dyXbv5KRGPapcF
mrESqKxyUgIdN4hsmxo07nMlU8aDG8WQrVpOOwhpOLuy7CBoijsfYdsy0qqVdykckainy+X09DdW
fIe8htBd6TlwsncW462pKWVybKH3lH/paEXSyXulbfYzVKY8weDeUiIRFXXT2V2qyV9K8/1g7tI/
WlcfJ3Tau66C2Ypl26VrrGSk+RfAdSXBpGWAZBiqJm+FA16LDdPwc/84DU4Yc17PWEo960h+JJlG
29lsxj8SizyGb5CCgG+mq0tFPsGkXE0OmCSINVasznFKd+dB/qdwVOP3nNTz9OVbi1YbUySvC5+x
nzmHiCXSEqqpxlFYRj+8vGMrRlWpA2qsGTEUhPrmfHv+RSyXtfVypU/6TAgZZ7VsBpLqQBClRc+f
j9CXsE2Ac7LH3CqecVPuFq8pPQIGon5OYS5EAaWL6BECw/sYM/feqheIU+QKbCclotg4cedWZjuP
R4bXQ3zYj7GAt8UiIMGn8yjfLX0YdMkpi+HWqfaL5xzU6j2+I8+mzbHYDVtRDtybrOzXlYjMJ8QK
/XUxEv5MIZv/mOSeCioSxJT2Fas9sQGY6Yv3CbL+/dcJBiDcp90HcEVzzNBHE/wwUXkP0/WkfX0J
/Z3vbdPpmKnaLP7OM3ad7leJ75KPTwpxJ3uuTRvpq4+u2oYssLbFuTvYzQ63SSBYlGcAM/4nH0OD
M1HDEqSzPObolLGUfdaJclncxhnOi8du6+DQJlo3/O3iRdS73BZw7deyDhnKHdrebjtMzHB2Re16
gbv0yvjL9D0X4ke8nPGqp17vy4VTS0zgr9rodYvwBTtW5wrzQdtfZTl6K0x3M+asymS7RsKgBdwh
QlEEzidFHcsSz+f5VSnJaVRCk385WhXtX3zgjQtNFSn9LKFgNl7SuhhzMVMeVfdsI9/iuCK0WXzy
RQtJRyRmYLxV7nEvrfDUoXZHZDM/jxB3ejhAIxmk/9HwOXy1TqWjhfbDlNunnErflkIAjzj2MKVe
rKhIOnxlc6YnW4wiya7O6VEPiRu/lsuBS2nbJTIZFWiC1WkjuNeNG4dTDfT4SlyfRV4jzoBy/kz/
nRfbSH88MeoOd1KbYAql1FM13UQEo5x4lxwnpIlsDU0YhjiJL2efyVztR60Kj2bhIfHh8qAeSeVT
bf1mGs8fImL+PeHRUptOfmS+GLuqnHc75iLkhYNYw3WBlIkpb5UQ3iFB4BcqqLc2dSvUiEmXkUzr
ickWyFb6bgUzP2d3c8lzU6tAvGUxIFxQyeEHCQUBxXS2F8gCDPEeBJd2dXKdwsSpT+fwq8qvK/FE
FwHIsORSjwWdagxS9Ft913OvNy7007UQTtdGRyM11iM6YxPU7iA9UwcfO6BEwU069eaXtBsFyJMr
7tZ4es2UbUEkNRZD3gUWVIsFph42LLM6pYKBNMAWl4wvaQDgY7ksMnD/RXfmOxV3xAn3o6r/wMID
CHYkvC7UnhuYAK3w/fSfWD6ukkSdbdWl0D9vELCZ0x4ShaVuaDOKrq4CViHYjqnZzARXk6ovHXsU
nMxrxzImd/GmLwBWI+Y1vWQTKVuALFjFhALmGtSOIFDKrbjiSd/9LVd0+UMOveo7x0CND7TjrJvB
ZoDAoXKk4OcJyO1qSrboljP7rU7Wk7ZX6nN/wW8faB16w1mc3/gB42gjf5Jy8RPBxNqDjh6m5qma
MjYtr3tg6z1HQG0hVnhK/Oo9Tu6Rb0+fwXvwc0GMgPb9Qb51h9zZdwrqGoM/MIOrfOo+QyYrRFkA
69/+obuGHDuCSQtnWDTyONHaSVr+fwukFqTh93PX56zI3bzO8P+tdUq/PIjqymWPhylcqRECUHjq
11UKqOsWolJgDCbJlYyqOWua8OaqwM0l21FHsGfaCxmFU8/DKzPjrTR0mFe7aTCIXVCVdFVYO4iz
nGhEjVtPl8hgWj4JVTG+HG3YQh4SlIuhLhU8r9gVxQEaRTyKrSLKKzNP00Z6nZAxh9iffskbo3Mm
jKfoGkCHj5x9bbGwCs+HbrlahMqmVWrA7gDkEZay/hj5XkgKIpkdNpuMX61ouBFNF3z6CedZtLCc
NdzV6apOOn1Nh7lFgwyrKow7oIj5ijy6OqJtXsFOTr+ZsJHY7vThs3cjUF/0pWqAt/GY5qwX/I5P
i/KCgv9g4N5Jqh6d8GdKIvCfo4kqXqY6XHGG3cCwwUGHzcBhzVkx3YJy+An8d8JfuLHkWjbzbHEx
kzCS4jHH2NNpMgadlsyUq8lZJNXfD6nL4K4KG4ceOFnkAtxRJQnkkyTwFTg7CpceIiRPn5p9/Iuq
YLzuWyCYbduwpnAFN1JWQEEP7+ZMDu77M6SL6NdtCbEvUM7LPsAFwFRwThLO3F+PEOOTi8DeoqXC
kaRxPkkF75mKNsixgqTb0+bJFQUEN/WxsLCrtpkMEMl0RkoZVn1yX14aelweSJtGltBZWLtwgg0W
SEex1m4No/pVF1HCsrD/V/Am0TPFkh7kbDTd8YIsFUldP7fFPwd5UubuFzoI+0wFHrUZpd/1Qx7H
B0vnaoJbEuRdMQxkVZqO1CnI9Shc336X4C/RF7X+/lJbB6bamvGkA+N92MS2sz6Yo4qHLtVZNGm3
SZaFqRIILjh+vdVojZBXTyIA7RHvNlcl1J2oDnb2trwXV0cfmmTsjFvaEdlJ/VRhZ+Fa1IBBWQdK
EFtIymMatSCtu+i3fOQWP78Yk1P4brG4XW4/Tyer8yx8RfUQ/teIOAk08YrPX7T0Z34XfZwAqYyo
pl5AFg2WRzj2zXC1Z0vuoUovN17OM6edBf1tJhacxdJ/4+NsRzQW6MpVXUVHg8KOJw2EOm2OhBBd
3oHGOWezcwejGeyvnYjCWM8XKd3C3oJzcMjKPsSXHHIwHHnvCUTGYaSK1BzmUXK0gfHFjo/a+hpo
05Mvb5pDjdVZU+xN7fyOECrA/rJc+5HozR0MNCN47JAKfm8l0c+YBEM9AK7KX++Sv2WllOeNU6AD
WZ5xeNQhwB/WkQyJNHGgJDlBmyPcSS0SyVgxETLWOSqyqIf+CelJL6G2bz6mwjkD7N4tbeh+gTOn
orvfYCmPJBoGqlwoRvvOIoaqzYrvqs0nRZsjX8KeNBDqzzVePCdBYWPBK5XoPTk7bGy5+Z01LvRc
RrPiihAJ/q3dOMg/XW0efEJ7vLJQMntAScHnl7oYwdYDz3GKWHjmrEkasVRActeHhJ2+2ZY2oTJx
61fucVRykM8U1ZpNl7vu37y04KeXPBuhbXUodH3vVDRp6abuyVK+9zyyZB25s2q8Rn2TVv++FNcc
KNRUZQwIiKqgBg619N4lw0nFqENTwkxF1HXG/jyMInbtaquAcReVGkSU16uUrgPOr5wzPZui+K2E
P14K0gba8DYcuRD4elsLY1yBRo5Yem4DKbSz7+f4rk29m660/ZcYJaQXFFXsf3U3IIGKmFDwxMyh
0cEpl8OLKmKeGY2DTMl94NRotzfPxBWXJl7KW1ItRGnqSIhVosm16lNhPTiV14ktvoWDutMXz+dD
rHIKqBDdo0D+hUMWa+CM0KUlktyZ+PyLiwUdZA4HuowofO7+YEGSfT4hf+U5HWVSNtwVhYpmq0nH
C/lwVN97yWgWBeu6JCs+LvG3BlnUd4Uzwb15ffqPcd/vutB1uEQtoZw6t8jEzGJfmySeoa5Vz1wz
irYx1B466D/qw00RR9OCxTI8vcQ+JWP5RcJPoU2+QTNruzqROwBxIhJxqFVtUNIZ+bhVU5ddXpHJ
ZwB3uaQHr/adjei/vbA5552IW/cy1idEAGQDw8UiCR2MVLJOYyvRiivPn8RsJy5NPiohMNON7j/6
pIoIa3aWthabDjf+yWGlob99xzH0usVYXCqmVQYjdYJ/HiPpAR2ZjZliXFPoAIdvAPlFslRBgZCl
Fzv+Qzu7YDD+hAOzBYlc8ac0aOtQrMgJm+16XlFeqIh4daOo6WZhoSWcNe5GUWw0mPf3dOnbzEqY
JUtckTCad4ap0x1zgSuxi7insae8/jGx59i1Dvcnoo6OFtD9mpBRErb4OwAEk2zh1qNekemDyoTg
TGaqCjo7Ox3yQ8ZyvJaGTZ9eoDnDzdlv5UorkMMXaUdlDaE4YjZyLEOmdGr7Kdzz0RUE096KPIIK
UmM5oPgm/XURK2jhlnx/w4v8yUjQl2mYk4sy55eK46W2Fdatqmlt8lApcWbf+htaEVT9fimdiZPj
dEIyTNc+RW0G2uGB8ytnefIavluBbt7pruNoIov5W6X0fF5B2fc6L1DKTl0GVQp2fE2Uja3BEoke
XruNfKzx8APbj1yXiToeXblRsiBNCpKoPQE8iRka04Ysxej9lY2y0bnJPPok9xTbzm8yNj75vlIV
KM2q0I7GKMW43+yPzZRL1QGhZkQ5Ns3X943q8fRP6QNahGDYtx+sAr88FQz/gV3hXFxE8qM0f37o
oGxKpekGp/sGCLs9196SBhBsqAwkiXf5HXLL93mKOxKfwckcfE5zzJuvqMW0/Sg5qrdxktye/rdG
heo3/6qqrgrdX99TEoiucG6P9EDEx/vrMFYafGgbYv7Z+WV/dDqFMPObGgP5yugOvtBlxYU5sOKu
pIZNnBI8Ny+bpNGVKD08qPaeRezYZgalKHXIGCJhht/MeVeSpNqNWeq4p3me6KWBMHVcJZUbB+mx
3LktMKsf+g+mI+q2tMjiATi9ygdVmHSeLZJaBsXcwLJHG2CjhOJ97G9oatqYWyvSnx7pmTbUNKDC
a+oQq/Gqcom7MRo+sfSo2PHpHTQkeocK4sHcDCdKB48nlbWTLF22RKCGFwzhiKNnIYxfb3qwAuSV
SB3jxYRv2cFFxz09I/VNYzdT/rC4daJD8lMLWePqSNPK/VsC14umb4tXX/T9TPc3MbKil0Ksy8v+
WVONDNQmCDniRVFcxp7bP1gwHZPPyMKrxNXafj5yk22oceyu3KeTubhDc0CWihRPZiqELiyt18VS
HTUZa7jThp2oVKE45WhzuQPwXdvgmyCbH0sm3z7YmUwilAKbpYT4MCtsYM3w3uVlgTCGlFAhGo8M
ApKxKvj4+RYpy1FxpYj7fiD9ZtiuO3jmYnZcHLq/qpU2lckWwPSQktxGlgBL0UB27QgkQVWTDCJb
b3OyfAE+fMr1dUrc7VMLZsp2xDFCbqwhPAOwQtkC0PszJP19rHKr1CacwfSZ5gF0VlOrWKG/X9SZ
fFeTw95xWLUyAADqbkyr3vvXG8Kuom1Di/abcC4cKPhW9bbd1HKJo7N3+NLHIR2FXDfY5z8NUHgC
ZlZ4DdXZmEqOWPKvKds9lvocVapU44UrtojR1P2C0RoM/A5mPj8ATjgCbC97tAHbaYasu57mlOoI
ujTi6SY5fu/qjOaeMZmKqvWZZo0raoa2V34g8KwYdsqfcfDAPObs7z9/TVU8g9LcxSSbVRntaftH
roJSgwcjnO9jf2kSQazu2OM80SsqUJVU8fNf390GeEeD8JZ8a1fzqvqcrVcrA8ItRB8rQoEg4NZd
TXs2p0DmN5OETEgtmJBLXVfq6FVsQW0P8Efoemr1kPgDFmnxHscKm1w3fiHkfDPy+NWgAda/ojxX
QPnd7G7X+nq4SFnvKQIez2VitWO14W7JnG88o7NepoM16AD9vPaqrxrnjAS6qWa0BTKzSA98sWqF
uZYSNjFNlvAmuZDkfC/0tphTSsTm3c4fkbtUZLry4DhHzw4hajp5FsJ6bXv8ZYEn0X1l6sAaxAI0
CQyt/hdSa/a0UGPBs1LcJQHpE7fpOv26eH/Q5bWbiHyDfBJiCMw+nXziJWVWsj+WAAvm2CtmnMpk
Syc6nwz4OGG4Tg67nzjCldTp1qVzl6nybHWS/YcT7bVNSjp4M0pJ6ZaREDbj0EW6R7F+kbQEDyU7
E/ENbA8Y3XAKgpAM1a5eS4nI/uDdjqneu5mCUlFv5hf6OuR3BF/AYS2LoLUcXBiPD6ESVDmvglZZ
EjAQx8M4qd+v2OfV/v9Xyf0YxENJc4Q/sw2isLIFqfT4FYClXCcgHWFUmepYfh9jdfQP8iUN8BbD
GQ+5dG5TMQv8+7nXGfp7psQCmYprJHWXylJxyBRB+V0zX+/e5iCIRTJTNPpJaSMtRJGP4lErZXqR
xj+/jC8wJzb93rKnJUERy/zoe9O6J6f7KhIal0XyE+vC45pto+/lJ+bSeAQVEoqvg2hI/PzghDuL
ivJJ2TshrWCPY5X7rRCfWiGU0PS/zIDZ0F5qHEUVlVJOXaAFs4pFIOmTLdUFfvzfdfSjIx734WhL
jcHGqZf6TjSKDqtNBAQjErUEF0tcrSCMvLAHy2cljiAkux7YnoRGxniOSrAdppR7xNA9qOO0oAhG
8HoEnNTgi2m5/rhfHBdtCjdETBeJm/5Um9NnRsPVuD7ONOV6yXIGIOWjTDuQwIgruXAKKg3ZjR2h
utf+RxXmsFiOt6XC+ilkKuwKcPHVYF6f1ToLdJoocOIbXOcxN3hsUCtSqhb9ecMv5XbaGhGWot3d
qi4iMIgAMSjvBbiJLNRJIWRXu/A0AJE4WpVSC2NNxSr70KH1EZx3z7zGYGmzH2XlWEatcrIYSbIz
wHwD7Dz2tCwIJR4rQa1FW19qcQgYRb4P5qXHUkt+k6XI+q1KuaQ6XyXrrQ+E7peafj+OXhlTmD81
FR3gSRn5/sj364NyrsHmUXfjpCuGquFlf7VFZj/KXUpUjW1UtsVwZZWHRmwpjNVyikwwOLeBtZKR
Q0FFKSuWFJC4rmfeyXgahJN6w4TVw49yCDUo0p/aLwqRjF29Ok7rZc7stINnRrdLcq+gOkylLAj2
mJJ1rNPXd2wbY4gA8CQqYbDOn+9NvPwZfFSjPoAtLj0/lgktPpJM2raebzUo3SOvjcMDJJtx/rDI
BWBw5FJ9ybxMh9X6RgnNtKYh6URR2H4whmjjvrX41U6KUTSwzPJGxqNIhMcfgAkHyUvsX/9mNv0J
d6JnsL/euiF3Tbo2KQ4m2L3NiuQgADfVYCqlA1HTUm2DbXgo4lQvjK7rYAGDHvef0GQycNfTlwR+
hCvxKnqsoNojavwzzIovBnKrYDwZH0vQ7CJ6niOGA3kFhNLsSn5e6WHlmLSrLGJlQuqt4DfjFZnn
GBe5nrS3hXMfKtH2zM3EgBIyQucq4HUT3Cf5aRTPXQtaZVG5TI6NUmlgOIsb6owqZac5dUgrJdvd
zPrSf3/MhJE4sD+5Teulqjkg/QxJGwv6ieyaKGt91P+jURd1nGTsPULV5pAF3U5mp+OHSKe8CF2I
HoCFClCFWleKpXlvR3lIZ6ugRCSUhrEPUQdXMQb9d4L8tA6aviB3IXIDFa7n2n3ygwD1pEAb9pTA
3RTLV58sFR0lsQU0+QIMVFrZWflQXzNMQ7kHi98aoPuEltf8UIbtgpPglsNcpWL7Nlklyst21vtm
LoLixU9Qr5BGt+a7bIyRB8w8b69mxpW7DhKwy5qmcmhhZtImxxfAEMzp0Ytm7+PYwmEne6aikH2y
8i6hEX/1+Q2MTbSxA3tMWNcdU9mkOfqLXdSFGFINj9C8z62i4exUTHFmHMWNPWmAjg8tjk3bI8dF
61XpScIP0OM7kXMqpJ+dyu3FMryRy2iKsBuVlsKaj7e5FN/CopfUTHyA2EDrp93BTOzGZFmGsuxt
FcvpDbXR2ibyBbX2/DC9ajVQq+dFWnsc2Ebskd++qNZTHt+zkLFvxmDECBjHTj+aQO8f6XngcS/d
qQK8QvOoJOqOvPo3BUCPJabpbN4gW4Xobzfzv59SsjM09DZ+JFRfcUwTICNMl2gPK4xnXYFAQGkA
xhC5su2LLX+gC3emnTTWFrZjpngpXRJUX4VxBFRZOGMlO7EOPgm3vuAffublb02ZRaMmKSTfRlgX
Y3h6OI0JUXqPwBYO8rBQ6RrgIA+PNxoDCH2zK/tovEgHa3zDr2GivrUqgEBVSHw65hMHFn052Bwo
cfgtatu5WsjqV05D2CO+UxMdOw2PV5XEnM10yCfdWSDGvTUxigjylgmbqfwHH1pDhWKrIKEK/Q0L
1JAF1HDiZtbvLLM1hAUOC5qpO5uiVBVfL0eymYDwd5CnSYhgz9MVNnnI6kTIf6qbf5VpuZgWl5hp
lHdDHMcsGRlLRU0GZCi+C2hA7qtQyg50PQEtAu4Gv+iIZgbk8BtdYNc5tLbR+49iArnb922aOgvG
VkviVfwvIn5zNWN3jYgzsDfwu1FbvmuBiL7PylJJ4wrE5eMW/f91AFWL1NZTXK1NnShg9O0UxlkX
o1a/xSTY4lz2eaA28tm6Q4sm6WYLh3110VvbzypPHhkEKATAbKovAPoay6Uh7iecT0IdJX3S2unP
sZWaiMByu7NRtTDfh7+z4ETGzKQjgBmbrrpOR1UzVs6UrOZlUlak+5rTl0Fa5GXWmkCSDhSSvr8N
d4K5heuDIvxsACjQpHpnF2mGVsp3jR+pEqnqAIfy+mtfyx9P3IxdQZBeY8aKAnQ84+hkJtJ2dP/W
i6m1z43M6ewKFoNQqxb5CQqhKGhvcRCOp1X+gq0NGfspu7rZf1NrKvMESvt9gshO4FDiwvZNpfNJ
yhUVQsblsu/E40r4se+w01fhAagaAS3Vot5uwlqLkpcO5JfW52QwJBJt2B56aQOZL8MwrX9YgPjK
zPG6LU/iOfNstNFJhvByBt3eDr32FTSZ8vwrW688G4KhHVCiLM/nQxDHL8FYsET+Du3aRMlYuboC
Usdjllp4h3q71VFcLnL2hmUDcQb9pzqLX1HdAsdI0tDbt/g2Da6VwdTImusO5iKfiH4WtrMtTrR4
/WGy1mR1Q1khNT8J9ygESFAvXhHflUMRrLV0YCGuCV1dNv7myvEwuLVn4TjjlyU8A2odw35XnndS
dP0Or8KYvlJF14QF3kNyP7wuzCGzuYJP+WIMBnCcoSU1a9qDzI+B/n5JVJekoh134/vyBSQkUr0N
oHYm9Q8CEElDVdOqUY51RijTTu0j39UPwm2B4aGwRiII/hEKfqK81Pk78hk44QnAhqDuMAyWW9De
blZQny59ltCXs04UtI9pbb9GcqqzM/Vk36UC2hEOmg+oaxLkboUMeaWqwYGIxiFTqriaeACwuEww
+b4ONJl36pp4TpbBM/3sITUnbwJyUvmu+cA5hI8s9xm0jsRNYyzSoNVksFlCIXBpAxc0HLiCigaQ
QTflNBFjAiOTAcgtBq67N29zTlPZuK6ndepnSt/R97vJ6vCjC54v2KsUt65PfGfZ7nx3AxsTgA83
lvsiSM/fQQqgZDN/R7OGznE5Cj2zOFB7K2m8K/sZQblNQAoX4Q1zN31Q244CzqDJJ+LjW7Dgh8R0
FWiXqwLfwyeyvYVKXfY4AXnOnrn1I4gpL+VbWDteyU9DUfaSjTCb49OtW/Ajj/XbGl/nnBzJ5ird
p04+fEKuB9JhS9UjWHlzb5cwohDNeaY4lmf5MHOGM5zonaX88VDL1h0/vK09sBlCQtTN3/iO/7GQ
h3MUyQQKdBVJtXU7aAfsfSzivve2BKxtZQgwTo85EPxZxtO9QYwBCl1VMaJD4PCqxhep3XLO/dv9
Gx6sw9qw/rNi1vQE09z4keyi7ZbTuQDPSx1Ua39304r6q3gU1GxjOe5zZlXgVFm8OUadji6HjXdV
NIIwH7ZVkhWnP8UcE4uIQiTLFKQwgk/gEN3UgjUx3x5A2myj1wk+CU/qBmG71buwofajyRgEwWgj
5z0uHGYRg/TyLNaHm1Jkdudr6AhEp6o39ocdNPTi7yDeDwbWsYmUR33iihnaTWODeA8yjEUmp4ZY
QLqJ6ytlaXGtrS5r8/jRdWp/WLJaPiMzLHkfK9/c1iLTqTTh/ibP+JI5SXv8cRBPrIo50XcPCJgf
PBevs8eMZgJM4FirNB83mqhRF8I5jcgF5F5IgU9BHNpRcpF+nTqXg2vcErB5zl3dx2eUB7v52/5T
mqW8aX5zrW8VWZYSejNe+EoE/z4+4PopcPopCnjPUKw4pK6ZGChMN5eX5KWOQH+HKc2Wxiv2dXPM
+9CaCW5agPFRlCqR1zCX78ui3RW0PU/6mmKDBz5ORH+5/TQwdSJd4tc/c07ClWX+Jdjrj0nM6mLg
h0tbxBJ1sDVfQiq3GDIKJyDpDlF3884D/7DdFQ1mAORl4clKpzfZCr8AmIs5InztWsQOL/YcNsW0
qgtO64gTbbVPBTvesIBzOLahH9aHXd4VisVGlAgzNCzamqq7hONNlt1uj8wZCcE/TqbX6VkZKqBl
99raFiFVMcD+k8NEWJC+BRIuNDtdB1TMNLqjqs9pM6+M91lR5JUq3m6A6kuDVChFIfqwm9zJfCms
GvA6omy0kuNUGmO16PdXtSZ9Q6QcYIijcmWo61f11kZSK5eogti7S8PVa0NQqyNso8pPPNc1eqOf
BGvynHIpKGhZbPh46QN6aPruiHsYuIWgppqe/wI69oRpYaXKaOFzCcgm4tKvxdrNCWlshv4RMEiR
YkI7Q0jcIwOXrEDJz6SooYLG7t1vbpoFUH2saRHQS7qdtnRm5RcVmmLMgkoBOeCWTBDWIIGvnRzv
E3em/1wubaYPCeSzsmkm0dTNx9Dc75hrEObhHnYqvq/0agdAvVK4rWblbK+Wvz1joeh8JmrsASvc
bRJ3/YdsC40F3UzrL+xVPiQtoMTg2gwhzEG8wOAVicOEir6IlyfChfuU+yHo+kJfwW5hqe4LMVaq
h4mtEmKYrt5JP0NaqNpYMVQOu0cf0igbx+IhVCdmK5donNuYxfC3qx6HmIIdMTcvadJA/K2tH1Lx
wZVooux869P63V1e3xSkl6MB/e1GQV/NI/Fr5n8mqI+DAGm0JToMWQIdr39Amf9LGoqS8QE2aHvB
j7844pDwW/m9/UKU0+NLITwZNCfkjCUAuoXukmdX1DffbW7+Cv+gSO7VOzNPCLe+Pt+MBnV8AzUe
TukGi2+KQPoZa41mfXG6KBIXS0g+gdcbjVh1+pKpM5Whj5asYB20qniWsXsIVb9bC6q8nq5LfLkU
4cz1rSCp+9RLxhLgPX4J8Y7q4G/cZv3vkixbiZL6tplSL/8mvwlHEdRKvc6AD1W+1A4R0s1m5O0m
+uayXAwMVDIcz8G2dWUYGdDOZ8GwEiGBoawe/iyfeDJFwyNdhRgr8qxQidLvzxeNPHG+jtN4CLa8
wDRrSs65S6Ae9eWcERfkLwXpvsDtHFaAhpRIC/WBm+2wUsOT/e9aSmcF2YqC5mFDYtS3hqomkNe5
nrxMgf08ELZUC57cg4Rbt788rnA1tkcLRD/buuFHpz5tMprGLlcOGPBL0UJfUlpzTOn/P2VBmM0+
k0hNzfFOg7N0hbIZln9ZcOEJRE4KeBGX2rn0xzeW81Mv13WBaQ7b078KLuONzh8pj13+Er2HExu5
nSPk3IdesY3LHdAsVsXm3/7u71N1Zlfx8eq0emVUForiUn8CCoQinpFTyYgd9Kpt5wk+aLxHmHDw
7iHNn2VTAfWCM6RvISSvZkxRnNqyrthncpQkwFLd2UTtMZh5e21fMOJadVoyK01u/mNoncx1/1ku
aIxppkj7weDWdt6H+5kz1RvYj5hOZtNxk2OAFTWTo7ll+f3/CdqtRGt+avaTcJOJrvVeqMEuL6qp
164IRL3K3f/N8j4z8rLmBlgWH6kVFLI6e0McjWGguPvkduQJuGDmqa449tihW24B1N1VcX/CMuxG
PIwBEyNvUwTcg1m4unJNPTrXEG0oEYRIMewc0y/VadWSlSNoa5msGyqRMIsRyBLFa9GsC/OAT/Pp
GIvaWrTocbGJI4EaG4reNVqaw0GfAklQaQGiiitIodPGt0BeAVFHCn2fyaxB2Ij5JbZms3LeVSFz
Ijf0KMMYtOWGidsXnYqy8LqXcHD0s8DGf9s4/WmXoE85fOtU8vcIUcbOrnOwTcJ+SDPao56z0jvs
s7qhNmDmfK90rzqXM0chhv/SoC7LppRNQdlTMHOV3T5lP2TvpNUoGBo62yJprJQoEfXxEHLZk+z7
3RxSNzMJGUfG49i2dVygsFXnCxUy6TIXxh0GzKvp1mAECiD4cnpbLMwKcO1cqDFsPYVHk99Rc6Qv
3LR3g2C2je+yRwoAWbjtxZ2n+QO+vFmMPue17OWTQ8xuGBH3mv05SrmNYHlKoG7MRn6P/9SZKfTI
n4nN1JheMeqIcijSpFPFg3Z0AyLWyE6CTcQm+TR06Oo8klwMni7d8Rk4bgLo9PRZAgI+2k/l3Vty
10HjlsBCs8IbmkgE71O+BFQfgkEV5o0iNcMf+ysk82bnhLPzyM+ZXImxJ2CMSiI07iK9Qm031gha
6fBI4x9ourWYiYl6Z7YU9VCeEG+PdhATsDFg34Q/9Lcv51w4Zc+C3HhYhLmna7Tnjo+JwLMefjaN
KHbdRRXc7GpGw9kVo+Gn33NfpzO+cPcbpfmcRf7GhNhwH0AiG+kS0vaEqpWAUuzgI3AbXV7J4twr
fLFdIE+j0O3sEJpyV7pUrCxtMcszaImLzLJbA4Sh2NKmVq6q37X5IJ0ntgP3Ywv4cbUli+tyPKim
am7HSaUOw6NVRa1mwizwxmlIdv5P0e3nm3Jq5ozGvZE4x6DiIYMfrJVJwImiE6xw6TPflD/QY4X/
V9QfnFOHz0djCS5HRKaXS24JdFU0vCtKFndwLVGKkJUtlzJfimUbb69VZOL1FerSC3n8kQNqkhTA
eY/vBDV02zAn/0jEi/9TAj1ncDtFsEFEw5dW0BWsSE/yhb27pFVeohjcr49pCO4b4+lQgx7aav4O
Bb4tUJM28hSbPrJCwM79b9po5T0nbUkLkGbodFQGkX17Wf2lpfJZpTC2seY4DusX71g3whkgORSk
D42hQjofzGomZBPz+4UYfvjnYbSgIRomlYSFPYQWtz3RMGF3NQC8gYVLnFV5t1s1wU2+mV5RzUBz
/nsoXGm0xzE8bXzhggxAPZaqZUt/d9ixNo5lauNsw0SGM8IrT/Jq+HETXdjQS1naBJqvxUKi7SSb
1Fxfb1cdgI0E8N6Lt4TCWwGqrSc3wq8gj2agdx3HFbkfExAnNM41htmewqxIxdaZboCWbOmdyP/h
npw3Dq3SjZn8hdmwO/Nzq+UqOwo1hV4p7UOZitVv9v2WnAi7vqK8ZSJGlvxPkjnKWDZOh72PfnWj
VtS5Lw9aiCLObBsyrvbW64UmCflCgcbqvHyDIupxnSqVlGl0sl4+RL4mI9j0vjfnjmEwMEalKRNc
2+8fBzhRt8Ci1z4nvRvF0oYpyuHlsEm1fYtAvqE+1akJTT9NLaDWjmHj/R6X8JL+B3MzYSH1b1tx
fQnt6MyoZEMyL/H4zeYbn+OvHwztvHH02oKeO8vxLzX6UTWpeT4iUS9omp6rx2UWPhLG9z9g76ch
cDrMdQUrkHMBTAZCNIKuduEGz1GTXxEkOHZPalGGXS1JTIi69LFRNlZ5sUvKIBbagYRsZuDfrBzg
Xr3Gkxvvvi9X4X+KLFCfB4Epf62lXP36o6wxOpkjiFUroUMWBnJSAmB7Mj/tPXPLVevJ67XmbjoW
T1GJUfTx+NEk7mAfVeGaBIm+HBXT6iVeKCa+prpiuIrPFtIyClJJlBQ3UOBb76mE5aw1ZeELv2cW
Xb32qJ3TARUchWhD7g0gXx6hUZ2gZe2Tvm2k4yW3dgTUdfz9WkNj4hnlCi2ILcQ0Hcpf7tInugHM
M+nVNivQyVrfeMcVJHyC/RM/yUOSEzrEJpi1enVJeNe3z/ihhHKi7PhBEHKsgI5O1FlhuR7JLK3n
gPxeGC71TZ9pL0RDmNVK8U4o9X7Dpn/seJ2QDsQM/lTxZq2CryBQi+q015gyCThjgbpJaU+DF04A
yG3nqPPQbLV7h79KjtTbj/UJVWnchf8LdS3Ir5uW3iPofl7yRUZz/dMVD3950UBwVv05p59A4fZf
A9/5ti9L37bUCkTWEmpDpSJAP/lRK2I24DJGmYemxxq/lAod1d1RF+2WOwfu1VFIhd+pbDEJbauY
MKVwyYz7rkALd/T6eO2qH8HWfZQlQt1jvTZhGhb5MIffD0TuCsluRPZd6CytuizCINCRx9DUPx/J
xyjZu0cPkNaKEFHOTZFUHOda1dOr76gNHMqc99zi9sPo0eB47j24Kwr3psmlxsZxKemBVI7QSXa0
cFfgmLtXG2VCyOJ22V9oDxiXTp3NVG9oI6t1Pr8YlGrqKdLDvM12pymj9TpnBZ/9nEVhKsdsDCeI
RxPGHWla9lgC4n6E3H/LlXY5pndHXCQq6/kxD8bnnEUrJUTTq/lc5X9+TcPGLT/aEvqH+zQH9xeP
b9qJqki3q8ecdVCxDoq/Ez9uXeE99+2c7P1s8HD8V6xfqDObdpIngvoG8lydWLaUPrwpdRLAVJi9
KkDQ/5kWqT6pJLtwXRnkVAxTVv0FoHc38zvqwNtFZSzSoUIGG7kjzEX3pa7ENBaghDB8pPzZ6zfC
wLXZhZ2MUidk7mLqoY39v+JQps6wb2EYAc6sRk1S8qC72E+oOe3wSd83mdZ5398R4mScRbBWQONN
/poI4X/F5f1lepGCIuUXyJ4wFo/LOm2YXhDW/F/nbjIUbiESHh4xsgKlGq90hMwA2vPuAFz9cP5i
Mp9KiLPeIjk1lddprogNtQrojIdgdy/60yG0BQhMxcpC0V8erqGXhIk4CV10ehmsdmrloDM/3agx
nNbE7YlBXmOYxwvjccgTx0OjL6bmAzUmFRDCWZ1GXJvsBBO7Wtsmc1HKcpvLlKXLbf8V3fhx9em9
UlAGr2dTdak//per/IRFTdTfq0DAUirjcza0UVNU/zQNaScKETStCOlO4z+LmzR3ZS5u5pDWGDe4
47vI0eH/w5urlISh/X7/IIyr6Y0TWglx9cTYxlq1D4yZ6mOfSCdTN8mbngf4fV9jPYNjaJ0+pwMv
J150jwhyUv5SsNuoNGIgR64O/C9DxKGbvouz0DByS9rwI2/1/KjpFtNpf36/nMlwfMpKac5zR1Jd
nVPdUuYolX8l4lSYPmT5phmZpx0uo0jf9dwia9P1LhA+KWOdFlQGuT2Ir98qSjnVBkn3KicpUeNk
PLFBZqzYU3MxtFWGIIwmVW5uuIF1MK2EV4yR1mun71kQgEwJwedkhkHXPER808Y2Q2aRGh2C6ZF0
hmJJqRc3ZSxwOOVas8c53NVZrcKs7h6jtT/G8LeOqBSflU2wpNVS0LQuABxnyO2qJiSAcZJpAlZk
ZanK9+lygbAbt1XLA7WdsPJ/97ojEnLNdgexXZRuwsSa1r40bFse7ZGy3YNYeqrBP9Ezxea6C3X4
pk9xFuO/FRxIxCuBu0If2J1C6jBWPhT4ZIVcaPx8D+7H9pHTPW+kxt9cBw0sMB+oeDkb3b+urgGB
HqTPMcAcfb8ot2LrUvDLOcVfyu77Cd0CtKgrFEcSnQfz+dy9jpivWvvg8BudkhLwrUM3JPArWt1b
6QZKK+B9oGg6MLbwKeiNCiXDMq9cDYHKAE5MUxhQHHnFt0TLE94n3cpW7EMg8plOnhVCKY/qBnaz
Y3IjF0LumrVch4eJPxQMGqR5eTlHGH64kBmalIsgPRHsueObFcPJXcuAgeKVQ+LI+VlPwOQYhEU5
JTGZAaDIeaXp9yLY6K+XWcgHdvuBnF/NYOz4fzey8jSGL9VqDNchf8H4KpmSyD0NzgOB9z16SHMR
l/xaDLkvnle9AiirZPGX/LKva+bZTEEoVNc8OvvYX4Lhvq4jv9wSWzdNxnxkjosF+sgTpzy7CqDe
8pLmVk93DZ34sPVTvB5EX7Eem3jLA4ge0aC+5EXvDaPuGFww1/YbwAvX1SxZKIT37JE38mJI5Omo
1NpaIVSjyx0kYRsuuO43f2r6UMMnO1X5bA1Ow1GMzWb1KG7FU5aUnQaUN+fNNWnX3XM3ClZSifux
NBIlDxw31txR/DOlOZwxZeUFvrG/y0OfMjdH76Qofyh1gSJLYTC5SG0YMABmgqZ/xrFvmsVaZyfO
6gw/2e/LEMFWQcDC35WX4obCnap6pCiO2DIklrmJcScFGknoPFkncjVutGxlCe/JcGYX2yuJkZfF
c5vdxGANXKlG9wwHpuLLP5tD+9qdtVPUcVm4VGD09giR8bWFmAzDrnaUQ9Tio6A6o/Iwfbv9L3Lb
daeELcV+wi3M/F4GcsA0/MnkgL/2K/dZZe872lA6w6zYxikVdCjBA6TXa9c2Z1tV2ZshOVrohgZT
jup/+Z9/6zeooaN1MpLXW9oX3FRh9k3VtySWhv9ZfYtSxVBFw7q9Yvkc4R0WPOjxJ11gjBuL5e6q
CdZAEGBmlM7ggvABgb8eAJ5jhl9CR3Q6RtgaB4nejmouDNrI30OsqvM4VL+nn4l9YYzAwNHsUQf/
m3AICitQRwxOQaVsS1utQYw/FxHuSObyzOZDRd+4Qw4gtzeGgfHhlJCJN82b3BecFEA/Fl7VVNU/
mj8qSpYH5l3u5PU6FJ+Tb6lggDp6i4nwpaJm6QNYhxz3HlWVbZAVRbbIcygpJE0RP3FEONrkQEhh
ijrH9x3iZ028A+632CHja8c7bL3ASLNSAnwmhUDU2jkISZ6Hx83FOdcUPXjtlPjpXFOeDATgBUYo
yzfx/qkSAiBhWsOJZLPTg9A49N/VHdvWMSCbNd8H0GQIeXmnIF+KwWo0pcFJM64Cp71y1JPhkaWx
GGnMdD6vSLxjdND60H7dwqNdZxeNd1x6ni1pYInC5YQAU+t1RlQTEwNr+9YorpdVMiZlSYcgftvP
RcDT+to6VEk3/M7s2i7j5rbKmYryAqiHBU1D/NXv7NMET9agdwvCuf8piHm5wEacgR9Y4jS8jXss
Pl9VDgdRVJW2e46Q9y6G4ekmIY0M8Der77vHK/7a/WdhAT46mBV18jlZSo81krGu13NRFsL1/osa
uEYsRy+Id09Kvn/K2Mo17703nIDirGt3a/6jynd4rcjKfa7/1NWhBLRPPUXrfNvX5sEz4q0aMIP+
6blqzX6uCL0teV5f+wjP9B8j1NbAzUO8U4sJTmsHcFysEfkk8TeJxzzbvuL/M8NApSE280x51peu
gp0P2/6R3zqTopIf8dErsAm06JKnmt8RyrNXKVsxKdRfxyYTzHGEQAUZkW5hEwk4KyZ4erWmQ9j8
KHPtmXfzq0aWdm9hnK83NGMrAA1uw4Kl5/vcUdRQTO8gYjHZQkfrxoCee/Jxag9a5M6XE1m887b0
ne2aOAkPkABa1hRSjAeoitbBZeEpidlK0eR+WIPl/jACkplb7j3ln+l5KnU5zIL/ez53BNWx4TM6
i8tU+OtAFHulGreoShJGIm86N+pTc+JLuvU2vZtn3p8aFL7RCX5lj21kxCyCzHmflONbmwdPNdvN
sdBByzdAqqCjCKRQOkWjsdg8OMwdWxIzqRoW31FIm6F62UaTmHlAiZaJhDFmnBoKFBlOT2HwkhMQ
aCJUrHZwVBYs3pCHZFFKzt/pGe4TvjINZDg5sZRcfyL0wSz+gTb8wXfVqQPFxIV4xSUo01mVzkwr
KrhfrEuScq6fcVVwCabKpfv1l8k0XbwA++7acs6WJ6Y+PCg/WJMoOrBduGhgZ7KYhJLEE4Ry9r6u
ChngfZaExgGmEKvRPiDqiaaIftq0S/Su4LHhdbkaNyc7erBsbXq26zwlXBMF9w666Itq0TLeGdfC
2xAfdItjXAOsPmgVJL2m7wJTkhlvIJngH6wtZXDs2YCbk72NzE16+ZmYPlvb58WzmZN5GTsljALu
CpzdjytpRjKlzTCgVfi8XhFigQan5dXApQzsp6aWDc3wsOsAERkyaIp9eR6w6VU+qU+5LugKvj0W
bkgyhRdljVcrSIOI96RdaWgHksVBRj5FnxAWBkYZlT0TZcdVG8nVKgRrIQBQ+6a2sffUXf49aL+U
sXv3HBjfTJ3K0yKMjUE1mmm4lZ8CMoOGcREiyaKtE7iTzFWBOgY+cAfKNkcOtXgRvzng2yYK6u1Q
/q57E9blv/21owpmuvAttQcF6Qoq2M4reZMelcm4yUP++Bn2aUOzjjASs7yllrrQJkMpQZxY4abz
zYuVIMMaQ4oCx5tXoDGuKaO6D3NFTK87L3h1Bj4rrxvMJuU4giXbvhKTWhFYdFv7SXMUnTHv3CaY
lURKzdDk4YUCImo72Hs+vwSwnNT8w20so2gUwzhUG8d0mNbglDrUprye1hlZKUS6shpTOmokHGwH
+KGKSVPAQcbGlPKsK8yXpzsOAI4DiXJ/fMgM73d1J7AF4cs2IhIsva2B1xiYh9yIQmh9yK+ir+FX
dqU4N36gW9c4b/6fOshgMT3yzk7MSMjeC2RkmXKnnkQNhAKcxLUIhR2+mNwEKXp21vXsHXM968jB
6EjDvGZ2aqkkUb/wu0epnqgtsc+RgTi3KlLwOQorTiHotiAVabP6BvP36VyXR1raSMDZcU2bv5vN
55Z77zW5Ga5S7FxXLbKkUrinWWpvSrxsJazifNb2iwTq8sQC5VpF/s2oJ7AstEo6AUhrguGqMoHE
Ufud0QSI9CHz6yLwEosW8Lnt0s8R7mQ/yf/uZti0NazOwsKW67UbNxQAvSSAHihX9zBQ0P02Ckac
6acTHntnUnogLsLnEUT33IZz/a13f7SM64B8qeWcj2zN2ADHl/PmfE9ZYBvU9AYgcmblgjbrHmWG
1AL5uY1LKaSB8rVk8jzDQpHO0cTUgOLcjSGZFOO95T5zqJfOcjORI4N5BIwsi2vC84vKjrXbp0NA
PgL8BKffEg+O4A/elKm1E8/y8hnlEUePTdPz2x7n+g5KYNzaQbA1nYgpUXCRLAisgXwT9uXlr2Xg
kMc0LGtlmO0C8Jb0zIHwYP1nN0nyoubBM0XDXk/bCkEqMTnuwGyWAh0O4Y5E2hhj6cU3IyKeF9LP
N0NoHS7DrKEldbny8qm9CgruWhLmt4Z54BAb1NjhGwGHCfXotfvaAFaF1Ge8NolwA4sgTvKsyqde
+yPd4P4V8ek1VB35TAk6ddROBquG3YvLGEVWY4GzpH41aMF7VVj/H6BxhDY+a41UxKyM7ThnDa0y
f+hlAXk9DwYjbTuNP30H42QIrmNtUxyAIQ0Z4ku2uYRO7bcD4phKBvxwsyx0oiKlBfE2wdQhFkIF
MqXgfB0CpfPD1zvAOJjssYJqxI6o07qGTpe0WWw+9AveowPLe4tTA+9T7fZiO3NXQcP2M0is8N5/
iMSj2iQQoHz6zG9kkFtZiPkQmRDfaJq8zuP5wexOC2OfMi/HZ13xv9iCxmKyEGr5vn+ZLGZAHbAr
v7AmopQqKhAt/b525LMULma6y2BcDVXIwvBVfG/ErOWbHGWeCs2OREHY61ML2RER/tM0GEAtP3b3
/hmqOBD0snq3f279LALN+AGAeRjuZoIS9NYvcIbCD2Y+hcwRpI4rzfAMRGY+tg9tl4/sfT1OSaK1
2zatklsSuyrgsj7MdeXDRtcruli1jkADY7U2i3shhiIl5/EjVwkZDq9SxZyzNMr6TVTnvhTVjeuJ
OktDRg69BcLpJt3XG7k98migz/vnTuJMUh5jJsV3xN/0LSRxArX1RNkN1VBiyH0rEoq7aChx7PR4
pxrm+Bg/hNPOPsYw76jF4puqbGztIwCYMdRE0jWD1DDS8a3J4RrEc5m9Bzx4sj7nml7pDy/A918S
8XM5fFTabubHVI3jQJY8mS/3ny9ppceVfod7jqR06QkjNCsoD/QtoMeX3BU4d8S4ns4C5sLhmK5V
yQBS7QDZEiQKj3+JUk2rf+MrFKDejjUwGRphbxGSHZs9UIfqes81Fgr+xAKWAommBpuJLpaVegiL
ZncQQ2qaLzLus2mVrVz/acduqLDTD4tdbGPgOAxI4+/V2nXk5wR4oiGeEjeMQpyXbD2nFTiwcXaQ
8xlJ6FK8KpSaabkYQNEB+gfUYmiPyedO/0fDHa7viT9UB/yZnkaAYwc7iXdcKSEoNV0bZuNK/2cz
2fWot0m8jzNBdXYWC6bMlAlXhYr27UDBzwn/mJITdmaMsrwD5OGbZS8sYutBB5UbmAk3g7J3oI+3
yUMqL4ebDmxYJK0tDsoiAMMw5602sgU01UHzurdtCJJ1BQjgbJcGkPOadmkKyZFmlzaLcfm7fp5u
81mQ1dQy9qaYM2ziuIOvKyy7yd3PPTV2OPuYKrdKKw5ag6qihwIqVEv3lqoJVqILrLKEOWmCLRS4
ccFhlLl/tocM//b/D1FHeKEJYmc+9/d18KU0+dpcxtMwky6NImV9qC2uSHymllmBq65mzRaS6l+l
jp9NzzOw3+IUAShymWrd7XbTNu3ep+I/Y/v+PMMndE5d034ycrm012c/S6Ow2Miw0CfCCzSDdGag
6+KifdDhJzBtR+XPKTirbpWVgp+NulzD5ks7MxZ5WRmn3/16GXAZuPGwLcQjRH+7YE6pb8sKJrPX
CNnOP4lxT92u8XCFQrSAlKTr0B2gOIqeIkcT++z2oTVSCk83lPr+0+nTZ+KUjVE65eD4rMTkiXRL
8XoOG+F9S2K6GpE+8rT4pC8V2743vJku/mKG/b829yA1zLhqcDrwO8uCZ4bqa+Qf3IInpG8mihVx
ZIhAsdrPbG5ym2SwF+8AKCCWEOPngbWDluU112UFvtHtAEOy/VwaSW7jt2oo6A0ejWwuzYZ950OU
rvzwjjvoSjyyRH6308DihUKTA6IacQq3YWF0sEJoAeyBjxRyzMhFW2faPuWKcjY7/3TChCAJOOWk
GcNRyl5ejmwKJRx7rFjbccirwPUKQZq1WwmR7qtllJeu1w6uHC//VdebfcZwwHrVVnGScIKO3SCt
df0xlZ5LlGhyYT56f3wB4UZAqxKGtk5nbgTuLLbCOm9dlaoTQSnxaWdVU+cUCYmekAy0ulKEkIbz
NNWYOi1valzTIU9nLwfg/SYH4DYD633IKxOEqIPllsSAXp/qSDYB/e7mmgAH+QaF3qoSX5MA7VUx
dosy9t0898MZH+jy/Isw0cmvVTHVOWbUUndwINURmXmfieuOmS1HEAirzEwfhczRsJIwxlsPXKJj
uxjHqCQU8tqvOqYBi0G++SYf9yHcphnpX///LWjvYHwxBhtXZ6kF/YHmN9mfUIlw6AC3yLxXptjN
Z4Pdspa89KoMaH+nba0LP2WiFqNLM9IcYQeGMD2towL3wJGv2VXsfRnxb4i4thY2yDARLk86YIz4
vkgj/RVe9YBqtCQrQw8jwYAqaX99j8BRaXkY/mhglqKgvPNUC3rO9ds5P/aXu0x/7KNwlgTkXrBe
awxaUU2M+88Dcp8BZKi8yn0idIg1cv30Ab63xVy/2KwDrI/237ahyZvwPUhV40iEd3DlvcW7W0mA
kYH7TnPld9IkPbL8YrHpPZu7u5S27ALWgdd5Jv5h/NGFTwna0r/R7b9/sJfOAUNZMbUNnq2OudCE
Gukm2jG3Uh4HLKIvg0V4sBht2batIA5yRgH5Fh56J/PNzdCJTUUuHUuTOrIDruTIEpduSoU48TuF
15A0Z9h+2s0la1G0FGmI+HsK75VY2jPUHEZd6BxEoaybrdm2CovQ+H73lk+97gJFj+R3Zzn89r4y
ZWUh1ldFEievILj4iDD2Qsq5vA0neQ+UfrNg5uklfn98GrltUJD6yvc/p3wyKYw+tNhEFPMklcAz
QlX9eRKpGlNdewoIKiuxKA9zvTnxsIrOBg4Fc5K5BFHJcG80/drN7OT8HQuerCc4DzrSaeLpqHm5
wk/6GpXiUpeJd2iydvQ+lkU3hXKYApqxN45TM7M3ukiZORV8dGEEsnwcLsJ45kGJxgZzy7FGnZ4K
S/b2PPB8hENJw8Tk0/AYv4LFPAhh+Ai2xGHzqCtN5A/dwoSjOGl4kMOkliCVUxPGcLdlzoZm848v
G7tX3wB4Q/lXAevKhjIhC70940vQ0qyYJi6Fhq8QbyqJZ9QRXBAB+aao5fSTI9gC5lOuimeEiTy6
vl5XLToofdWG6Vs5wsUK9GaNPqBzLcgLSJn6cIaTsXPcuAH6Idgt6x/OXB3bevP4++HSjsq+hryV
reCikGAtY9MOvqby6V4VRz+T6TcAu5vCi4I61LOO85ul8hfek5f3fyjGSMsSJ42R8NvTisraPofd
dv6CdZaTFOgHLjVY9BkdP6ODCOsxtm+YoRTWz2TCw2fJpl3iohBk3TbWQyYxg3LYUiGLwSh4Cg4Q
mM0pHMpXSswY7yzG4H4BhbMFa9tiRZsGPpFYb+GSnqf4yEDVxEXUFR8UHYdsEbuPjMh1BIwHKCpf
P6Wi84HYBXJ/rSgqA8kengJSQ+teJlUV9buCNU89UAZEswvQufUwHORRKJeDR8ZseanMACIcbZbU
IeRNJzipF/4HiyMIRVPfzZigzy18gBNlOHlzV2PJ67JbB1sIFfFZK5zV/gy4llawnhJxTSVFt+a2
FsfWG8uGI0XmUsjMUnfAL+aI/1byiyxnO1Odvo40qWxVhRpOyBWTju/DhMuLNQmyT2jL2MZGKX7H
fccoE1o2zPQqIF8WSTQiFA7gwMNLFdmBAjlUcQqfFAt06zqm8m89louci0pR1u1X/KsNEXQFEVd/
+hinU3uSUzllpZcs7Ov0vZdvh7IBXbSHMHvpuSql7+pK2Hg2ML1c9ECIIVcXJ38e2UTnUTERrSZZ
5TdfGDrGxJ04yWMw8NvTc8uTKt8Taguu/NzpJfukmaZmAp4IiK826QcKdnl6uUPBPpl2hKWasKT4
Jkopi+FljaeHAEwxiNFKJrbhdhzPTQUTP107hcK3xv+64vPdz0EpfnGY3KTb35xuYavmnGQlzK77
elOYCpFtLURKtWr63kkC7SihGp2YminDyNf7Rzx0tdNYk18OvyBiNVR/nB1I6s7qu8BsHfgAOtQF
L85AXz3u+D6aE9E2nSexmEO6KGSBrpvsHuTKEMSAV1cXT08GO3yTFfTpuPTpzu0dpLWMREbtOqxC
Ji9gQ6Plu1ydWoUSuMVl9JjXHOpt7K8AIEqEOOH9kuyRZau+dOoD6Xvg9gZy94Pqk+qnkDUEtjaq
sxf7NrjB5Nn4K86d5w4hg9uvdo/vlBWLgKFYy0R4gYijtYsXau0oaUVqXHXwG6xRvlw/G7g3Qoto
ap5Sb66fU2yHP81cgdxa3qMXoY+V+PQOnmIDR7ic2RewxnHMNVZvu+1rbRqubL7hKdzgcx5p+eYD
JjqdnSFSxFfFMM7+eLWohDhFt3kkBb89nwsDp2/zDf5gdGJ1cf7UIVmTrZt2LHizz7Kw+W46q944
2v9aEn+rrnyHbKxzTjRkilW6XmlZVGaBtGN0QdzttjR6ROklL3XLXzV+gBLkxqaznSgg80gRpGMj
kt/q57M2weRC1mbq6Lbjyq5qxTgihu+82smYUfYBcawuUeYjesWfBfkkFN1nOYj3lkONbRYevwe9
+W3U4Cy0bcj5BOhODJxcpsQ33W6/fwSQYmdgp4xAlBPqe/DlxcftR5Vy8DW8CzFdxrEbe6SGzZ1u
mHZS3mPxWduPXszvqhrHa2Ohp4YmG5m2KC3E9+SzkqqxxJAHs+qGlidk0LcoBIVp2mBZ0U55xdon
GvzdQPnYXA/XRtDU4RGnZWu6OZRwvRDrkOisnavuGUJNmkCCiixWWP0k49Rhdul/M0KwXb2Q3Shn
Z6RK0dTVL0UpxyNk3LgwB5s2ooMNy2LNijCi+YpCbgKGfYn3/fKmNevdwHsZFP5WMSXpsPtAsqqJ
yPq+AZVL9jrpbpX+1QiX+WbTEzu8rswKBLB9d8R/HS/Bo7UPeUMUZNsWV4eYIGvxZxP4AqExB8mL
1n0L1lb+icaQuMZn66FMOan4+hv3VM/N7Z0Pm1JeFGBuLW5OrH0Buj34lt2HXTD4loKdQx/j+O0K
5icEG8vz/SycwlG+0uSXDe3xU3gWpCj1vbijP2KirHS7HcPAzMGhq3YoEvk2BP7f0KN1JT0Rotxd
PD+ecerV7J3tUWfctLnh71a0o+QSeE5NLHfHTFzyaycRHZM/EEKKmAjk5HAOe4NQBH/NX+9RJjV2
VGoXAnYEP9Vt0O5psgjW8WP8KT0/u+ch/cUGv/i4he02md1cdoN/yqm+F7/IJWZ9Hzj5dFFVKw+s
+Xn2BRoPNSOaJVKp3E57zKe8t2P+CrPujmGkHvIwK2zCMUP9VKbz61MalYgkoCjKshkHJBXtiHq5
enBj+xtZ56+SRAL4Pe34Dh4ThFW/oNtOZhmyelvFca75yq06yxFWXJwrftw2wftubwJyLnJjlpWa
Cblzg8H2p2A83zeCNS1+JyDH9fwrnz/CS+PjJGnlCMnO0Du8AtKn2r9Qv3vQKJxGNEkPGBNKIl6e
ilvt7fzn7tgzaKkgbn3C3pKIAqRKjuifMbfkmvDOVXK9NiBDQFRZYHJDkwyJf2tAvXnOfbFVBfAA
n1bvuo+UcQnaqljhai5vtRY1+YxaJ7LChImGm+1u6aB7dnUwufZrSlN0D4OvJaRQQYJHTT598dhn
xbGQmESp1MHh3B0fjE41rM8MCOLKaReAARoCfuUAm98GESQFujp0b/ftIEVirqjpJH6q0g5tXUmA
oVD5EyVtPcQ3jkTLUHwPpnXFBEopsCMHRUcgK46gsjafv2leGNU2hR3jT3HKStiRObHjuFvtSUNK
Os49l3e4zsEZ5OyWYLaSHFnZlXDqcmzkmbIIIWN4blRJJgRnFINjc9TzHVrvqOy1UUcVnVEWh/gW
GzFVrPAIcqNOdwciSRgvyLjebk5jazzGuBx+xnuC8RjBoU+KR5gqGh0+N+ixnCC8JWW3k3+gbqdb
0CD5Fjs9AgLjHvYQd0GQnuHrS4PWfcepHS/8gNaHJDEdbwIxp8/x9L4Rw4s8A6nNJCUArrMaylJJ
eipjCL1IFBel2Kk1sJz9JRIqr08mBRC7aFAER8Q6uY4tl6jskboMdUa8eC/JI9IE0n9PlCpIAk1D
FoInJ9SXg2ybG1aVZM7PspLEQStzAjjQ6pWpWk7sT3XFA/SMIWt4Ib9+awTnDmk8AT7pI61fdS+m
Cwtvyl3anGwch0n5SxZTFywV4MSvzIYucP4ZxZH53v5WfvFn17WHrgZHryJrhkdphUMTt0CNHPdx
o5wd3qgAAPy6kOMsRpTNbILF9dId0j37G026lDAfUu0cbO6pMn9EgN4kf6NBIRqk9KzT3JlcFO8e
XcSSyZgLEKRZHoWM2ttavBRtDKgG9VwGp5eCe6kG2X0kiVf1LI1vMoub5gr2PzitNPdAjbDcRKSs
T0lv6mge81KbtycjL0Mj8We76pzL7fPhMCG5eeuGn6Bii1jhZ/C77rc955pPnhKrRrZBxqDaoZgW
7jhlZAgVTb1y27Ns0Z1ymS7BpDFMiTZWsC+nRDLKfRxH/eJsJ9skiTyLnD2akjqcEoAo3hpKcg9n
stQ/zqw29vSG7SLm7OSvGGSRISC0/ZoasxlfIWs2m/WsEQmTh32SfabmQXGWy0LEtpf9BMRPuDP8
2ZPkofpBx7COS0EaiWksbyEVvEXj42C4eBBrgaM2Vr0Uj0glOzp27zSaSHm/OXzZp9Q9zeru8rCy
1FHd9U/UQaX/Y7vDrb/Ptcbfeh68y6HnPkm26a2B1iBvmwBkcMpA5/x8H8SLzh/7TAPRiaIbffvM
rscR3+1Sque8Og2Yk78tTQHP/c77yLhekMQanoE1FhF/d+N6Vz7upNvTl5XqXm4m2IF0zSBaxKTU
dmgEJaC2ffWCajwSr3vrcvFK8WnUYsCwycjwKye1gCBn7nslg9JN/4YGLtO8THEjW6zZCiAS8fGW
mViyWqeW2bT4l3vqCTh5BIxx3ns/CTrWm6trJEHCy82AHzP3/GBrO6QI2A1N03t2H8mgoeLP7PoK
lcJJXN/KsHJaAZB7rrG8Wx5XH2EJMrOV+hc/CfSnuloubBu1RhNDV4KQ3TuKgqcc/NDeNTxCnFm/
Y2XFdlJSr+GdusxPfWGPL8MiYzsfK1m2z3pSB9dohEnMx8w6Jp05s0UGqSk3dU+TaND/lcw9T1vX
5Hkm8CIvkpCoJeXvtaFnA9l1CEC4UOrtwKITqc1pEp3KG62rxLKwN72E5HEq+unNuVEyVb2Z8XHE
APRIAyWrB+wr1/NoLDvH3BVVxN/COZNRfsXBxUCmFV1b4H+bW4nEBJTDZCv/1/HLLqoZGQBvL4wG
GNbiVdTBeNJiitOgpvWYaeogvBcUUC1Ol1XHJh/JhwfznF0wh58pc2Xi0X9ARZqurla5/V1NYUAw
BnnzWQ1VzJ4waQPltTmmKwfms/p3/+Wtr38d19y7MPrDoyN4K2QLrkBXcacTjii9Kn/56scWg3Vc
7h7h0j3wM+vo+L/LOLVsUXRw1/mksz6m90BkYsgAjRFA5vU8vpPXfANqhvSxnEFZRDkeAAU41UCJ
FniV6raT26NG8P/lNDInphNBulMuS/V0VpkhLkO//epzDtCT579lazjiFSIqo7GlFCYx6piOrX0u
Lr2B6jEIuXGeFFXdfN6OC2vOvc2oJLvqZwQHMLM7OfMihsdBWEWzyeabtLC3VodhJPAxDDc0IR44
n1yLSz0+nfL5y12ccHNGq7lVJ5n5pbjLj2s+rUfyDwdVpZaqWIeGdr0676Caw3IjmFLew8YCyH0x
c0Pu0XEFJLkWLOTU9sEXDqYNBJfmy+Cp7iy1O6Rb5ic0RJpooQWUB4/pjUAkoleBiSBKnJ+Z+/3l
K+Vu9LMxDCYV8RfXuxxexJEYiMfFenKC1WuhYfA+hgUzPYU2OnSg1WvRRApF9lHC84VSIq+ILLYJ
E0J7FMLArp4rSqIvojpfNTBQ6BxfJBeye9xR9rSXjWXCjWluCitDUNiKxXyxP9jG+EEnYZHH2kzi
0Q3i3dUt1WMSn1LPv9vXovWiKa0vEzGyXAPpg7RM29m+VvdF+bnXLEnW6DQ4vkiiWHjTsL7Vij8e
18/p3bDr5TT4owrWFzeqr52gjWYW8f/ftSVDNr6aWDkV+HZ2ZL8YFBUUxJLEywwhmzKaGE5Erndn
kOiOxBFh4n14bAqUcdZ3kl4Wo7B+ysJV7r9JwP6DNJGDHakdlqSetCWaifMf36DeO4lVpuYBAEk4
y8uaM5bd5tnhYD4vOrUr8qed6h0hEgPHOG73stwbqL7t3fcerqn0ISUOb4g7whMiI6ziaNL8iqdR
kdf4fFMWL/RjAhWBil/Yj/dxZsIbTS0S41R2PGP6Zz8zpySjvXhC+hD3bwUwh/60OWbVs8XC7SLN
Z67pP5fXFVENrfpWhvaTU1rV+ZFtIYIdSdiKRjA0eav840yJnqrdIRqmHjR/UqQwRXtlobhxRKse
4D4rH1p0iCDU7iazejt5MetNBU+9sINUHJwxzFpCx1jnSz6CD0NaIaMo9lydvWcQVYvCd/zEu5yb
EvBQQuHY/hxWV1Ry1e/eILNf5E345q4w+3Dv25ACi14/7oYg/Vm8FHwAP2oxN8d8ZnKnaulYHkG/
nUxhDRxHRRkNhkn5zvuhepC1Of/nD9H80cEniXYdLAntAhpBkHvalRFTAsKPaZJrUWjVXqbktUun
+m/WaKIhV1vwXqEryzLp+YNk7lOwPrHGhJISgoYVRh1E/aEyCVA06RvxpNox7bgAqRUJA5WBkkKM
eNXwJ7FBlQtDlXNg2ALcnENSAw/Wrtu6Z7XM55ljBqzwudaYaDHt/oA7el2OsQU4dT12w0OzDHxQ
rN0yVhg6LLw2GGTvgHBUf4zss4bdbyJHN3xTHMj/Ke+K6yIkw1SJvtl8jfvc3y81kQ6JQsp5xUWd
053MlURp08Rm6V9SQB7hHFErbMYChCuTcftrfmF7JuJ1tHtvXPbWBqnQueZEsAq6lYxGntQ5W9KJ
lJ+zWeFw3DI54bxRTF41ROSl6HNCcYLDXUiMvTD27vzLEGzpKMRMed05A/XcLvPMvhUif5/JVUE9
wGicbNtVdsqBMO4liymeSZZc0qGg3ibrEzpsIyrdXWNLIFFpZmDTY+T99Zxh/O3dC6ihYX9jJJ1t
yS8Ra/q56woxAKV5GNKX/pOI/fKVn0db83iLCoHZveCJ3gjCbn5dvjLRksEAPnaWsr1qLAsdKjxk
98C1Nr1H7Eh+AqmJR+LvzxNicvNi6gflg5M4fiRFHlqWMe+HiiFwYgjaLAjQW893h/8PnIPyjybl
8DD3+ZDfABUQxxEH5Nxq6I12Uf4pIsvy11MXQru2YvkgexK27kytDryqGcZ+igYtRr7vsZJ7jfJ7
n3KS3uFIiPcaePSv7p9KFv8np02wpv/HPQiobMKp3DCO4oeYmOa9bxGj3RcZmveRr4rvzrsH4+rs
rHRuYWETTvNcYtOHlsv/d0r9g526m0cIp0LApWnntooMgC9bSEfNXypkLzKhlDxF7mo/5mccjbPx
cbKopknslLoTNk8Ws1fATYgdBV8Kll9N6fxJCoc70MfUEK2JrYh0v3CJZXT4rbxuO+vsxN8SVAyk
+um7ZpoHyat6nF4yEn0OeJl8G8KvMKH9d3EQyqxxDRp584oF4RBixWyaKANTBmefFTOYuvQVSJDY
zxJkrIVlneYERZyJp1cZlyjP9VZsO56Ianrc2o9OB8j8rIGqOwS0ruZg4mTvEY68l/sZW2XPZ2XM
PdhgjCevSn56rw7RQbUZUPkb0U2tnbrHbRsvz+v1sHC08z7rjIMIZuwuwXSviVmqiBwkITEPAwWT
iG0IutKSTYCK5EwVeTHen9iSweqvYFrN+DCsQI7IEKBjAWp7VXWQFnEifpaEGUZi41rKaJAaUx+A
8kdb8X3xBSloDp1Vr9QTq10WDiVgFSX41ERTigUa5ftfQi75+G1sFwrN7SB1gWWlgZmC2ZnDQglj
mpGKl7CQwrcXQfLEmhAe7KqSy7qHQCiJ1ueS4LWTfVbMtzsDe1Cw4bpeSb0bP0o/EHdis/pPt2jJ
bLVd2UP5BXzaYvOtfrI3qQxTB+JnOF+xowm+1lEOmw+mvbBDSisKq6x1rFVplWkmKi872AtnNttg
PMy8Vi7WC6vMF8fUKJm7kKTISqn52Hixt4oa9YyAQklWeghCwjq6i8VoZGNgsORLpK3aTnWD1uXt
dLK1atYZvYxilBxX57EBviu1ZXUm395h54cOo6N8EdKcnxAf4bN+g9Um5iK8yCnBYvKZiYHQLq4k
PgOEwOm9zF6pse+NlQZH9k5Zr/+6b3uUOmOrRWTT8PgqJeECFn8tvp79UwyHBFAgm6DHUG1DUFz+
pBBIxrPjFMMQQFEEtd+WbBi3LZ4gWkI8iNh1Ye+wUwwHwLzCzWq467TqXJ2kPXH++kKSQ5XS8Eyn
ojOTs204Ra6O+g8QI3KrA4pVsY4UPYv5V/qoiEwsqBZ/4Fswdv25iXa6JlRCs36OGVvvERlE9Sq3
1MI1o60LSm7g883CIsBu23B0CPztwTaK3z9nM+MXeTdtJFoicO1JcWiijU19lEaHwA7XAeXkpZnM
M6neHq2fnpsTYOdNWczUrpmV3vQVXJvjz0qYQkqdvwDp5IzF9ax3f7QfjRmd3aYyq8iucT0ybLYv
/jKJ/veNOWAsoXoJLd7xLBAHhMM8sI85sCgKciKzKag7qc9L4HJN3SrDtNJQMM8VatyMXrySvH0R
soBMOqYO4tUSE1jnDEAipuwzJHGdD7/ojGcCGS24kv5D39O4MZYLfKVi03Bjx7FBReRIGtlRcL7C
NXWi4YF3C7k5W13I53+EoKel0CbM6sCgYJfNl/hDnfecfOhOSVELUzBaRGTSxxqtOWbelHIfGwPw
uhBE66ZLaUW7uj3ettU9weGgBNORkt1Ih2MQK7MIyPferOHo5cmgn1Jvnv8KXUbUS8DjfbxhDhZR
e+hO6enzC4Mownxvzhv27sX2E2cKxowMNUx0TrRDO74gIoeK6BlgDRzV25dw1umdm8JpsUnhx2VO
NYwfMDW2fKES1Y+bepO++0ld04pF5Q2V7cEj3sSOYdQD3RBgllRjjOHZOsxM9/jRJN+NfSAsFBX4
7lDy7n7EZEODcV9aZgcde3mVjDzRMawQeY8U2mZqGrGd5J5IE3zqaZ48U1vyXh2u7S8BDs1StPFB
bjeMLbZzplyhYmiM1RJ+/FxJKkMfauHrTe9vi7w+gPGqMUbd/eICH1T/YjTJ/aVvJbgLxXKZ3P0D
gmoXc33FpMZ+FTI88pgY3c5qeYAXX4sbkq2KTpCXudEx/D8dFVvQcpIh8AWww9ATCQvSwoPKFJMN
J6D0GOCKxoTNvz7jKVFQrApJwuZBO6VxwDYEdThki71VjhhCsyVGsA3fTpxa8DjP6v7W7+CEKRha
TlR2gFqnnQrImlpw5uShsN4okTTNXWgpxcYkJce2UwKZ2xyRvl475ww87m0i4P4ZpNhXmTzO8QvH
xMDzOWkB4BTv78DrUcahQpHfcgj9+yRfGOUbdaz6Ia17j5gA5vBT1aySw6yaTXXfl4QkHFfyAfHr
eF+FnZd52rnWH5qg/xgSuO1q9qd2oubfBFx/nk2IK7H7/S7y2yQjL0QHGuEa0rZqqdNIIcGGgQCD
o44ZPZpir8DKwsAnJQCgkeEDhxar0stbn/SWNXgeNRuL9FYAfu/J/qfIZIH0/j3onvYiHs77/Qhs
ZV4c1jA6O376hMnTa1JYHOitF9xetta3ae48vdor2MDQRFZu5gUNFrRAXrbwyw+HPMKw6Ke0zPWJ
NyJdESbG68l7zBwrhMTkjO1Kky4D8ux5CxilcV1oNTRfL+ncQWCAcZlecOMZ3ME1z0UgPT3I8xeM
6+BIVhVPkjd25NOW1a58GYMRVsIqxJ/tNQfHJDqSb1KsULGMtva47FbKtR36Xljnyvw7KZhn9DMO
ww0SfCx7b/A6zDWnJa+ByKKtOmbAidjhZ2M1bsqGmo9b1iwkgFbU7FFtmmMelEyClqDbMcnKWsE4
Icgy7XA5LDoOtW+j7ElIImTzlqk2vmdYObI7MIeuwn+9heuXWWW6sWZHQuPQ5S2JRe2EbbmeNnps
hGz6ATUIx98oFy1iyGxMlGsHnvR+Nb6s5rJKw4xaTahrYbpKCWJ7Z4Y1Srxaj8mzHbKPJYMB2exK
qVcBXI1TITABuBSObzlPiZEQkKyNa0ewgEBk9dDT5Smez9ZfE1zTbd/sRnjGhswW3W+doZ97paKY
kA5K5C1bDvCK+P8nNw45ruxi8d9dZaalajSKJMyUhsg/RrcylJjhazUb5nKh7CLTDs67k3qrOirV
uJLcQ09533NesWfVK0ymZ82hxKwELnMa3N+q4YNYafMDAlmRg2SpqmIyRmzMBPySpWrHAJgXeV9f
1sb/PUTLSfQVLTJvv5mVkMVlDdcQ92EmgLtudmKghChnJW1fptIFJjU/9KmJQdRXsXd3RuDUXaFE
X/zEicS1Z9Nrn2wivPJ1Ar+CoJeLnMenbAtAicI4CsPZ7qfNyiVKszUzIhflSN+qKmSgV/oZF8wD
hJny7sTf0dsd7P6IPklUWnNa1z0CH8eyq8mNncHNJp0HSuaxnnIPYEAfEJrXGH6yHlr/QuzUPF/1
OkcS8K7RcZcquttb52Pd2WkYf5CnuJI3Dq435gN8FkXg2WcAnvyMrrnYO7uJjDCX0Awxk3B5jxtf
yS44bw5Pn6s3o7sQ9/5vuWQ2XDa23XelLnm+c6z0Cs0Hcet/agv+c5yN0wvhv7X9VkTdZnm0mlqZ
vP5PkbvpyWQ2cWcwGER76M5f8AWcMMoT7X4MfxAcSEe61DcXVF1gU7SsTfD4a6+WOuXdyCXP27FU
t6WCEfU3ZKF/XxZlzzbQrcchhHPMEN85L2GzxRQaXSfRvJE1i46APWyIojJHFhWW99+/2YFVBvVS
CaEVMh4D2kYYHU0/7WYX4y7hKoFrIlUSNBn8i24ik+hgfL8OXqsBDTVVKprPsi9rqFDlvTLj1oYV
nbfVDITXD4iQzkJZQkUEdmvOVhAR8vQUACvXoikpeRBF/ceSmhPPUxq2ZQeHs8x5X52je11AbWRo
kJd7NHNJhoRZx8QI/oy4rLqvFNQ3SinGbuDtK8UM0Kn8FRUpoouLpDlG/lfEN157VeAaJFvIAP3Q
ZZc7IHmNr6DWs6OvCzRkDXJ+aM6W2LdBUQgxToy9kdcCZU9luEdnDaYeA6drscsL4tX4epTrdulj
IlTati44FR4BL14ic40DFc1Duv0o+IWmpeKVkVXz7bNHurQcL5ECBstSYUVwGNWlI3WnVaPy6gy9
aF30MIgAiiR3RXiLmSwEgo55Ghc7Y2nx6qXodr3pj/+b/0LagxuhqQYdePeAr9F5aCEPG3KDtsYh
Zcpz8k7fCpBL219dmaqwu2KoFpp9mImZnjIqFot7HPa8iT8JhD1MeNO0vqg+7W4p8rIeIg0k8BGA
GdSeMCPxYvjWnaSsscLx+zA/VOtZ8bS/MusfyE9ZvSc1F3gcipzT/qFOFE8pbD/UTg4tZc46cFHJ
ug7lM6wrA4Lg+3vM9OoAXZ0AGIIytGBpfWQ1bHRNSsl8MBma739fklrmJGZRwoxtNepXBebprr41
9NP7L9Zg125/OYsNdc8uny7fWAJp+y0i3PLOXDiqStsXqYn6QxIP17jOmgflfy/euvYAhIU8e+Wl
bPfWAjnC9NPH/nkjOnhosniLocvhMidC1ZSo2Zrn/mVmmGJDAABzNHPAh+1iAc8pPFobUbT7FPFs
V3MSTN+DJ8BJoipwJAYj/8AbExP3oZ4Vu4AmreO+Y5mh5Tr/W78Uvus4IpRTWN9jKrdmR6fXLq7L
kK0N+slReGc1DMKx9vweTCbyFniKBpQuKaZCR/zG6hmd0VpfKDjJ4mzGC99fcTQiSKMuWPkyv8Lh
klofjoPd1h8tlwutJhVU/ecvdFmBeIaDieB9loI5xqXDryRq68fQ6ivfbufYS7hwDlczogBGRCFm
cpsQQPMvVipfX+n6AcieLiIsILC2C29mIo3JTO1w5+disl7CMvcu2J1vJrkFM+BgBvZUSePBZEwr
OZQ619xNM84Pk7AAzhgN/EYIEp1xxuCYnBWYiajZq6ti1eGE0LyveidOHoOeggKK0ByzXdvxM47s
28lctQ+6a/Y72TrS48Xy2Iti24CpprmqKtAC4ht56AafhH0lU4cYXMd3TcqvpQ7vfo1UsLu8fhWt
cvW67zED6vcgFbxROmF9TUypdxgJKhbpaCORwCx5HZIYyecmBUScpV+kG1AvAiHgc6U0FchTD5v9
ymF3mMyPI8J1EOuQnMmTKcJ6zT10j8v/L539p9Izbl8+rNwTzH5Alm1fDYx/wKBGYfkBZ0hlJJJm
wImaEMiz0oS7Ef38LY3DVsdBy9362dyyM6HsXAKDTaMjDOY/jik8Uqu0nwcORSb9DV5kpRInM0AT
quOVbG1HXgMUe8jXeWPsZRAn7lVAGYrL/JZEJgnfqLrhGseGPRqPQi9/1312+thMSg7ifvIgnUSF
SuoQj7nk6dKhFidHBFVtNeCuQC6jhcF3X6NH+Z8X2uP5QUGPugRMq0Wi5EKq3uPoWOYpcA5JFika
cDdhfiFIQLeKrnbtS3KvkbxMNPw2IBDHbqNgMknSWgl9hp0P4AKoR++JbzcH1lB4S8O+8Uw9Laqq
Li2bjlytL2pys+7P12KmH88QslRJAemmhTQawbQcTYqLWEbNkYmhNhvLOXGp2cuQj9r3YCjml1sc
9b578DiA7Ia/Tn06I8lpR+YwRIx2t0vRbp9e70EBxibvPcBa+z4TVofPqO7xP9ixSdCNVquwDs3C
5I6Ox/occQrjJcZzijsSuGkOyPnAtJPVgD8/Gr3tbYKYhzTEa6/flit2UX1IQXb89UCutnuKOqdq
dIxIFlEeFuv19oMt5WlcsT1CgMtj8HTN1dZktoQEBQe+lCPlzS5mKoZGZ7s9QKawyqW/c4lwQNON
hLKDmspBnW7KSRm99bQ0Enbs02aoBaAuM0kMtCrfNQIKP4mN2YKep7JA9qvEL7EHyaSqsHHmQHNF
fMrz35FAN26zqWHPL/VUZAdwbpOLfjU1i5fzw8fqsobfqWbTeUjHkUni28DUqZ1c6PG74HWOqa20
P6Nu+ygr3+CQW4KIaZgmcWMI4F07oqzCP2cbpNf4CZi9nte6cvXukZSMA5x7nSwqmjNemXSIfT9u
ZBVDgqqLAxINwveEWNsPCm1NwNdySxI78maYaUFrkr15p2eomeesAnI7CcUF3PjTH4sLKpbByEHv
X0QbqfmXkTpQSh2SbkW2s876memKtp7EwxLvKU0W39Qkq6coiXVlx6GO3TIYk6TKLH1O0DKKWLxT
lEf0PBoZUzjrE3nrpFY3i2jN66tHN1ha/D4rmmk0cVVZmTCEK5Gmfbh/j2067/CRvL3n+wEVODbc
L2cyrSBpjuQM6ZehGdXG354sKiKxDkozhhrgcz2MslIcI3QZx45ySBUrUUHu11ZYZyCEYDztIF0o
AIT+TAAXQKEYlczT237N+qyLBO4Y4Ih4FQIbMlPRlgB3YVR1uq3p1FAkE/KlHx9Qo4ZbsYUSeQjM
RrzewfXAAkKxc/NQ8tIumBlMOdebncC9Y/HTURU7eRHDoF8swkbQqkxNx2o+rwfXIXZUtditGNYW
FGMZoYg8z5WofIxJusBEMd53McATnDysHjJh7wj0iRc44j9a7UK05HOlGF6pvTK7iIh6D+QoBkaa
HxZ9ErtNnYQeM0Y53jRsUHDxPJ4EcuLREOxdpNPj4npmwjZCoIqpY9VymAR2QEqUN4cDgUkgzy+c
dXMOhcn2mPq1A2RLkLdi+Fvyx4D59wit5u6/wMiEBzScwQNXe44Tcvn1DGAGi//e8kVFC5tmq2dg
Eqbd9HfghLYnm74ZixkgNbkXqaomI73AdkRe12utEO0KteiBBm5FIsym3kNMqdBOneqROkXlGY/z
Q+4nJ0CncLC/NkD2XO94/6FYu0v/JhwrpAxCBtEy9YSRG6LopaUWLqBnzXmwgOorjOWFuPBtFaWu
TG3pU1DT3LohaunUVHA2iqihdpbwNRFsb4KAbOSFwCRcE9FGMgaWUgZ0MhzIEnLEyBBzDlnSt8Ko
rm2EYwwVPnfhd2Ki8wK/FVh50E2+f7JSSRDnl9w3jyfiRH+PAfb8xKHDkAf+iFJaicZcj4jkWjkl
xb/R1N/IMG1uTrg+UM1455mHV03A/d9Xo9I9P+uEbNu2RzVi4ZCKgHB/GOKgZlz4yfOJNcIs6cVn
n5HzOfH3v2BK29ySiXsFszKdd1bRQJ5QM53/AzDhcVgW/S6j0Hz0Q1/5AQ9D8EVxs8vHrmLXD2C7
893t8XdwhDvkoX/yVtanLBuDbwhdsEWDqklJS25tLkGZF14pZrCK5kQhrUc8HCt44pSVNmxrE6fT
3BITv01mq843k4bSwRotemH/kEQcwD6Zb5RV+fs8k4/qFlqDbK2y0hSmkhkBBvai0Gq1VWUS8KdD
k1Trxm7iy+0iYZFi8PS1/3KmRW6WYXf0zwCgZMYICDYTtiY57nj0+CXsAOEWAyOdtjQQ5bfBhOIK
35z2L3gThYYm75UhXMekTOPQcX5B7ZVTC/RNghcubjiFLqpKfdyRodrqsidy8BOJ0ZxCFzGYj8tx
oD4leh+Bf4rQgERGDZbXLSiraYBuIyX1A7gJNLwyr7vk0rWuyHHJpe+cUy5m6zvBJakvsqswIiYI
XNBgkIYNQhnKaaqhrqnW+zU63LAmVb6d3PAyWfdug+FxM0diCAFrywRXMVZ9U1Sb5BdXLWecxZXO
hG3sTwa5wkOmqgQBbyDbEG/ESWyWpzeE0g4NRGjQnNQ0jkRdrO0TbTlM4mwcNn+3fhrhh/9lRLAd
MW6G2MQq588jik0PCDySNhECghDypxB4rUHhNKybOM/HHxXIJEwE2p67fdYl1CdHycPdAyjT2iyl
9IQc60tKzJKpCv/64u0NR+/fEZVPvzJa+3q84N/gsClQj8VnXOSxpN8m6mMGZNKFn4b6OBCC6bod
V2uFZQzRYrLHIe9RcGZENQlnp4RAR1AKgHsfQRpxTF43sk1VV8oDJfCJrTnMTiK+GPxmQo/kC22u
I2cLbKollMxXkhwoRnZw7wdWCjJjzRMveXrnUMbll6pwoVsBp4TIGVJGyLX/IrDh92+cvR0S0oRJ
/OTlh2m7VIuwSxar46k034eorzZw28In2KatgndE5aYTvRfjg0VOmvbC/y6VdXRBBDVilHJj74b0
/u6VFtwUpW5B3XbmgWoLazXgLSoXA5C+k5rqHFd6DpxDnXQ8pdrQWC0qH2mHUD7cHEci00NOJNo/
484IO3zYaYOPVZ5a76uMU5gfw1HFlNpWU1qYrQu/tmF3gUzI93Ir0wA8o2TH25bxC6TfD7eY2jL5
Qj+ztN2HS/HxyxDJYZ5XGb1fUIAn07NHOC0j48PbN9b/fZHOumeqhn+0E/Ic2cq9OEaFjETF6RW8
j0To+s/4HMs4rjzbUyBZ7ybuNhMqaYUCRpFctoz3KcjzZEf+Lpc32kCrimH1WSs5dpmbCgC4UMHP
PGVbCUFNTDyUZSEoeWGyjtjXsqFYIbaWBvxr2lLnRfTQwTmojXodLhk67+QeIUvRGDg0bF7d69wX
mwhmgcMCDNg0m9xIWq3U0C0NXHPHZMsbBA4BtAsZDmLEgah1kSbH+UaAuCfMv1uo5jP/sqr+Gfjx
wWwukdcbj0r8M8CtSvbHwcvNLzR634bexgitykZ5BotAeiuKTFBoFJxF91ZwghYSxXDNd/fiqAsm
sowhzIcsHuJNX/9GruZoDjnLqUgiQIQYhHxSji2Qhs/J2Va8n3e9m/2DKxTaWPguSYyVJWmxRAsV
0bqgTk33gvxRiTz1FXVEBmAZ12W+bvtiVGRJ9kTNm4CQMbzQ1N+XZJ+lN/kl95OoB2njoUfhLIWU
Qsw6vfdBkCd+t0jM8Hgd0Ga6/kODImsWSGDKRyA/tXogwh8GAjoPi78XHBpm57N8+sg4o/W9LtgU
vixvfdatY8vzdkFYcUDgxXlQre65QGauU4xmKYfAmbAFHpHxhNt8TJFTa7cdvc9pEp7k15kiR+s5
O/RwR20F23UjkcIQFSycrNtnsgS8IMMjll0k7M5yD+18pqws+7VpFhp824STNdZha3GY5UFcUweZ
dEhhJy7E7YbNeOz1/a8V0gzxcTynkaMcpIVDvd6Gvt5NLbaPggb+2+guQlNaz6CgubTUlypwioj2
5GjA84W9XwIUlHBPaPyQa4dMStScxSrEKlz3BEP+n45IwmrDTMsHOOtfjkwwI3RAiN0NSAa8b+kR
hOAJsHAr3Okpbtlw+buMJVTJLWqMaFvMZfyavzSZIQfNFNsvWX0qMSn6+iwH8/dE/QCnD0U4Z5mW
R/93HhMn+BbbJj7PxN3bQl6DOcrwZPVEYYgeyuHkVPxEwWuBt3rdVYr09NkOU2laTEZJYM2yYrXs
BWY2UP9UGIgemBRMocOkfH7rXJu46crm7aZ6iGvPF0NYietQzIcZvU7thZgzI77zMfILHJxyYlaf
xxCi+r8pT1hXgy8z3VQ3kessylVLJ2VYXi9abgO6z8IYYnUh5mKOt4bHTMnfuF9e4Mm7O7SIXiOb
VUOiug4wehAJ7rAllvUlSApmpUY4bSceTX33+TDy1nj9BvkpXCNr+cQDVn6+5JBtHJaqN4eMYgZt
cbDHQDPSOerYb/CBurD6fTtHWcgrR90VHidMOQiYgO4cWZUhP0c6CUodSiUfN5D0SkuSlCVFae1X
sOS3f5SJzC0di7QJxSAXF8UQX2Kp7zPRqNJpCg3QDpVumvsvVt1OYI0ORIqEGsp6UqNAxlTku5gN
vrgR42adHTzV8uOO1ATCqaOXzl2tjdrTK1EZTq4DejfPUtAcRcxDhx1ZzYVB+fA/4qgyteAleazS
FqdtvqnjJY2HF6GuveJJXoM7OxWGxiFEXsrP83smRmpZbN4Zlxu4ValgESf3MMEvtTRnGCbMJEGt
wvMPqxrxVVRbheOtGLN3AYrBLq0k7nYH7R2CefIXVvn8UlD/ZhlbwmcLhV49YcURYxYRq7rHRziH
sOSIqLEoaoJAVn4peJp1fFd02ZeOeDepKpVdphbVeJ5cv0VCkbSpXGQtaNYuhEdzP70Ovs3LEvQl
x43udUMbbMWoCbPk1OH3LIcaiubraaVEcNiDvxlDKZg/0xw3G1VwaLVtKpJ6dYmcnlGhvTTXLK6g
1XBRl9cFCEh7vHKBXx07u32ZrRDknf1C1r5iCkgr7rpWKWaVmHKeCaB/m4jC8R+qFJpJU9HCvIBF
yWBL/vA3bmjsyIm0B2rdynHGx4JFz4PTkd4m4QJAtMRqt1X0YGw2A3U+Ns9lNc6KJRp0gYb2kqtD
Ya1GEs+gJxDld1cuXlQnn/LJ53ff9wHG4U3/sVYH9aRbYYERZIVWr09UweTfn+2Lyo5uKVD/ARm8
Eq8lT9y4FO687gfuGk36nFbVB1DhxE9+cXNgjSLRmiE8hg8TdMRC5zLMYeoG1JMjKBm4BWLIe4qu
BPrAyYedUQy0yqSWPqyMNckn8ggGP5qFhoensfx470x+yQmbyNHWLBydfguKVtLpuYmngcOvLbBL
Z+cPnQQlJvc/EIuQNeaOXvi/Yn83O86+2h8S9jbAj9ijIh7+nEU6OTsIOl6jvn273ZWCwGjZeYM7
pKp7z78W1TCg8elOI1GUQZg7A2oOScVwVLO9nnoVzSiE8lMdMWbkSiz4nfH+DwTVjP++kmezI4R+
nCUXkk0O9Xn4BFWd7qOxo4lPiIkzPlJE6bW7ui2ykqqY+L6gRlpnKQHijkv3CL722iSwTWjHQnNh
oxd0qVfWlDyZSOG4cLXYWVf0/fb02XW37UtcUG/jr8P0tFmOvQKDF8E7GnNItr1LguCj5LV+vpjT
aVJXOO3DLabrl7MUQVWMHqBsCE6eHOYEyDqM21TisPwuoDdnOjLMrsdsaPphwc4LYi6fKZ3lrFol
W0UG6rRAt5P6AcmYec8tkUieQB6yk/sRwe8MdchKTpMNBpLyu6M+s2YvF5gJ2UA4HXqrnOwhUPmT
3K2q7+ib7asKan3kVdgys4w6O5GofVgMOoxx10M4MvPrUaHsCPBywgzobSMDMnETaWSKP+pX8QN2
DMc2fInVQ0in2lfdcqS356hjXh1Eatcolo9+vO8GH3ijPrGzLLTjE2PECUB5vVZFUe/i25/Eswq5
cGmj+4/mXjSOe0LzGoP8i+EnDaj68s9Ll+EMfqOx5vSdacQuz6pqaKLGNn+LCE233nH45g3/XlVd
8LdAHdTdGVwymD7blGR1Da2Kn6PNbuyklkn/mFIP+YUW3qKDfoIAk2d6vsbTIBvWw+J1SAZqNrGY
1+OWZPK5mByWkGVS3WrsXvtevwan/uQ8qy0SyALmUR0OxmF/TeFK+NYP8/hm6iK9VzON34sAl2GP
1YUj2MW6jkI/pHIIr7KGX2sYovOcGaWrPeWj6cW8QNPdPSvXFINn593WyuzTLPLn9ksMOUb0fefJ
jzc4CkfiBCX9idPoskQCBGaN2vv+gVcGfy6Sxjb2b1WugMRyASBSMSNtMTpMmTktyvu+gEBjlnWI
yn189e40Q3O7D/mDV65HS5/eUaaekuTSFCo8+bBsa0uYSfy9FIl2CXed8ihdcnIr9w6SGvoozYbn
v7k5pUC88mITxiv7sywlyeG44XRp2wHIS2y4vwsBPCkr45rexTON//rq8vyZJCWqFIBPfVEU+BLZ
BI/9pM9UBWOZweCON9wAu4LEGLo5Apobz+C2xF9YFIr/hRRH9uGCs/qQoL1iMDvBZAwyw0Uli8lu
urD2LbUmbu0WYfzbOQYH7KESkOH1WR2xFqSA2+anhxekJYep5rUEAPQc4OGJE8P69Tu6Cj8Axq8Q
Oi+/WMKZ2zsw1zi/eyij1m2iBtX+e6qta4rKfCQFupnOnHiLChZtSTyfeHcXernFT0pZgFdlsUe3
Z+8ATH2yxtark96Tih0zznVol2rLnDqC+RNZGLeGGYbrcmFsuzupn7Ws4OdSpS9r5K/uXzoUEotp
VOTVD4s66h3FdZlgb9C+rlNQCii4fJ3uoANolU5uWjx8OJEV4lrHeDydvBr8l5y6pavlzADLolNg
xKPKp06PdHHGysAJSuDiX++FxEqDwfeQTs/Li/v8mtxXiKXAiU9vtrmHTHofqaEOCZGp33eEzi4W
OMLtfL0FYk+h/93h87YAEldnKx8m7rWUJOI7OhyojWu7xypxQlsQagR+U3WYmzXS7vRAXI4JuuHz
GjvFyyjcbUBdP6Oq78jYlnhyGZ9HuNolhApBFckByGw/HW8vFnOy9dAeqecMhAlzKRBMhGXdRXvm
48dLsb/Z0ut0thyI59g+2/kBwWH52Wfmw5+1QHQK1ScYrgQArgt2arT8qVBmzyhW7Si9mcLz27+H
HXN/oHWqlZ4K1uqg5Xfup4Xd2b+jUdhrMMMiYVeCN03EqY2F5iNFatB2YdlN4YhBDqjQ3BgrF8KZ
ddQjGbBQ57Bni1KhJIsdUtB8cm+n4hEe1OsrlgJsRcXdPSwXCEaWxbwgrRdDJJC4dN0X1M2/I14/
b7+k8qtWKrJThpLQ1T5gJJcWPTlyRqA33qNmYcsokoJ/7iYJSMf6x8nmXp6D53GY0rV8O4Z4rVD/
tqoJEN6FHD+uvl54TQZAETwlCKAImpkazHe0BIUfKdUxzItDr3CnfVkh5BPfHsYwH9A4jJi/KrZv
mGPxu53jLgfGpoGy8y7vg95a37GOlPdFZ+uFRhUGFv3m20O5+Ltd5GilkgO7o+EUy33xAr/SnYGX
5ZNebBIpIUZKYKvHGozMqJ7Qq9mmFLSkST8VmunJop9WctFO8UcyuKr4OyCxi1UgSq3vn/C3hV6q
DvucndFdI3ib1NMt1V/e5U67iHq9AEdkyjS952R/0rRMDWXuPmyq5jPNEV4oabwCNO0FfzZ3vb/o
8AuiWFfm65p4qxdOSjFSr1HtPbnZiSR7HNyVvslsLFm1YOPrzozLkSAj6JCmUjEcn513KgU/qWiG
Rejsaoc71jV+nXBbpBtUyxFXNtnGU241XHS4fEiP9X2MlBsAniChsEx2Am/UZPIPxAezuc0TQDsI
AJR98HLXePSb1h03w5isajR1QnUIExtXJO1P291DPv+A/LfEHkn7E8Jzjv6gR6Z+5UNui1jJXWuN
7Onz/FcCVxWSnfH6WMFoj1w2k0Vb9PyO1GXf7uzlM9pIsy3dcwE6iinExViUIV/+bWJ+pbYXDQJW
WKKfQtBOmMrcYe/LoxAaVgCJAMxokuPFIyqxhYgDsPtttQ0QlQJS1Qki/H6I1R3rWgHjzitS6l1N
Y9wtlGtTR7P8AjWepqYlf2aELu7IXYo1CxTcktOeBzcp4QJyb9/jUeZrBscPiQyVfjH6sCvsrr/8
hnc1t9YadPWd4fMLELm2wsRRsynHC1g1XRvT/nW2cVegwKCfOvvhKVKNxYoGRrxbdJ6Pg/dalv0v
1niRisfFZzYRBuBG9m6Sc4z6MmgLXkqDvj4ui1qZa6UZlonNLTPa7S8JXLEV4MiEMoLuzP0oXxMO
vh+p//QgdqjUcu55h2IoaQjf8xqNt1I1nFbOgKM3WKP1SWHHSwojgZe7E5WBP+njKIY5wOddOl/H
IHtkz/hNfHiXi9I0FubzMiPtXXcjKN2CUeekaLSWlP1k736JadML4EHffgsAA8Remq9qeEDnUXph
8RQMJH2EYuP2a69P0AArBOkBpp5VD0U+Nm+Hed7OiyT22rJDaJyNItz1QXR8kd8/avRynh1o1o4v
k6Cs3iqM1v8j8hiqMunCnJAq2uNstCAk/sgZpbzT6+YKNV2XaiigKeq2E4NsfG/h4bDonTOSlkpf
Acera173/qbwj+KDHzDrNUdsNDesJXlsDD/8qS7eppmRodIAQNnJ/1aNwWejpxHukDICdjJ0/vRo
gvsdqG2fU3FXpYf64ORyozG/xTh55JHCE1u+QKd7vX9etjPBMMpNzpfP4V8b8tD6TNOBB3nvQMDl
KemJqm0vaVTJDQsGiy9t65yV1QhiA7MFHHqtLMq2fTQEh8zQyc5+ZrtVwuUNqHvPjiYO3FewfEfo
Jh5mMRwkhsiq7weUC+0pU6q/yt5WDXtIoekamsrhA4w3uuUaJShDxq0W8y9q5bBzr/xaYNPrwL43
73iLA8g69BS5hspQDF6e76Axj5e+Ya2ku3HWRWhWAS0JT/P+nY1bo7VEYPx3ivgaoExJhhOVe+BG
Qr20lCBNV4jM0RKPFFhRTCjYeFty3e1lvXZ42o00/E6JxVjpj5LWcx0z9dS2YbS+ghZSyhovAWtv
VGV73wFPVcV04zZc774akIaK7OMEeUs8kFUKqhF2cCL3G/jVh9zxQYCDRkqz01OHBH6WObCJTNSp
i3yw/BwtOQxu2Ne2wAMLvyK/SpBFlMUOHAY9yCkwXj8jHTX8HORYJELHHR4nmfa2GbijNVQy8EK3
FlQfZEu6t2DXK9QSXemdt6SmTZrxDK3R6Rkp/lO97ftOo6eJOBiH5DlXlH46qkJzjxEPvChJHGjq
naPBPjjhm2epeLEt/kZdDxU9evYoN26fn42hogRANnru8FQjtNGtQzzL+oVo7A3m9EDmm3oqfYyx
oCAMq3uOu5SIMmMXZ58Hn4q19ZDFScp9g7eDSTOKfSLAjFIboTsbqnxJapyqydP0HuZAdUXbRWyD
SmjC+KN7hd+U3hXsLvD5LQsaaoBWOLToGgVSfW3oXN99bZq8PoTnq0RC9QbHhKQnl/1UIuwb4MsH
waLNkAZ7aSr3eR6yLOZ276WIpZbAtsDOPFWCX4gVR02Lyt03yJUledvBLMbn0oUPr0IIVkNJOljD
vYF2/yaBptxQlQELP50mofyGLBeI6p2ygPyxuycCuQtngQZLTKYzJiGQR+U9Pc0gEAz+LWBXVD4X
9IvaNJE9jNaJnXAxUXD9x/3r6US8p+hiuFPvZKdbNEFUYDFW3HJz03dI+htLVpPu4bggDxy5jJMO
m4K4UtzchH32FE35nP34vygaq57KogvuABFG2EsmsIB/c9R1BN0pE8goLATmKbkAFezyCTxjdVXS
grNAxS0Zf1Mz3chWqbFFyu2zdngFVKkXSZBzTQmPmDuAovqmCVsNR3KQyRFcUbh1qF91XTKqiA0M
uOIQMD495qqGuC9WYfGg6cMkj/F8vGhRrPuE4c7+eO+B+RJr1I2Yh71DQcnzJ+MjvO/PgSGYBw7H
s4JPkR7Y60EMZf7rXdkHhuNsHMTcYyQs9jdsUhawB/J1jYEM68PdnUHfAEYctNL3yAlTGN8Hm/Zj
JTSQHFh9LTxryxCx3UWGCyly8I7MNTeIgRXLjSU8QXEw0SvhTFoP0tZDSlD3ZYDsERGECznzp5pX
z6OJqHoYmSm87vuZYltFfzEi2cjsPOmeQ0g4v8U2/z0AbLKZp/n3RBw7lUp2r8kl0ir8Zur6qzds
I5b4N1N+HmlUXvUn6Zt9HqFKpRNDRvZwAuLiKlg/yz0ENy8TNpAbVoFJOVyKmB6jrpHH4NNejIIT
/3dm+/qVdC/VsWhKRcHNqWL7/QXwSLQjRG5f0BYFjEZ4AZ4UnpbXURA3/hwUf03ugR/EnwrBBJk/
PKvciVhqMNNxM0rnAj73JOSoQ/zphqwlS2GV99Sfr0N3yPZDeVY3JbGzONVsGpbatzJG8ex51eIl
Gtlvo29ID7HeS5A4mGk3e368QPaXohs305o0abTAyn+xYcp6QCg9JmSHan0qIrTWwLVmbdOCxO7G
OYbpeiQhMXZAP8QbssYNS+0P2wha3UseEAXDtt6f9XLa8DQFz/uAuQBPaNTZQBbMr2f8gZLIiioH
0cV5C1ipdNbO6+bg4Q6EOKXOyY8f4JmeS/bODyrsorKCc/y/bV9iSli6teif/3nud2VtVeyAJ0sT
9FE/LW/hbUynpHu4cju355Dw+B7UcwSg7xJh6D9D4pVq3cda+K3qZNxK9UdjWnKL5gd0oPfQ2/EJ
8sRWp83HLWT9XCe0bdpXmqPje5ieMNA71ob8BBuCr6mXKpZJQVV5k+kYRk3h4fP8Njo/f4dZqRMv
5YK0LmxfBCYYnejH1qLBTQljdS0tB7N93pM3KmrgdVqL3+Q8wmYvV8IAvwDKMYFIhNzRBfZSAC6n
+ASu8ogb3dt18C2k3MQVJJZTKXYYagZ29aCloFOMhoynbDjBv2zmpuW4nxVdbEIN2aL7p5vCaDCp
y7ZfedWIdOVylhZ9DlJ+ldwvCKl17tMcouMvRi0+byr2NaIIIrbV6XKZsNzgjEsxJ2+bSGrKNalJ
V1p66lVWc/J7FejM/de0m4qojUTTVfFKDgi83OuryP9bxa1wkkdmTSA4jBy1DA8Td8ZNtalMUIQY
eDaF/+SVZWzYPxjUkgsPjkKzAZVb75FqXZEIJuGnHIKQz+d7n+hDnexRrxmhMmLHA7uunnxsHXa7
ubIAi9OGTq5p5YDNCwlfw2s/mZyTOrc2EfC33SLWOuk5wcIw7sYvlZv5TOmzj095bnHXWrbI7/aP
WsaplTobTnsg+4nzIBQfXJrtG8uizE3i2JIml6HjfrpnqqGaontO1qlnCLHLxi0IvzmugVXSJvUP
w2Rh9F8dmgFi4iSh5HtjKFfIq+aEVSPfrwl5OSMxfEupkkIYjWiEyq+x3/1A86wjZdThFmzDGF+S
pLzyCKpdkA+i1CZtO3xBZr/djNIH8JFFXEDuQwZ6fI0WYVdU+CaonRL6YR6iG0EnzNzd+dYT0elA
CwDm6R1YuRoRP88yovxZTeFGjWwwVZeEb8AAAVv4gQmXAWXoBOGM7MXy9bov85vlb6QYbmuYdi2a
ZvZ7LMMfCTbn4sGh/Z0SQuMggmo4xyRGF+iCx7uoyYpAvlXFleqcr+xfbKeIMU43qpVd3Bqqpv2G
LPv0D3CWrr50zEAsq/t4A0fSz/L6fFgAjjACO2dG4vdKR2+f9asBfLAoIScQV1HLOUFf17G5VFpq
CT1wkMBpJJGqylr+j2QWWkVwNLmoqIdp5LfFlEbq1w+lH07NKhwleNE/FJ2OSKgJI/FuSE+vyhku
lMjcCSL1fCPeOjU5Gc74sNSPPHG89yx7T3qoqZBi22We5difjxG4v+5BNB/kHGzXHIrGiiReB91Y
VTPnBeSwWOChi0lXWRcSBzuuhHLHBdNOuVDZi3qhP04hH27cpozEnnfpUi1UFM1PV7d5VR7hcFU5
wx072Z13XCO9wUgpo6wU7n4ABdu/Oks0ma5OYrHZWc5V6cL6bixROnwGA/01luiMZ8j30UKfHYhm
LD3NhglHDxCWuifAfS8lSFYelW/UtY6AKIYyUCZgaVuv+tZhYllaaKq7M7UMpMfNwtlxeXIjkQKS
RuI1lNuY6mmNbvLUzBKYO1Abp5+CYUKDbWKcjmZ/6vyaT4sYKSKivu60sUe8h+PlterN73GEhR4Z
R8cLuRf0OYf3sLKocZ64XpBsB473nPbzhXsiufQ7Bj4JEjx1qCW3zscYF3JO0bdqZcWdR9n43tYY
/HE6ysOVwG/t97bOAZ5ppBhmjkW/n+WMwu/xotW4YXGX4S3BUpdVm0vS6fKSwY+LNZa028T65CMX
6qARzU1dfuWaEovvaYL0fUNVtG98D42YLNUmjuYWtEuxtybNnMnNcoBMdeOiz2BudfAEglrOMeSp
+TUylr/1dD2qY9SAqWsJRRF2aSKu3bWg4we4fnM2tTmhajP1fbMX65+pdZL57knEQZtvE8W0v86B
l/89s0Re0PNQsxPkfc1ikPuWUS559YCrG7SjIl0PinpLZxOqx1dY13s3yXOrRn1RgHYrEcEShVFK
gOA8guGSXzhrorbenSWI7THYYWfmaI1E4gg0uZyha9sJ2D31f6hQIIjRo4WVVtDjpT2WYrBJnL9z
oITPr7yGf4hNK0ENRpHxTz5aqzx9ByC027tiTpquHsMAcLaRzUA7yl3ZySqP0ySX3T1Mu60KrOnw
OejxaqMN5529mgSi9oeLbcxC13GlnFVTOv8Xn5XN6+x+d8Z3NBTSUqyY8Z4/fzBaEbx+1FFh4MV2
9e1DNBY0pmif/KJ0OJjCDKU+1kKj6R7OVbBBcx9WJLG3ZaokFz8RjgXuRYPHt7lXk4HY7XiSd53T
3Wbbe1zCDDb6BdwkPax0acvti839OErURSwBoh0BoiDizASFemZ5A+Mau5uR1EQ6jJqvyBp1wbd3
Yka/1+dnzQXMmioGNz1SDhCWP4Cb/HpSpEGkBKt/yOB7Tgrm/cfZ7EAQVoYAvA+nRKYrDZAiPLds
0RzBlfahjlqxHh8OgK++tsRJC820g+myvAXUPw0VQJ8uJvTRHmiNxWtXFUi/zZVzzyo2ASCB2Lfk
X/Mbgaf+4oJR9pHR+xIPS2z3BJHp4hPXUeOAW41KgMBKtpiK9lSoq4rJcVyynA+VP94SM2pjOVEa
yK4u5+LqUNdS4O1svAGik2veHz5sIVnK3wZ5UflGB2flHaga9M0a8QkL0lCwmyuyJr16EmOAca4n
pjXq+c1Ac8QWYjtYT39ry4lCMQE4wvRpsszyd18pjxlUrynxFM43x2bTK2kpS2c1Jv98Gx2cqoRe
NTG6a4iuHgvhgrz5ZJQwUsUP52/foMfg6ecdbQqDKr4NaI/HTVcPAxxnBiLWRjeOqLHLy3lkeu3L
5w87yFhpAw/NHvDF2wZ4ROoRYI77rja6SoGn6M50Gav4twOKeSmBHx/ftghuoFzM95cVsViwRqyb
LCbfmEs+sSfHqBBkiTUeStHRbvLfOM7cfS4mwdHycMYX0lCngMBI5ESohY92Htl0EHXizahJG/vn
jm6InP6qipf7BkiholQZYJ2BNCU6UwvHBVQTgOBHLj9ZwybAplmRlJkVqE1ivHhD0m+bOmBM8zLF
+v8oYB+MDE/m2EjqwhvIFhRhMBJhhbHf7iRs0cc0wJgn9v5pTsQz6dbCHnJr6/E00AROWqs9Pq4c
kn1rUZ96Pjd7qGry/sepgEnxqaMFylYrCxG63SavQe70v92ZzEBZL4W+wkT97Mhgj4NtLsrXww+y
Z6rRLtluv+keoxkqHOCMkEF3rbhZMrGuwPwGYJki02ytpkFT9YlxatHGh5b3BLytkHTCIgqdQgXJ
WJQn1K+PQLO4Jp2XsdaoH91EBzS5HQN7J+ww3TtSkTOhGA/KDUd+b81/q15fj16ixPNFoQxvRGzs
qOf1Z1RADZKX5v9+4iWqNgfJciBcSZB0eJgNzR0jSheZPfvJjGjEVQ37STLIAQobYvEi4jFINx7E
skJHUSf2we/FrzWRvWtqMvIXNLPL31dAEfE16/yDNceJGbnG8efiO5foApJexHaHBSzK0OhuV/k2
KJhsPTERv1W3qHJPWtcDwf5Ad9HaYHhxVj/2g3utu30QxTn4OiRhuRHRd+CFh7psLVFQDqpYNbWB
FGWz8zspZzTdvFOIJleS9Qve+eGRnCX7iXhfk1x6miC5mKHWgUWDqStXqxRPL2Ta6STPIRBTat41
E0h2AJ019s7b0aMbzGsB0mkuXvbN+apk6rn6rkd5yqEJ0BbdgVWsCOQLRJWJqT9VBtz3SWuum2fo
Lrp8VPgyX8cHc98oLGt6155IrlRT2flRm4uDwP8qMP93NOzJwXRZBby8u4/GsqZt7XYniX79OjKU
pRdPCoYsREfXELhdsPxn7rgJ5Y8JhRAxdmTUg1QoLfBbqCBNEzo8vHlQJqkIl1JXhvMGWv7vafSg
e6KkFyWZ6P0OO+It0D0UPfRWuqwjtunI3VUAnBx4oE5bjwo5C/TlXU5t+kEvryL4X0Jbu4/N9tZR
hhIYAhn/Sn5GZifuoc1gdBwZDkV8p884BkVwPl1gpKwmRYl0H162RyO8KiPNFpPLt9IZwVy4lchE
2cnMWcUhqenpIMIQyE4rprs2U2OKSPom2ay0WR8VWqMYKu8Cb+n0vdKkFFMwO+of3rkV2YpbBbhV
SI+7fqOhcL7M3TYDvqSw20sv4EHSbMTgOkbxnmUqbsS1O0jjZjTTO+c36xMxWyPapefPy7N1sagM
jeceaWAWbDR1zLo0YPRJNvSqW8x3t9xFEBfDW8t99h80np29PqHosKC4YF4t20/nLIPndyEMiDkF
tc9BRszn83NnIE/pDRGtTBDYRBngSKwTrOxaiQ1L7tgW8O+pw6/dwUQKs555pLbncXMPlhLvlj7w
jk4Mzq+VUZo78iMdmOZkNQZK89e7/ZatP90p8AUOM5e/XOc+8TGhpzh4YSYZQeHM6WRNhGL1p4P7
wvCfL3s9ULYh6VoEOdgKK54CbXAgxCGkbR+rkYPBTorQefcGCa+46hG+bs9Z9kplSu1smjhNkr+2
nVhZfgyw+Uv0C57yK1WfzedbH6v92A45HJHoUu/Y3TfugERugoXarJdKypT6jcIHSwVTjZV/lrF5
H4sBUHMnwAfJbPusnP8oXAVm43S+iGoIAllsekbJs2aHbFyFnYw5+tjU/hKIw4/n0s00+qQc/+iO
vZFz8OCyl9ljQ/95Hwjr9WDT1WWZv/mKwAorm3c/NDZM0TY6n4K/ocfYSzokfB3ODSZ9hPWEnQbi
vIYq3UWCbVpG8efEhl6GbP8vofVkdEsLAJqymo1a8Uirpmax7gTaX2GveO5DGINV2HUpSPgp6wJa
201WvA3o1MU0oDVFphnwNmCCu2h5oo2iqdKeOYmF2edv/nlfWFLail0DKVhD2kFj1JHEEa6niGSj
wVCCY1L7xhHkK+To34OpUnqXjZa9JG9wIrU2RFcZkrZ6fTmav+cxyrFF8Eo0yF9jNM46Jpr8evTe
bKCO19Wk3LgPvDJr2CDjfLe/FRnhw19KllY8deqeZppW4iFN8GFNPvQwS4S45YyeoKMBx3yhs1ht
9jPjmO1DDEvjiYb73/uyxYLq0+f3IPxKhmOwfQVdOYSKIFucayv5iPw2mUYDFfaPyWdciklHjdMo
9qHD5iIRNXSeHJu7aMC/PVcPWcSqUFZbA5VAf4pUNrUvN+23AMOBPqh6hN+uQ3kBPfYoNuAgvV9P
Zg/AyrtIewXEBxYPXAslEoeZhPHTGhYPxSjmoXVmMMUqtDxumxcH1OMxZko/ePnogkvyRfcieFOj
+yEKHd+79DyC/uHMDmMAhSRr9Ckwpz5v4DvjjJYBPAdM5X6hs45mqoGzchN80t6EthEr/J6qUl2l
BVpo92VekdVuvD7V6NtUNcaQaw2hnD3BdWp+JUTdMPN39NlwTW6O9t+lIT00ZHSGHutjJbwPIOMB
ZuW5IMDFIk/p/M7jtCXkxHQJm4wlPrsRlrYN/wFEDn75yIWsBoCEwCJpSYOVs107anMshSf6ppm5
fCtHwqT+cZMGWArSeSh5/QNth8ma8ou54q5OukgTzK1Txx/5z1uzn1MvpMooQ8U2Pcon+xIFq1pO
Mc9l9cBJnfDKtZzMSbWnFfo+4mxKdDd8suYMvuUtZ1nG4JGy4pHoNC8m0qbvCW86ekOOXjCh/lca
lXUoF4iggpL6ApoiN0cvt8lDjgavEGtK/Wwnh7PfeoyTE/uQMxqFQE58+NDLhgQBraOl/QLtmNwg
ji68k7NxKBv4o7oXAh8YXXhQZmBisRz6QsMrTjiC6a9Nin1K5T7mhCqdO6SVBx3L6qDouXd1Cbmf
4qnCAnKB7ZyRehaFAbHO4ZjuDO0uAORN+q7vRxBqnxl4n7O5sSevlslOepvLSKxg6P1Wk8n92X6T
hIOIIhvClD/zZDY5bZbzgLAbHvqAGU2tjhKMyyet4j8sIYxdyozGkmNoqS4prCsv9dSsMKN02YQf
9LW/bxQvaMOobLctkHYHc6DHdeuVVGBU67mfCgFUzB3Mj2bn0DJZ4AWiV2xewmJUmCueURwC9D1W
uWFLfLB/CstZq86wnSqlYfIlGTre/ksVvqgOXx0x77qrh6v24JHtao9XLnx5rW5LjZvk5/PKjVbf
BJEMfYFIk006ssQtqZRkqcZIyyiI+aJ+oWt9KzvIqkjg0CTaVJtUi7oufqZ0zZiIYH1JRbUXzb4Z
B9IvZjbtyO7tTvBN7/7R4NhIIMuSHDKtQ4J7fU58oqXeWK1+ijHyfHKQ4ahNYoPEf4iRChJD977y
Bt+GWsEMpQLsHjQwPYMmSMpzprQzbklO1VNhEectCTHjvSmbCdKAie0UolIBtsmonroZ/8FmfmxM
VfPqHMk6hnPCN+s1wRGy1pl3hiOTf+Z+cJWv1vLjoCx6Q5vIJh+bI2yXTl8maJiypsnDDnaSntkv
+/s91e8DLQ6Dz/4u0q0UVeznqEEEhg//hZGhFV5gmCvKr0+gfORAEpRpwUC6DLM35/FK9pug48sg
nCMQmB9cmfq2X8VUX0mT3cqUHShFgEal8HTHspmbGGIDZK/sHkYXn2R/9jKF1RAaSqJEAV/G4Niz
TswerFIsimcE7CYbJwNlmMSm4NCKUeoSrUe33OKWOsjuDsMpz2ytgeZLNlWM5GScs9k2gcaDcq+M
CHdwdwY4Lp6Vo5xJGZb8tQRQFXf3ZEisSfJt2C2Mgik/5MtjWjNiDPt6SKRLRKk5zR47EJpB6US4
S3tmI1Swy15Gn7lTZ1ZUYyJGTjD3zgDalHsY9uM1L9YaEyAF2NoqeENnMksQE9hsbUGWpKTxhz38
rxKLm5kdwpmNpouXfOiy5vN7FrgAJzQMR2HyJuqq1KBO2S56Ols9D32/bxAFuWx2bciRUlUwAeVv
la0hACw7yLTlkevuj22CQ4K9ORp6H71K640oJc0X1vexwPz2ysu7UpxBkTB0afTF1qcTQwldtg1M
X+0IfnYpHMusi5n/9ok3kK+XlAvI9RT04jfoDjH7gxwoakJ1rRzmHlwNk0KaNVygNXVHdxoquh6B
iTXeT5cthhoLuf3OobG2AcSraP8z7OWCYq2ZjoTsN7G1J09+WLcp1YFRsLiRnAzB7i/rvMbwIoPA
9u1wuENyaFyXwzN0giq4fDurVNEdsZ0+PlZf3RLAxb77JRiCduS+hO+e9YsgejxSvhq1YZUpohjI
S5SN/zoQpyqJ/d1nXhfdUeA9sVN5WpwZFfFyqH7fj2vvfmLFPJ3Yk1TKlEUSuaf/MH9KB9VKmZR4
mBvwSI3VYlIPa3nFQ21KHm02E0S/cyLT6xet0jod/FiCxJZPwMxJDZmnbOcAGytOjNQfy8fQeVsN
DoR/PQROMXrOhxl0p62b5I16kn7HkmYFpXrPJCriFThAW7sRop10bsYad6wgvuUZAVWqEyUBPjRb
iUEsaShCWGZSwx9dmx8E1j5myT5VDKUYjAgPgKAxNmGkP5d3zxhHxSmVecQPiOKl1U/7rNHuOw0i
pQj0MJcNMmqNekSf4tixQA67I4O02KAWCa3Zy2Z3N8zY1dwnW9S6LZ3xBsxHNcIe0XDQl74udCT6
Gpj40y1wzvIYU1aT15ldjKTM0s/Ojh6YOy6h32E84Z0NEEFK+xIJyAslnEdwLltgQ6tS5goOYeEt
Rx0qOQ6ic5zdAW2wzl1qHsgtg62AaDVd8z/Hw2NfeN9reEMY3FEWweFr7BtoEhd/UaCCw/Vd4US7
BYYopZF4cCBmcULxN41LPnGwCK2VNUcW8rSmaA1IGzH035cl2OWXN80FhpgiENLMTTvUW3zT5cbO
5KypygWykt9BSj5OrPA07ss5kaFA8P2E/23sO/6bMx6AOpfpiV3r63VE+ysBVkNYAl4dqN8HMRwv
bmScnVU6V28dbbla4gXYKVGr7+PG7ryaQKyse8KJaCMzQhOYzECpKZ2Wipg7VIPCr9q7L4AAluty
U88GKBj/oTwV+ZwKze9PNOuFzdZW2sri3p/IXdWzuUnamviTLZo9Ft8rZBqqkmuSOrjZAIkw1/S7
ThG3EbvbzN0n+t7n8DKHCwW6wym0lqErbuhy6ByjWhheOfSrc9hg0RKJKbkxaD+Sy5vHrpZffe+K
fRjAIonaxo3Y1vhrnceZaYVYyRsQFZOxv2bVHnPgBQn5aKfN4cQCSiGwQPoOkz+34yz26yfdhQ/V
gDJnC0/8n6yRLfkjhv6bHPptg450Ei/rnWfHvxzFvkQar0lr6NXJffBBjR4Dw7ERq1PNuqG59SMN
YAjZToQl1hdMLA5igInsHkIOM+LX3mv+SHVXLx21kdMD+CSyYTwXxQhCu5AZjpPZ+RcJeaQQCe26
h+zn/lgFcFrchVuyaKxTviqKyb7ctjj+euIu2AqEheizY+iEq3on23p4Mn0ui5u0UjHzFQViXGkT
QpjmbFuJbL7UaZKIXoY4pXBYZ7IFPZ8lyW4CAUu31YP7oI8BeS7P5BhnjflHC76vqHRDlL30yXNq
TDN/RpXnj/QsUPMUMUpcHtU80CvGMK3HVTRR0Cs7xk24vINcsur3mi3i4Rb55v9+KmxMH3BjkQSi
+JQkI8B15Vhl8ziQmnwQ5MqwQExrLcAq9ySSnMF2vlUos6CufkCibnEUH4Maj/F8Z6ShsgAS8lTH
T9aMSAWwyInoeJ5NFb6q2xaso1OQrpVKBkI87EVEuaPI9VWO0gUz9ilfNPK6Y6DPCKTMI92am08k
h2tZ1RqO9t9To2+3bYWtW6aFPwku77WTLFfwZz4TbvccYEqcQNqouBu+MzLRTAv9QZEVjBmoP9uF
4QY/M7GDhWlHu0aiIm+8EE9scvk3RcmdUwqy3NWa/xuPgPi4kakBf9yvExszq42DXOHXB23hdVMO
yzPLpcO9IvQjPaPWWwsmO48N+vyoiWPSC3qz7FnLq3mW2a5jYlYVjIWeZE2JZBffhgUbczkvD1wM
y6hZwrQhxGlKo87t4H2AwQ2xO9nF02wiKqjHHYaNNZ6vlyk4xbWjH0LRZNMDvuTudtP7d6gMIPVj
t3YW6/C9r3popZDzp7agFxiTxbODBdfhlvsVde1Oq6k18HPeZSb2ZZDqaAv7PNyPJmHba5WXGDKS
TNjc5LRpAKyK8wOi7UJ1I7b73Fb0McTXdiuDb3DpRQrTI+xVAUDx3UoD7ijAcZRcXbS7DNFksTqj
Gd1FqeXFj+qJpu5kbZGReZWrikHpyPVKAc7GwJLXIhcy19RDgin0000Wa3T1CPt0CPxTO+q2bp9W
XoHgjAEYxqt7fS5XcxsyhUj3fLQvWSE6mKDtxRS6JLWfkqHp6p6VUhteqMiXIDQtOiDcknyqAsTQ
nacelb6eUW1pAJV+URWPlf8U+Ssr7a2OYdlZk7koxdViPvkd3otPx5q6qsTzQRbUVrrQbC691NOu
8Ue5hHUF6OGd4k6HD3NyeaFGHLjfUs60bSek1ejc9CULsuDEXkAorZEfAvrmG8vCbF+kXhxaHN0n
smFeuow5yUVF96lyeITl0b9bdNgZz4BMw3tg6Gswyc69Y1uUJhKSxkKtSJAbk0tjVEUi4Jzmw1ik
cQEbqcOYP37NJtZcowgp/28c9oB8lKnazsq4xDUsALc0m8m6jPIRl7g10CzGhWH41poLMoI0jSQ/
xg8L0jvh11SRYHzrd4IE3SduPz6ea1sn0hB7mL+3969MfRAoreUCwCXBPL+DrO4J8qBPJnWteguz
FWC3b741kxbKNatZdD4/wC8lQ5sKcW1NitS+u5+wd4DOM3vwOBLys+iQRdP26vX3t9Dm7UxME5zJ
T2hlRSFwG59BPj8E9urti4Q35Aot4jlcBwvAc9y9FBR3A/KpH/dkbRZkt8RF4fQ5BhVfKxfB8wdU
oclZBpxfvB4rM6vDQSMgy1HOxIbMdN8PxrdmZxOJTr5E58xTWPn/JgOF47tem0rX6b6SZ5qHlnND
aakMltqMWqB/tpKITLizIMbQMPAwEfBLckDtHO49RmxtRLwA1sB79BrqwgmLlxgXk26u0qT2o4B5
etS8b4XodAHa4m8f2Xs0gScXqSMK5REQ3IK3enBIw1HgXhzf7u/hjjb3LWb5isOoKVnGIY7672Lw
OmCJsLPyGYLIMxdyUTR66WzuXavnbdwkxv/iL9gF95QZWoeXfscYqifJqaIaRCqUJfuZuZM2/ww6
KbUmAqYP5tJUbZ/FH3pFgQsCaaJT2Ui4GBOJ2+QeAzEQ+udxq7vCVGYfC4E+tO1pmv3NrMtdBCUA
nQbayRxzqs0YQVCuYN1E2GuzXKC9NrNI/CflKFu8tiahph6/qTDiskldTMYNUkmWPLy6ReP7cY4F
1bt/jo89qzGjOxGkZysiHHjDyhAh7Qz4uGFeFXAlHaC0Sd5lolKDwmuECKGnlYI0kUxFpV8gV2nv
s2ZilwXdOfxXlPQNXf9sDMhU6bQQ1Hd+k4UD7zDOKN9OGYpYzWk2PuU7KZSsOqb+ER109+sPxD9v
65CEsJPX8sv/jIjNP+MBxUI+PSea1Moxwuth3K9k0wF44my02qmCKAvjB4IJoMl4zzO4GX01YSw+
u8jKer5CDjK41pwbjPNa6JptIpkFeAc26FUVsPNwvcd0ClkqQXx6wlzQzf7suvM6GZAJwFvBIjGy
Ry4pvDZODfqTTdrEEa1wcuGLGwCRzLx4pC7n8xZmxZXAsQ09W2r8TErON/ZX6FTLdLJgMyDxXWZL
wwt06EnkR25RJbDxaVwVM1KCpViInEscbueD6Vq81DSwmMNQZVA53izIRS4dEs5WKlkF2El389m4
vyfilEgHwbMMrrOQOr6kgKpfieeMzmTl6dIhQVu4xrYrpuTSQsh5id+TPUr7FQtaEhkaC/V6RFdh
d2Ur+RpR921FURM4eAeZaNpcoWLKPy/6v4Mw4EphShjcYtkWunmuBqFWu/JsYB+R6Ou+yIySNNLq
K7M0rr3ix24/wXc46c8zmVrYYbcA9bwYdednArdaZzI+trA9tLRdxTWjRfExnkwjC/mDF22dci5k
jfGlvFkURrtpc0bzBc1AlWSlq2dJqp6wuJyNqpEeS6/nKvkWD3Zoq3XiZBnCASjJzcuOndCCd3bt
K/EkEI4drMChocGJUxB6Wxs+GFLDBfnxvk3LbWJzeR1iebbGj1bhbSiRMerBDtT59at7dX6eX1t8
U4Jd0keHex+WZeSOV0RB5tLpUS0G/bUHTqtfLVkPXRPnqyvEOOyynrIAgTDVkOaQkD6zH6kC2eYu
HkUeIzJtz6rtlRTHaRLPn+n+08F6duzrvUnQp0q2NUCv0o0gzlk46b42EC5J56Wj6W6NyrcPkhIf
Xasws0a+9IU2wl2bZ5lBnF3Ntg8N2V226QNlKmRG3mkcqS0I//PkNrZ5zz6U6kA2ryUoEZlf+3D+
VRH4pGKIPOTNLZUc44DDqDl5fWhIdZY85HbJl7V/Dna9A/vnTWWqy4L0KxcIrleJ2h+B5ilRMn9B
04GCoLXw973dhRcFIED0oSfc3Omf213ctF398ynPGgVq3bazSoYA/jvtHn63Zvea9k8Hl9Tixt49
5+1eKn2v7dUAcGjy86gqgpdeSNheKDWs5zxYqYrIYerKfQPIIJCuhs+v6Asa4QCrkmzGrGz4NNfz
7sx6pVy+HK4eDTNmzDDvIqLT7iqcX/FkLvleQqUyLTOcL15wQiTcebnIdJPcYQOJ7u1yLOc9/MMy
YJkt1IdHypD2EdrRoW77lKiIjRQQmIVOeq3gsvHc99g2TtT/yoZo/Nqq2kuvbgutIcqgefxCVu6K
Dz5lugX9BgU5lPBRl5aiAMnCGqEXSrhtQXiFrTHQKYeKbUdVH5Si8DrwlHMQANYAhYYTcOh/GAwu
ue40jBD7lFt2Jgloe/GPpeSdz00kzhBHNT1rJbcWNixOjJv7qlvPo/YQ11w+fNlXrwq7+eCvNB/0
ladcAOcreIDiryM0MjIxL85t/ohpHOaybNa6zIIZtyQZM0cfHp+lquKiiqtjr+GOmPwYfI60J6i9
jVX4sRa+4sCG38X+UERBWjSfhvp8b8FF/TRywbjqisI4Spp2gbAXi/Cpu4AZxlE6p5BhQbJdJ7ZF
j+LCDXpP+TVKEoaU71Z2gD8IRuqk0XatmhXqOqaoJM+JXwjPPl7SxSCtSqZe2yGJ+dQNphBaFRFs
teHIeC7rIkKRkXjJsb6On2Qv8X7U96lYhM7zsODodd+PcWxiHioswsncwSzabK/IdqUMaM3q2OpL
Zu9V0yImlSs04ycQN6OCSUQ0HKuMOqo4MbxYdY7Akt5ClN0ebRJcLru8HzfONEVqplZ3p3KhVE+H
+MH6DWoF8hU506p3u41rsH2Skp7rSwEOuriF+8s3ovPo7pSRtLgJOoRTBj/FOj5Emxf6fRxzLLck
qlRPSee8AXlcDCUfBXD610X2zQoV6D7+mnCg8283EiBv8y+R6PELF961gW6viCLIeLNGcomRW9db
229X6e7a2D1yQS0phv0NWKetyMaV5DKjqKMqO4oNFPkK5z2QbgNRKXM4LM7lUwaJ/78eA83UygU8
H/r6CUMx4UArXcoq1e1KBCw8v7LbgeLChVTLODs8+fB3Rfl4sJ1HJ+EaOLcRP97J1MQTKBvLeGxG
Io/8qn2wg2pkpmK8KOOLAATfH7npNlDJKKDQltbFgspTBWbQ3zCu1XLA8PE+xZOvsb6VFeFJUKQE
aSJzYzkQQeuxmzi7ARcviyGPiG1YjIELFMz1TxcgLhk5RMy5CLJLdszFFj5bfyrEIR9XN+/s5VBf
pjtEISlT2yRzgb7g7wa3stTAjQHAIDnGriK08nfxa6iSWCAxNO96X5WtWerqvsgx2y14RhMoaNS6
WXw6LJdaoFUFsNt04aGVuEN/lfEPy0gbWO/6Qc23EEkLSait9nIC8kO6+DhMylBW5HMX79H/a7L5
Y413Jj75ymPz1d/R1V3BOJ6SOUrIUZKi/e8+n+94C81eFSo7AHMTuD6+4BFjjpjNq3AsndL74/14
UjG6BgLSKSQHz5O3/ivH02mfOgrFVShnPYihLFuv1Zmyd+sM0dPKrGUwx5NEM5SAB6fAoT1nWqs7
6svty8zcxnV01qLURG3eHnH3HjXMEYRkjIXp4jizy3wVLEDpY1ooF1DnT8FftcV9Un0zzUnavcXW
HLAwNzmV1FT2Mcdr0pwWeWBQequii+GDzEVa725n6NxAC/gApoNOKB2uCb0gUM3SjJ94E1+ShgrV
xyZDr3hbrNFZRk7xiL8+5WZbi0f2nK1qXTp2iQVloLlIuHiKMib1qS5dIybIMBL7D3XpqVEtZN2B
99QdF+wzC+eNEiomjwirSf2PG+6ZAFpHwBYjVKx1VrVoSk0znLnvgtEae0dV+qEkOxgleUJsqyAX
KgIb624kcor4XmQGRYolBr5ohK5C9/VrxVwKY9v36DsA0EP8W5OGzYiwj2qcnWcbTbbcQ6beY9/v
VAvGaVGBqKZfj0A9zs1cHvhv+cEjG4N7s34gDqFw87a2ONrGUt3+2sae2QIdLznaFaEXF6eejOH8
1NdI37I4+c9ceFpnpDcIIKh5fQ0mhUgAy1hqzP9h0un6PnYTg7RrbVEwE+tTFVH9QH9v7qDOkNFY
qR/pQbeSLpTVK660iPZ6Yf4jY7TdKpbJsP67u1UitWnu2bzU/O/BeoPl3DNjUbtwZQ0LxWbnwZFt
dpPK+bnZNXrCqv9ImIJnb+aQGIxch7pSNyW8PXRPVu/OCazEOt2c0CRsgPrvG7rpUa63XKuonjg/
hYWczr9boqQ+6hs5D3qItBsnWF4U+MJ64y9GxS8GHXI49KISArlY7Ej/U/4mP2XfPIQjGr/RRPH5
rn62g41OmXfj9BEJcDxx9KjRCjDXQ9bU2PxDYwP51NFFCzIfSMuVXVS6CxAhzAx3MGhHmMJGqNNE
Hs2VVbC8h7xuoWMnYY3YP8zYOQIF5EHtd2hzyrTdSwI6D36nTaSTd5biZVr/FBCdmJg9gMVAf55f
lY19UQUwh1cgLGb8AhS/R06NLZ1xIYAD4nFYEGgWIHmrZBTQCUtKfRHzNT2vm89BoROYs1dXSI51
ItiGy3V/EFCkn1SKH7MIoEw5t3i+js2dkX0J2JaAtXkzbpSE4XyvgP3tUCkFp+hKvZfonEIqyK50
yGAKboooDENBxzUeu8/H/U12oUM5nmeqfVSDMOIhVGYdpsHPNa2qzPt0A/RS6A+rWKcMZM1Qw9xN
6ulVaE9RQT4uXcKAS/POp3Sz0XZ7SCf1LNAwQP2u/M3i3n+/XrT5+c/OJsQ3Ex0ZqmiZqJpeK7KQ
tZeNL7hCALe0n7pe8z07O9YjD2xiJVm5y/XtWcIxnLwvPuU6tOp03QHNyj2E9yQojjQtx5lYKLz3
PJW40N4s2WvxCc9B8oJq5/bmjr3C4SUuLve6Djh34eIGvipEH2A1I7mj236uBSuOpNjIkyGRP5/i
3a5e0LSFijbLUxwazPIyu3PE3Jzp0f/UF97qofODoNCcRqnxhu1zIiOiVZNb4Qxue/UIQR3obSeI
vM8BAv4V7CeiYFRsIb/fzE/DtYDS4ylATy5QdhSFlm3uY3kBCukL9v8djP6QLOrgftSWWHGoxixB
e6NMQlbzh1deHAw+ap1fNKlGBV6fhk3+y8NTfU5jZNzmsKi+DCkQhYIrDgOwjILgn9OQ/m9b4tqF
bQUeIbe9N54kJ56PIMd7P3gWBRHAPrqh2NfnBU0HsR1QTbwPylozAu62RikEkAmX6JiqVGOucZy+
oZ4uLVDukNv2c+FJ8miYVoHvSPxUqWq4Xk28naY5Isc5/O9dW2G2r/fUD6xbG2g0zXB+qL4fcKyW
fy/0V8V7yEnIUgBWDRL5GDSJdCerQrv3hTXRWQpR44+j522PhzIQT9vLkLL8G7+ZhaJ8exItYmYZ
gp2AJE6RcsSrT1OQd+4SOpja0tIF4lSd1G6rFBoT2Ap6Lgd7oTWo5iN4YkfZetn1VCDjdVM0SIIl
CjJgacRXNOFHQpDqSlXEaYh/uKEyH5qAHLXjgWLGQXHJVndCnZl7GLnXyGj1Rp5SkCdUFk7DJbcm
yqX8vosZzhjGAw6yiS9KCJyz/lcmdzBLJZOABf3ZDJ88VOSvVNBbwkAE+sU6CGtvy7xQcPjR5PXx
o+IwR5fnisqlMqcn/KiqqLXuxKd+HgtovaKBS7tEb1sVoT4/Q3cEQy84QlQAZBjs2nWtKcupLtYf
tJyroaTAVpc+y7j2UlisxGNwxMINgfBeiCenChlnZATzjVx2dPHXVBoPlmds1g72Qkk6gFAgD+ks
z1X5t+lCgFBAGSS+CD08Zi1BIln1mkKb7kJBQz3AyrBZxrmC8cTrwNERVL+Zd7GFbmawdwnXmkIz
Ctt8YpvGKRr9bCeZALUgIQAWh+jUY9d6wTdj0VMizKsy4zBorG38TYV/e2C/yi9uFoKBboF72+9N
7ph9hGPn1jHrLM9w1xKtXK7h+w85IG3BZ/kPW3jk5C8jXec4gvOLLOkeBeXuiRuKvZ9yUqYysXT5
ykguhysMU60GLhnFB3gGlVdKPG3YTfYFu0XJqMkihfsJzoE7+VeOyXWMl7GcnqImWds8hPPDgtZl
P4YfsNtBKJylXzLdCFoXtNsisHdOF3QS2WyVMNHElzo1f44mnF2ovvUs5EBa1vUrOnuFicQ350Ev
XmR//NbJCGW0dC1PASyWgg/zDv/mwhlBrEYKf1bVbOy/deyI8OpK93fY9gh3ojFKwpuNigOytM9H
0VdnJVBevjTs+R45ZjkVyYJUboya2t91JBlgDUE1rhTht9FiKcPbueFLHFhHVzDgM36SLKoP3yKB
vQw7iwSoNhDC0iqHkc1jpviLrz4phuT5v+zluT2bnV7DlImhRQwlO6dkVIgFTvvx/urB/2Anzvr7
2rBRWuqBDv6g4LR/Uf8Wa0/wKyhEJc+uYBcO4XiL6691zPEd4JbyCIhBYOqqb5J1D4mfxeFtd9pP
jc+T9uzfjJqDvWPfVUqYK7/wrCRzxFC0twviFaWnIjhWiRUxR9Nq0CQmDYasDWlK1l8u+7Rl1tAU
Q/6dEyNVvq05M8OYy+pizTybpLj7nroHaJFSdjEPVmYBEYdfk3nqz+qr58OghTC0fvMoByw4Sqh3
pIydq02gDbOCi3feqrhzh8P225MOWVgVLNoql5FSYD6KhrP6qn5cMwH//v0lDKJAbFbbW6bEaPOL
+sBkwnCnHGARQEbXXRyl21GqpLdd7+P2LfRVfAfkOiaKnSYpdauQIZ6gqtgmWXi/YdOnkY6LUX4o
8N378Uv0Cvna0LwnnfPyC/z21FN9+YsA0pu6OJDftaZXPQ8sQ/a1Vp5Q5HwHfzr0MlpLbCTZxhwc
5DC9CjOlxvesLHcMVPUd5qnzu1gtqLH/PKsK3qE8y987jbDrtMr/OdfC3lXLplD27qihhNmKjKAL
CfizSISvMdKHHJERPLiDH5Jcxt0ZZKrOclO75skIt6vNoUeUGQfXBB9tWTYjWolcuSYxxd57ImDM
x/zUwljmy0JsVWQnXhwMAh19+8AIUlkQ33nf8xFQgb+cmwKXo5apZwXOFNDZhqITGiCBnsF4UVTx
ahsYs0bxCP8Yk/NJSpzzq4HdfWgfCcT4jdGcjAQm45Rqlk62UYFWUJZN4jIVO3yy5hrCO7c4gbzM
fIsjGts0kmrkX0EnEuJO/7kpjjXEe8DK1SMzrjNh/ZHL1wBzQckYMFbofa+KBAcB3DcDS10ZyVHV
waekPBBIx99yrdACGrd2gwsHtbrAAPMF9gyUKBrjx0gRNDOCjr5t7Y1W/W6hxeywmh9+Ri3cdVq0
1Kp20sjqep9Az1CsOIjjtVBayPJ8w8TQd1Mj/MOOdnC/w0y1MgvxiYE5XVO4EcMvyTBPwm6+tlhV
Bbrga5YyzxuPTeA3Ol7mPNl2D1zKQwDU8H/jkkSV6VmTLltRuzBUEFE8pHsQ0suYulJ1jLNT/X2X
7mDlWL+jyMqZI2o+5x6TfFEveexQfP77Z5cFESpSijZ3YIZlZjTyOjSg5bsFBByW04VCb0A3RcFr
/fWVBHYeRM0hHD7BnAPFAArqvC9yc02PvMw4VhRhT3jAxyhmbC2MZLj+eUHqo781PtoP88Y3UX8m
jYBHFydU3hcX7YaP3CrP0enT6Ht//8RHLASOlxoCwslg3NEWSyf5wVkQLaEyPqz276PEuC7f+cMJ
+IYIycZEPe3kpHwCOC5Ry0XCwdYuL6teNGjgAUdlx8Sx5DIO8o31TewADYNDHvLmK3WiOyeILcAq
Ee8erKFyDPeCN2do65YjjLXfa2WsDILH48dAQRZ74UeCHJ2qud6zL5G5MMohL9Hxo0QYud9Kn+fd
WvdEkYPzsgKS929IBBJX4Or/xwQ9zvh8D4Oms+CMaftjzq5tJTLehbv/xexngO3JqzGkPVPcPtYa
Stmgi1DCfUsVILotjv81knSdXkvNSesHm3Gn7Z4/yotdgwvvZb0W2zLSPXCXOOKUBkiH289mrQqS
m0FRvFK/Q0sZyjfXMF84bmEfZKpkZ6apNOoqtsGws8TFSjITsodOup6XbgBCz8R2NVfFz6FELzBp
Xb1PyA3bDCysWGQv78rEUh+kRM8pzjG2t7TrjQ3sJgoO/RW4h0u48sb8Ux1qyZMAfANJS5VRwbWu
5jbXKcbwfBQHXi4Ut4/5nl9E9r+xGIi07l15eK0mD82CIhXsFCtUmrO9+PU99VtdE7JgCfYCQqEE
6RW35doFwdI/TYfr17ASZn2Bxjd6SjXSPBGpq5vK6uDfSm3oaR0YQ3I2/dBk7hGsjkhPSQMQs89C
qemsTOhL3+T/zJ4JVi5fSXdBLOFJzOCAo9W938xThfkUOpBs8BJk80KeiBk8Pw4P0RsF00LE+Y4f
yvVHKH7gAZ3jSyJ5YEG9pdlRX5OUA75w2p03jFkURGWh0j6bFrcB1qiuSDsG45hjs72ZGBFyXJnn
dhlk1qoucx21AcaAd/T9HfmduaqJJ28C1GMq7xL70pj4RplCTpa9Vm6EXNppRJClL677DatjOBKu
dZyWSOTN6j0uNXZ/vWbD2M5njCUU40GEadN9zRpg/FiF+XD9Ji5flUOzwO00WpL7g9nHcctVvPto
qYVR1a66ZwmKHNdzxjISi4LkIFUukNUwOxB3mXwsQ+96Ye1qyPXqWIWXT8wr8EHwOPy0pKZKagfT
OLchREMsQIzT2FHP1R2hWdT5ekXbFEzUOujT3QKH+z0/EHCcg5beGsXZM9o+niNPcfCr+gpXj4VJ
U+MYUnWAIm/yQORU+uu2hL7qyuNvvsnX07Q/ZTWliuiRBnZSO5EhciB1JAfJlXcr8KhSu6wUofDt
/gkhj66NA/FcNxb9BW4gfY7afz7tpBd9j6h7ynNpm6pMq8xGvOIcjmTJgkYm7wH2Nnsv1+utmxNw
AE6ugSPJ1Wot+s6+oFi+yCIN4EDW425ACKgnDTo/O13uyfIzRdGEJltoyvw5akQD+b3lxaUiG6kl
G1vNuNiQ4Xtw6y+mBC/A/4VDt3g4CtWWb6banWgS0m0LXRCs7OpP4mIe8/eo5YVofXwix/kdyz7k
lnxwKpIiNOfKnivI7bQGUfziRGtpmu0ABV+C8ovUeUrhYNnTAemyTwlXJtfyQPocLEtBAX9HvQjA
MwK3jCh9x+zbTFsuokyjVhoWEySbqfO/7m0439D7iIW68z4X+6AjsoFDIYZDn3RAnr1imqqaC9bw
kB8s+SiFemWHQVvjgklqUYqcnKtt1lGPBE4JaB2GuKNSr87Zc7VCWs6iw+BGPLAa69sbIp8BFJuU
ErkUSB2thmpOl7OtJ0rS6+FiUI1AGGk8c7yPxnaAZIq1zUkg3b+x8joj8c5BzzRJidcFQmyfy0+W
OSDerw0Mgin3XTT+/WFitGhP1tg/v/apMX+1c2VJPhzDB2esvFqW9mZ1KL5xJ93ETUU/h7RjXMbS
hfMcw/0kz5kENSgwievFGJOkoR47fcwA10LaiqSRbp3d7O9jZ79oFKidIJzgiAy1LyUIs7f+T5PV
591J5r+VrIPX5B+j8Mh565S2M7+LlSLRSfdXsrbxk76SiUsWPUxABwdSeYGIwTwlqxtbAvG8ZnIk
WRUlbIX4OXTanOdW8CMJMP02/H+tdMSZ/c1ZN2EfppQIGWMy47SyzL3v6xP7teG+cXfcbntd7sgs
rGPP3IPoSNXVsg8S7+TRR8lMz/AT/tFq4wtvUmfYLc2NnjfEtO8zxFwsVxjOtvSGD9MpZrVy2Nlb
W5y8e74DEZjE3qa0+EZ1BT1EiCVIucPjw8MkQdeGIA+VL7taPilhZTkfc2IVv97QeUCt5DCi3p1r
Xxy/SRdWlFqMl48g1GrGbotB0I9rS/ETQJaoKo7swu55axd2E1tzo2dqxNKCEe+rd0+4CCv3eh7Q
C7CsK2hXI1/2I3khqfYspgkLtZSQaPdgh7aE+OcBd3eT5vd70a9LMgKHmX6fHZRGBgjy/ctvy36o
g0OjDzMUT1GmwknDy2+JPwz/kwGgcqQD7qGWuVDqdxhCFpRjlaJapBraBYRpoGSGxFI56f7cstKT
6RWmbtLH3ZTF6Sn76ps7WMI7TJivovC5TUlRHsVsaC+eqox7UEnVgvGeEGjY2CdsJcd3mlyZcdu7
3RIu4mMq+lCV7UdFKscTibIHspeXp7zGdqHi8jl0aebmdaPp1bHNoZ58oOWJS+dUAPn8ClXOwLSC
FWhODy9mkNwXDUrH8wz2ShURAcmsI7dJNe6dBeFG7wetRt5qPFS3m8//gjBgDMqU6956sZkowUgn
uzWzLxC5qFqBykkbnfbNnckOzqeEeH737HVzhq9p1SB7p7otuw4igw8izLythnWgvUsQyDDt3JMf
/AyVYpOHHQvQDudKS7l27D4xiKxG0FgH69MjqOl+ALCtVqfvxPob6cFJOokBgqXnjR0M/33YpSOh
wXCqGY13rXLhOi0gfQhd//P/3/NLiGXZLWduGT5h4hUa1wBVwYKCjEeKwZGyvO9pa8fQSPw/L3m1
LhLecGFC7vFbd7GbQVbxjwOQsK50tYOu81BAInL05JNLm0IzjhxsDF2jRNAapZUW+N0Va3qwQgOv
zulZXKCqdxBNQUawLWi965MbMvFc4oioWVIiQiyOs73kHHljRFCO/7pop1ckQNTnkTKfqY57gPKX
5gQ2Zb/sjwaTBibkfW+Ko56unmybwfBl/0d6A7z1QQlMaZnWnP9iwecLwUViQmCRPEqUQNC9mcUh
rtSC/CoXPZ/y1SOwX+1rsa/j8YxkLp7CYVZl11e92n3p8h67jT5shAcduk4tNe4OtAe5eOozbano
hkLyJAbJoVIucFJ7suwwwBT9zc1SM6IaM5bdL7KRicgFj59OLAnKLraSQqbLdd8p2nQGPauE5XXO
t9VPlGYzG6qHifVtPqNMqjdAvICGVvWutd5Vso01Ywam33JQU/NcJtjrp0+r6BKPE7PDu9Aor9CF
6g9gN2tUhTWFQq0YvMp0D+R0ZM+d/qi3zvsLiKdHg1HWCb5yfGWCH6dyuYB7JAWmR2c8wSvhlIo7
4b8h3XgX5gfjVfXpgvJ9KYuc83ZDr3Swq05JqZ5SrBThLOdDad9pAqmfwKUkv1A+CaBR+zhSKZDL
/kHXcVSrm33C2q8jPbijdKHmUxBobEt1ZowjLSIf3HEMxPOo7DsHSjgIhnX/+GT0AzsAIVxlMwud
TXoJO8gYePBaFAJHPDvu6HQvn8K/5tupIkRmqFd2EuwzokJhVByH9VUCHRKlHqESnTts0aAHcAwK
ea+7JKm7Yny/ESzAMl+tbk2NTvtwhrMLzXUd35ZfgvAGuwZmRwJAX/B6ngJb7CKRql3GLlpnJQPq
QJ8nXi8XHyQXex9VDKnqzT3pAIXEPBsacfFO9wCPgqW0kV4nBwLcU4LyvqyYUnc6kSIwH1O8kuWU
SYeXzauEMfkPsydH8di/Fy2MTj0uktYDDTPS0h/R1Pe3baJ5+clEpoHPxkahRAsr9in506xiC9au
XJD5+HI203iolvsakMm+blxoLZ5M9qxXjAJw52S5vlFk1Vim+kjHF4SvMNDleta0o+aCbDydjbru
+h2XAxkvmSGagpAzmy2pntVTVjcu0F+JlAv/y+IFe+loM3qn/kgkDKgdatg9ZSNcUazStLMfUTJt
61s5/W2XXcs0pw8Jchnk5+W+DGtlQLWGrW8FF0oYjYLqAgiqfbZtnOvORI76qrwSXNYI5i8Uo08y
4HehFKiuWToT+gKwSnxYxtd9dBsq4pygQ1NSVYdxkmbb0bUNmJrPG+P8VT3rqtPiGTbwuaUvPpkm
2jYlZmj66stoqmIkqFNYlu0I8xWtmVIWLI1JlNVTIIfnhanBeSrXojxc2lTWaGgGyVg5ielukNxM
iJEYtlnXUMbtbZCMXw32Re5PmDBfuFnU7RFfJaBt7rC/scwNLsAILRPMI5UNBazrm1MBUihIYOpf
dF5MWsrG6F5s1Mi7ViXCqDTt6hEAtUs9ZN9gMEgOACnZ09fDQ0qi5+B5vWGPXNJnfv9utQQpIZe2
d6OOMLx2SrKMwXHSbmMiPk7a4Cr710FK2wPA3d4SpyPsG9/Ef/HWrUopAeKJd3HZ+T8snIdebxSl
p+OI6U79Ws1AmwpT2qjB9OZuFMfvl1zJFldyiJsmd8B6N/g9dhzHhzyEueHVBnV/uZNtdZ4pPNoJ
hQBa+5vBdyx2Ay9wej2iHG4a8KQeBPDZeZjloWRxNEHtK7LCUF+FNpALo3CfcFjVYtwxfU7pMlK8
BDqoMKvb3oGDwIhCVaKnBd35fjwd66GRg+WTpJ0MPCxrlYLi+0OKCbMEPhc70UY68bUDUexgu39L
jjAcd2NF4m8rIhek5imfV/zwdQCu55XzQW8c3tGHCO/ZfZQiMnH8o1nSitTB8XZNnW4OB52MbY92
jYAgu/RSpIMRGN9rSiPV+GP+K4B/cQjRGOS4rWWtG0cDeDO4+7i0tbvLmx8alR4OBSpigy888b4x
RlWee5jrOZye4eHeC9h8jEe1NBBfYCcBB02O6Uo3pbS9FciCtMJZ/9St7CbyP+fbArief96gIHkk
SPix27ePKBQkDBQ96ezHiymvvtmw+D3h0Q+dPIsjrhei4qyI9rgt7xbG/RvcgN/rF5MzmbAOHjWf
KU+Sjl50faIPFfjWXDkM1JsXeFg2vmLhquqJ5eC2RRwKq5SL9fuLbTzxSW5C2VU1FxMAFkYliF9m
7vXszvFyn4h1aegLikX02I/HuaxYtcb9kjSexLmC+dZqzmOwfuN9WxeNGqvqClNI4jFve7Oqy6hB
1vIXzNsD/V31IbDKoNpCzPjHRb/afRH8unMXlEhEreZGdcXv+wVHk/WWOypPVbboibvKuqx/un1Q
ymMJKbIboUyCWKhUPGLCmZR8RCA2kHLfNuOmq7CVHzfpgxuEk3/jJthiAK6cNFe2IpGaQVS5c8n8
XKtcK1o39+RZXn5HcvDAuWFXeUJziwqE3nRWmKPzGUQSybJyaRM3YGegjZpRNRCncvEfIYnVsdYn
kSRK/YRshsBYIiuf1oifl69XbeNEwXz0sBWA/a0FjeI5TNx4RjDXYZHG1TEsFI5cEUpI9WQouaRr
6A8PIHFwqa2XXxLYeufuBk3+SOxrvevnFGWoclrgQrfwN6pGrdRZE0imki7a5NV8A5SxBzGNgNoG
JFdDWH28TkmIMh/f2TNf3y2O28cHqOXGWAeMLicrKEYITYPV92GwOx2GXK7Hs0yMa03qhYBhL5QC
ci7q8t4x9IdSldkajl/ZbIXrtTQOG82P29DkkFgaRpescNYSkYPECBsj9S0CUqv0Z/rZ4qOsxCgy
AZkhPSRnhI5CJxsJRGwZl+P8jggGvHppjNitU+vNOwPPhsIbjDD07jlthD4LTk/yVfjoH4s3hXKW
xH5OjPEq6qIWoGK4BT4MEonKyVD74OK9rJkLswUkuFD94B39TYMRVL7RLkoXwaA4S0OfW7scifUy
5fND0ipeTPFnRhroRI76W9/g4WL5Tiea0A3ZLYhM3psPzjQDBsIDCgao0aTWshYDS70YFoaquZ+q
HFvHlWN6NdR1Xs+KY+9bh73qfg6eNMREDj1udy7SnRk3s0mW/DPLmpQf27dcQY6TGyIYG/GrcwXM
UlZ249H4VRXDI29eEE6eqqTx+HoO+8NFX0o/80qm/PwVUz+qUoAZPOt9rQ4KoLlcPHw4UJOTfzpO
mFmiX1oc05apcnSBBfEvsKryA+/xRgS6YYUl9I5a+jPYrJn3JG2w2rO1Y56+ngJ9gGphsOePHXit
h5RD3Aues4NKBZmQTbg68e+BiTHWWZ4v+oHftU8cYjD+H0Lf5ox8xn23TgYMcGgF+EbF2i7S0Amz
S/lZq79M/m7YraxFFaivFdS2ifs+0qupNSy+3nrjb8uS6h40dAk16BtiDYnz6KW7ylHkQrOp8W1M
v4x660rdGa7UV/nPx9mSHcPyZVMygw3RGgC0RvTsOa5OxIYFcwG0OHgWpAX5jh6+s7UbZRoCCwSJ
Msox5l+xAZyMq2+4WCf/fPA9tKNp1qTmPc4QIVGPUXFCw+JldaTOnJQFEZBA3Z88Ka0jaYbCyxDm
KsNM17+WrhZbz4EvyYSWMNV4ujGL8fbuz8+oqNGIz//S67CinGyJvV6o45KOH59IFGg0GS1M2awo
IbT1dkYe9NygtkzCy0iddD+rrMAhzm/W0YVF+ZxGedOX/X2ujX+nBOuGeaxPJKB0SoHNSF6MPs0h
c4oltaW6JJ8PlTl/u6hZrGVhtrEYQP3+oYsNqXMey6eKPNVd7J5BYJ80ICVlf8WzBBXiYpODq5Km
IKbpWKIAPi0+8/SNhD3t8T/Ox7R4tlQAG+LLVZB7JdtTBVPAd6d3a8M21+QljwKes5yR7jganWci
FT6+dKG4INVVuI2WcElpNrYqVURQRoLm3DkJyUmnhC1yPnsj2MGDrTyQ1oH4PjtWrrSqsVVttoLj
61OyCs4MAd8zszKfYFHGK7+BbNs0iHd+4RnehK8Mlby0BB/F55mSUptvUevVSmBceA+eVKounZLu
ZlfNDYg44h7dtND9V/jl4jJ8RnJZIEOdP42Nc8JTRhSF3l0xl01Ms5OytrE80xu08Hzo/nHCrZ1x
Fwy/yZyB2zXrxwu1J8FstA3GFbeOxnL606ulsvrRwXXIWJSOZkED7KaAb9a4njLWcneUptMpocKH
9xCGEQfx+81/+p/t1WEvpLxDH9hTZe05mobrBlyPEqEcKIuasOQu9i9PXKTwOVsHWYycCTS4svKH
x4MZAmFYZrADCIFoC2p603QW34NrDfQjlYC6e3kiRMH+U4XjwAWoQKP3qxW9rujUjUiheDyLbZ4t
9J9LRUx7QLHiZvR5hZ30UiHDP7W+HwVXWu4OE3vIGO24Ih60SHJ0CrezZ6qksol9esTcIadXB+3l
20TTgto2uwDpFeMueoiNByXVfUJR6VgD4T5FPNxbR67w5ZlRiYKR4iSQgWmZ6zj56+t8DXkGfkU8
wBzWoupijTWHluu9oliOK0nRqC31htPO2TH5xqPjpwogH/94EKW6LZTw+x6UDn60ULpXcyOCYhuL
bHpLf1GVFBfbF6tfei7pv1SgCOf+sRFb6DFl9OBMm5xnCpCHg48AfYi8GafzyAwvGIPLPApOyx4r
VqZ+/oZhDyGGgukEHYtl+phP6YtW74ajRx0I26Z6LIWhfgz/ESe+mR75k5rOU+Q76KKmtf1Or+mI
yUrXaFRpxkOqVCJ/Klwontw4e4Oo1Sxh680r03jOUB/K67vYsnvRT43EtfEsA/gkX9Pc6D8xwTVC
cru9Zb2r4z5If7utteaUF3x++seEzSSi9Dg+5Hlq501ToIh6/NvFntHP2zpbaVcWCk9RvCYjmzsj
a25S5oDGudqEFsM3DNenQUwTwwGB6Il6HTu/xFf7bufi5nUbl1Z0YH4ZHlQHy13475Y1wkVLrkOk
ZfiO0VEaSZRgb0GS5FM2dBYgojk793GiWtz7bwJfU8AfW4Rq2tXXKtYUk5uHPhBe0a6lxA3nJPqp
is28ACrq1RknlNxXgMjy9qrC3XwOacvhH71z6cMvGA/59exeriIh+AC/IsUq4lvfKI+7MtOFqQ9E
WV74YdbmE4jHUZg2bAIdYTNSLpKD9AuZ4Wt2aAilsR7d11bVYZXrUvm9sgAwRUoBGQw94Tr13Hdb
BCOr+I7gh9hv1Fit0TLZXayuA3vAskodRr/eZQceg5ckz6GTe1qSDi9iZDRGFC8Yd2XIa1tai1xg
sYO04pKGrMj8udOuR5wAJj0NaoXv06RWvXp8L14l+BPLmu+ayCm9Q/wU2pB0kaZW9jCyt7KsYjEC
VM8+VLNbmV+DsQpG7bowk4dQVUUPC+mJPmYe12vVS9qZMsyfHd8M6OifmD6iEfCuTbuW/2p20wmG
ri+fa/nnsRdO3p1T1UZbbXjuZxccjEl/3Wph9cobNlXYdT/KrIDtxxSGn/U8V7KUqNrUmWRDhmno
fDK72sLIRiMA/GcE2071Bn9CcZb1XFh/6MTXxS3SvEmf66IsZBT8tP+6LV6AUvGCtekd6owbEtnn
+uXcFetGErZ5+NBA4Agih0gNeCLGEWLPuMwKK81Zxw7qPsPqPWK2Lfuu9fHUvgBybI3toAslJjPb
GnjaUoYHIbV0GPEL/mCqy6GE7Gn/6cQykmxxMOAwwmmVqsXpTEgrUlGqNDJuwvAumdE/Vxb2lqIJ
LLtd9IHEDe1ltv8G/lWEfp/SLZyJRixkV6IPupEMq/0rtopGYevREPFzimU+B66f150pK+Y1yC8s
YqC1wltTHcfhxiW7lIITez/Xkyp1tW1vYlZoDVso23jAlSkaJvbFjmcPw5qZ2iEANqBWUuqspMSq
CbaQpqR8xdmTIuPJgVeiTFaffZekBwMYJzgw0ZNn+8mhSzi1CW1hAAQSkySZT/M1nWuXJMMOrtPs
VH9hzRfGBHhJ3v0RllsboeL56DT2iG1GDkiLPwPHArRIo1+GzRNEGdNXEsn6O6FaITAiIneEeTQ4
uaFR6DqV537Fko8cNJt6wzAChdN1soXMyxTgc1vlAwAhijdWBAxfsmTSxe42G/GyZyo4I9tXajGq
qlW+RlU4jg9iYbI+69FeIO7wEDAodfEHknyBBYULbdV+z1mOZLWX7IUQWkdbj5ohIn39IGqrhh1J
zHAgCQwN1aSbHlRBRfnpJWNpW+x5ucyUfVMKo+pyV0tWfSZPJAtYIFZWOpmya3bbNAJVP8gTVlHz
YEluyNeAWdkY8bnvjganXh1nasrFkwN5OuEOYl4dzbuh8mWTs64jGSW1PLhDn1W5HzpYUoUMwJGb
e64LAdC0WLE5wZ2mJLos44/GrYDba4rCwyWkKDFpB/6p63xoFilaaF/ldakpKDrJlrzsF7iGX38n
xygMSPAgetDTdCnjPwUcxx+y4Ie2ert3jvrpdJq/ttHPh/K5T5cxnbvYwE3vTsrwCh8PntH+3Eli
+SQTnLr7sQG6/9DO0nTrWV09bqtw5R7j9sVq8o4C6+gixDVT6oHx7cRL6nvpIJaWoLw2SzIrWd95
m/0U/DpS5s3343+0R1vKbPDaSrB+Ku50vaAVXMJ5I4SAuU+UzKMxu/ntojI3ekq+ssn80f+RENDK
5PgdxVyOKj0FyKcnXCxopGz5dttmXRXe4Sj6wzw1cDphCuboJGOyJBMfKhpOmVINOnj5glV1It+v
1aQHXOX/XZvYLD7JrruOYd7ejqVo08U6IWbzeOcCG958XNEw+snNNnf8NhVQgpD4rWjcx4CbsG22
53d6UBqrKOe4Kw5JTkMiiQ7/RRD9D4TO3tlIi8ui2BaLY9SxbLPqPCjBFTwyW4qdjd5cZQ9Zjyl2
+RUg5yq6rz93PLm0FEnOwYl0c/tkxq9R2vEejT3LefD58X329FuEpzu/gl7zkvH8PV1I+WeuYfgS
ArZbDxz/7BiOMU/ZVSQBNlCEnX2tqVxMMUZEy3Q10RaHRzo+KgvkBY/daaY66y4lUVJL26PGFpVI
BqkKNuKy8FffjfRDVRqs5aMysHifUl1I0QGHLdOERjGEPUmIwp/LdIm/otTl2J1oU54XGKQ67nqh
IxMOQGhpbrUo9uotIvMs6E4l/d/XoHyt/31pxhkLlow8HstBPiAOcYUxx3u+ugZ3YB5iGALou39S
1tO/Av3txtZ+ig7OLISLfpUL504ebA6sfEDOhRtK+5dbpJkAs2WCZtlUMdm6g1k5hMh96BtApd1E
lvxcPbJjYOKeNVNyJ9WNHAh6ZFszDBMAtRvoyXjes7ZnfBlHg11c1Dduuq9nbPDGw5GT5ifmu9M9
trHAIuUZ95RS9jPnLklGOPSwFlkfxofajoT/L7CGLJs0nZcBL6S0FrVxM1tHzwC1050Z8irfQc6E
hOBbXjIPLm5YR6+l1/OlZvyOk4wj7g5QtLGek/X1Q4CVJEbWeP0n7Nbcj1qJAwQv5lprVCyRBWPF
9bSwZ8dxNhvp7oyVYsQrybnlTzklkLmEJxddTu/he11WkTpdLigIu8h6VnrQrhB/XSs5coOxhG9n
1gnjSOrIfDfcTVk7TdJ5EJbHGdbFnRRB58lFXeBbMJWuZCPV2azRzXrZGQxC6VpuE8Hbe7+Ge98W
e2bXHSMfGjqTlqOMJJx/YaCufh0amqrTdqgGPCyjZt/H569U5duQ7GtPXmH/UQAWUmCmEUGG3JsW
J9i4VGAxBM3biw2lmjLMRY1Ch0C6+QuQTiQTpAJi6PoC11y01JuLX6NS/iBmTXff+Aag3rFiq2Xt
cYMpiTomHR0R50IYVFmif+e3Kfh8rZVyH+VWtJE9ni4qZlP8v78JGJjAISLTSATbS3GI6nNVL7Mq
iq0QtYEoplleVKGpM/C/gb5I4SaBrGm0HB50VSrEUXEut5nIlP/vld5INolfP3Tc1pnaZTLp7qBH
O3PXcIominvS2RzIPpOYwD7SI2V5nrFS6USH3CBmkJNRDBzDqJ8iKfeifISSqXAViJWzU0CerCCo
pBIKvHIWn8hu0B0DIGV8peyT2k2yzExFIXmMNyslff0lbslk58huEzKP97sW5RKlQeTd7Q2D5GGt
nJDkgujLrE5tBQfFxZZF8sajINvxAgOoYUyCaxysAXSI1uum5Muu8uGFlmNfNlfwwVDn0e4p8Aid
qIugtoQsrkTFQ46ZPYGOGxW3q5RTdt6kTVBLgm/Ey2M6C2qF+z/tVvu6L9T42EutwOebuPM/7EJn
EP2QdEaJ+KOsCRm6+D0MQ0jXgNF9V0PPDVGcavErJWhiu+sv3dd10FRi8bXSMwDlWu2tmnxcCHV8
eIrAvSSL6lFwz2bYdN8i0ZFVu2EmVd14zDKmscFe/0ln8uf3GV9rJMstcLq4DfIOratZyKpTAZ5l
NvjtUvGdbgs2r7m4oMdrjeDDf+rkdiUC3X/4sAbOl2O3+prHLIc3TXvhPYHsapE9XKH4Gx+Zu2YF
mILGL3S95W4bjhT0KMguKL9fIIMPqHh5Tpyyb91EMzLAl89Zvt0GA1wirmBp9mwRzU1vZ9JKgU/6
Rci0Xbbsyb2yOBsrwjLpUy589/LlDOx3QBnOuVxscou6jbA54wbQm//lRLwakLxNRJQZyJtOHovD
BHDCSmQ+wMwCwoODP/0NrTA6oRZu7SrPqHJtMzjI9TIFk5ixcUrJv40s/m1ENob/sTb6q22PLKRD
f7nSUbJaZ0zXfi7+a59oQNHZdoSaaCUk3UFry/y10DkF+//6ewykpE2OIJMnfckRAVuJO0Wfa3Tc
hm7zAvy7E20lAwaZZf46r4exwnqhVpsBgNAhoCGz3fMnS5qb13U2SFyVY3uKCbxvKRsTexGHyDjp
buhyzZTMUleP0HiaIEnx8jXLBAWvEv1EvYbXiOom/+SyYrtSFJlR0uSYPnwiQWn0LF3Kr9yUqgMO
Pa1PsOFEKBuZ5qCrEin/GnsNwxcErGto59YHM7SwWA/88Vam1/NUtk7q0OMfxSdcQv8oaFL7DVb/
kXA+8COebBdl3jNP31nidNai6yuZAqcy9E4nCZAELdHBU9dhdzJr6vQo+HMDKHQwrTuaf0m2SA0B
upOVd0rqDIaTK+sgLJOKJ+s1XFltgg+UW6pI9u6ZYZpOYIVUDoi+RdX4FHMfu7NLwFrSJlAKaV1w
vy8TsblO7Pga2oLIyoaeO+OBuLK4nYjJ3RUcQmZ2p6A9Rl/qhJALJg+ACu1WLuxTOtz4jN3KTCxD
lPqONLzS9nb0V/U7C5FfRWnDr9aJ+b92VrxIc4btXrU18HYSgM2kgGDdDONPKwzJ9j6/6T5UW9vG
JIJEJXP8AZDJxRxA2ibY1FVfYz1C8wj31xLkFbViUr9tgrkPVuxmworZnEKCNae9ydTWbO5lLj31
1jBPv4DVF8rI1U7cR1Y4fclKqOsYPP3kFxI9VNfJVhKEG33Pi3lKkdDHMZOtiasIvd2GAt8KsClS
JguiCOhVC6icJjGcviMr8u6aUYZ6Kzai5UPqiyVnK3kQ85FuCLP/wxJb1Zh7PpRhtg3buSv8eQk+
dXtczorqUgQOkxdzwuVYY/Dbg+jNdMe5zbHGSLi8umhMifhK+w3FAWSSUWJzA03KqQnQefkyL7pJ
GGfqNuLIpRUX+lVO9Twa+li2B50PbryGTWdQKREohYSM5EDSKHmW/9U3sj8PBtAk5TBs/f0bw+Ab
WcDjlQ8DKJWax2fqj8wgsgE24mXKVCk/axK/jWZp2hO7y49xn15/IssL+/L8gIYf10JltvGKLp6k
jZ2KDaI6/x2+NrZSTF70VJ5c+SRUSviulbcA1UAPl8/H515XRsvZuBH7GbND2ybLEKdvJrOqsJ4T
EQ5po4FHVKWUX9xypZM6N46ZrCl9DNVn3t18jJaGjhjXUYz4ljMfrwQ2l42mrN5E+WR3xQqGoyyp
sxE7+lJlSIsdw5Y7Gs75UEfUMu2pqueQPUzfrCf/+NRhOO2qN3pMy9I0wepYAdt9tXan+tnCvsC+
mK5DNemmryhZ8OgCbMV5UGDbF637ZLbRQUC9/Ncck9il14dNbVS2uM1cRPfIN0PEPqWbE28OngG5
UC8RiwASOU2CNaYPn6Jw2vVOcD0GgM6taCjaekYtXZV4sPFdB8PIb/rtdIGZj0OqvDn+BBUn9mlz
RCYrEdY+ocRWwc8xz4mfv/eu5NtD7EVE4XsfuKs9Az8TpngYwoyUAcQpHawXjmrCs0Qeblh53sET
XLhCd2MaKMGPRTQEAw+cSy0gGRSfQz5ZUG+WSJFmiSs/Sk8xti8plheyNEVl7y0uj5umxTRpsvdy
s+f5W1obkIvcEtC5QzGCogbAWLyz3XivaDQ4BM7MIlVUUK2enAqrm14D+845mDrnKnePbKsggsYC
A5kNpE2Ojb/TZCgEi2m4cLJr1BqEGBQ+IzA/0dT0D2ZZJY0/wLkApyxIQSOWlYtfzJnBMu7+9qPD
vbW9taFRxOCrSIcNxOhf2qZTVzeGnc7CHkmsBC7HuCq7yHDjSAg8LdwRcWN6n9rWUwutjOJJ8hsR
4+6cmDcpMzJie+BqvAcxS85NEt33+rLTxuF5hLUg5D0i49pSHIwf68DjbNUg9jZKazB8u3B0K5R3
xIEZ3J4/+6O/CUACC+Lkh/NH3nDW+ZHf4cXuupMwIdEUeBQrjVJCa/83E3Rb0t0fQc2wLIHyES5j
GyRgEtb8RpGKCzPRFpeYKJfF7Gf7/NQPEisp4W6C7cqfm9uTtUUEtTymJ+j26vYGs9rVNKR9b39h
56On2AEwmnxWV6zzOa574/xgk6p5A0ZStOzutJKc0AEnYmpjX1CPGv0tHUDTVyslJgawGDp797s8
g9fYuLtUFGWMf2CnAWicvpzfsuWKvKPWtcOfozSlGrQFRLaxHPHXcUU9P/ZVAeZWrwbwWkL+3N+j
j8JsbNoRocmf9tMbOgsCqmaC1rsnATh5BIHD6bKkZZAzPTOyj4sKS5vvFT0riRumiDJxvaO+2aZh
bnNi2gZp4TolsIWeWRlpFq6xhtTs4Dibf82/gPt0jWgY01zNPq94h/wSCwhPny+MVSdnTD9lKox3
dfCmdx2ElvIG0Q34TnxY6keyisGSq1uTOY5X1L1PMFAm0yqCcCAr2z3/NlUoWS3OFfhaNDQslWrj
GXcZpzEa3nHqvhaYSoIWa/szNjtrcCYFcoprRXUSise1U6P+c2+mcDZsYDDJ5kL6jVtgE9ioaUIL
bYcyeGV3zqFdSSCSTMJu0e9YlOGgkglwdXPtMnDU1WwvuSmdiNcqcn/++GO8mJLNeVWqPPwQKvN6
Fs2ZVPebfLjaB3XiJQf6iC6jBqRhwcsmTtv0tV3Ht9T3VUxOGUBBhR4UGGb7ZTYaxaqlS51VeGtE
CcFhkkon0Ng5UZJLv6idVJTPA0ublAgHlXPYFcfvYmD/5cpKC8h+Rbyc96FlVP4Wu6E2dwgD2YVJ
4zDYdSUCXtB5kd1r1jQKGCVSRxTEo6VQ3utzOSzMgJf2ICB/AFjG5qzgxsN+gwVVDc0qZGFwUMZe
40dNmM1a9KX+bCT4rKphfRNJ/+2DRmM4vKrusIIVqgLTiurvg8hpjmQnbPKt/ZpEglHvz7uuCOkh
eOQ52TotcItNHjTOP2BbOyJdpZysr/zPpDeKn3YTlguheImVBuvnQIHu4+uMx0Uo8H3IggiEHv8t
TE0447IGOpJqC3bi0NQ3iG9iOubzu5EBmhS4n5NEvl4wPSq+oGIBR9fC4We9QoYsO9CZ6e7/++iD
NNDTDiOK2mCkJtz3jiPJowr2RvF3h4o6Mc8vvDCqCCqDCg5XUnxo+OBHlWih/J7rgZYL3+jMldbr
yPOblULhR7efult3vxj5IkCROqSv/ouuPzNLunKOVDuRc9k2s1DNyl4J6k9fKbRJ7ubUNTpxAO70
wQ30jNEN2GielVRrjmc5HIJ7cBtM0D1rQFnh4tRuGiWbc4cIMUaSOpcnFpWmYqDaVwb3UTpPUu5B
ESUXXuWneQKHeMAaV0y3ycYrnoWxzdk8TT41Q6+pjrgTc/NBVFbI5bzGuLuHdRIwMUbYDIMR96Ap
ISADHpI2fMP/cgTrFezBmSGNu44Vu7ZJ8a56e8Nb24hypLhDHzBpTKi+O4wJp7ro9WMGjdLgTLPi
GA2EPNcTFffWoY/BmUUCTLfZ6GKrQvwxIRlBCy80WiD7iq5YRrkcNAUt+ICsQ/ckZDLNVQVNdlic
DAoUDKZCmKRBUfckYpeGFHxqrqZNiRv+eXVugnQczg4THd4tuKb8dxkF56ucqgI+cWa0tTICMB/H
56tWretbndpPYJKB5CvXIONBUzrMJeFzSV68zMJRCZu0JNDX8uHRQL8tvkvgRe3JxTNiDdlrxqeZ
IfcgW+6fpNGBezl1Nbg7iFiDCPiMbW/3wYxR7+r3UO6gr31QRORLnpab1b+7cf9OTGLXFEAHLF9b
vJ0SFK/c3VvQYvFWt57YG5/2XX9p9F+g04IkJ2TKvQxJPixd4XECo3N25Yd3rluuQpKpuRNG0uyG
DIPSS6Q9YvuUaxPJGA5CI41GaLil0BdgLnTF56NprZiCdp29REsBc3JuO4s+I7E1rQE7SM9yMHIC
aoRxg/w1jr5sonDnx8i0Pur2+IY+o+SGhBhccX6KHZ/P5aDYDdxDDN0yq2ci9A8OfCubYV2j73Ej
Lruf3vUNakTi2vvxFiBP8WEV8cOpN9qxGaze+ClmR8MO4BUUvMosEDdAFQF+eaSaYDHa5OTSno6U
B3AX8fxYdsWq6GHY62ThWyfDrcLbPP8raQEt4RBB7eR3bRxIQQF1QHU1bY71pMBZEBc5NwqtPkdp
UALzKFVYPgOJXAgdIWZqcZumQi732QHJR1wZgu5TmbFYc9anQZGdYUciwsv0nlrKqMTn0HLFUC3V
ZSYW6Zd/AG1cHeONzwQ1v671zeL4HSZwR1YqHUzKP8wqjsy063rtjSHnWmq94UWZtY/Z6WuxEFGJ
CmMl0jg8SQWF7JivU3k4T81FP4Buak3j8fhbz01NwcdM/Sb3LzmEhPrxor5SaWi75HiK23+3r6y/
LCopGxHK4HJQi+GpTv+wlkzJ1hMVzxDqWEq1TQh5i3u6eQyknhecQlNWWvQCftIml90BmcjfmWWY
l2w3dRdmxKanf7j6BlNPTvRjlfCMm4IDEdUxw8Qt48FvqU1YUcJGuJ77ztqzcTc7tknlq7lVXoR0
QV7jZBSbtLMg5WGnsTaz5kesgchv46svAbdMPUI8j5Exhq7nfMdk7CB6eOiwZlM1ZhKDW7vo73jP
KhQjJ6G7vG7D/ez8n6hpGKlUAg/+le8NbkvNBD9EnptKP8A3vWpzAGrc5Tp3O0iVgg9SrTCakxW+
HHQo50oGsFhGUz+HPM+XrV1huvhMKSRBL9RkcsdimPAoMKhjR0el3qlXggQTlxPAUuMo6VOEJ2h3
HWR2H3Ldj4RJ5J7cttDOgE24kn6meIF9+ALLCyKIaO5zcyzZNoYjs1dIMPJlfDhfuGAZ89jmH9Zl
lbUGIfkTjqkdOQv980JphqcLZE7t4YUpDsAqAN6bcAS6n9MFsjXWZBAOqOZ9QWYTSHHYaVeqtm3y
gJXNrB4mOOZiYf/Nt69H/fzI8tErqAbgkuIZLbY8MqDvG2C5sTsrMcTl2todPfybF3mHJt6vN6oE
mXg6+DigebyK5qH3AiY4XG/3HMo/RyvEDHrdC5lYkV8dWZ8kws+jdYajRLZbcGsvaRdvjH1qPbZZ
ACEoPVpbkbM1JYVkhk7ODF4C22/80SJp/ZDb/8yWiuLh8xtDIulJrCnK1GK/k3AfJfPkhSXBWunI
kgrrb/3rwAsg/yy9aQDoqDHTv6D/unLv0MAlLFo7DxWB4HkKRSyFkQsAWG1k/0E95lQdqJHWVjwv
X/uYPnKE+jgdKpHlZSnrkx0s9xv88m1SRu5j9hYk1kg28cu0q3u8sS4Mc1FfcgUXHNAqjVfEki2r
8v36Y5Dr3Yt/Sxv5I59igWWBLZInroc2ju3vsM5YJyLM0L1l+Y2m89Xny8kgASaC+TYBf7rEPW9U
1OZI2qql2r/eVH/0ie0hX+PPL5eNE+E4tArUhwfQ7h5VtLd+vOM1Hw43egDiUyfN/jM2W2sL/I8V
EgKpwNEHpDfYh7hfFqiU0JNNFcEVFHI1CTrg7JGmQcGCYCwWoAVf4ZQfJOhz/6XaX6IZBSVIH9Me
SfDw+pSo1bO4315bFaz0pXgEFUM93FAlOccXVBKXNxkbmskGRUij0yo6IIXBKgmPvyUq1Y/28r5A
0DOR8nqF/U7vxxd9+GjqtMM56km+JwLYWn4dmDDwKKILu0Z3tLpdbCzeEFzEam1/5PKyNDxPOyLQ
6yhoYvhiujhKQ5/XxClFde4SSwzpWlZU+qKxLbN+sxpqUwpq0yIOlM+VZSSWvT3NhUjbj2wj3LaL
RSOMmq+dlLO0/f/IwCzjJPWp41jBYtpakz0Pikr4Q5QLXOb+7eA6bHS9WJzWYq72bogG4hpaROHC
iQjPO3GHn9xKep+zPhsPRjeyJRIatYpu285pcWO15z/UwohBz1xMV6ma4uSk8/NpaU9Vv6xHcQVc
Td6JI0lGP9Fa0nlXdkEPSyP45mSa1ymwmfV0Hl06mW5/8zivgbxoFl6+Jsw3enKj3DhNqfS5rkZd
Et1XGBBRKOxS+NxyePpjAlo7mxHSDZY6dmSHOOyeo/S6btv4KxqLIsHdi6ydjWDyLZtEM1PpK+md
6RfF1gg3XJCBWhIqdidiCghdtJhNyvbLcSb+8SwhHltzmNim9AP42qEhU1yR/euApzpGL3Kh2Evc
c+K1766+IJRi1PN8ONDmxdnvz3aoko8yL4gRUBF8eGZvER5ZmeMGaxEor9PdReEGQ7JO32yI3lSf
rbaF6dI5h6AZc6ZT8ga8qeYkTebM5aYWAoEjpDORUqPmq/s6dmkBXb5hctfVJA+ayTj0ikraP68n
UD4hsbWpq/Y6HKcYr8GIXav8+DSmBS7KIuI6kk2yl7brVS/Eh/OPSjvD1ZuImZGr/S0I7PNxcyUo
FVlTNT3fMKXLK15/ffyEMSOGGe/KJTMaHYFSdHeBVTZnNkm5OhdyE9pjuoXdpRtHGqPkPbkArFt3
Ht8PTI6ytdM5Fh6PsH+Dr+jtiFQZW0HQnR8ETNcxFEQIunk27paArKoOeN+pIPrML/vIRNhqhx91
2rd7il9u/fZCDHZ1Uo5vTRO0KpIC1ESvzB8TV7lYjUiGGfL2mBzFKqzLcuC7IuLTs8E+4H8nzrhH
Jfi9mqKaieGeuJRI1+21+ivSnOGrNDdBLy+AegzkSKjmp1hUdPY8u7Vb9BB7YhYc5Ag9YMm/Zf+9
146qGnWW7R3Zr4Xnr5SUumYHNC7Xsp2o6lJb3ivZMWZBJJL8WX63yJ4rjpPVw2d72bZVnFNGNtlE
7EHQMMniVBmcmZfGAufAga8xgDnNO738l0RV24ZncNxzghr84kmFRpLD028rwrk9NEMvZHlfERUK
FOvPwSfg5ywupvrjoX4adBe6ziFjccqC8dUBavsbkqvcI2cYxoBvIIgbSpl6ccSHGTSaOMwAXJIY
smRf4YSOAHVvgFczwGTc3OmCq8JlyTpG0FhHDIjOlhHCdSHDpj6JY3seBo61JbvrvDJHN6uCcCxZ
wbI0Mwf3TGr3CmeT20ysgz2ge9fWNVywman9Uz8NMMWx6wrDUVJ8up426vGlSQerdt39iXy6gBZ1
WrTxGaoSzFtfGlTJXw4lzE1CArMT1TIHm+LVyJvCxipL3bOun0/TE1gQC22ytDi3PQpT9bjC+8J2
6N2GDjk18ZzxndktvM48crgptcOEz0cBXBXPnq+V6XCyt0VtCm3JYn45x9Ku+xwMHeT4P5syhk4S
8L/pJ/XxetRlCJp/6sDqAKtvLAkmiYTLrebU4vVbn559FdumSB+NDFOKoGMfCab0PS5qmz+I1DG5
ZigrfvvaoppPtEnChQ1YAzlHa790SO6yV3eCaBQ0/V7KOA7wHu6UdrdnoH8z1bxih4Kz/INBePYl
erdpgNGZL+Se/4QPQ7LNrXUr/4w4ft83WcX8v0VQiZuudfIxrW//c50RxENWk8AL4BcqheUjTv/k
JPEkDPpacHFm/cGcO7X17YfhZAF9I9VaMcNvo1qx1go4g9yhLa42hklqFrnrpLDHKnGa7EOfalyf
Zd8rxLGRjBWA4PAepOsO5ojXw6Jq251ZFampL0ALqbdWdEWt7nq/BHMW0mvLH0VHqoF939JXrDAh
eVvwc7lU7LvQlGDgf0wRYI2XCPChsxL0IdDx8PJzcHDeWdPl68EVSoFNYR9X30CRWYWbgyNeLB80
DyrQIF41AFuAODIBXTNYNRP1CvcoaRCQpwgn6COk9W9t/Ao6uHDqr7zcUOKSLo2f8EEL0tLIZrRl
rhzN1+8tVRl1Gj7BcdvvlugzVLO98asIoX70S1k9hNyg6R9MzFIIPwnuijVKT+IS5GUANxEqxsA6
PJ1iOW81Mf0XpQBVZMBEpCKoZE+1ZWLrMdhNWcXJkf+ydvSHEfo5r8SLt0idpWFrZfJ3VQXHtdvY
rVBqt1J2fo9D7DCagTjadL87T/+9lQ44iV+UmJBoi6ILChxKMvpM47D2BOVGqsELxEpRAajiMDnv
zwv3FmOe5R1rNA8IjZevFYMHTU2ETX53vWEZL/rr4DnX5pakQ6QRl7E5nCBBXjzZiaAvSZAnvjc1
+CGHru1STYtQFWfzxaHVdR6RktONg5M5pLmjukwiZBro5HeCwd/plxXmfpUnBjSo8BZoiUB1j6Da
FxzvHzJhd8siIyCe/NPHFBL7Gg12PUng/XVbgOM6XiHkf9X05RZ8hDUCT+V2BwE69Vpev8xKqkiY
MlORn28syPHJnPtgvMJyn3Jqzyw2TEOQd5WW7LLBCHTL+rcLQf0oRwiZj16aV5EHJkqzoQxMUiT1
FbifdtZaIUgWPnXuFv0fMd+UXYV1HacmVyIyM/bVao20JUjSB6IYw9LHVhVDYQ9Iw4tNLU+8Fg7A
wrMmSppBwL9sy/ps5RzvIbpCyUGAYIIhHp9jUet+mSW39IBn6yH0+UYBR42n4FbTRw7rQao5uJFy
Ae/8dss55DCT2o+RUR7Z2AegKg4aEj+NqXua8mkvxPdiyK6NKvB4IbIlEkjDd3tMn5rhgYLGFC2P
A+SpwsORfIpHU8oUaRxXla5LNmg6Nk9KM30IzHArpMeIAaIXZlT/pMvtLRoy3NDE6+z7AQNgxVo0
BHfLCoSC0wDSb6GZa0rZ3DlpgtWPKjQYvbUSEMEYs4Ey/UXYFsFXWDXb1xP67vITqT/o1qdAtb4n
s78/Hrjy1tWzAQ9JckvFYvrOmDnGeYXcCSeH8tETKDbS66fB89lRWYAu0mh9yP+g4c+49Srnbcpa
TNk813arSHVfsOmniiAKoYTybIM6h07eBTIaZSEr5mWcEZE1db9QdmL45HPYOo+L6dDYHmSjgBUz
rrloqE7CJP4wapR/fTY09gTgC0l+ZV0Gq1g1AHrI/sF6qe6BEa2QKd6ZeI/+hXk4DsxfTvuZWzRd
hwq66cwRPHhKnFWLDyWvv5wbJScZgWH1nDO4jpzL0Jy5BB3Vq0Fztn9zqMDV8V66CzJLJW9tJ9Oj
TEQFGQki8QIr5uR2i3PNcDgCEiBPIYVU8uAFygMedH6ZgSdAK/mvsTiCTOlsayCtpJQnLltRh82Q
XbhFytfAuOY/f9TPl3CvMW5fjUwlYI63wWSnc5Szq+8MO3Ft0qmBHXLyNogtPuBFMDerF66muANy
G8Cc6H+8Vxbysj6udIPDT7vC4jmEhw9EY3RpJwL6onippUMCutcBxNCGIBfDQTerKeIFkkN95YIi
sql2KJneMGe8ZYlbzmpM9DxXRJ9N/fduW2zJbdR6ia9X8as3Q3wTrzPuN+DV1DL8M2rup4EPBSkZ
6hiFQpz7hAFc8qWwBzBXzzsjyFJR/9rpLhj12pWLR2MzyFwhGkjRP/4D7HtyHMoQ40v3ARxdMkCv
Mt1TtIsYq8H7W5w6nJ8jC/uMfPnIy+VRxFt0Lwjh5o8OSwwfgOWKYzmSBk5Vw5lKsn0tEoC44uQ+
LOIOQq2D1bqUhdJ64UVTTc7Raj4NGKP04YqnldTVhnKxrTXZo6vFm1RshJjsDzlWSVN2VtGzJHxH
yxYIlpdX1ItHsInWeE592aNtyHnlhGqgsuoc9pNQtVspFozPy1iEWBeFzpGEMYxVOeg1tan9idwb
f+JS4wveByEiEaGY31jCrHClU4uKM38xRm1TC3++CV8wyY6zNMk2jzb1ayShHEUqwfo7LA59jkJU
Wa0pLkxGUvlhHLMOvR4YWK976zjYSthGo9ldnFZrr8urdKdDv/NqGNVtqWC0cyeSWopfYtpeOED7
6El5m6vLUtLbNEHbcCiy8qZHZNxPBe/y7dAS/nWvqaStKll4EqTeo0i4paaVZnYNxzRkA8c7ouVf
CT+A6e3BnI59h6NPorv8VGYdePC7mzzhhJc53CatEAJbOuVHJd/RMOVcaTbOpxBriwh89guOdINU
AoCFwh8hOBH4mMAPDIFsRTgty7UPG4h2ZECUmwIl4qwB4b/oIKM6zQLyz/sOQx4+vsVmmJk+exqp
lgqdgMtSrrf6lRBTzsSeFLRDAmQ2C5na/Y07W/wCu3vrfnjk79ee5pu4KNPMJpQPN9xsPV113F74
pgsYmaLiFq+D3F8OOHyOzbtztp1QmUuFrf7E41KPU3ATH0b9Yl50P3h/WeIJSAjj2PuZp3VI66VI
L/bZb/qDPJkvqdJnW3GBlqTr/WD6PWf7ZU5xTJJkov9vIugBpg4BV2LM9MHbq+CyyeCS5zBSDlrg
3YkOeGxzEjQEsmFgZI8dqltPxk5jAQOG01IHZyzMC5KVoumeyT8swJzpuF0jSJjWqTqA06JAcxSA
kJiKXfgb3eHNmHo70AFrzzP1nYF+i6OaUJ4rtp+oqhft2r4M9YOSjx+GjqSOygfUJIB40a3iq8t1
X7qstMAJwyFXwDH1hKboRWHPATBqcWvDvSwwtWIyrXEc+MOLkSMRzne4yZSgKKSUhEcU2JFFXa/b
KETpSN207c4gKwACuaDRXUpKtD3XIPkrCYquVwyr/bdwLnBMQ9frjeEfBB4XFpfjcErb1YTv75d8
zRCwAm1OP0yA2G+6YqfChxFwUoO+mMJ+/BxEOvHeRMOjG7nvwzauRM8l93kbryN1RxePEGpc3As+
vrqR1SjWgu2XejOCDkOSFi2CjgiaIx8hpcoYqH/EHGBZaBO1C62rR1fojxuOvKHMZPMqjkTs6GDj
fv8xPCRGh2MRJJ0rdhENSGGvVwZNURZQQ92BXAdXOANOpGRdL2O8d9gJhvjaHKzAGpE01ntwMb3I
32XyMQlY14GkSGnfu2Rim3QkbqOABehycNpa16kn5pAQ6oP+HkCE9KPLiiBmZPU/5xG2cannB8ca
ax2KXsc9+lRLBpC5UXalyrOb/7ReDSvkOf3jEWL2nqzbdO1fus06B5wmsv0Z4QeQMt34y0ILczaI
dOpdpNU+IWABb0mpR1OuWvRKh3PYMNfox/Ws5KDzjI7qVulDvq6ajpvFm35slY3LOYgDR3Q4h3e2
afy8i1bbf2px/tH6V6q/BZZahPICbABrKtoiyIOQLhsUOopsXTEmBEHiPpN8+snYidtqFlDydlUE
pBBDn/hYXP/r2MCkHKgvdokTZEMOio9IlaKSKV0nCpsF1W0i55B3aBeMiLsQeoPY2lQof5H+zcE5
QsItmF+WlhPnS3TH61YXOJ80u+Cax8s4AK5wISHBxk5lukzs81lCsFHaXi+dSpxqkR09EIRhPtKk
pujJ60U9mYHQh+GbaCbWr6w/viVYxtj9dlV3uPxtR85oGUbq8vsDMxdjbfFLimITaqjprh/7IaDw
t8Du56i6iGBEMQo/1/DSE+2VUbjfHFJVA+72W9hq8Po4BtnX9qO/urfyRvmATIqvTjNFOaNTsSZy
XM++5nCeu1rZvHyRT0kJoKkj6Hnd1MDnQDwsbKOb4U3ye7vFQ1XcRQSLGox29pjDrU5dd/BHGdyI
9G2rDrwO00Cj4nWwMTO9rHJ9vhbfSmAhpdPgqWDW35p8UyIaLb0bKv4tRiMru6nmWg2mAKHrD37c
msf8z9rBq6FmDLJJKOWyPjenpFoPa2FPMFzNA8IneWDL73MQxCNhuDN6KaSDm+3NEnakVLI08wu+
FpK/Kb+dqBIbuEosaQBmCTASQ+6uoV09y5khwJ+BZXzMMLm5awjUr2O6pIaKU3OCVbYG0FqhTuxi
mvdvf1/JD/UKJdDSEtjTewRPuJ111ir6TNasg7lVjQgfEqreZWJmzFpfLFw+sV8Utbtq8FWSNgi+
1QcrE4hExavjl4EfF4++Xs3sjGbT7Zf011L8VL7V4i2BH2Df7YfXzbSRqcqYlcW8Jy8cYHI6rb5Z
rn7yJsMjguXz49Roh0MWNseEcGQtAiaiEDMkc39bKQX0kjtc+YaEqSPWU5eoeOgMQkWe5Go5ClqF
EHW6TKA7lO1yicJ9CNQl4DyTX/JQ4v3OCeJIi8k5xW+ArhCJHv9EIpLd80vuEXfBWknnUyLRDlpJ
HdgOHwjDrQbUoR/QnYTZgvIa1EOGkaWwKmBfrI0VZj/ppp0g+B9zeYwrv2AQBt3KS7vcjXWmxoIa
xAEWSeVdYeBS40/kQYVrrc6wW/0SwvUyC4FWDfhVNRu/iGka00IF8e56dkMxSqpFeCAVJn9x6GCD
3PBfu/AvLk7af2gR+bRM3qHZvnu57GKiJhrq8R8PN4TGNvAAdB0KlfgrSgx6k6QBjKFFAi9RItmf
3sB5w1RvdfrMSoMXWITDEYRan2KzBQD00q0uZqdwuof2KeYJl3cHTdJAjqrVKRUzgiDOX+Df+7W5
UYkJmuo553XR0FCGYAM2UPbYHT4sL/Krlhqoz9SL/debq/jY8fyY0CDvaUU0p7fXOQ9fRemNDTQ6
q4DGCOOhvZTT0/bxd68xwHJwns3yUUDS4SW3E9WFZvOZK1uj8y836+kfRrPhg58Xq3lvFfCDanZk
tSdefy46yhyoP9r1W4vyt75RTSNSxHXLLAJ1u/mOsKskupiHxdQkNAX0zagmQU3AIIV98bNAG6Dk
3vmstSlY/+ubBcwZsomPDOUsPdMExvW16ztfeaX/HLYspqELkEbEAEBdRFtgacbBKV1Ir7k4yYdc
HK1P+I3/cGBtB1KJmuMp0ifaIuBJO/AsiHC1LYeZ7DZt/bqlFiLwI7/lLRS1oAT8yTc2LdliXbN5
ipuFEfUwqxL5BZ+f/PyzxFrbsoc/8DNLVtiRHQZiEbiLF2+RNZEbETMLJzZfqWQnN9guHfmVyrEI
/tISpr/FafXmWwLZw9lae6pPO4iJ3gRTt/eokXPdu5tqXdkJlJR0oF8I5koD1qO84W9CNmO1SYq4
DDjIWH+oRMupzPFBXcZEbyIlyqZkDwEYFMcqasM2misBbxupFETpu9XXIkhTKj/h2/Lgzf2dnxvz
VLC4/2q2hbfw6MN6OxlcIxshQxKO+zQ6t7nnsP55MEm82JDqzzh3fRGCJ8+t1VBQjg/DE5lz4x+p
Z3T6OdI4vlr1cvQ4+3VdOJCspZyTZTF6d1eHSSHxgTAsE7mfB7rzjpZf3n2fBlm06dpv2XXcpaEj
LNBkjLD+kkA4HW6VY1WMJA2iezzrGPB7ULGxKEwkouDRJKrr3te51E5BgNUTfnOg6L7YGcy4BoC8
t2I6zj8rYjPGbVdY9Hs4U0piVxachG3UPlFcQqjZPrMuk6k2hlmym83dRHoo2oUazfEqjAtZ2wFf
ZyYmnocG778LPqNDwKrzZ2hCbR46xFwtQr9zE7aUrMPoRsIkFi5WCAoM8HcYo3RQawOyOrwEqn3x
EpxWFeEFtLnyPg8foA+6sdjK+NujmsuleSja4qTHOEeuXTZfx/Vba0oZ6F9AhYnLkM5Pv7nGmBTc
93IbgXGosTTg/2J+ovELqcbzlpP2d8TC2h3zX2ZLHbx1HUtzNZ9KEn7YtMbhUCTh+ewHeTUD1pHC
K9cqCZv7q9n2nW1FYLm547Y/5eot2ispoHJ2TlUq6yKTp3Je/IOULBaNG8BwloyPYGUuDtPDBy8v
R1WbY6TPlpxHqA1jZqR/gWRJYVftAHGWgqFCK7qHSz1BE1fE5w1byGpDdGiUvbGqwIXcAVBbYYzl
AAdKIiyXr/GwB+Rx62T7SViyz2noFQ89M93eXObvqw3NzTnaehwLZyU2KL8F4YFhL+cF4b1HsXhl
AahV7pBAq34YPnZ+ShyV4aJxlWrijAJ/kBxbblITpx4z2qctgpjxjVtb9Wkdg977BBYmdJn9h2Jy
Vcfi9YvrEvaPoNEIOVrFefQJ/j9BNB/2zrKtEUGpfPwtxP0aTSbnMQf6Bp5UOMBfruwD39RHnXke
T256MF7hf3MDt5J4pGETEQbNYDz9CjnNtnLXnWuOL1rT4jdal34rFew1wkPU8Wqi8xfLheOp5V3H
UcLcNzH0Lyv5N9vhVTkUegxhkihpqL6NSXBviRpmMk7eIYrhFhXSoC6mjM78l0/d9NEAuRhlF+o9
vxxKMzrfFBBGp3qKuAK1X4nWCBynv2z0zT38dsiZmcfQVxe9i1DqpMKN1qKRQ0cEBIJF6w6iBTtW
HpK6edgeZSr7EMXarGdlvvCAWuwZRrsd7CKVk0DkKsCuAJnAngE3tPTUA7jNxUAT/ZR2OX/MLbEo
4jXnmo530gbRWfa3W8SEUZSouotvcXzi2tiE7zSdDeAjnvXPnaRXVU1gUQPIIfmYHnBz0J9k9Xat
sqAg6vqDmR4GamRjwIUs+AQELrPB1LQLoyCCzKYDfmALOmn3/Jeif4BpHMIuWK+7kWwpb11Y5ohe
3r9Ac104QyIy90vSUVWHjQeM2j2jpr+H4oKZpW/o/dUlEZuJmZHKhtPmGSpVrUVDkVP3puMdnar3
3WsUNXQCxvtZbxBp5rn3yyrgJm0OyjY1CFpCPaIebUA9CBviiun7Nc0AGJJG4sujofA8rJz9s766
P/KRr9jn5McRuhw/kOrKXii7uz0+/+XPfHq9g0dYeB9R13X2oKBmr+jo00oRrVbP1pTexq+LfKu5
5+1rbFGO61LosWXROLotPbBluqd81EJTmqdgzqmGMhVA2K8CelxuuNXOVERL8xW/62hA/0mtW5mr
cpAdaw7ILcrT49RY648cYI21slcHxgh7QrIk6fnLIW6tRwI0duG3U5LKkB2I6osJhcS+zilbWu46
CAJHOZZ5dSXTirT6W13aZSpgRJLpCPQfKdHAKeV/e4xoEVkPXUCy64/CWDCa0vxoCpNKFxIPuyHQ
B2PsafbxCIjSRT+qBaKgefwV+ciLGdnaTO1e/QWIHN73OK7oq4SMHa/9LPoIcO5f5QyHZl+zxXgu
CpDLcQXXf6gCOc9GiOAfQqNMY2lKiNsMHEPVon1DWXYuTDdXOtZj/hhf6ckbyeLzikDv/OaHvXbo
SVx0U0JXu/0T6wU8EuVzQbv92Cv4UUgWOrUrCzrvXTw4qNz+1obVYAH4dq2CqEwdq6/nKuZ8x4Bj
WJmLigEljZXq5uN5b7iQ6pQgsmZCnFMwyBwipAWHmtAoUASW2oHB3lCAgLbBNLIwXCoJjA0/YOjx
AHga1BoaYIa40COnxrHr9WNuyVCsfX13txiDLOsRYbpSNoA6v+6wWpZBdoAk5knSjS4jForm2AZf
frZCpdzJOwKNksM4vQZw6EZGcH6SKFVmfxW04lKtA6SiZyJobSodqXvqJzxQBKMHWQjFVdIVtcnW
YA9pBUKjIVxBXI5Vm7ywTtQzpVQuXLvEFkAmMKhuYHXlKX3HmHsZRAHhUqChmhiQlzwULX3IJ4+W
3scFFf2NNn+oUG6ooLISr7QOmxL3TKKck/t0w74U6aREMEOQnr327o1xneq70NSJaUBVdw0ixZD5
VstzatEkJmBJR+kMzujR1yhlpbZlEfCXFoTaZxoUEIy9T7CyM8essggUK922euQVFWV01OdSQ3Q1
zWovRsMeiLKcd9l2Rbj6S3GTRtrnTWfIHscAdmWKhBDtH/vz0xPSVtiAcUTAJTR1I6PspaQQEhlR
fLIJ4wMPXQfbIOdgGc89IHTmLsifXGsBH+6ON4qTZOAFqf+ddzgfUwQ0HqdfDFyMSTIjVXjlUzw9
AhvYE5QnG4DSgqkuX2PC3rNj3IbleUyR4J+Hnzt04TQ/Ox7cgHn0Ru/LomtNkDkFFXgsQ4XTPkmQ
t6Fkh3RTWdlD19ziFPHcHIzSKI1y+8Z3/R5mFq1+1YCXJsguUvRgq7xpuLAYg4wFs+qLGPH/tqpf
1yTTBFoFY75NPhwicXHtPUAdomzGa3NnbzURYcA/m8gvOwk6B8CEEg450Ma49hrzE0S5waSDkAvj
OBN2QFl3L6G5UC6jPPP2DEG2sMh9z2G43D+zWT8jdznr3KnQmEp+EqRKG3vacphXPR2ZAi7ffgAm
lJg//DrC2cOKVSdh0C2C32FcTToosJb/c0taAVUv7rnlT5FwdgmT4Rg7ieEH2kqBJnqSvpFdZScH
vZN8rZIsPnpeBGrqymcUlQXUHXPzR9ojP/46tovrpNhnCeq3g1CTNuSqgfjdNaux4wmOV1BBVaeM
rPZrqVvOYLF2OlEVprnNoQqJij/isXWfu9kGZJAXbXzCZ38gi8DGwGzno4VJkuMhQftik+naJiCv
2Mp/HYxMH70yRF1yrhuFyzoA3PysK/xwp1D5DLcgjvvKpDmRIVEwrVyIHH0HE9kShVwhH8PC3D6B
ezU0V9H5zB1uBQifbMPnnESd26clNATfABbscAMQOEFVmmyajkwscGxr9PnH2vy1ipBkr4STM471
1W0g+U7zSIDWvwL0jWqiQdZzHzby9lyxcAa6Wew4WkaAW1MpSnhOAhss+PBu2yQD791ZKZU2Tiuo
YlBBWZ7SC7p/lIDX0HpCSjQiiDRr1fyZ4C2+zuCbAkNncJpGUR2qNBcz30lbWQjBcaemCJ40rK1k
q9Jm+BdmMqg7naS50yO+uy/W73CojBj5ts5Ik21DN3+zS9g6w+bELg4O9bUoRTGcN45m9hAoi83W
cs4C1491vgQc5EQZ4EFSXrTUHseLWf5owcYH8GHDO+ugQlfiBhPUJuK/jORYhbf3Ee2VpVy8nhZs
jxhHANKzXMTuVEPIY7akecCAJLW3D7Cocdovy0PrNQFz/LlDf7qlagaC50OJEoiYD5py/Qm1QtOe
KnZLT1gFPOzXmM1O4ymlEBUqkMxTmov7d3/3cyG0ic+oHB2v4zZERyCPLxA2gL4c3N5pUS8Egr2O
FPsWxpeGT60WGbdThVUyNZmqqzMaxfx8rmaLRTt2Wh+rG68zzkgqojQYJWXj7g1SP20FliUsYfUi
5Tyxg0ovo9qvMs0oA7S/DuE0u1/BZ48rhga8TU8CJxFD+L8Gkvqr1bHCj3C79YFpCgPiNIL6iKSD
vrmTCOZWGJVqruOwFfdudNBjfTfNAnmoO49Bt02ii2zOMB+7HO1oxJ3D0tWSy2b8SiWSwnvy5w9J
XeM1mdi5PB3CBslRzi5RVVfTETPGK5vLqXLIuOcak/YyKkNaJW+FYW+3N1qzrMs1eLVp4hYvFPLY
lHknnEtU+gjC9lvYRe/SanZXTI7z7+XxPa6HyQWAGmKQy2QovClu2pZapvQMP1eN2wZgw6UCB57E
zqOCpqvoxbCMdWoHOj8ttx+iQVShBitW3bzbo1MP0O+54+KUkcE7yglIuk8DkEozgA0wcM4X/e83
CQKK6L3JHP0UD84nzh5GhQGu/cvRnQtPOsZ0amOv1h623/LORtegbRIM3cKCPTDA97hxTKN/bITH
AbIbI8uwMtD9OGUubfp1Y+uUQgrep2l/EeZeDadz7wzEkTLWcbZ6/p65qmp/NqiJfFGvRC7hEScj
MoeRgw/yRQmrrNddpWfAHtOe2+pBB+piCSpwwXnCkNIenCf8C0XXWQfd9GJ8YiuMJeDrxrWVo0LA
fFsOjvXn2XyLr6BIHNFp1FM9QvJZLyXbWwr7/pmjI2rb/b/jouKUfxXt1y4ehG0OG8NEF9ubr6cR
LvTahV0p3xTms7/aLLk/5smwLFmw0L/L9pIUSqNAckoAlyqgnzxm8fDTSUzb7l7tBYDQkBVEsLtE
ZeuCC0mzu8CYhX0rMF89hB/yS7uvK8WD2ihVg1E6k+OskexKbLFHeHGGF3E3YGKXzMbBNVejOM2X
yMCHDHLWIC9vOP0jt0of/7MbojkOaIuJDskyY31B3I8urh6f9gjz+ZnFAw9CClk4+zDuvBCqazxM
67BM0hvH4NNyGMG3pMlf5mofdzoJvM04Z5McHfNqzSvFjrmK1E+glqwLq1JcMH7cj0Gb92XFUpP5
E5quA5EiH3jhYdOS8bYbSwfJk77tTpP2ltICbmSMt/1wLA7vHn9QTm4U+bDIWF/lrCZcBbISnda/
Y8bSWVd1qMcvUAhoB5Y5h5VQa3cdkYeWbls1uBubXbmjzQxGgCbNfNAhJkMAJJxF1btK62W2njeq
fACcB/dcZtEbfU7diLPNqGu5fLBFN/OQ4utT9QPhgSN1XReIUNxb2XiL1XcM25wFQdBS14BW7jjf
8dcqv0j497slBBa2I1AFHGj9UMk3hYvHjizUs581CVzqeeEzCKBBBcxYvcAytELckohxJN9QpusK
VO1hYn+ic6tZrIhYvmkX3BKl3Y2gkHvROyUEhvgG+gXdZoxUijW07y94BvBtobFRqyFu/8HdO81k
I/mUF4fn9lPxBGeoi3JrXoOVFVxA7jlz1zh+RDHxiqVcbQOyRJfVSXShctIZMl2oMV//SA+L67Sp
aDAcjbua8qj/S0TDejBwlwHUj96O7SQKb0/Kik/siHqu5SYai0onS4reHogRhpzdHBE/qhrxv7sv
QQ6LA7Cff0E/0+B7fc+J7lQ6b8YdCjzutr7RU8w1qHqwnh9jM6VvWqVeHe3pmxdAffscSlrTVG1g
HqXzd9WRsmBBMjAAAT6LD2KLYTppFWQ/ewoWTYr0M4ddvku49kdHU6iOcnDoH4L/iXvZE3MOkKCQ
sWvptbo9IfX8jn3u2peOINev/tO55/G9jBAfqZzVY3JgkkPOmRi+QcBhOhBv5YCQubXFVUEZi11T
EAyYRJIRobCzk+OOoTFNa2FCGkG8TqCFv5D5uvvUx6mLrkhaLYOgcxLkyS25+n2kmOwwKr2Bjp3B
6HcDr/rQjJUKXS0uYhbMygE2M1PESYa9VM5lWPYFlmvi2epV+ADLt86xn4OG5FDjCN0i0l3FCTEa
KbENY14VEE7dnpNp1wsKfVmfXOI7ESxQJdFD3scBq6mRuwZo5AkVh1CpkDrnxw3iwN8iD7ghOdcb
3zgn2PCOfxGwOyjAoPsQr8iO0Lcz36dc1L2+xcSRokUUHbwbpL9jF5NUWW7eppSKOVK4qC+Nh0s2
YiYltCJucSjqW1UwHjYctCaTv/biOPXzHQc72KZGtQmx5enLpZCUF8pQzJWwxyzh17rfmkw72rWJ
B3nPriOzgnzJgzUd2Arl9jpf+yE5FHwXTY0tVVLLe5Ekh+iFa43HUEbQbCGj7Z9RBHlEkomS5y+J
NPOWj/NCqm0FT7qtlO8xq0ayY3+jZaGZUFZxhy7tycOjFjmLCUrJXXtiAC4agzXH6kXeh/xgwye/
QfWTDZq0BY/B4aHzILLjr1OBWXte1fOSf0uxv+T/HzXMMwdxAoLGnPlc9WLyoD+GtzdLBPb9lmc2
2Ck75sN58cDVwCKLhTcUKkR2S/v0hQMuD3rljig8avFNxiN+D2UzIpWRqTN2gvN92YEZd2PLrSKJ
P48QO64J1aI4H5HCxoeMcH43SIeXlxDnHR4LuHw5EN3xfSkL+2cXPFYk+YK5V9aNCESlvTdS6xOa
kEmX/9rReew/FrzO5xQ+TlZz+PISO6Et7sIRSoStpg/oeuM5IAJXgZzJMtqESFUYqrj/4s5OxpxU
0xSAxKdJrHMBmsuLLf219WQzP3Jj3t+n7xCUEuC8sUB4i0RF8piZQNMBoH029k7My/mW73e1Aqeq
T56Tonh1DLAaj06USFuOxjgff0OV0G99daMbAE0ODG0nmtlsOA8N0SUy02BmUl7K2KHb/GVqsvu6
muynLCZAD5RBDEtqy3NTwQT8eoNprNuMjpKKglwxmgLy1MGDlOK0DFPHmbpyqPs92mqnvGbYkqsb
e9ZUt8IOkfX7labInW3yCiA+z17R/onom+6mPq8DTkowcJ2Q77vSRqHlUogPCa2CKEgTrSc2tMTX
muWjR92p/kW62OCKY4MsHlLFEkLQPBo8R3m8dmwfAvAQVJVAkxrWUyCNpWr4YG17p/DnMV0JdKy6
kUeps5G5r6AyOBD1WB+eJgK62UT6vj25uGrxng/Q39WV7YYKYHoUp3+FbHy2U5xZoIPuRz2CY1oT
wL4VBaCbY2119Fo/i+2O4uqGeCwnNO7UQPQEGNfs7pvggOV/szgzcJBe7RjoYEdfhOECJXu01t6L
CBOGlGQWjLSSKdsAZA+V7jD17YyH/KWOw728ZjSKnbkes868K/Hbf6n9veejIGKSD980ZBLjESJa
mZej8TPxXQF1cAJzNCx4lz17O8+P/GUmtsXDtKO4uDMVxGWAiWX6u3lVs/QZKTMFVSmkoB1F8lph
YHExwB4GV6e11UZYkvvwRtfwpgHVkCYnCUHT4uGWPl5zlklFms/W+BJIhlTcb8Sd5YSgBBBH0LFh
SqRcs0iMw8nwBc6dKopvyJGxVGrSjDugK9A+t/85NXfBCy7ZroVpm8C6yZFyR+6Rszrw7sd3bPvX
5N1LrXBbN8H2FtU8mpclXZdsf4JluxMxBO35GNYkyHXEJRt0mZBvQ6LvjSWRyVTRswSzO+/tQeGQ
JaiinUoEHFsh7aspUvUTZkokZiCSkuKwvYQcnPjX98V4BA9vIYN4WBF77FSZ2TdZlFLt2lS4AxVM
XB6LTe7Eutfr/Ql8Zap1jXrYt9RU2g3ZksHzVKYteWhD7RjXXcr1Y63ZPSyJHGm1vcuOnSPZqZjb
pwNPnCVvnO2i+qxg59yydYbTkmBnFr4vWeA7LfvGuiAOPTBOFXnmG9qzr02j5AcKE7157vHAKSMZ
0dlmFLk38bGUvvpdRlX0+IvM//Yl3iV+Nfle546KS9SZhlvCeWN8b5oUw6KLDw5t1L6Qc9X3lUSM
+eac/wOW/2HFjzfSAjpatF9oARqYssVkbXWiJT69+NOpbBgeueDe/kUrJ4tS4oQHGozUnpyccjx7
aLGFw7azF84lGRVj7HZD9h67b3XbrMw0NIr/PLxuHiXREYUrjKcGHfcORysAcKZvwJBHHbzHnHTB
2TvWYC9w3Wlh67I7odGXNsBOdIrTqXMbyCr/vnk7DFXRgiVInExVUSK9Fzw/yixb3Iu6e9wQaT9r
j9v1/VFmetFWfSBmwFjI3QhxaFDRo2z/jp46jptPFnYfTMIeY4329Nu0QieL4L88d0KRxJkv+0AZ
R63uSOxjyIG4fRRCCGmyjm2jLI2hsfdujwgPDyTCzcg3QJ+PKQo73qDg7BMjrYrfIBceori/RaEh
0KjVHDQq1vP0+BQklFRt2Khu6NdlGy0qdxbuQbYmrAc92kWhaM6xwnQARws/pd7MJO4DFZlPffcF
9IecaINYVKmPWyn/sqSQhwLJgKtCXWScq4BgmZQxV9wMt5R5AitXk+FboAhlKhAta0tJLP9pGiSq
bQAAeB0IpDbJ1SR1X7/pyB7xOXMe2coQ7v0IfO//buFQZd7Jk3J+YE1913OdSliNXS3lNML73yGa
OmbVnvkYMea6cBph+43x9OZlPSCI42YLzhZkId9h7dnPI1n0wJ/J727/f5lDwo4nVkqVFxIQWvc0
xvvoBl16ditJblbSlNVumG9Zvt7KhXCHm3E73lwiXFaBEvpPNhXvYXniYYOZ+YV/ECrs4suI3aTv
nVdRdgu1Hj8Ow21bTWsL4LXGfhgm2gRzvcUZ6bw58ZoqRSMjLdOBv63cbRwYZAwHljGQ+hWXP+72
hz0KXR4pnau/rapvT2f3trcebtgDEXDLK5gNBsEKn8F8YuFheMQzOAmmn0R5xVK2kAhlgIY6aiYP
BQyAnJHKQ5VF12ohVLHgOfIgLSOkibCbpVgydETUKOQaY0jZrvfffsBVEsc4OTgDymmvh3KfibFC
kyz6Pr/q+rDi2eSY9WRJVks9E0Kf2TQZsqSUV2PehWL9xyHfLUyis+UHXgs+WwM3TDyi8/5iQuOt
6hUmNJCqZOGMS2+G7EYfKwjLDZVUKLEQlpzQQH7zIpTaD4649EfLRLRDrprsumw14dP0yawcCN7E
5lWg4sUq/psl5+9DF0JpJ2Na+kFC1eNxxZYT3giFadOoYf88lHpUsN82F6sz/xM+V5u82TRKBxR8
LOvxgeQqs+vXf3bHjaRsXpUWmQFLqCXlu6K3Vug6UF6yAuFK045J98GsefeeRishqFqbFKtrd2Xb
+woX01t5n7ArlUg1So4s8MsdhgU5aX0dysEcT8Ss93cKHVkiMTYYC+JMJ0BHBOZ8c3FE4yl3rUdh
FcIDQ5hXiN3MaeJBMJEaOAGm9D9oKjI7tkSqWtcbvv/iclYB855S4KluDhJUBxrOjHNCtIOc4j3f
o15L19vu8c+JFfwGT/3ZTGEHV6McpU0suBUHDdVtUC5Q7zynF21ttAcZuQm40CpFTNa+RV0CYFAm
kM03Szb9B2DWHTxHUgLIghCBBNYz11A1mGCTwZcQ0B8Ikde0pJFDGGkSjnJioci3VDwvxspRYPKZ
wwaxRA6OI9cBl3lv/NsimyWeaMgW9SG5onW72ILdPmkL7nEVRYS1oZEOZ8CTY73dp/gGtj4MsAVe
DaqcLLBH8V3A2Q+NnpwIiaGRDdqy4xn/vvXcIgjAaMV4Zg/sFuCxOIZ1YdG4k9DI20seDyz9Eei+
cgNL/o1mzCBcjZdjhZN1TyMdB7mroAC9WhwGMNR0c8hPMJc7YuA/V4CHa6fvHGU+jLo68iEWTod7
OzHi1FAXB3fD4g8ZlxjVF7ee42zWNfIulu/FFKYmIKDclyDkvb6h5pupN7AhmxuZt0VpnsA2edfO
oJvqoMr3sI5+3g3B5EjLdV3GAHD/OKDJqRQzWLoRoMYhb181PlIs/6miv8dgorAYvI93gvAAY2Bd
NojWt/miDp2lOx6imzIjQa10clnY9RiiXDWVKLB2MQYXpGREkwRwEpy1OKAaUSkr1+gcqm8iyZ53
i8Qd3Ldc+R9YBO/Oo9xUeHZxAfpvK1nwt3mwPrHpgi0IdngOXmVrlspCc6UDvzs3WndAG71UmvrW
gxgtW4qsD9r5TxS7ziDOpfc97sJ0G046U1PMXKJfiIE66Ou6wTfCCjw4x/5RiGX3J2GO9Feb693C
45WfNMlP6ojKJE5UJ2UcmV/FUTfVIhoIG1XjUNdRAfDrUttMaAbBFakBfIxs1SFCGT1JAUmhLo6M
/O3Cdo3/9yM0QLsBj9nu9H0FoSPWqDK5L9if95sp1+Y8hTQ7ODuqAWyct58n3v3iX3yUmybqDa9T
oEcqkgcayzu3MjCiGKISudewIh9+0BreJ6Wep7FusKGLZcN2LEI/+yFNp0YX0kHUquGqOJ2WWDKn
uac+VPsig4iGJtnQqTB3DpM/RJwD+bN8xUtMfqZ90mGUCU8neduLlH6n93CYeTFSbyQmj//ZShbJ
K/+4T9IOcjAGisBu8AF1abQBcZRq33+sULjoU5Iq9whheR51Bpo/7egL5/VIgucatbRFyh0k7qf6
wJ+RM9rG72bBoi1YD4Og0Hv7/+89pcHlfrTNakpMeHHgGepAAfC38QmPV/EPkxWQR9YJLzyJXZ7f
qCS91avpM8gQLD5uqBsbTLtHwD3hds1ufbjSQYAZjCWUZHhD136XNnGNkP7E1VzwWy5PJU5g/VPe
D6rgc5VOmhyosDftZD+hrLFz1W+uMxR3ZMfVtAcC+z/NE69rrWFTG45A1KlfW/860lnAWtad9U/H
6c4lI9okHc1gEgK33TNDBM2IXIAe+WVbCik/2va3ESXdgtsoSztI7aUZD21fjA5dlL5T1PVR4fJ2
7nk/rFGD51Bvb2f25VoMpzT9wE8c5t5GHbTt60poJHAIEGI/l+RHsEuvn9EMhnTIwXtfJAhTF+v0
cPH/7eZXQ/UpgiiTFqzbIRYdkaVBvL73KhCMLn39EsAfqSxhqyiIr+aaIDhjfnIbCn7x7DZyg0F/
rpa0FRuX7uNVbLa6+l1MeY8o29OReYLCTCO7IqeeuZKDrTlCmd4W4dlLLss09sBpdffvu6hNBndy
fYX1dHr8yiPO8hq18VIeAxhukdJ2Ds0/ehnf94Q9R2lv5RgSfXdb+fTpkAspnhuh5h41ujLrLffE
eM57s1INkDLUp6mUrIIXoVKlK+tDpmMmEXWe6spL4TBVhok0/ZApVSUeAK2eo3GhmWOJe7wncGsS
jjBEWKtxlqZjjs79eCTY+GLe2nIZACPmP+L4MFJvOEqyPo7Dj5RKS6b44oKfIGCo8voZSbKHsdBa
DKD/Frj1iGf4nsqUdNq8jprmR64Y86sD3TLpgw8lHu8aBowcTk9qs9bglpk8qF49KuY70bFrp0cE
TpvR6VPHPqN1nINQAoyPiSUslpyHkphrf/4SuWXTm/YnhHf5EenXtJ3YKweXG9csTk0oeLVX40/A
PIMCPchCMy8TOTxUNZzSiWlSZC/UnQl5RtNzFs6rqucRFQWerXE2f0ZIevpsrO4HXlcjVXCAQkHb
Djs3zvmBpDYMmaxrZ2AVYHyKgz5NCV/8iK1EYDAJ8Q02Sn0VwzgkwKazoSfM513lRNkndtPplCAy
fO2fhMhec9wyJ5z37uRtKVpuKrsFSt7KCmv46DClaFT6XaIKLSfhf2IK3xf2mXMbj+yGW1v/kekI
IIPKxFaa4h5ROPUd2eoPErTrcJe8+SRFghs8Zumquyxr7NzIAyrp+x97wjOZwbNTZNYVDZ+Kpim2
ACF3TUUZgn7sKIusPFZypkLoR+lp7T2Sfy71cTR8Nuwm3bZjLl5zLqabNo36J1phHgwmepipNIgT
e0ga6pgRt4MrlglBGKFm88luEDBmrtNmAMwykra9oDQ0n05RGnimfkJiT75nQVSENIzbZVrSGDki
edMEYbQ/25It2tee2ZmPWzfpM0Yfv6YubPuSizEYdoZMCeUEps5sIqO6u7o9AAHi/mHlSLkRNJ8H
1Dce4fqj7UhiFA9FWwzmUqfAmjfLNzPmSdE2HRAE7qUZT78P3wKbtIVlj0flVKFoTJ18E/PPYg69
zHBKD8BxqzSGHJccluju4/GTz23w+2buOgaqdG4iyl0GuNzYgc4db9duHVLjP8h0XypBSKDVRMA/
PXjq0bOSchh9VwBw1OaV/f5bNVZ6+HjfYuGniYAIW5PLdn3mdzr3fxhrMWPEz5UaWRSiLuONyOcd
E1OKZ3mVVe8tyOQI8yqq/jCUH1WkDwLq/mwsH/qYzJDLkE6rsV51ohP3PReTfqGtQjHyWUnVMjol
6imDyyKfpKXdw7q2dmO9YI1uc0kJJYkstHlkwdSs9UXao/HHlgr/XB4BjRS/yeSxZE4oJ0LA6JjK
kp/jQa56qM02LNvzATnBeUs2bFqWNVsPS3/+hB3lqP3Nazt0/VDTddbeHkb/wxYSkD9xuL2yfMEs
oR7YkCm6uCwclgB4pCy4zjDkUGCrycCBaENwuNm9gfOMLjjVcFR3T7+mvd3aYRnBIMYNxc6ZiBCO
Aks/8Cx6cZJURk6/QKSRYaI3ehHMFCuYb3zHzomUUVHN/PRNqnN3d7M7kR/ZFpYoKtS+tmpfl0IL
dXPooS15VxLxm9EhAk8CH/1YqB6aTPaeC03SswuJ10HyFF1yDFRd7MJ5e+J90IWli6yTCiEkdOLa
pq93eXBoZU5G4HozgvUPBZbd+kkoC1cfmRvcYv9cVw9+mDRMpCNP8X8gn1xEmf8RlEUiWTAqLtnQ
Wls/nkG7Bap/1Oeat0qyj3yWRuPgunfwZm9/ytqtdSXI9B3xIhr5rWXL4BqSCqPn/6cOQokJWQr1
h/BEZvSsVtMnAGwZzEU+IqHeWq18ixGkmPYch5qDpv3MQG/sIT2Xv4Tn8kNZ04qSJ7J6g9NT5xT5
BOkGM/HtbFiTG9Zo0qB7nEl6y1h9ZJ2r0kourcEqVQum0P0cDBCnmBDVjhjeciaZ1cU+XB3pbCUT
f8+arCdetjF4DVFVmK9TbKLX3xtQccx08ESeQQs7m/0KKFMV6PzScfNsXqzo9/ZVP0ukyWecIqO5
ztKrC56B/Z+2smGRjLES+1/AXGR9lSU1Pp43otEYn4MjzFDEFuOnOcqYWvE4tGe4X436RVJmQww3
4zIdDA7pxWjXn/1lFSi1T7P/ZKogz0iOKgSDkf4cauRa+7cTkYPb8d8Va3Tkd5ZgFJWNQYtK6DTf
yQ4BwpuleV/sTwgYNUct9e3knH19GLgOTBr0eSo9d4pfTLXnMzxX0OjfG1eFQMv7AB+TKTveY0JD
n1LkvryB4vhZZqRAke6eNbsU/VOblqPvdgRhlqLbZK9FNzsEEM2TEVbcbord7FfLuPdFl4iDbi3n
iH78mWSdk3WS35M5FjocKqOGFb2vUwxnzJeen6i1osdrKQ++d3YcRyBe6TMbzj+Ek7Finl/oXvRq
La2xXk7lBOv8mh1WaHZuffxHd9pj/xE9hglizfV+6VRSoZUHHn0xJAParrEvlCeCb4VjGABMeYR7
gvIldkPXBK+4x9K0OQSFSlP++ubZeQ3LITQwN/7JSqdytrsOXCUx2tAvct5V9g7Oj+nFkCMZ/aM4
qm5MfDTVEz2RNup4FBcZu+yDKYgBFzVO4v/KLUfy48UtplNXR0QpD7ObSzVmitbd6IXPTZrgW0W7
nLG45FNMUUoOCSozZzR/wq2ga2YaRdGPHOJWKLwY48Q3ybkpRCe5NxKWs28Kc/Wr68oPwPC0CDYO
CVGWl/C6IOgWXzyliPu7mERTgKsM65B4awxu3qVWWXa/ZuPGFasQqomcQlccEpMLkqeX03+4HBzg
PcBl7HIWlXeGqNdTchSMUMXLxgc5oZRBEGIr8kuxBneKI1a8Y26wrANGFCcGnzT36uQdjB0J0o1X
TSJKyL16+ptKHfnri+ZeHkNQRgGGKJidbdM6AKHy08CJUwphQCBA3/RKJKKCWwxMspvLT4hdshF8
QxfR2dXo4p54550U4NZ1KZs0id1cG0EkIkOfwvm4fAAZ8WuhHMSvT6OIGGc0jEEFU/V4nGsIXA4J
iNdP+tHlrqfj/0sBYQx7m2gWQ4OvF/YrfU4qIWV72gY/25S0JUpHcUA5XjotLWcqzDzthFHHq99h
MWDlCm62hj3TAi6gmVnmv2NWjXMy1kP5ZW94mPwdjbx1y457XhgzLyycmOXiW9Wk5Aru3A0oQLVk
9/G2/VUhpvZOUjDKhC/whwAmm6PEF8jpGyzUl4aq9CiJxL6wo0cuzXHtzFsVQJkZMGejdzdg4d2Q
rYOPKPVmcA1ukWJ6gLq+DsTVeIzaksIqkkbUu6xKIbDodwkETcjL+gN8n1rYkYTche/OaczSSnNS
I/eO+Pc9MNWjS2g9nGAPXMNTs8HIi3nmkvFjFmvAibbNySZN8SbPNolHxIgJCXpADzmQX2QOHS3P
71FzQYHe9jfLo1A5tO8aVvxSfWdLmTAd+CUdFmRnfy0l63zVfykm/BQ7E2fabyP9t75S89mXlB5q
lNUmq+TJQliloFDmBwo85YEmLvmRE1yXUlRQjVSJlUvy7vhZ+6AY9rFolyHrEFvbPsf7jw8PYuk1
ViEK2ThVKYDVZgKt157krUFlE2/J6CAbW4j49UJZDs0ugW6/1jrQjw4kJ+x5B7cIBKTn7X265b2g
eW78T7vzQ9W9KJOq8O6P3bpBJHu+k0xC10SYfYZhkXx7akolNq1B4+ZN/NCmfPWf5DidcjG7UFI7
7ROew4Qtwcg96fevvgAhWHYYGGZnZvwtfbwPBH1iFeB243TIeUd9VR6UYdhfyNBrwbdUWWJMvXHu
zlOPo+07OaxAuvFDvK4dHFaS4S23qB2hpU8jPWFxRRQCFLNBozqn3Yffst0Q1nBT7tAU3C7u6Z/S
nSLmhkMxpV5fs1q2srJRC7CCBngN0NSXoFzI0Nq/PIuqDWCPdK0SxEv0vWxt7DLoh3PRj84GVIln
/+0Omjlty1KR0ti/prnnMIErtR5JPjV4KsWUEhzzRtbmwMve/vcEhCQ7eKR36ga7dnfcGhxlCceO
AnQ4bOR8qrTv8OD7lM5EEcoece/aOu+DGlpA+y2wmEz296TIERQozLCtTeh4Cg10VhOTZYrXPV7a
31z4LkWOWFw0YIby7YhlBYjF8LuxcTIkZKLRTJjsJdGb2tqxyIL9oJWXxYSeSelEkUfQ1pFzaPbY
IMZTpvGyKnYR4jok/HHLRWzOQUmycsl95JFfAcji4b43YyGBjIt2DvVmMhE5dwoljXvUhPkrRRuf
IrlHpWKSJB4tX7zxEtDoQe0X47kWbQmxy6obqYTpJipsxD+Q+pGqA/+6qBlGbz1loxoEfs3dcFd1
7IwJ771rzbGTDiKGPt4clfFB9UA5Rys9aURRUJPLtxUYGtL+3PsttUu+UtTEEK2oLDi1n4PCU9uo
5BPOmVIGNCnOhbH3/zg5U5u0v4VTieTNhJ8h7N1t8jm78ES2hUoMDqAewwKTdSBc4HSoKIozPR9y
rJd4Ub9VSbcvc84tlj9fLS9NCnKBK3Ne2p+Syvxgwbzfls2Nj5FKohyk1Edr0BzIubw0IGVQX4dS
4jnxSMX4TMBWR5SLbib27KjMPdpMGCq6ZP7oWAF4qQ/t0gRsNA9EUfRsmsJZPNzL5BKjgpeeHGJC
rhFExGvSaMGxmu6IN3KYE1MY7NcKXwHHOXo67nDv4YXGu4wCEoromjOcgDq4pQ7X5IBMWygb7Q1f
vtj6XEExNw8TsMBHO1SFwrUx13c1ovYnGirJXKnZK4bCdIVykGhX3RyU9s1YuimPPfvYiMWBKDxb
yxGFrg6QR07Ohb7Vw2QWxGZB5EeEIjJ0qKhrDP3YcWqIZz/riWM42AQHpuqyt85pC0phaprePkT9
CTsw63/itcPCun+jEws+W57U8WXUury/ZncM+UiRA1PyTr//1lSNVdYo1hhx3BbcYJjXkHaa+ndL
sJ/rNU/q39rb97jIfBcYACo56PW+NV1rFvN+C0EwmF14S0YMO68rp9Nzy7H3xE0dYz5GqRf/jUjT
lX5PyPOQuWfKglR+xr8ZhKFtRM+OL652B/9W2h1p6+qh418srChDvA2I0O75UA/MhThiJ0XgCT9k
hAKTbhs/PDWLwBpOAXypfF5Q8hvHfTLe9SmmmPWE6RQi//qrF2esKZTtH0rT+mguwvEyGMt2GPZS
10BJ4VU9a4bUgpz7PEw5qL6N/GyTqUgAjyrDIhVKkdC3j15uk6KYtrHAvkm4uwajQVfBtTMHzdz4
xfytnA2+kD4mTQT8eIfoEEdG1EG1QxfpWVXaU+rBDG0IQx5Ge3DEzGOOKj9JxLlk3851n+6tTtKs
WmSeWPxdlInMvyAv85FfPbJnLCyrKVP4AcmKknASb5ediiSwM7k5RgY/88Sez2pEllBV4TRo2qac
qNGifgXIUZr2rK7od6gqwYb0ifFvQ0VUOaNOcr3xDrWmjID49hcPpPF3VRsahfVYbWS9hoVQspkJ
SeHoKGjRFHR+GtTHYvv1XKPgvR8Qf+ECut/cdje0dSRhj3HOHKi+h+ZPWtmP7M+RgkxpLhHLc9aQ
iNnh3VhltF4bdTMrbmZ6Buq2Wivb9y+TbGuyLTRUnVX7jsnzQO765872KqPz5bWj2Gmjjez+qYig
hX/hPZrGXFwe5KCpXq2H+ZyB4ZE0snMgYq0bA8jF3zeXtIwxzTjcGsAGfo4A3ctStOsmuTrg3gU2
JAeqmPuulwFX2on1obzgpJF1Y9tQf56PwShU2l/vUwMBkfY7NQI1GZymdyJLHViZh3/HH5DybcUJ
TxZUZ0H7c1xCnp7thrgiYI585fcx2SACRAw/FLmRtXgA3Ns+bAqaVJqc7vV4h62KIz2OXZMlUVjC
CswFWc3woRQq+XwOvRDZm1lweOcxltZicfZfy+43RCHRLMNEHkAp86C5rOPyVcOa/oC2oQE/u2xv
1mACt54OdplxH3GWHmIRd8gxshw4fUBcszztOLVlrwa61g6n1p/Lbr4aBXhfaMZQr5dPCbWXBEoD
BusgC4BrRtY+RA47MGAHEJnaKFlZdK8uSsgHFUcgkknvdtgDnm6t/ircDBXp1j7LtZvhKzEm4P3K
Nob/Ygv/F5onDwicFBeME5yiST6Ek+Nh0tBLSaLnIk+38AsaTJDXxP0lRUhRgUF+Jw02Fwd/5+aK
QA20G8E9FzRIkhBritNNu2ikxS5H/VLfRd+BnPd8FtkVOVlWek8UBxDTZ5b7oLxTTLc0tv1DWh0Q
E+VQs5QT48DWt7fXmr0iLGYoicP/Hx8ciqFTs/TsiYJumqv5adcSjbe5+C2HcUBu9l5TNyOGIK95
qUNsCqXJN4f8MvvrlG5VQTHeoNzhh0/LGRpNn604R3mnBSKrkl5WwFvVxZOb2ncNAozmNnzkuOwW
UavhUIfIBt42XQn9JX+xEMa2IVlYNGUe49QuFwc3XoMZm/W6BaRP7Cp8s5AoOKGgvuWijxgfDLTO
lNLKDHIFcqEINZRtc2IBWARICpKdhRc+TKyCNGbnzFk7EBQcVNofi3oGyqYD4gK9RrSm65qeLK3H
bMTICkTygMAJdsRnyzjlfbvJc4JfQcrEDrCynFQWRBO18+Q3+mL5HUj0gs5IFRS2/KQh8c8wHSIG
I2LtKUKnoGFGsVyz7sHeX60YMpqEcZfZPE4jJLaTF94LSHRFzdd9SLGKiZJd9t3xsxIQI1BsYbjM
4m9rbwmfewEeZ36wJRDe5BGbWpSaqIyExAGpLJ3Mu5rxBqM3ZAOaplday7gh5YQfEpsR5+0p4ple
ZrxQbCQdA7RuslqHorOfsYO7rbjVKhDY7s3xZgX8fTA9C6wCJXnrOVtKoWMHtASBWvo+wrEkPZXW
h83iYxQX1zuurhizZ5SbgM1d1tCP+su/xRfv4YfZpVSuSr9+4wdAatQ08HFDTSS8pBLIxkq/V81K
Ilhu3yt6uPZbZQAiGF5mGJZinqbpFw9mfYDPw8BMo7qfQuSEndLdxDPeQf8abSB4vZyL8FeWRVfU
UsknmAhWO2x/SRbnXyAS0b+FiYKUmD8ZkxQqY9S1EnTkHwfDdiZJPXmhGRTQFdbguw+vjiMwfP3x
yfAS6oUQ+UzETUbyLmYzkaKeO3Emoc4WAqQi5FFVEEumO4OhC1UhPXusO3xACHCVZYZE0lDOUJQq
BQBeM0h8Ml1s7pkJBlMrTW5Lkq9I7eToaotfbbCbFVApjjwt/BsD7ROy61MApHD/Mc6FZJSwYBJz
lDjqNi1EPFjzNAvd0y60Pgh1HgaU7JJNao0urbBgk9LgHcHpVb0MjukC2GYm75SReY8spY06NwJM
BGxk/wiLoQ6HK8ngwlS4nGXUeKx29qW15udLNIHGp0NItj09jd/e1MskN+e6wA9nd/zNdxj8zb6/
XOBWeWOu2MxwMePDOl2SYrdyqlImSvPUJjRa1TlSRW7uBPZ90+okX/PjSh172N16BOm0Lf1Wsid9
Sf8jDj7Elq20XqE0aYLjqmxNC4bjhyMcKcDHDkIYnR7SO8jKohKcuEsz1IMRg2nVifeFzKyNn39q
23KxEU+pkVSQHkjNwfCvrEXUxBKMaHSw2pYi0wT8koFzrcHOVCjIknRCBux745SXHdIj6d+tWshv
NFH/eXycQ/8jiMZ4NMOUyGAdWoXEeJg+IR+YefkDIt3C4LDKIxeI0bIHHvZBsUqeclCVR0aR5D4Q
cvmwMPCHqn3nWUc5fGokGmtTMCOc3SyKKI1SuVzKynjvPf9CGQfYInQWH5nMQlvqM/6uDady4F6Z
of63zMzffnBtNjg0aSFSvT+dHgz60iLrHX56u/IvWlL0pWG3EJ3xDOmDokeh6s1Xj+WnxqvmXC4q
ynWYw+bc4hwT58ijbX1X5wsLiIRWMoiPlMkLWjshIQLWp65WSERcDsFhCf6xLELjhqCXaV5vV2nY
JKeqkYEU9Euo5O0tbazSpGlsFtp+wC+xZd6tkkvlYaBS9aEC5YJuTnVl366VJPVqCODoFjAWuGPj
n037zXDmcs6x9bLAffkHwJ8/98fzBwEp0rWBnWN3SrA6GdkKRtSJ2Jxpy4dYt4hd1VxbwqUfv8mt
pYHS3DSVf4mrBc4lbtcb7JxFPrbWMkf3kGH1GBOv0i/VDszous8mkhyjMFh9DA/bpaOOHiskaOFu
pni8KM7rjZHtaMZ54mgO+1b5YcUHDSlhzjiI+LxL4TX/HGMBQD8qV3z1U2P9qnHbQMj+8ajEfRky
oUrFqolbfC6qzFQTOfmslp619sxzByh5bFjpEY0UAnU4hll8ObdoscxV5F/PyALJuakZOH+Uz4tn
sUCwmlJMW1SiA+rQ+Uxweoh0IFNuD2FzDgvYpn6B5NOW6z7iLJ6ZnXLmZgec1DR/ua17ELjprhnN
hvtwfRK9u7xfsTHnEbppgUD7kSMDVqU/rui3HuHc9niwCTMUXfurSdPsHdtd4YWmCg5CIEflHZtd
MnU8qnSl0FseJP2ot+UVT99uVq6pQQoM7e0SwB8Q/JeTLTXQwECBUSInROY2zm84zwRIgCQxcVOP
ARXB072ve3LNi8g3ddcsJ8ESlwusP1igEnD3AB/5+cy2bXXz8zrkDMv5+AHmBOLIylTmvjAd1Yf0
qbDpPioefW0VRK/taK/69hur+DWV7oSzRLq2zo4NSZkv+C0Z4KgQ4ITWoGLQpG/SHrxe/NK9w/Yb
NcOa+zfaV7Yh1EmuuPzooi6eJ78cHHa1qIDob44750cOUerqhigHAkvkmbSxTNwE5PXm6/1E4N0a
kox8h1vfvMxCozUw+mj9TlmGRbFu97bwV/Nmi4sYiU07R8DT16sdaB/s2MkGhkdCOneswv/ibuZB
wxEJWLEAUieyVbYHVEZTHHBHnUdzIaruR1aXxxbs/jxH8KNfRRYH0dgVQgi8NgsF7YRosIjqdpLh
Oux8blFcGWSx84CYGh09PRytmOfqLcK5510MFXnDI266vDMlswe1yjo/hOEDZapVD/2oZV5G+v+N
tqrajjUga4IF1xe9fRaNIfibeJuhf7cDI5swzEM9bGyrOWROJc89HMvSINLQC/pPpdSa1IdxB4BA
CbjRRNe/2xahU7Dom4SDqExQ71Hf2jFXQ2cd9lxHjecWWt6od3qStWj/pbG4+1RoXac3kAMwFIVy
uBNf0f2HLkZTcP4GUPYH3zQih4WyS4AYvaJNPZC+8DEbW1Tituog7WeLHJUEu/Kh2G74I4LKNKLk
RiB09KTrlZCQDXOr+7FKKBPNXj5u8y+Mg+1xI1y0JqISTFEqQVCIYHFxjn3qPrF2E8MamGHZEl/Y
ww41VSNqoqWY+ejlacSbdmmU19HvngWRL00tcOAFAMGPfau7lGc8mkS0qQRxXYf9HDXzVhvN2E3g
3Wx77XaRwVjWEcYhs6vCYcsFIzW/NOTEeX/37cO/dySPcnQEeYeOuIWkPZM+A+somZZAqIRvLwAT
xkY2UbXoGe5Rlt/zI0653PjF2FG4dEorap9wgPhV2zqIJArAA9XVZxBrpO08o4Q52c2wzIUda5Yp
HqDzg9dM6/IQ7kctO4OZkhedRuh7emTc8RIJmBK/tJHXXz3uvzfMAFsIXxpjtO16w6aYvxgpQA0I
dJvinfMdoqRprtSV29Jdmqs/gxIj0E2cgTAwLchj01pjel21rqTmgaOoNCTAoErTqRLWUErYyLrp
3wPKbvIY8waYtK1c0E8k27Xg06xsi/XUzKqqFhhV6+JMjRL6dXdkFNH4lhMOTn05h58mNaJVCNbf
Ep5Zz1Rn+V5N8dsjxECzsUWrxuI39P5sPATe6xq+Rksj0B2uveKT4FJEOGxC20Z4jwCvcZu/7kgV
eC5L8tSn3khrhCjGYQYz3nwWDMnj23SioE/QLoGv2fQyFYrXDe/9LAVqfoo3RAI7b1eeVPNlCO0t
iAJpyXFDtl/694N1kzvX3cms8TQ69+fqmQSIdV0xyYE240JPGKAMPBqFVW4IH8LK14mQHbmTDC56
30mCJkTlZl1NFOx4KidVO42XXsyPMyV4Jd9kENarq2pHq7NTNM9qVpAxYJMbn6tQPqodCb+9K1wI
b7rUaSyQq5grVGCUM3xEXyqenW6LLrsdh7pRk/YHMDBF0B2OFzlR8JJj8zuKvZ+gbnP27TTzhTyk
pfONZ+8RproMKGmHkHsiqw1Mlx7V9A+rWUGID12Nx+upQ0Am8Vy9QcjG3+evV+asusYmeALjqmXx
PSfHn/bZH3FUHK6FM2tkhQdLB5PhQ7edA/SGzGT8rtlDemPgIk+Dpm++6qHzxZM/+zYFNgt6PsSo
/5wQKUXeyxiT5D0HfsJYXOayfe/YINMW0msL1bR7xji1VQZNX9ez+7lMQMVo6O4WbUBpcF2s6KE5
/3QcHUiNfx9B4qSoXXAjtBzYBIar5agpvEaacqLtUVjgiAFhozgJI0b9QXtuXu13t78keP4/uGCq
tDbNL5bSI7P+361WRdksAg0IH41DLzT5HhJugdnBA2UWmPAOlUSKSILvoRGkZLiVWOtT5YPvo24I
9xZx8c5F/9kJomUQBxno0YKX479+KcXECi4b0ZLI0fl7aeOZ4mF/1VDwmkBGgzXmY1BJ6XE+X6Sj
TSCqbzkRy/SX0g9KgYNooPpzp8FyiksEpG+bTPS0/kVmM6t3ZYl+yA89CFcmY/4Sz60zkw1Ll8Qx
6ul14ekSNlQPuvu5h7vph44bv1ZSXm6Ha+QmNeio3VATm/kYuMESqzgwSW+usbxsT0XpHkihtSI7
09laXbFomb76eBRByidpyLOGwE9db+gVcxS1z/8UEcFHUYUimfHNWTh+1vs5X0LAiR/6ap1YTSH1
cSYIkHJwSBwPecfNUviyVmt9uBlV/qqrl9NTiPT2tv3V8OBSYJHq5C3LY5qZTpvI0wXXBry8HfKx
N9KeuwJdcf08KuhjwLUJxsW/r9uAN/R+WS8r2dzq+0q/CnFqkRq3xb5qcH4174S8PoV7jdGsf2oZ
aBnmuVzaYotBnuChr83DgxyDpOfyEka9jscZuwJ0Fsd0S/mb4PXVHjiNTGlJs865ArTQAdMQ82kN
qWVa5ncVA9fsPQOfYCozmbxdbLbCrRewTI5975wZX+8vxHCkV18PoH/q14n7oZ+dx9FfEor1eoAh
ikV/lUsoXC3Oewe7kTdNs6qblmnshx2tUCodYS1WeT04ozUjp3jKFwGPKqrbKa7e9Uou29DSw0fS
j8cXrDI3GLb+DbARntgKQoctDbvJGy6WUw0HRXJSwweNowbLbhI7rtLtCRhSThHLKuEypy9F9fG/
4KJ9tp/TEFz6lu/r/JblH7riuQjoqjH9pLXtglX/xhXWD3kzrJFr+CuqZTtSPpL4EM1Jqwhuypku
Ks/WWcZZYbpPQmH8HlyN/sF6ALdONtui+luvGn5Bxio8pT/B9D/iyTlVz+J88IU48i6qyUTfiksD
MuekqHIosT95NLqR5fP/y48F+txvUceB4dYn6JvcWeqltXacFY9el4y8qPV/ITgaV8rvpzxEL+4X
OWP4+/9mWqR70HPiur0NbJwiRZF7ypRRQkT+//0a3ELdHsF0bqSNg7eZu5uhGvxA7F7+opMCobcJ
32dMQN/+GSLqbMQlsm+7d4ZvY3iU8/2/G9EcltvEngX7Xm/sEiQ9ahUqmekjMmZ0BAebSoLR14EK
4IBIQAGAibHxOJjk6xaaLwX3MG4moRM00Z/pSIy4Htcq+BWm++ewheFYEO1gZUB7/wuq/9T9Gl9W
QCYc5IynBZeBz8hEZOdSi8lrwtZsmUZ7FVhbMKi5RKzik/ZHc3rJZL1AKjYhes2mQR6uacqSCqeQ
DOP/bYBqaCmHbnGqF5y/VSEQRoXGKfgJupq2qyR6A02ocAoN+D2Q2CnkiW+0mMmRjlCMmJhl4Ey2
tYmVkWo1ZJmv/Kejrl1p50wYd4XCNtA7lrCMIZSPW0ercyVZ39ZxmmjJdVpOMrvEf3w5zNYOIvx3
H1qAOyy3Dbanq+poRuUPjY1FalywxdW+Qtdi8SuCAGLqieI6v1QS2S/XWiXy2nQq7vsdkZPqsDK1
XAtRBP9rl1HI8tHZ+7WTFineWHkoh8TDk6Q22ZXbbdLLbDL+NsMxYWECJo5TNvRi2dDZojW0LRK4
QO3deKlSAwkjOQT9kAxag6jAYCw2W5GoERNNyZ8yP6jGfhMo6AXIisnxZ/1ulvTvLmWGU1k5TPDZ
zVsC38HoR5F9tR5SW42FNQbq1JrfaMnClt9Kf2AOsYFmD7qlK+GYS+Oq63n+LvTKsJV+Eh3zVj2n
B3TjXUayN1Z4fKxKXVBggvvElnijX7j1ME5j671JnBxMUhQo+ebae0CnHAmsiUhzs5LS2eXnjh7C
Cml+be+YoFichXfsYnHWgaSrddO4G5wNKKULEJAIo/GJyf/W0GViySTc9RqfvUF9J88Fc3lvpaqq
dsSWYvkTSAb6xE+cj5UrrXYEL8f48HmmUiGnQfFkBSjjQq+htF+7UAJ0ERNvKySYQRmP5QI4KxY/
TzVs2Tw7VkMGtGXgyDSnzEeU2cgLlLWy6szeQUa29aymkdJh/H04qkKcmP9MjXCyDPKZRIK7AZN3
k3EXIHawFKxHm1SG4TxpLuUuY7naO8xmJED4b8058CmseY3jzQR96TeC79AnB0eK5yiRCPOseARO
0rxJzUcN/xi/cub66VjGnpu3ZAKshj9C4ZdPamju2JeLzM2q/1h4N/88Kdpc5i6jO3/fdc9wLS3y
Zo1v8ZgY/eNlAq3d1zE4e4ULZBbtdpd1Kdy6iBy1h7xtOsb45Vs0cVPP6NJ1Bt6f4hDASurSD5Nq
a0A7t9B9+/xFsxqCw2bzZ1QFRvF9wVSLcjwqgJM4v4kGLUA1r89w1sAX1icAz4E4Gp0HMHoH3BGa
T1MiP9Npu0vRAO6s4hSUUm5TWvuBXm38WJQEF0zSnqJbi2TiaPE9EDX+rcdtPFDLteBthBKweTgM
fzKGAG/XYEAJ7WMpXnxzR+BGzndUd4q6nuTmzrVaVKdBk9IU4Amq7QLWWbTwH/CaW+89myGEdGab
c+uAUUIXmDc/C9Melb1WCNyC4NJkPqsdCx1Sa6kbJTkdKty55cT6Vcsxdt1gHXVQ7l0PO0SWeDzg
5B4zRu4kzPHsUGRdXXy9Z0Z2UKyw/uTY2adxXOgP94jglNU0nzzHzXKDQftzfh/0NjxWzxRjkjze
pXweQphZyp+ZdgabX/ie8Qo0ZZCgyJoxeYICooDJi5G5bqUif26QklobnN6BygG3ImOvvEtfq0Wz
hvPolqCdfFtadv6PYwJwYqoIuyd9gwom7EHnv/vwr/Pp6sQRH95IiRu/rX8hakVtS4Bko9SiTs79
WdDNX0qCbYuo9XjdDfb3If2Kk6KaBpPgA4Xv4bJhirXjbxqRgz13hImqkxGp2kQ+H9abCP9ojOfO
Ira9jHpL87tp+oEaorGpPcSVcznCdFipqT3P7cYOToWVQ9HYVxe5q8lu8DkgAm780CiZAS6zTNKv
jJMQcwTPbxHyZBa5EMeuhU8tXNkoNIdQoGTBZYa3HPJmZbtus8c9xTQmnZT2PAvnWaNdPj5lChPo
sgJxIKO9vYU/GYqFfsyq65e9Nw9vy6x4MyfIIc7paE1E6jZLcBaSA0SaeE91Sj+awr+vF8W8PMAD
BVZSIvaiOtmcO0vFhdo3VL6STxo3EIp+XBrcVVGiGwBl8JOIBJ2xJVX9z7NuwIYjoj0QRuOSmvkj
+hFot/PxjwrtYAK++eHpUePDoeelMFBG2CIsTivZiXSrRYvyyjsfG4TxMxK1fUOttXqGYYJU8WoA
hI6GkVgAergYzfs1UpFMVfCPKk5o+Phxyq0xatM6Whr94ennguW7RM0lF7DJJeOeaaExTQZ1/Z/D
eFoW26XUN66dsPWx8Ggpz9QVm6X0Pc6mBeZsl/0hkEXrx/uWjMb2aL4MwMQNxxMSdQFf+lxgjmnT
dCVsFbeCFBPBJ599NhC0VhGlwrId+92jgtxct9JISZ4CtmnBwcqvFSIh8EpO8kLqZk18zkwLIWwJ
K8n8ka94B5rJDutKHQE0M+jpt9b6IMf7ZMrLt0Xnnt43GMtOuTn/QW1o90ObpJTlPo/2z5f3QbQU
AgSN4tEnqbr9a6HNrTTeBJ2ZHXEI+8MmHuNDu+U0cAVOL3dCCUMvde2YIcFuf3fFkrkj8S9tCfmP
3zWTzJR3kt1Wf0oIiytMQ+6+ixrTpl8/gkeorhWoEL2OHMLMXUXmczU+HxSePA0w98BKnlUd3ofm
r8ArcoXl0NgkhIxtb9JQMHMGrO8vP8TYWh7AnIqEud61/2HiGbQyHL2DVbQWmISBykvkurm4FiQI
gow5gpe4Nru8S3FVjpISHAuugvW2cjoFD0IfY7rdK3HTBWJCNx0FrSiwgjGf9QnIBL3YXyUOlntx
rH6w0V2Em1uR+30+xd5x7zt3i4IEy1zIk5GTdmc3QJmyJDsbLSIP9bIgybqIFAgHlEnSpDC+xdFo
j81XL8pw3R8PNULwnd2es2WJAb7MjL9I1a4lxWwer12tZEXg5UNeVoDGAvqkLOFzcF6DV06F+ugo
7/Yk+m+tUpriY/IZ1QCYY6xQHWdSgA/hWDH/O85cHoSmn9xNTg9K98YxWYlPJrkONRQaF7yR7iGU
9wAWneA4VMS1WF18J0VBcV25JEHIOlB93Zhtc73WUJJe8G/IBir8SaWqhi/LiFMKHvuVZZyC5LCs
5bkOGoqKcEiFrqRBcwfIl5wIMFfbwU0/jP5SlMUWVXL+vHl570Pk6WCpeflZyWirTdySis55TNA1
qsk0ZccfWy6fOqYYxackNl2o2u5SqSXBKcB/8pTh1ls+3Z1wO81lzYBcaQmogqByxzkjW6eEUuJ3
bqjLHl2sx6Wc2cfiuQCEqPLehzFIVkta0M1TOYxwheGC0JtmX/nQURMjbIb+tjvAmSzwGWjY14Mn
9A7DBrKVe3GW87rPtZAp6ngUaKGdpc5SlH0Qr07J4ohJwqSP94Ja79UOKSmhgAW3z60H/g4S4l30
wL31L9Z5iofMVlAMFcAxAnjZrp4jwep80JBRWjQoNVboLDqxDYhp4qknPJZYdd0tVJQ+p+iD/JaZ
tVA0Awe1zX9IWCEq8TaR2NVi7BtXBkoieevUr40F3K3YpBJwdUQJolKIgCzi+vaxbytcvU6AnTto
XHFeMF2dLxl0yRcEX7RRoMBGP2WmzPu9M/Ni3mZLn01LMA1mluf/FlAkB15escXqL0PuVeo9h66e
ywB2Nzb5cbcYKeDPKRe8I0YZ2WWd34fwbuJGGSe2YvY0o/kZN+s8qvy8vig9m+UQ3T5ioVuj2FsU
40fKDRowl6hsKOpk4Hak0dTAwDhFRJQ9zYLWbmibRw0V33WEnin4y8jge7KuIDCOAGqlRYX6Bhk3
hvauEAjVz3sEIDPh3HeurYGizgSGib17AX2PoGvUYOEynmH9P6VUEbRnZzfr5tW9vvd8sXNm3iA6
hj5IuV5I5Pb8emXXUihD+pAc+JGkhNwDgEKT+8AnF2YI2qU3+bYnBdAa197c1DoVHeyrLhzmUp4g
lnhcRIPSkwKzYLxmjHoUbkJTwhu7Ky5x49M6RLc8q8ljryJDDn61oknNIhl8pvdpXtC6ntbx+Yuc
Y9o5lRZkqScC8c8UU/BYFziIRKTkZx9Zrph0827vK0nCi3B1L17LTq0Xxj+QahVWX2FCWNlA3Pst
F5VZluSp1T4+cd8lrcb2Zbo6mH3VdSQMXLJ5JJSPQUSAs0KTYu/EIul8/tsXe/L22VZHrPyVVH3Q
07Gmng/qgCIw5Yk3HEWkEL2h3svdwdyJDMzQBklUoWVotqydykOTiMPyUhKF2fAT3hRDGHTQMW+W
OHegBZSUUMAGGtCwFYNw9ATCgVlWgnHRgkDvkK6G5iM1fSFSe4q5H/tRSBJZxDcjuQZ1VafjxG8t
8kmbconOcYK6MDVPox0vcR/iewM8iqNndBtqp5/CmXGqDJjTXYxh3LUKxtgOxTxrHBgE9Ajakdku
wCHkXTTyWEX6Ve0kBGnx5QJb4MU7p7hAI/ovZYZYbW4DX2nd508RpflefmUw2wpMZd4C3VgFWodd
JAu0eRxlm0gUpY8Zd8h01cSxEXoLuFl7onXaeG14p8J5BtvSwFYxC5W8o1zaHKRwklNMwiLQmGFR
aDh+ItfIdsw4MDfhmgDOOaENIevECyKxfQ7X363axWWj8xmQlvhxfFOicE3K5bBdJ7oo/zTrLoiW
bmYizX87jG0h4T85f9VObSiYHFAeF7WEFwJ1jRY7nv+3po5PLagpqhp/tUZzFkqU0bT3cHVDMOom
RSWtnbn9CdcCadarV2EKvN0G9imgZ6OW6NKU4/DpGvJKIvpFzaPRbyIrM0BdzpafKHJFkUXwxpbA
C2Pb0Vm+Phn0V6vhfOucIFV9sD06pBSXAaCqEJlgnp4CEAbFg6wNhDmAVdodmCMEd5zj4XfIlMEQ
m1jE0Ba5gfd9dNQowXFIKsWaARXGgvQou7P7dCYHDrhursLg0qQF2CWJblyyER66UrSVPV+Hb/7d
cdnHoh/yyyieRc67m7i/Uk0Cit8qSPxLDl7SbeZ3oX3uYPXxoKV+ztg7e1JytcxriFA5WgrGLr7a
w6dQZCXsPRXXDZK73jBBxa+DrpSI/T0oGKu3LDI59oeZDbR9Ellr7g3F7C9CmMHOFqa1mBq9qgT/
DUTZsjghQwEo3M/id644f4aYZTgLHw+vEcgGrCy3cQWZSJR66NnvrwztXNuL0/Cd4TsLn+ENumlH
N8Wh3ZiJryRAY8qJTkqWvvsREAt2Ai6EbvxMZtki2jJekyc3bEyERl098HvM7B5HbpSZ4E8Q0oyr
P+/IBdSxhHAX3tg8wNWnlZQr+97qa0kuQ6AgL8L5pVnZ6ZWUVfWWwCPu/8BnN0HVSjjVQIuaOrhZ
F7H9fVLeAuKI9PhQokZsjhNUDiZXeRDemMg4c6hZ4Oj83FmNzbmZadV1Ld458hgmiDeYK8A/19/c
Sjj5bYZ24YeLPuDa/D+rmq+P3pJi/VFH9rOXkPW6Bxh1+K82FmpioDkpXlSp+K4euselStivqPNg
fTuBU11lyF6bhmPVsmtQLZRaXEy4MyD5/rNht7Yyj1gxyfQKNbn8+4Bz8Y+NFNNDGyfLjAnJy1mS
usFAP8TWF9qdVlfELWJDBZ1AkZoC/koG9SgFwdQT9uS3BsdJ+dOGu+xvlOnIk7b40RGk+6dI0vI9
CBB4ouCZcoysxJOnhHYzdUGTrjCkVS6kMzfv+AaA6vfYs0e+8KmZTxn4r2zcynp3Vu1HJoqx0kk5
b9BgsqV2VcHbiuKHjHg5n5QbmH2eGq95KDJG7nOZtjQR2bTR2sAdZ+Zu1xJ1O/4/3yKjh2rfLgsq
o9cq/4DUHWnOz61gTE3cN1WcRAcPIJ7E9EMoZECTXaNqqOGH+ADl9pyxAQgXMiSuHA+AELoNzh0i
3BZul63/vN3aXoZeMU1pzET9aNHyrmkaOPzCQ/KwZhrwvnd9GK3PPVFVGleSj+hYtmvYPCqQvXdO
8gnPN8DRERos9tW/JocRasmKtj6R1TcwgkHuqnXECtj9JyUl6yvavwqoQCQfCHAOfy33mXC0u2jZ
tQPK2q3R9k6c6bWDiIjuhHgmEQyUO1OeQDXlYWRTui1FduCl5i2+Y2R6XN/EFteou4clLTkXPDWo
OuXo7bPVTKl5VXIv0haqXJEDx3oIHt4PiLN3oYjDjs9gHX8lFh3D2SqVw2Beg2m1c8KlOl3AMr4D
zPw1qR40d9Lu9hapVrmJZjPTGnycYb4lO266jG8alDV6RXdPhYGENxmg18/FliVuE3GsLFFTc+iv
FP1iQyvM6cQv5KzlGr4YkTWxa+L4u9eZnoAqfhj70orwNKktEDLlDDE5JvQhQdE1JfZe7zl0McGV
4XyD+6NchTrDx4tIRKnfCVvsIdD91Sjyjz2Z+yg7vh2j5VUPdyz3BuD7Ohfgtue73bv9aRRFEk/B
iCmoWm92ShKSik6QHnpJ/cdiAzLnQAe7gYg/S/SwQlIDRNrpaOAJE9S3cXixwCM00KoBTXNzZ1K1
xEU8kqxo2bQdu8v1HTO17oI0mSX/4zgUzA510nV7N0tx5GsdkZaz92+SUVN02MNTtWY5XawZkNDc
VgListqxrFJZ2D1p1qvOphMZghixMcPUK1VW8Fdz0TIxGmd+InAr26i0U7Ph4nE1jD5lZBYQU97H
n0Ex2H4LQAI4k7IwvG1prAy322tbCglrrSU+TGxsvdPbPqf4fkxrLUMFkDdU7CdbRNva4/CIZE8y
0DXyqxpDtbQuPo6o7PSD0oN0ZbW4ypwbLXGMT9QvuBBnYxRqzLFtcsN0n5LJlWyhn00369uKnv6p
bzyfKHVnWEmVwY//eEO/3GKV8dbuVdintZWiT2aWw5beSND6LlQPYNxoDsRNmLBOPbduSj/YMje6
oryi+DS1d8q7GncxIyKaaTyN/p0xGNvQx4U7GbPDVvcz7EYoEdPzVpg1Q0fkE7+rTpRyYpsME48w
RfwNXRnskdmmZogFcsJyHlXJF2agnyzyiB0OTgqD7G6GfBciZiSf0e24d+C5wzwQT5LWQhNFsIIC
Ydi+HQDtEC7g6hpR1UwgTUfIg9C03dQj3W8w5a+p7xHpgMIx+j/nMctFupmcVqZ08Baf6tbN4EJ0
YVUAO7tr8idk0iUUaNIx8IECwyGHtjxrSae0zgWYAqNw0GILS4+WSI7VcP+PvQTYqmb8RptaRBkG
4rB5DurTgBn6y0QqaRJANwnzEES3GbG1m47qv+bo4/lXLPJk5r76WEge22iRDABEpjhAMqUlf0pv
5Hgvg+ROW+yd63aitL4ph3LVC3pI+Re1ujW9T1NVrvNMA/zDsi2eGuWrft/fi+qF4b7KcJs7GTbt
GjluQVe6qpum/IuQuZLdoEBe9O96ZbCGLVc2f5mDpf/STX9PqVgIAJEGQa1kT/wctmCT6QdDjgbs
AYOHd5d6NgKXXyOlfKhbRgKqWQUbiGPsl0Cd+roWMy7Wm0fxXrcauXCUw6zWZOXykQywkQs+XdNy
ZF3h2gegzu+V/EslUgy8cWngmjtQlaQLyuNnhIvf35NL7UXcocTcw0qHrc1dMTnOY4Pk3SGQZvn2
9PIY/OJYkKFbAVfk2MGVHGRSOPq7aQqABXLO9hcVDEEyWpkuvaerUrlkXwMITkIhJtLcqFAZMNsR
VlFavcfoOKw9eh55Yv3H03PMX4YzLiF31ErpI9qeYIJ+ZSNYelyQcVmm7vSDApWZs5+FwptKGPBE
OpljL71LcE0e+ttNbRAWDcg+wOzYHDWtL2A5xZ6euf3/MMrmKq7T+ZuNNDdOC3JbZlUOVFxRWbFE
4j++7148qdrN0AUrvjx1ELny+MzwXo58KB1JQmoJ1yvV1dwM8ABSIgMbWCJIqgDAc7o98w33lPys
BkBWl3UNAX0gzcKLEhBt+rAW0tzSTw4rGgykMEU7RVQQuyYoitGuuVICHJD5fxtaVM4IGCeP/LMd
jofeX/5PuJXTsZM5jLtJmUkUfyBj1MvvaFiDGcLtqrfdSWdBv/Fgq2NvSH3SwwJgdiscpN3Gnzo8
F7hNHwDCV00SP9PjyCgDAowYQ3J/ZPZUqRUyn24/aF2wCxgQsB1Y4Sij0+xTrkMdlMcAkabQbxmy
UpgeUq5BX6QhOYzNONQDejpVRHFHYQT0vm1iJe4VEpkte0RMxPJ+NUNrgmjE8hPj1FVifqyXL1xA
xj86j2qibj79ZfDv+Zb6MtYHHGTsdkEmQxsKYxtR8jtn1OFlU2+KMHiXFqHqg/M7TrVTVuUeGMZg
gMYEswxEjFGqfpnicYFQysuCLslyQc1v8zwFEv2jNePLNzkJoJSWXCjq+YSC0+JiXPD419WeLbR0
YaayXSxTw09sks2Zc0gEJ47l4LBxgP+YKcF7ydhlQut7gKTeMZR2SlhbJad0RYbwXhzYJs2zlWUU
5aZDRao4ReqbxozfpS/P0jw7Wa3AFC+Dv7DlSqjEw3v5XE7EioneTR4DdD3tQmCshrpcgEvzQeR4
TiuKmhDy2Ig4mt4gipRC1g9X23cf9uLz3xLCZWuYgtdHW1F7n9enZHW0LTJZZ/iW8O0WWLYpA/NL
RrK6JXTyX0+5KwbqBjwzWKeThivhkThmVtiPDJFrZFXrnYrdtBKohG07DLEgZE8Qmn4T52s1qfpx
nBT6PAXoKVqv0zfgBHVqq/h+Ws2SZkfx5UykGiSlU81FpFF2DDyoEg/a5Y0EXJnIQ/9paCzmVlX7
iraXS5n9vlyqhBzl8QxNXN30vkedy6+Dd43jKKcihDs2/SS979aQYnwPpIiSAQkJ7o2PXV2ZBVAG
9bDnByz7sHVCrnBbvvp5lnOH9YRKsrfUAJRGx3dPvU7uhbbNRQg8u6OzQzTy5GH43rVLytWZ/JiP
TeWPtNO0gFyWGZV74HKt1mOhD7GbMCiluwfNAqBLFMSukqHUcnaKSwrKak8LgssjYdKcJ4OowAew
0foaTtfL2lEQNw+Wjb8XQec5mYRQ1uXVfIhTOrFBz5nmaQQieFU9YjJ/YiAu3H+u3gPa9L6pTBSq
9quLF12zYD0Ko6x18t3rJdmiJIPBs2TpM+0Br2ydLY8XmL63nQALQxxiFVEEVkrpaKF83iRwcUYs
p66TzplAJxVRsQe72sPwJJ6Ok79qyZH/VO4IMgTypzZTuDISnFg2vtoZNPUtPMD8FqEplTzIO8po
IvuitMuDWIQC087woU5XrDGdCdrFhWt5DWWL9yNsq4Hp0Bl7nxuVA5xIPc2PLoUSLQU3QxkTsTvB
743ZOs3MSM3TIxKHj5c0yfNKyCLGNxbiHAQS4RFi2UJJIolA5Q16T3FDFQDXLXZ4SG5JXYNOaRrg
BmEOiilkILMXwACq2O4x8qaoJYzguOCGBy2RDc7VH9rYJIlihvMgZAQT2MlWdI1wOvEfy5Hp/dzs
25Lko+HBN2yki9m0EjwtcTGP4GEAki7bEvcNAtE0u9jnRsEYomfRLTTqwZ6u/CZp7Eu7bVAEEqzI
cyEgNDSr6/CAtlj5tIDCQQnuN0NwYoTsNrmtdC26JK7X1wdQEHDUysWT4Mt3iE5Ue4fIYTzqH/2E
IQWViGqo3Pj1EH47CKG4AlFxHIk4d6g3doRHOARlhZyRQzikDXUYnmFA4XPZngVV5KW2Abnc1Cow
fz3t4SUWVqnL4r0aljIFXTrQ6Ml6T24AQU7QpQkaTawS8BKEY3IFygOyJJCGM3Jg8jvz069JhcNt
9OTzpCzgU3jOsgc5huCG6SnnyISL+lANBpGtdLN9Gycjg5pdbH4vXloSx2+nSuFEiKVckFsGV13e
wwqOMeraJrMprdPcvmK9DAtMVXielnXdRNYT5kSj3aBSJ4qocczPAvcWE0VZyFHMTfvgpIyVo5uL
5oHM+kRh3Rdj104TnicPq4dZW3tCStxop2bxltVZ+ev7Bfx1lT4tMAqg/X17poXeG1RxaSJRj9YJ
tqwSS71EQxWilXpJoTWtMgQKw1DRZMoQS4PucVUN5yOQ5KQLYICUk0ep2XzyKmWT7wjuriJWZYhV
ffYd/pabXpEjF35oOyV3+Q/onTg6pDl7+VK2zKZu64uoqy3SK7WDBu8kkfxlh9QAtEZ3RsqlYNRV
J84gAIQocCFDo4nasL5abEEZfEqCzoftb91ljhedMk+E2Srd8+BiZ+Hu8Gqt/KfBPW6Hoj4kgQ1d
5QpXNmkiH48kYj/8/e5V+G01UCmIm3g2ZKmgrSmUauwW2Gq4recv5avUYHk5fExSwpU6YLk61qdP
1wWBF27+i7wYGJQMZcMQXCbrwzi0i6gvq01U5nxNdjd7OpG3OwlWpLDXY8YkM0b6Z+Maj8ecShEZ
ixlZ0ydoVBob4BjKUK8pEPOBKOqW076Q6uvyGOTvYMVGBHpiR/X0UQrAt7ckSEk4xUHNb+kH/mDZ
w1NtQiIsKZPGBcSZ+LhHtBf+CelFpNZF/fw1QjrfmqZzXoSQN9GAOsQyXlm/cpAd/Ej7Tjvjnr4F
JhTYm+jXBL3MWWD8r/s88XRhXokrqMaON9S0t6o71ktmMi107EFDV14oBp44S4AAvTv0xglDlZ7D
XUYydp3QeYBPdSjIeCmTqavsPwMkC7Vy39ih0nmlQUr9Py+NOgVBQRHc3JCnJTp+jNBqH9XTmvHw
7i3d7yJ2KYTkeFcxKZvMVSTBU3MNoBI+kkHsm3ndOza26l5LrVDlPs4BHw7/dFdjrt+nMH0bJhox
L4wzB4NSh/AqzV3Q/diuYpZ0K1ZEGuqVYT/lNWPRjkQ8pmxbVzWt/vlfF6uRi4G03aW8SBNEkQ+t
YO/nVPhX38bxCCMoRjI8zThyhX54EO2iYIMu67pPRUrFVKdXY5eAuneZA6wLlKv3794IPFOwzgGF
OqIYS0lHiw2v+Vxy23KPLyep6yMUu9EhLPpVVNipLA3ieGENaHoQMzuu1cqRy+BxhPLS0dLJEnKS
OIo7+QZ4VJh+nj7Dx/lJYPz8hrHsPd7dfr7j8t1PLjnDzUt/sPdrUWgNwTXMpSiA1Hv8bb9ZBNib
4miB7Mwx3yun2DhjGMo5L4FqDOMmpd7EKj82kBHh32Rj6RAwmSvu5VlSrsW+O/yZSRSrzl1jgzRC
I33Yy0U2RyqN0Ly0mSKn5PAI9MVinEHOvdP4TSWe2plSVRAyly6NlsMg+sv3q1fqNcJXx6S7hxPZ
krXgr0HoZ2M0/TDq7AinYpF0PwjQqKztRLMod2ogx9ONt48Y7rYZg/nohrTGnoIDkjTffxwriAs/
PiAGrnL91fzKmmtu5sz9TyLcfbBdTOPRlvO6IgDy2ql1q/lQ+aVeQRx77FWU58ZdVjQyeXAxLTP6
b6dP43cX5C4h94oVk9jo8sqWpoN+r+0HQCkjoiSuS6cscj3PWLvyNak2YLhH00FSxiXhhDSWb6b6
ZGs8bsO4O0hvGkaIkbFH/6z4jZ/ZxtQM2cQkqleOKliWG/y11964eQWcYmoCJRO3rArmYoMjlu7R
pPANTNDfJuDDDhm0pu+tWB01Ki+3iwH3LjHHWdDwsBNh8Y+e0U5stxsMNkeFYpz95vQMOOZ6SlmF
zL/AFu54CeJFEf9gqzd57Ke/SHfF2Jd88IyuZvAefLiAvSE+g+lSNoAuV6gDb1vypmMZ1Mo88qr3
HxqUU+ZooJY9ELEwmBFiC8VUWnLBa21i/455uw80Q504+iEi+hBW+kUv49nRdfe2eA0Eg5cU4ZyI
8Dsxt5yKH9Pz/1zaDmLsGV0KPdd/gGkYSycdK7wybuirImcTYkDlAQd9/hUxoieWocGuypgExbMA
Lx8mstSIu4b7quS48O52u1tI+bPdz/D+LtzKWtyNwNv3M0ih2xiTW57sA00PZTtEH6skAxLmhz+M
B4TaCF35Pnh+AxxLj4zpF/jWkkA9meJVBWdMhzsCC6wiqD3afaSV1DuSXY8zErPOavELEu8PLLTD
2gGqr/Bv43sn5PLivnEKfZwEeSLY3lYLs4VaWk0wb3pc4kOmbu2aG396bTTNJUEb2lIVAG5rVWUj
f+C5ezYCHzoNwT8m0BKQHg6KIjt1sA76K2ZBhLNXNBq5gWRPUZAYlVtbp9NGbNE2tBVEN7cPeXF4
24nr4npVLfqi8s3RPbkS+EFjYwtclmRNR2NkmGRZZnvgpZaMo2TVBe1IzmjxNqJtLlWU3lhmX6Vm
mUEnDmTRZVJmKPYDH10nv6cvIMWwNqM62jponCK6iagf6tcIKX+zF/1979OruX8LNbw3/ZCtXzy6
cg4v1EpZ/MfmvqnvjubTgsS79CX+OMzbjhv41NlkQmonSdSRUvTuMxZccCpaxXJyBn1Lo9WOAyVY
1KY9ac6LEoFRCeEgFRfL1ojH95Bn2zz74VzzzgduGmqwt1iX3XXY+H9Jrbs/1g46TKaXVFRX62gc
Wh9W6lHZeH2Y0UwUc0qhNapBkvZ++Out7TL7PpViwAv8SqXW1NPCxdI83q4CNpluaxKMLJGAtg6J
+2HAp8jj1+q9FAk1lwbvjem2tmfJA8XD8tIIOzIGVaknLueHxtOXvYwFn971O5Sa18CjZrG8IsJL
+oYfQQ3F9v+fJ5K3TmYDliX7VHbknvqj+BM7BPhO6+8jT5wc/Kq2+FCfLSNQA9HloOeOwOd/Tfv0
aU3BfEcGRIf/0KhHEpcdL4ZT69xkQXszmKOhqZ6PsFBM+VJB0nf1QE4ECJLMw2rWGZgIG/OXFquN
bxavK0d9AbN+AubsUq3zcc/fpm7/pdyKfjTsnKRHqPwLgGhqLNZLbSxj+Nm7wv6/DpccTDm6WPgF
qtGtuFYjWrDviquNovX/r+uwN3+92aYInzMeI3afma5eL3+9Exl4Y/7Wzo2vevNhymWclTUDXRf2
VWG3QlDaPPT6l5Vaq8Xq6PZ/lV49PfFvbKf5OVTYNwRpKnKDhdeQHFIyTQNuSMxnSNHkKE8fEVhg
iuWsPC0WBRCL7yQA6TblB2JpXMwhaOYqZ4s9T3cGsY0ADERT7dks61aYX3rcWLJ6Ve4EcBplBOHD
P5j2daIYq0samm8Vd4MC5Mks4r/15MthJdSfwzW/W6K+zx2lv6K2LuNSTCicLJssePzC570XfUaW
qdfORWOPpydFene7LKG0R7LO31Bb2kmGFMNofQ19gp5XeMkW/6Cpm1FVcSqHhCVf2mWySWPM2PEZ
CViw8vJuTmH2l+/q/gebhkriVeOzfa6yWryu6EtKJSmD21ht+rT1w1TLGpgQu6YpoOFayYCLsM+Z
Z3DNRmy2lIsu8ok66+IocVpTcm0S5GK6RTziMfbbjCaXm8In9cmOGb4IciEJR2t6VO6hHowp4Ep8
AfI/jARSOblcl7gNT7PaR+Y8nB6/72tkykBmTgbtif2mQP6b600orIgVggYkkdCKHOgEje/fa65C
b0ejdR/AzQpeTAUNq1Y60Hrw8eXrKcJf5XHQVTE5gNXwhjtU9XmSJE7FLBp7kriDoAMdlO3Y0yKX
6F02eRFJLPbxlu39r0I3XtKRxz3sdD0aKS1/LK7F/BsT6LviT40OtBBRQu/hmZopk0M/deSMLt5y
FJCefbsQ2iKDjG5c7mSf0qOhJGkJZAanqzHzrK2zoYtUt7jHXXcUjPcUbhBOkpmoFCyCWecsQRaz
Q46RlDJ3kRkofLAGL2TlMMps6CCF5oEysNRnL/a3+dr9Tl6tK0xTQLLG0U0/MBolcr0nk768ZYBO
KAXzSdxuCaAEJBJ+sRNnAjLoDPN3w04MhEF3DWUiAWtJrjQfmQo3jd+0+42lHq7Gkopi2+jCykiu
vM7i/AgRvsdQ/fPyitQ46+ev1sR+1MRW3SVERhHWB2gIBKWvZR0BYHRFz8gE+K8zlnf7ckU3r1Ok
uPG7pdzXV+Tx9M9S0WxdXygmcxDK8riqHMAhpXPKIcGKtyxQ/Vj/rac+b/g3UjIydO1KrlsY25Nw
d2N6Hbx2BYLaU94wyCe1XrPxlyMrROpEGxw6sDER4ol3S66FPPWhtag3BmJhIl7rxLP+w5pI0RVi
1oReLeMlZLDUafqnniUWr+Kh/5Y+NEoMgh+mEGGyL/fffAUEVEcheUx79yUfhGUq5pn5EtOsk2ym
nT3sjb70DM68nuutSLFg0wrCQeIXhkYD814cgiAOKMI6fNF1oQrUgdUsIfcX193agh6kSGp4t2Zu
LR/6/+IGAA07/oOUkNS06rCvrGSBWeCz3faucjRyA4x/2ZIFZnBkZMQiCC9t96pvG8/p9lcG0ysR
1rqtyXKhfo1H236LvuzRn1z3EJdvGmW54jSOzQzcrz8soOI7O1/FnVXNcgiUrSlmUbTH7niR1z3x
vzlImaTW9/RHatYNb/Tc2Lx0XyUoQrzl2Ctwy0NDYSZOxz++TODjLhvltMrrzWme6Gk3SLfEoUOt
ROAT1QvIslt6/MTFuvOa2Nh17Xc9dBeOPIp9kQ0lsaXhd7d5q2FEVa59asdBev8xCK2geDZeiPvt
hQ9FahkFMpGWFVPGHCpLoKuPLxS7uZQjKAa0Oe7BaUkJzL4kNu62TuNgRu1c5iSf9141o2YpOzWx
2HcMSkkq13RKYc2NnXzHAXhm3EHHkMuLD5Ri6JRL00fvaCX/vRHjxfNgJw8kXvlbUAUSEWcEPaOX
qIFnW1mfhPhZIPs4i6q+inku03oTumqPKcb5eGUGtcoUI4sv6qCC+WEf5hVIhHFWkxdYvtoy3uLW
ehIhVWf3NXDptaWcwvsLSm6gvgqnfa/BAJqKw8+DJcOQWoCSDFxnJJiEda0Fwp5HdQnWqJQOZUKJ
GKa14gFz+WxZTPvYBIogZ9p+EdhParuj6A9mDFQ4pbP5bdkz3+wpqr4jFdpPgup31es0HiIIUBNJ
4j5K9LLsetLF43ZAzK83sAPWpK3XaZsn4CEAhqHcfg0owWFpr5pnbECWbjXDBCEmHscuj22JP4b+
3DzCm/we9zpIGz92eDHC3PxBznvpetm8mqiz8YtXaiDvplFM4yAQ7C0/862aZrbOQ1R0fsREbFJl
NyUgQOtEfW+XaRjISmYYTd8jFxyeJmFUt+WoMMtEK1jjDKWziPAImSeioDQ8587ofwmUxYnF9taW
N5i100gNEX4LkHK2h83DrCKZ0xQ0kI+H9O5R5P47Kv9PP7VOCfMRATrwqAwXN9hIpwEt2CnZbMDb
4mMZHXulyKPoeGmUtc4I47TmHKFAqbuk24TeGjAZm1upk5CNq7ELO1s2pKq9kgToMO8JOWZj0rrf
dPMptHr5oDNhayBeJP7XtYbEk99BJ+ym0Ltmxjcj+Fio8DdnZT8OvNQICuZEt5lZWorLN2xmiNsK
0erJumxfQtzbmgvDAKSzdO/BA2WFmaYdilrCrDVMB/WS5lvrv93zVVxuH92Lk2uKJ2TZl3blUhDM
9oOioIFW9r+kZfk5utfDBZpkZzhSjIC1K0J7uQcjvv5ZyFUJc+BEMnX8gtZtYiOlhFSJhiUVt1GW
Q6hnzlmMw5JqJ27Dv+eCDvocSqKz9EAlyUjPQIGyla05WAjbwi2O+OEYC84Ju6FSbqaB9KvncMc+
jFxcYAfVTtD+ooOPJOfLU4R/zMOFzsQO69EPJOlQczT+IRsQknfH+4SUv9Q8SqKrkQQUjkli3yI8
gtUXJatov89I/R7ENbzfXVV9GyX5DCd4EGYcEC3oJ1oeDdkxPy4gfk93OYP5te1pXsUDTIxlVRCr
I3w+z1fND16cFg6EGA2XIbN89gcEQB/ssOk2s/D97Zn1kEeiV3ajSQJ9arlSyWsWJTBp+Zwk6R02
qK+xtLM9xsAySO49HLADYK7ZLLcW20iVznLPw2Sf7bSXcHqpw2ZuvEG00nm//+hvkxvOJ1oBa9Uw
F8hD+HC1pRBMxgFK3vXf4nF5XXZO4z0ZvFakRC10VvqtXHOH9rRSHIHLTwvX1RhafV7cHHQYkw3k
EMcx6oMdgTXL5EQQ97zQXtuCD3Ev2YZQCDgAq7pD5y7KWcWJpz8EErWvUTgpZx+Mh46ytUumUHi9
iAzRFqTey5Mg2SoE8cSkdMWXCswOO6Cgm8ATQPhoGKQ/5FNXuXvssdSDDoLvvXhoDZyN7Uk5ZLJ1
Xp2f7+1VCpUGyjMPBwhUNDBgCBcEl1jClGVjycWqU0DIOUIiwRtFbElquSbQowske1z+h89HVQwq
Mvp28ubluA2RTPltF5XMpjqs8dFmo7ywhMb+cXTtsPW3qKJ+9Zmgd3PD2oNdTP7RLlHpdB0fsHwg
rQI5yWed2MxEFjSl9GopH9utiTsAu5/liz6EFDmnsbAkEvGAIbIBF9++yTDn2RqnlmTveFbjOFPJ
HF9ArJX5uid9dxeIvzqPC3Ku0s6fvRVhOzK/3T5EFSjtAQtNOF2vhpnw2JdpJTkSbYv5SaRkX45H
So+ZS1xeR4i/PjTsF4afivnZD4MLNT44yiH3j3roT4UJBMG3HmcQoym3xPv56hBhnojfcwLwoqGE
KgjUO1jhi1Sv96jtcLUC3Sp7o4WOZW8Bo6FPGnzLam5b2kDMxp5KPVKi9e6v5Ow6TemBBv+p2Ou1
qooP8zcyGFIrNApVKpGqtnyMa8Z7FrovE3/jY9SIxThWfvYQVPSsNwJRXVfcUjRfnVktGvlXjtL/
+vJO6ZB3jO1RxWiLRJlnd+K7707G6ENDeoFgvrNP+Bi3c3wcPFOSIodiZNJlIB4791sGlS5L561L
njtQBJIB1vgWTtBxBdN0IM7d8QA6Fx2uRr8uVji0HChJu+Y5pbrU5Tu/1Fy906DAEQogZcfWkQSJ
zM/zjg1zOFHr76MEFt+jMiU1AhOunFT1FHLCuSTCkC5ZVd8vebcBRUd1e/qky7dE9UPBTswZ/VPu
/7ZdaZWyYuNpQW8TlwqFsaROPTCQio2ONSHhwz9XB46ktDpgMNZc1LIrGKTEJRTUQn0giYeoGU9g
KWMbkYTIwJExJL4CIq5lyjfqlcHCNZboApSvBDULZ0581XpIxTzGQwY+CdKERfPysnaXgMWwUH1x
/deGoaDmOnET0O83ejdHySTAiVXUlMb7FwPgaNF3qV2GOV5hL0ZhcRfnJS2cTJ4yZ2wY4OH/QVkd
kIF1vajySaClR+foe9VWH2T9LtAYNG23bOUtgQIGRsnV7pPbpiO605WK8wdWDpQk1MSN2qIrKz4l
eh+OeSEdaZya2fW4aoyhhLOw6A1A+fqWv7ubsgNf6A77RX+wrSBH2GOPPsv0c1GTna51a2ykMH4H
6miHW8xMJsd3mCnYFGibAlwSDk7bsaoU8C7HFEk7q5nBHdiIPvRgz8kdon4rlDAxbqUWMVMnXzFA
PX7A1rAa3Gsk4U8+ddKr2wZD7cuqVKKNAhu7K+mA7RcYKn2xAjUt10/IA9Qt9yJWdV76LTDbnP1D
ADgRCASLN9RtEUjauqTQecoO1MKFQRVY1NHqvBSaAycSPT3Dia/pjZg2LW3gw40dB/MRsbk6jwVH
G9mTSx2lVob9X1NB9XNhI+8LeOkooYwlX+vSoiXEEpuKehcJhUd0XzjbQQQL5zHSVsjzpWqP03/y
wqGFri/oFyELl83Dtkd9zNuMzP8HXHGRLUIiRO4JqWKQabrZpJ5H3Vmfx2hnzjYNPf2bgv5j8V+a
7W1PWcMd4IVcnJXti/srVS6YQZEl75U7NTuVqiSYxuHWdkkH7ilFS0+UuwndfpWfU1SLbVgDTlSd
3eC+PYXojJb1oYmF5b7d3OXkxCW2+YW/B00r7jzCtOQGZ7xO3qvQAdC0yr/eW1CzYjSdanBq11Pd
CwfkgjPZhZQC181BJeSeQH7Ly6wbRHshjUOsklfgVfACLVXWuIr/s6G+Ws1fYGdUXAOA06e0hL2i
MVV2TpS0+wPxhTB63ErCipbyudk20xl+QoAZdaAax/SNlrIx1eVv9/4FfZeV7CkGmf0nSg8fwSEH
mlT8mt4e6iw62J0D0ysjRY+XSm5HL+moRIbeeYaz3E/M4h/SRMhS2AnH48kC551WmFKAw1AIJmdo
aaskndKoJyqFFv4bWIx/WPvzIatgMO4lGTB00FWFLg1/78CW7V5anr20jXgyh0XPZLsi51KEbI3G
Ij9GAdCi73uYZUi2WCOv7tw9y0XQPRBPKqx7/kSFc1oi9MqhJtj54cqFqJvK0B0WurXzhfSfhC5q
ixTg2yYcMja50YEwNqCzfCCpmJqhtPA0Gatt+0K96LdXi84Le+vQVUmo1pj7a0SwufXGYHmkJkLT
Svywe66epDM8MdUjG9KCCUeonOTzOqMgLcWaNP50HQgsCrXuv/BH+Eis0GqyXQNzLpwFluhOPpGo
rwL87cz3j4yxmh+cQXsEhL2b/3UlwM/K7TpzOQkwQMgz8XIHXWbf3Y/uBu/zsr8ys/Ym5TfcXNAW
wWLGUpJMTBfZpCcyxat3XdlQFTu/+SiXGETaIiL3R1iOndkN1gz6LXMECE1FVNQV0CitRlMfBDMX
JsV/mnuLIoyyUCJPEJ2/HBSPgnYIFrV++a4hWq5DoPfwL0uXVMc2Qc3RaijpMIMza5GZ6miNrh91
P2WHgc4c4ly2VmFx1tgWH8edxg3AYXU11pospw1a8N1u5smy/a+37KaxSAIggydhK0XJnUvje27r
plQTa96LGvwsH2iy6cel4jAjST26k5HzkemUklOEg2h22TYV/TX8xzm78Gc05sm04c8wzSI1dvFX
8/NlzUdOko+Ln1HCJd8lN/fXM57/9doN5+RHpT5zjMObqFGs3p88iLF9yw22g28ns7KA/IdJ+xo4
73H9Q6fzmywzBtMDXLHO5R5aAd7jyEyh1kaa7uVBOhlSDaoj7EvOExkC5Hyijzto+GmYRJUjiStQ
oH8w+0RniSW2G1dRrsIGOwiKrA+kL27k27ZnYcPu71thIXwHmzXPoRBeHSuNyJS5+7APo21EMOUy
mATv9BdxNc4XP0ViOpTqWFwpphahOzKgFW2OEwQzvoIngp/S1SQTb+4O5N24ca5IqgTx94Ib8xlS
ygBz7PTtMAldGjG7d1y7REZPmtFCkxFL4iciV/quqVAwJmqAaQa0EtlVnUd1ifuC0g8rL1PJUk5V
563WJxEUM4cpDJtB84CRaGaZMNPve+SpPhpd4UeSFvj7B7qCphcrKLhZs9MVAQXZKfqwMQ8XekO5
nLxE6BPtu82fwnXJa4LSOR2D70u2U6EzAtl2Nso7jbK8qYw/KCLYGJuNDcD01kDuu+qp+XuNWLOP
JihxmJxgPyaEyrRZjJ6uaKBSwmPpm2H20XxDy6sq4wSzmblmTO0L47AqBpkHcm7G0BfG7uTadZxE
p+Vjt1Ap1b7FI5SfK3wVF1JnLzMU0Ky586ngABg7ZmLMQ++VRHqXtWJIO/1O6kKEKW5WoItyTAME
m84TpTjfVWKvbfCir9l1Q6bHhIl0o4uRU+eWR4wfYjnTFZFFvDJQ2Ojjgq8bmCRDRLJvdrgQouxF
BaA018icDNEFdYfRlXHXKBCY2UG9FF7vxljFa/8UlsM1rrjQmTbTPYYkgB1X6EZtxCGsVc+vcjta
JifLwoEsi0vR6zasgIYiDNkPsA9tV9oH9kfMcfHMurIVxU3L0uV2jLfu7ai+ldmSnl5t5u6MVy2N
jkGbxFEKqAnnOciaIkbRtsAGB8/I2VtygoUN1rT2+pUGosONC3E4CSRsi6/KuGUQjXQFXdtD05Wt
Wwub2z3R+MolY+cnWQBxG8l9q6HtktX7CLt7vm0GoXf6iUKVLjB+B2ArCRl0/k+ybFDhMaRcRy1Y
jaWvIh3sclAM7SZ58fd8EUGaHPWADHq0CvPE4qKmBPp/3s9O5kYYqlYNe7s7UK1Lhv3PYu/DktH9
RRr1ONiEsko8aHLOYEH66MdWBr0qODaeYPDrJ68D9I5/8jhgboKW85Pxaph3chxjN7LEqXy5v3cg
aGeABk9R8aQGFuXMAIzABj7x9lcun7HxfPEAU6x6HqDfBRSa4WBPpuscJlpYyFanSQ3XSTf+CtCo
7V4FcXPs1Hb9Ur4CUhA7ccCjyuroIS6UiSoKmpvcOBqdXhg1vooiURfkgf7MBwIzS9RKZPiBEqTe
dL+EiZwAG5WiJn4Au8Lr+s8dvSad+7FMSd4XyXnLzenfY4w+n2l69iBN4dDB2sGWcfOCs/axXaK4
1IhPoHHu/AzvVtFpsewH+RCKdvF/a+CiBaYLE8Jn/Wb/z0n7ZM5ZAmDSKf8xyOLYZ0RHAx4cCAL0
votiZWBu0+G3tWsxUEAq6RfLyHJeyuPuo7VVAiHDpcH7OBb1B6ky48yONSfRf45er2Yo1S9SRl4/
lC5TLTqX+X533HrPWFk71XEod8HS40DIXr2v+3PJcW3L7aRaR/q3jkRAvNm7mO/2kGyfOTvjTW2a
RqM85EIbvbURqU91RLzBskVSN+5U7XSlFVf0pCFdHptaHbJBI+WVwlapof5X4V0cp+lvU+8zhi+Z
QvZnEs4Z4vtdLlGNGwiT59ybJ6QmCaQ4DScbVDlWEDJRgKA7dyc/PrMKhu/QSUhh8bP51HNMOWUK
BHT7TH8e/BJ3BfJNTdfvCKGlTocIKQHQpKV5cRzudh8OwCbJaJpboVT29FFox6I0ikbAs+lZkX35
xh8MaJcMOKECT9dj66D+fmLioT/US9W0KREtgxd9RgpgRtBV3f9ae2VFqEo3ZCRSb4wv0I5/LRNb
MgNMJouHE8fF7sca9GIQGCHnp6LMr3IPexiNOdG3t9xVYq8WnpvgX+kHNQh4M9Ec0ZM9vya2t0uF
Wo8VX4sF2ixQh8QJSNK6+CsDEo3l6SNZ95KQZd0qFU63AbkQGWdnckMpLBC+2gOYsPieJwgIBQDy
29Bn2hbaKDZBQJyReohqBE2DAx5I51IHd5fApirejVIm5RomGnsNCawyHLnrDtdH0T6NexItA0Cv
hTgAOzNV5hiy8ufkD8y9BavMYuCI35MscX9Ba5POKRuSGdMkqawGh9Ztpd19aak8U3Ms6CwswR8D
mxZAFF+Eqqssdy17Et7OQnzBM8uKmX2G6vsoFfTrm4FXfEFDrx8RlBxTVWLHF1EkElDhHLcmDVsh
t4lTblbeGQq6/SczCqbcy22aUVl6p2/NS/TyIVymhidQNHr5bz2a7auXRaSo+99oQOIxxQClCU6D
P/i9vN+Ezz58loXd+k1q9rQMfV0OQShzaApd8mEUvI7alEeOB/QhPqxpoewk/0YUBimZaVLdIR4Z
PU1tnuiT/QbD5Pnl9yXfiKNdkjk2DPzLorm10ZhHqCtx69QTHP3LEP063j8FUuWuSYCPzZksoBnw
TBvu3RnBKVLh1c+hyztOGhX/OeV1KCGvSeFKL5otbMGwMZPxUOZQkduR08mtcFD+US4DVXF8tZI0
MHyghx9VYSINeq9fi8FYB5/bUFzm+Jv+om/7DAyMGo8Fu7LZCL30EvbEE23G06/y8PU2FnasB2ZF
td9331EInUxoACP4bvDFhpDjbEu3HBChKmMP1oxAMMn1cfWnxjRqOeSMHwK1B6tDD2qYUwnihvsl
O2BouQWAHKSGididYm/CQGtsneMXaopvfck0Afb+lQXPWFVu5/IeJwT7C7T8Bhyc52VjiOPyqwnR
kim3VOSUgQax5lidkRr52s7g18ImeQ7A5mvh0y1umIOsUjtLDeI2klmbbASslhYfiwmYE2IcKcB5
GlRQQbHIsaSYW7hvD41WXjXUerttnl6iepvmKY9iAAJruBwdgN9ViN0fkc1X7+IkmSE7UbXOolCX
nwqfMlkMqH2M3/LvTBg+CVSfmhzLU6dVQKCzWelmgwxce2fyUafCVBf39XF6Id+3txnN/Ikdtbfj
HwKW42yUbRLmiQ6UKcaX8NQtTn8xzFXVjUvm7OGiYPOHpDHml3Arhm2Dxx7D76hJxPttHPBzPk8K
bOPVUDkgo/4RjEt31DE9m8Ri0twSecAxXCDutOh02bQ2LRbPF+O3Q8GKHJqYcvy7Ews1r7svUGJx
ydgSsMYxZLNx0rkxIFk498VCGI2wKeBDrb7+MMz4H+ZeMteyfJUTggDAIolJPWa055Ym0h/x7yT3
3ZLM5Ha7CLllR93fpWFKE5dCSxs8KUhxNjFNC7VEtHa1YJ6Q4736Kbe5vwIv5s5mkVWc1b0uO2sg
qk8IBsSBW5jmd/gXGH6LDpUNPGaUdPjgLuMo4FrSLPPtxwHkK/83eB/63s7TZXUXmg7ZRhmQdbsu
Jy6nTRNLPRgsIdgRr2WeH6028KLvcFvLSOo9TyRZ+JvQWRpk7RjWKNCuFVV2PXeOYyplOT16ibxj
8QTLv+QR83PNKK5qp2/uparAHzpOzAueHh/Eluo3x1qbhHdDMT7HZyuVl5AekErR5JZDpia/qf5L
CuD5yN9Tu7Xtiw60ueWqBiX791MTRwupU9FvKBiZ447nzkSfVLUGMNOVa9gUYQfiRw8QR3leTLU0
O/eidC1o1ZZxaCtl3NOfe2/YgJKM6j/soYUu4+4h2rHigm29saaZ7RZD72urGo4W8QdvOyO2nWeh
jHArfl2XhUHBygxHfkFjlwDyQjWcmlszPeUDZOpPN25lwJnkCC1uygkjuWf13zEliHrtqgv8PGmp
bSWgkW1wU7FRFiI8ySHtE0c8Jgrriui+TGS2zxsXPagbhX1DNTwLO5rXqHfrL+/fgZa7oneAPf6d
bBUBGHfNcQPbNprgSfSJpYCz8xg9BRgjwJsVwwMui0k4Uhl/fZUh3cTDr4lCK/YWlLDkK9RKkqGc
IO2GJjlwBrfJhAcNJP63HmNTogG6+eJdaluMSygoZAZ5sQC3Q/F+5pXGleWV9TqcSiUsuli2iFLc
H2pAEj5iXDdp+yWk94E3rye3qBvHS9dNW7oWwRa3TGzIqu3woTW1JoT+waKJ+sdVSxiFyJLdCISx
XWsD/XmSvZBM36sVtfK3SZkjP/j3rBY2xIHI+95SIobokzDzFm2UyRYL0IMduMghOLchY/ijsSy+
jipgBhG12CcDYJkwilYVgTlEo4qFEeew1CK6YL9hdY96UH7LHLvF5/ggn7LJjgiKe+kmNgC/+vdA
UZYEn/DJknsCSWZUbMfXzNa6y9NBKTYAFWTHHkt3xvsw/VUOmtGiLnNEp3RXhI95Crn6NWL2QO7R
j6r/wU6Guf4CILq3oRk5sOw0uez8mms3FHQZG67M/HMJj+HN9ZeK6tV4xdcPAz1lOhu7RRBuAN6B
Q4SnQ8RKa1OkqSmh28lJslE172MrtJ37lNfTkmIRIgUQr+OKWEJjzaAhQ04+l3UfB3tZNzZBJjyD
EolmC0cDHIL4/3JADmk9VnGRmjBDZ9Jpa1gRuK7q05M0B/i71EIjNYTyX40hDaJ70rCp93XOBs0Z
0RxKYTKD0DUmnBqag1lAjDRpGke4zbMT5+Nepl9fH7BWj7ihmtBy3+rmTXqwbKRbO5pqN2KTfKM5
4RvSP+Zt6UbyltEYs2R5xVmfH1tGwW6zOHPPMearXQR6pMFr/QtXQhUAmdMPoieaNc5cMt+zPEIe
NRA5tuNSy87VsJsGGFtBn7iUYQc+9BdkjhVEObw278C1XPoE/DJ88tJW//i8tUaBoItrf20Sr/mo
loRyH0KrNJ5Wg79scWQFJ0wKIjZKWRqdsScgsoqPoXhtBeYJ9DpDfbq9jKKxqqjRIVi5dZlHC7DF
0FTD1D1fMuOebaYxM+OpBVpf1qCZH1i6kFbyg1bLYQQc1BTuK7vmRJcZd42Rj+sTma1Y4k2XjJo+
BHuFlcw8ro8YscG0jOW1SRVdOqA5SXwnEHocrluRjm19bOJ3qIL3Ck/T37202aMIH4cQkFlQ0SbC
g5qDiJBl0YT1hQsS96RUJqWw0fqv9KBZ+AMU9cb3Ff6MdcYV7n9wFEl005jS+aq1XkKm3VmfLuuw
6gBmC4K6I4oyFjwcOkK1P+G6XxdGR47HEmyVvFBM2G/50HN+qRYqD93ZH5m/1cb/AcPNUdYuFciJ
uHp3puZ44TD4P57KEbPfIEfQXFVcHqn7EId8dvWnBui7UcMVRs8nshcsTdUkgqD/Qz+/09SaVUrr
9f6sxAe6h0N/MOMlPrgXeeuRlvBHZXCp0F5CGc8bxu7N+yM3h8UlrppxHd/+uJ/YitAtdiwmvSIB
Zp0tJMfEzn2+k+6BNx5/NBbR4C5rB1NDX1ox+D4zfgCF3gw/kIFQgewk0VgpFfDxbB90+eJk+cbM
1OZL+QGD5cC7RbNZEZz3Ro9Uc1/VlqMs8KtC/O0O/0L6Qsj+DE1FSNDckukmLCn0MyrK1fnbAJWv
Mt9AJ/xN0c17kI3UoZVcmrLzIL+9pf42I6y5zeV3Ti5ehpsuvSAruAWAOqFfcy/6T2f2Iz8LZ9iZ
JhSwVC6ij4LW4efrzK4ZJSYsKP0RappP6CzBRAxVLK7iNnEJmTD81uhDdsKQHmz9RFrzyl+VW7kp
juQI1WchT84CNfucoPCIlv9jRiF7eCLQtR6xgSRxXVqURiDvXIsN8dHYSbhSJrn5qDxSRjllxkwS
1gsNt3CqXQiYcVI3i1TgX9xZYLW5aqVCeWGd5iKdvRDlh7dZJHIuabok+jmE5xpWf0yhlReC3MOY
BsBOwLSnRihuj/oeFMV7qhCAQrzRuWrJO8/cajewDNrk9UOAq+8cV/1IFkgf2F0nKJ8RSr6cu8Dc
pKEVPbtyCTOuEZuG9dv21VIfLmfqGF815X/R/7zEc2onWvsJwBeqBrFIO53lSbfKlUtaShNn7WzX
GXebuyaD4YNmM+/oUAgDRlANuMkHf7ChbG+xuv5hx7Yanz8tdcPd52a8gdsyEqVmmAVMejS963ie
fwBFj3CNrJbUS36IXSrF2psYaSMWAV+27bwz7VJkK9vdDJHzrFgKtaLNWVBUy80yPHHSiQ91dG8/
f7tZSWJsVr0HRlZLMosSbxZiQ33Bj0lTk6ruvoSL0M5kEkAc6f+t01litYMVGsgwVWmXgSdbeL1X
52QPI/AVY8esyaBW3dgJizoywfsLGiIZhGEHn49f5Mzyv5eZ38a9KuHL3aO3k5aMmQAJp+4t3ux1
qaUY0h8dSUSuzYic3CtnA4osr5c5oSh1GwVXQ+NCs0sekLUAFHTIuJbN8h7zSWfUcIFhWyX0LjQR
o1d4WuS2+4yROvnRNqbrWubn2lUKuk2tgPZmacg+oQ5+qDZIk4LjW9PmXWavlaxE6obRY6D7mLJx
VnjPUljYbFiI/DwK9erhcr6wzJZ8k17hpstbxa5x9Nf8nsU2dyAMPSUlClZdvZkJC5IxS40wfqTv
kSfvCmS8F7aPaYI+9ATtdelZEQc0z4b7a9dpd7wQ8pLWQXYYSqUUL5n6waPk5qQYf+JWntPoEstD
oAhKSKmnRmCVlfAyipjqPzXkdjGf9jsUPc0Joknb1VHm2WwXPprwQcDG+R4G3QaawOsS8+rClNoi
RBPqlfecGhBl70GUQ4l5eVXiMJk0WLEGgAhX85pcEqV/bCOUe4veUtGwwnfaQkX9PZjq8plFvv7s
lNTCCXW785zqh/9NekqtHqZj4iouH8aemslp3hu7g5zGW5mXP0RkdDTj/+rLGy/Pt72gVg5SHZPU
SdXY/BXzRNzT1gLqFqkdPCS1UPxkuFtmjx603RawCoy8oRTeMgB9+LE1jY+Gdcv0fuHFH5CPRfUi
frzt7Xl99PrmKH82FgMNE/B1v38fu5k5R/yRT3vqG92Ne4JoDtgzYB9uBceH2GkwppN4kzrTYw/O
/fGoA6+h0/TAu2j3UWEwHYVunEgm5IRPm08CAaUHzaeb71og6m2tTttvE991v4VvRmWCz9Swr1IJ
WRQBSyltcAOWlgVN2xLQ6hmRunGYP0m2eHsgrXcGlVZsgeq+vqDwrOGj9/h6c+D7sfgHGyeGSJ13
ZjnkrIGy/GwGLMQz5x8xHvQy9z7mWlCG7cqaZEVKkEmMOnSAnWHrRNpcxkimeX0uwizzIpfNh/wW
NgQr7eDr13dPRy8Vaav1x+f4xevwsFEKhdE28NT2QFlwzXFooxrOtaivbWenjeC1dhg8dCgU7Opq
KJZuYZp1TlxKb+pZjjg2GbDm5fCExDy1m6mXr+ztQ7BzXTWulnvVesSgEfB4OhRPTGDK6zBb3Abq
OMA35fQTHP96wsiCINM5L0feUN7wOE4KuJ2ZszBr+HGrlcJqKZ7fnFqUrZ2h44TviHzsvptpBXLO
m9IKML0c8l5ZQv5czreCLxlqpqtugr+Tc0EiXk1WKtEGtwk58A65CX0m7K7fhUSGuoL7c1KkSjDv
vPxrE+UrAUHF3Ypoyuf4bshxqi7346Hv9b7u6dOQ4DcGkAo+apIN0YfbSWxHEMS45CMHeRCHL6rL
lqEF9IfICNi0cP4yD44BD23ESIL8KkPOU7gCxYjuewxXRiiQpz6PSk3mLKJ8eL1rBiAJhBSVdZEc
JpzQTn6yYKm9fRDszDVZ5za3X6n08+E4D5uaP9JL3mfsZnzW/jWe3X9cf2Pyj52+ZpbRSTvWp/FO
4fG368DhXWPu3J/SBc3niGjy65JbvV+6k/6t3DpuBO6Lr8G8v7+ps+p1jAdboZuHs9WyGB0E8v8f
og24t4VxmqwlLlSDN213m6hsUmoKa6TKDUc9tb+AzG9p7BDO5axWUE/WgPhNVn5TbaJ67Gui/RDk
sB/WIcLOoHSq+XauN3BywnogfEFHUayJm/tL5XX4I4KZTZc+JaErIH+C+ONOPVbUmimsy7N+UJAB
7EKpwiZLhheo/wC3RO9ps3J2mUBhXnHCm3/MYA/dXEso7Cm353Wp97ZS+6QIfT2dEGxKkTICeGBp
EMkyZvpJVTMCivX+hkWW4kUg0gdqePpoAxj79xKZLB9dpK0nYxnjQtHUSxPwcGESh8gsl71rJSF7
qvOxw6iwhNiE8SYCpfK/gQ9AXdqf8e1q1ApbeD5SHzS0fq0kob7jm9MjX43QzLJUsQ8m/9AsyWDf
4Kk1YABkItRlxrh1I1cyEahQIuSKNnlx0gvyEMLqSQFnRwBoS3QPNWfTPY8ALqyqieZTgAxAY+5g
eTMfDtkg6+GhyA77SvnXZvn67j66l4nc0rQFfIQFqiz/2Bj4ATYw8+C1AibOattRc+xI44pvLXgN
6b5/JhHwa0KVOCJHMO7ZySYu+IvMryWR5Sb5lSEBUhOZJUQANMT/ZeRF6KbyQIAIg7ZnNHoNs1Br
mXnys/2x70RO+dJJI+KqR1DxHqd1q/DaSM+4mMV5iUsqOilQFXFhGzIhBvL4yKX1RpeYjHGLg1UJ
YFlGTqxo7io8cEk1CL5eJQ6l86lv9oVfGAj4Gav+ULGH1VNwQcsgYXzmWBMdq5p5FmgK18XJLvjv
kVDS0J5p7ePLNPCADUr2xJCF5UUVvr5RcoXNazY7q9Nve7LTMNXlOQEYEW2FEmVZVs77dSKROtBT
6VbQeczHz0ekeElE8wdDy4GpL634Vhl8HcgHnEjvMA+OnxXkQiCtXWCeqDoPWIAGHptFyskbYV5Z
yAgEho3s8mkbvtDKmLEx7vb4tNqahS+gH4eekWWs/p0/pO/1rh0iz1B0n8fj3PQP/U6kuBYvmrzX
sqng768gIcdPInzCezzj+2N0oEALxJQruOz3m7NaBi5UD18mkh4A6epvAJT+wTjqq2zOjp6M+DuJ
Ko1VsM87pvFmW3uaGOGOkNAnXPY3KGYp5rf3wUN5xzGlMXUb7zZqDugx676ZyA6v97DkSEi7JsBg
4eirDtuA3Zt0Pq5n5FsTt9+rF5AReuZYji/eKLOJfB1rgIJXL9lcjgPoKoAi9615Ie6H+X1FbNZ8
jdYYr4sdzo73tjPZrSCmVyBoVtamR/3ASri8YIsK0Il8khzezFQR9IikvPhWSoOUuxUhMC0ikQys
ZZn2GZA4vZSzLezRCRBt5vMgTtSYJOouEHRXSrCCQ9NL1NKoNuWYCXTr6tvVxXYcKVWU3NEZdT4s
i7OhKbtCAwF+Lwt0fquEKW9/Ynmoz+bGhPZM7jG/x/aBh8/3mEl75R7/cESPjBTWGs4LEiY2R6iw
yt1etjsvRt69VwngUC3PrQNIULYxGzeczeFQdLyLgIwgOOMT95Ir4aU1ESXKJnhFODMSCL1KGa/b
PBKZc9Bf4arphcAdt7msIS5EHRY82kuGGEdXbvOAc8skjj3gQLVT7lKgaFMe3aSniNXviuNcL13S
H3Yo1r/A9vl6KfPPkOAvMSb8nVjI49Gv2RIYG3jRs1UHIGB/s9JkP4f+SV1okbbVSuFzvwg5AvWM
E+juLA2C7tvYg4NJ0NlbA1VasqmR/NB+eJp6913ajCD3vjbXvfyAN6Mn9LaMKOyMX3qlhEcYGeHg
go8R2KeRxu3Gs3DMwZ2cVM/lYbTUfBFKbZSKRjAlQ8HF83Zq4cFwP/sYAr+5NdTML3FW3QCBjpxj
vXl9G+T8NYL6Zi8e4K2VMbjUaW223wlePVdI1aB7qz9v6ToAaQhD+xYgwdKZJQVlGV494HsY4yw/
uNnB12PHGThtq/Z7XontsS3NBZQASP87LdhAduAcv4JOjsp6kNyN+zprUUVYlQgQM2Nhy/3JQsZB
v2ANTbTsIwFLAqzreRKPrJVTsXmBJy71eDWeuKYhpmw+BgFAayunV7lmkyQo24PQkvNz1BAdOZYQ
e0swH1zGGZmKy00bzRmdL5YDCBBw/3bPTW2EPR6kNx7Tvh1vxZKs7yi1AxJ9zzSbBCxCSEIqyl75
zYN4EUbU1Jp9I0tkpBuTmfDr/R912LGwAE7vgs0aW+dk9bgP7zeihCME/gQqwAQMDys/ySBNsBfg
nResISrujgJ9ahnpnFlm5U9Ekjy9IP8dgfWcVjzFnoGfNercB0T51oxM5YUOv6m5pT9m1cbMKAfh
AAfKqD2ae+iOIHHPAFsI+wWrDZDSVw8DFmtXmcX9PT6g8F/paw/baRAWMsue3lp4R3O+nT1NaLiA
oQFwyjYP5EagtWLUN7tCRcdduUBrgfSomQAWMCs+PNiyhdhGvG13AsaQkwjCOPubBu/DX+rgZvfJ
D7iFcUD50zRJIlTY8e2CrzfhlppmsL6Ocr5BcDlKykgr54VZmWCtaH4qpNb+R4fq5nK7c/vgVr10
h+8agfiQ4CXkkz+KHo5eqPmD2US/tGQWZnCFE1vLql8Qt8vlCltN/owbNkZLjOFHdxhwTcVxGusE
9468a0AkqJYjNmOZEcZObXbFOT2HfFTp1qEMJNT/AlkTjvg+HYwqhfW43gZZEbZW5kc7lWW2/nux
5EXhVIyB01qez1NFHJepicmdHFwMVc3k8Nb4QV2Vn6EyWV3UCgN9J8Ik5KvZOaCRYjvtINIQHLUQ
mlbga1Leo+YtbjoVPGkIjs8HhD2GYKOnUz1jw534csrZJRcSzE5N9c0nJbyR+8EeWXES/bUp+O5C
uHzaA0gSIZv9/YqfzHkv2j7b0CVQMO2r7UtFtLnsU9gMtfiO2zHpFWFcvBwb2XWUGz6tsdF5lzUV
NUqZ70SB7eI4GdxZdJwVoD7DmHhPQtwlQW6tRVC99BbQOsOKzk/Z1Vrapp90kyt5C8cRT6CVYdA2
8kvEEHTclY7foyojX1qxNzsPK2t8mmCdnrtIu9vWftZNtfnvUPLYLq1Fvk+UBBzraFHvpHTc8QyF
hZ/fnlPrmXTXC2XZBavJZGkNEFpEPpq2YbmtrWVhi/oFwT0S+XCT0i/Z7agTALdES23wMhksrz2k
cswaUXN4oGSacf19qv0Ji4N5GTuwi2ulOq6O5svdy0A0TJKao63p5GGMuGBmksGRo13lAundG82r
jXyFZZy25NfBl0LWsQgz3yYzS6ThhA2bGkTzKEv1UQlr++GEG7siry7R9nJEyy7TnXNNJ9R+cVtE
xmvN6EtpIOCmVABeaiOPSKTFJGyHbAQp/gEqplaf2Pqp1/GW+fYwSW8/yH/SKo46xGLfx4JtBI3k
gkHrt2pnqdQPu2s47aiibOo1QE0qQrhPJH8d3LubnJ2qolCCSLJPGaCe8PuLBUiffip+7uu8OHBV
1PjyFsnorWVMJGYaHzp1F6EzUlB8PgP9BvWNnBq7GExIKPOjI3xvuCJE8pgLy8inSTsWqpUv4aEr
IWcq+p+hQmWwyqEHbTy5ZbL9GwHuYPnrdgBNK2ei3lqGCKJgeGgybHZl3+ymH0tdMtzzbuiDvTwi
BITr7KnmxQD8m7dAUFhPfud69ATn6aTEzBN0f+95ldRBuYf18Cq4ek83QVEgoL8VeohcmyUDM1p+
PMoWZxou6cGiZ2ZVX3BNDJeTleeYsLLVIKl91cksX8zRjdkCOh9B1X1qsaS+lX6UsdhNfq2OYyqg
iMqYQoWegz10uJQ3V9uLwHoDOvytLN8DLxwczBHKoI6AMVtG6klCAkap3JOEFSnq/AWLlu2gEKh1
3XweQJiud3e5Ci77kMXwWIbLVj6TXcY8iPCb4ZjjJBvGFURZobifceH4F+L3CSE54HLcBJvxLEHg
2ibEQ8OGSVUpdmFKlVSoqBVVI5K4jCGcD9nQE7w/t0cAsABH++72+q3Kenm4msm3680kI94b0FZk
eC0CPdqrxDnrlvFAz8tFfNWL9CCyjqlPL5Tb0XPKkODItqn6PdldKprA11fkms9kNVF3Lmz+l54b
1hgPmaAe0LknMFf24rNHj16NrfjC5kaJxAlkLRJWR2iISsrJrb6jY3bxeD42/Tm0cgXKAbrYAjP/
5QKn7Fx3CxKr+IKbqnA3D5hu9tzdmfTvqD2LXQw4LYNW968cm57D8LhsaGwJwbC6Bje5HCOrGOtp
MOx0OcoDhYLPXorzoNlzvddex5ivthBDdnHQoHDW6hWwsMRVUp9Y4+Mu5/ZRL8wLk8vxR+lfZOAS
LpxoCQkp5pqdg00gb64rjKxfN+h8ST8Tg/I9ahV1HFROaORHNh6AIpqLfHeaGKgW/rmfYAjoawaW
AGqmmZDILD9i5Lj02UCZOF11zYdV5uhewIKKnJYBooiOnp/pQuJZ6IJna3EhEnmcnHLRR56vZhwY
n38FeIC+dZRYY/WV4kFfVEEDvxKHWhbWx+R5ueBDQmF8/5c9MPngoLlgX8bW7f+Gled3ScQp1Jms
ujCBDnVGwKWxsGmx6iB1R9+A4vAjCH6SQy7a4Ml9JWXaSn9bQIAbJbpiKPBTvgb752Wy/WZH0zKJ
ppGpB6dS812uZwC0V5xzaP+Im2D/ff64ENCfe9OJqkqcMGwlWRFvYHCVrBfDeJTc+b/1eu1a5sbW
uie69lxVOWdBRrMRkoOnB8kZvyz1bk/4Vz1vRGgoVL9D/8PYIYI7kk9f4AfuxvB441MOU3xf0Ty/
XKFkd4nJPGEDAUEN9hKxuuv96mLWIdFFO4U30Omsh383rqpacHtNvyqAtHyouYUQfQXVcHM5Jbju
1WoG/dBm14xWQaAWmOosRN7zvkCkHh6ViJ5x+WS3raijERUQT/rzTCNPQPri1pT33UEUxh5BBSvL
pSSxI7co7UR8gY0zQTncGW8PE8SrKjKXzvDSeiPmSJv2CzayNMDv+yFo2LbYVPMYaY0F4yU2bosT
8on4pZECa19a4HKL+ZtuiNR1eald/m5p+w+QKlnqVNZFzbTvpODkFJOeus5tdqy2stei+v+wDeIY
Gu1pxfteN/GuWmiBONoMjD1BrqAKvU6oEITqnv7KKX/PczFQXjnI1da2Dt0KY4cq431uH0QUmNvg
YFoJVniJpmiLjIDFGfEYe7UuaAnYJFlZJqYiqfXGL0Da9QqdtmQWWkPzcQ+ZMsU+EXPliFh4s7sL
WH67xLxD5ihBYWcgcaEO0FMObdl2/rpjQM8GOLqHl+APAlyxkgKpkl9CAi5xclC3jkhoA7v+QsgL
1klv8Aw6z92zNJ3qMqLjFrBkGo1/QkH3YcqbE9IJXGCdZ8THD48jM9fQinQ5ODhMKNpvcLS0eUeA
Ki0uMHS4lbaLw1ucfbBF1jR6OWZnWI/UtfJMv1rOMp2Pc8Se+mqIsPebrpvyqdD71R7boqesbrne
rDbA3cZqG+fMnB/ycSWacp4d9cmQeCRqG+9M5Zi9A6Z5YDILxwAPdv0/+xYcSPTDTp2lFc3+R5RZ
vFzs0VQW/ey+FQeqnFxhP4K92+XJUkNowT4DTvr4vO2w15YDGuV/p8zhqc++9PlHK28vsCoLIjFh
XGs93b6fzkO+8rdV/RYbTWzEJNsMhRazYe7QPKQFiIQL8wFDrxKCSffWpTYVCGxBqxhyS7alwOry
Vqv532gmQ5QT/nZVsXrbi5ToiIP/Ju7vuzkovR7xsEGr0pVLtbipL5zNNllNKyKGhVniYCMV6uvX
OfzapgDqBGx3vJImo6XUGpixleEJ/mOjt3N16d69EohA6yEB4xEI6hsZ9xg40pVOYjPU4hAIMnzO
a7jVx3OC5T5jrVqErwOXp0pzgpxSlTM7n+q9KNhB4aWL1+OJ/XTmZ7BOrN72XuY5+ad43lL0paGc
27rZ1JTB1PlJk6m8+U3L2bRWGF4CljqT+B/WUVVefA8X1dTaesBX7rZmkJMLl2qkEKtKQnWlYdR5
BDwEYadg2FaoRbH3yyAFUzgzPt8we3AIGKOfcybmn0lR4u0dfNLC1KikJxM7l7As/ef6kR3dDzGR
cGNeTtbLx8vGRIdfXdKgks2k5YC6MnD2NqepW+dMHz1zCuN9XoOosU7Q86EBePIhjHSqcJZ5TCr6
auqgN9nRZy12AZYBFPI2BE3qvCsavl2AWXML4UHI0mWVLVvtlObr1M5TZkBoebk/SO26dUA/8fMq
qGlmOxEdU5wvFza8FH3K6h1WuB5cUrm9bJaWQJlo5kJklqSbtU3RdOYj0XcTZzUPAdjMsyDyn7Us
UjDcyIWr+kb7ZSQK60KWrgnVLavfqUWYMVz2AIwOEcEJXRzu8iNDu+dNVck1Sir9r4MBPFffBSEC
dcnyh6wAopv0X2f7ZgNZjwJ2J4iuVvY37Bz3YRHr975n2KW056lwgrH8nPB6cBSTAvK7pjEoORky
+UvsKWJ4hg7IY1wxUB+BuTtoCoYEMhcztst3EeF3juUh4IaFGkKPT/Gqyld4M3+aHjTJ0FcxltWd
Dco1SheVTxDtrbhqUsSt+hMk3oAe/VdYLCOg3htAMjKYcZglKWIV2FTbzE/5Lk3ld2jaDGQEOCF7
vR6I0ePuWq6Y9Rw+zKFlbnBFUxnc4jAwsUbgr7FgOliNlRoIYcMFKYoqTbrbM2NzDsOqd2XpnDQV
Dce6GO4Gzm8RhWHBpmko1LJ4dsJwWaBBFDjQi40D306ciP3JXa4jvbfARlq5XECfq44MXOB539CJ
4NXFcgOU5m0mGTxxPcvXS+K+RxdK/4Jr2Dj0MJM3H5G91Eh5U9NEW35SXuTsPFak0/AJw5mrQbXW
XfxYER7svZz47VDFVaes/u0whIAHlpJ5J2h6ayw4xxo8J+iZkxaZ1iiwfEv1bn2Ti+9K78SrRdVW
UT4NRZJfukL4fLr/YgO8ai7991tmzyazdT/LPWa936v0c37/2hlxQS9FX/OhgRkff4IXJ0pZFJLE
lJKBWgYUaDeVPKjIE7y3XVk/Di95FNJmWQXYTR+wtFG6WOLTXZlaJWUXnZe1RDz07DYkPAx33QzW
YN9wj3l9ZLaK8hYY++kwvxXsQFl0rOMUDZwYzt+qKAu3bJT9KZ6shdsdtjDrIVkoriOeSAy4msuB
3osITIyaB8lLLjWgBsp05MArtOzfbtuSsSBnaPoTd6ES9HOBfF+3KuwGBtx6sxPiY56P2aS9pcOt
ygz0pFUCPetJc0fieXNkUBkYn1/5Uz6/W82dwM0XEK5I1J3RikRoe4Bl8+2AOZFX4Zs4m9ZjKWxQ
ntyWfkSxniRq9/0OBIV9X5uA5uWTzLD9yaHKTLy24H61k4FY8u0QQXOLjMEkd08c/z8mZUnz349s
LwdxPB1tUuEVyfVLK35hZn4jh+kGtpcy30cekTDIrQJh+1IndvDQg7/Mxxq+ma94eZAmTqerVLzF
iSk+dCZDtvCKFYdQzXfiKuokkH5YZ3Qmttb3Xu57fjppUZrPSXwGu/oCzQxuV095uz+egsJvRDUR
K+aBb65hiRe5N86FQ9FyEGmUkKq5VhDWivJRlVzoee90ABaS19fOTJQ3US0TtrzipCy2EHCRH4Qq
CaKaYPUGN8ERzS+quyetVM1lXCMpHDje5E3xQ/yza/Q36jfqxpe42+sBew3S9kKCjsayLqbjJnkC
12izGyxhqZz2F1E887/k/x8ofX3PG/lx3buiu094BlGvzsUnTQ9mW/MhzwCwMfUyDwBT/+b+lWrE
kRuAE0f4ehYBE/rQXkCjgEyfiK07MEv8FEJDrmV+94fE+Hjvw5Xh0mGM6vnrTXFu9TDAcfG7jT3q
egLYoGRHUJIBJGhWdw9Lwv2txEOV/NvyUDqYHhLudR+gtztku2V06m/z+GAtMo8vdY15zSgccNr8
du6PjUpSOC0z3fzgE5CvDA46EySlS0sn3gKWRDkIif32UYu9PTxqf/Z5yQK8JCX0Vw5Z2YGcTdO/
pGxFP7A95ZrW//JND2Fjz69Caf3dLUDVHccJUGHJZckHf1dVq17j6UMdeS0aa4PuFXwxqgrVVfXH
Tzh9mjDRSsjNGMgCy3TawmB7PrAKW4kSc5jgFSaxMshv+Bav5zE0nvpAFoinwYOb133uTX1i5zeN
nI6ew9fp/lsurENyOb/LPWMNt8h86x1qRx68jO3c38POnEVFwY5YTFXxTzPqh64NWGEt0krFiNRB
7J65yrDLySNtiMrRyJyErre8KcUe912J1i1YQI8Mxj3E6lA6JagEq1DM/1fQscmdjco0A4txEZ7g
ZUPbR/lgs0RxJhBMJY4jGB+e1oLDCV4hLqSd+i82EXMmIZ0g4CWspqlnL8bdsnrDh5eR2A9BqjLG
83kWrrZxhu7N1z4C2pUR98OADX75dmTPkt0X8+LZjdzo6suaKxao2wk1S6wK7dlxs9k31TtgUZxO
xU8ZxrLoKy0ltmofeP2Oeu1t7iNSlayQR/8G9fTuW4Xj0OQyDXpBEDkKf+KDDs74YNW2pqylSxBP
dvv5KZbFXd7RQg2OTW+0IKboATkRQp39c8cT4huhhi/UrJxQP509wF0AuBLAqq5HTjrcME1zJzVx
p+6rMeusI7urzOfz2spO4D+BZ1vYmrOsO82jpXbzfBIgeXAZ2QaBW6kb2klOPzjMBJy74XwWadSG
XfR6rxZ9Ofu6Uj/hjl6IxAItDkw1NZjcC6++c5i2PDWOBYSK03r7/PQX//BPY64kid6kU35sKKAy
TTK1MB/gzcRnUUGb1ivzfb9tdOG+KJVD/ekharxEEOKqvCIlnigfqbKcTKobCdGtc4n98ozTmlpe
xhZglqJPEeTVEkw7Wn6HTJdon3K5OY7KAdhuZx5832xk3GRuacVpyzDbxEm8UZIGjSDd0eRlp0Rm
h40455khKMHLSex/fgZ1C/i2tM1Ui+K2vkWkc+EWUeJG7r5OWAWqdB2NBnp8h3cOP5om9xG/GpEr
s9KETcvcaSv4NKF/kmIAlhsTowiWH1sV/X2v95DLp2CSG1o49LFNDgQt0rfNR8t/AOY2JYj0l1O3
/QTDUfNcYMWCe06aLwml14t6gKFFJm194asqyZvbDhPtWHZaIaoAt1vrqgAI0zELHpD/EVEG+WFp
lrtGjXizFHgS5pTUcQeJyWKk5QPeYDckL+kfvBllKUP/R9crTNNazwq25n7nB9ZC4PIPVNER1w05
hxnQthnV7peVycEAlo3a9dPSUDIU+vKAw5vbqco4LSUVRPp23KNUG26+hCaUNPv95rslIcFOod9C
SBrpbUyvtkxfp14mWdVLNQ8HZ5zcP6kXl3JZ2kRGLJykqkKERoN4jrr5UqVQcYc5KqSaKi9bezkC
jumInZ8Ssb9TE38rUyRX1OHR92XuUJSeau6+U6FFxlF4fRB0qhHZLvAVgFrqEcQUuUYvnf/KoEQ0
tPPZvA4EE2SIxWnn3fwUrI3KQdV0jOLGiRrI6AbTTiMEA/FqHzPL0K+/Emsags1MWg14/wJoiy9+
T74uJ6KULAVHRfuavxXkePmk42DT2qdTrpiv49/SEk3WhPH7c6+/+/CIJG53HzBc55dYyNTgI/hm
vbjuysmEdKDSKxeC7TsUbRvpVP7/nMWYTm16n+U/xfq/OlU64J2SriChwxkwCTa4Ku9hyBPotI1U
y8+B47Eu/Wie77/zpwoh5XtnCCYrcMptIUHlTHfwZ30zBnt/+r+KlT3nCy5AYhAiu0iB/Rzl48lo
nWaGFiJMoyd76uKLQOSuUdTJYORoDEVkcuyJpuvnowGpVro9GCPbzYY/d2aPtkCL6o4uHJHVO0zA
4Zdy80uE4x94fDj+bR06v8yWitzpjEgHnmBuFWSERgIKAcS6d3uvDX5NFT1TYIaQF1ezCINtbuQj
JYUTyJWvUx6f5CbTmgvBvfC8AbPcn84eAYxD6C9ZteSvvtiSalesvjqay2ycU4NfuvNIWJxJJQT9
eQ9onHsrDDHzqO3t+L3FEVqfiFA+qJa5mDVQ5MygA6rok4Zng45WSmQzbUZdczWAQaXTVenA9nTY
mCKHq6uRzNGuOsxk9y1LSopSAbVROry+tG9HYHJGiZaVHS+y1oDaEojSnGHgKWc8IGczQxQ27UPv
VkURZs3zJNh5brwtpguTpRZRW56k5+s4z38hdz/IvVVMHPnHG+J0P4EjMI0ChVimrIEn4JSmyCPU
jTX3yiiKs6Khn9JmMknpXwjfMZ0Lst8raJ81ESHI2X5NPDyRNeTzrXbznb/m5MScOf+iQ24rbUHn
IwFirJohrujYFA3MRignWi4+0rPAd8KShm9WpqdpN+S4PU4VQ0+wQu41FoOweM4iKWw4tZvd4buY
9NRXNbseT1W+YoS9C6uyZ5LZK0jQMbY8aiy+NVE+GSh9XDFhAL97D6jeZYu0q+vUisVt3vr5JYS2
cuI8Pl2zwJSJNFjYIE2ik0nx0VZdSyZtwowrd8CSy66bYhy/W0Fcwdd4zGkrDFE6aVZp/8KQrluH
+xuGAhAGRyumP3+GaxlT9L6tur8yiLe782PyBcAsS3NJEgvEQn5nd+N6ibKJ5NQGHtjXpPJeXZXy
B5EL9nE9d1+ZCjcy+EHnnaEVaSlpMHZXPwbwrpvU0F1eiwSzmyPyo6SDA3QdSWOuPA5jtLMl2PZS
IVd1qLw11jce9o23rB8gX/UMWM0hM/NDJD+eK8kVTvXUD17YZHDArhAUrXkAZDGBCJ4ky2MoRk7G
JGh71KfWjR05SXApgLnC7yzh368aouTrvA8TYTRM5mQ+qv4g4qO1AKr5sDow6AT83nmg6uKXmL2P
9zp0QTzxRqtW1x1CavO7tY0XKgd+pYbTSajTj8Z+iJAAyXlg7SoS5lhM07RwdTK+fgmnLoMee+F2
cv+nOSUevkpyn9IznzRxQ3y6ZztGTzbpfwhy3mKIuVweLtOcqOd/pIWx3n6twE4EFC62p/IgnH0O
B/QHrSQI/6z+519AScTP6LDL96pX8xFALKvaxWfqCNlFwhfESHK167HJNy4hCrbzLT/LZlhRMkZO
CQwMZ8nAC8go+8oy3wfo41J7CFXv6sk2YehwQDtKs8Zvw+A5hiuuIddw/MhlT4CK/Vygi7Jjt2xt
N4gwtdGB/hy2GL+gORqeeYNVXWn54oB3Jc932lwg90GlXjUZLzlHTDA1wycBa6hp8IlI+qEmCkCe
PI8umkYhP71xjLk0gRI8owlESVnf/ZrqQlxWfVTAHNWR5LNVhq2wgMdLdPqHO4joWSjNd8UuUseX
HAbwmUP4iQs4Ak76NVgXZb2gmE/rkXQzA/WBI743jkzp5tiGmvOZQQ7N/iUdak66jT4d4BKiMzmK
yeaEj9Zr/4OFjvq8PXtZQfV2Q85HfJOmfXxPKl8Tcbrnz9MbITIqp92Rvsm7/MnUAyaTSaTDKaP8
FoZJZOnntA6gAvnJVOrgjpZdVs0bA8la2Qw5kwRG2df/C/mntoyX5e+mDdfQboE+O5wCq2ENkFqB
QxvgnNi9OoDZXRacPnGiq3yshxrwsb/MKX0xNr3RZcFXY/qBVIXeCw5mSiUoqiWO4y+pf6WuDtKS
vPonYgYx47Jv+I9TedR0R50VhM8OromwdZvW/MQuTv4CxDwNQRMLR00jE3iuPP2Z//fhu28nrFlI
0pIAb/cEWt3uBaXy+xYWTUNXX7WYiJREyEJ/a9NhRaZA6Rjmms6yQA4lw5mPjl5uwhGp0dSPiYkk
vl+tecFVdPyYG1T5hgSnAYV6RIJyKmKyNZMTt1CYwxwI5TPT8pPfsIg2WglC8kwj3uNDLiR8m83z
m1nK1WFEDxrvRjQSGMru1whI0RBp2vyYAVhEJNMQHCs8dAvQyJWlDfsChjr4n+qXaKJvqHAEf7Ke
5S4hlCYuZquGHYLCBv7nHF84GcLYH2fWbbIMAhRG0Eup8hfgxzbYzPv1m6k0rTlODQVSEI/4Hwrq
Lut3NVdnamrStAA8ANUzpPyZJMEq5Lb0EhifLJDOZ7rJTMU424qvSOupVpQj73JLn0y8tYWDIK8v
0FAoFwTAsdFe5w6VSzIJsmrCObcCjndX9LNPsu9eF2w98f8X8uDYNCRrSki/yCA01nhDsqR/h8NX
Humsg6JXEtaltplT/gNZwVAPXdybCQSrccITq79tTOY7LWHRVuCHl1k4rqzOdNAcFvziWKdzJ+ET
UiC+LjQi6lM/qQc9n1Q6/aP6C11Y7nwYkEaAg5ICQtOyqvlKhRwr8HrzhlBho0Q4iPiM5Ez3F5c8
rjpyX8dWqzl2w15h6oGtl6SzLeZz5JRiEmd0AlQGFjQFTIqdV/8RRfZL17dqmjYf7GqW/xPPEUz6
Kidw4PCaWheAJKUUJQxtgetClo4dCT2hc7sDJjA3IRf7d50PTvqBarlXBx/aZxgdKjE7joYTH4KX
b7+KEinTqfJxGY6lFnKBe2O7z8uMRyuJrEwgeDsrvxoGEyfy7hAjlA5ce+ElfipOWGFcN+tbRCCo
8AlNTjYNSwVw6xc5bjdxHRM4VJUNo5xH0Lc72r/CJA0JBMh0tGN9oNufxazBA6qIXRezK5Xl67VE
NTJ1s/0YVR2e/e0f8lupRiNY587HDxcu5UNb19JbFkzYnK5wZP/19ij4B9shaQpQpu8pP/rnd6rk
BA5P/lgzsVCAMDLoi3Dv2fNurqOTUmozOpJh/IJKP3br/RKtmSLOHPAUulUseHN2edGItXcwnNbS
FCE63T/Swkr4fVv47OkLEPDZAzG2ZmCGrxgAfPtdNFJuvDbW+9ebQaeJyN/od3DUjVb3hTjJc2qy
MDreOMtCxzFSs/mSCXzaVl6lq3qA66ykMQVUt1O8wgL7AxyhQp7Uda4M3X0glJG2Ogx2PJymVpRd
Xaih4ethXgMAh5c69koaMTTDcLLMBm43a9u31HpsWkXdKoxiCuv1fiFy8gqoIKTSDpCFbNNVH3qB
mgWQBR+x1+fDQ5fIJOgb+LorHzWGgqdNkCaFlS21AWq7/vNk50LaxR/H0tsKqWs7xcwQ11Y/BSUp
GOJ+pRkq1nZQ3gzoq9FOS+sbGAtpAqR5TepYPXzbxJDzEkVZ19SAj7PWlyZhfuNPax1HHLpCIh2U
LP+eyIjx3nurJhGdY8IK+wDjgAEbVQ8Fyqv2bvWgkP/YIZ8Zu7klHwt7BfS72NvWgG5ltCuN3ihG
oETSQjunxD0i1aayqKH7nh0Ab2X5h6eWO1jLM6RsrCibkNszupgIR9xw/h08nT1zsChFPsaE1aTM
wXToCh6o5mZX+3d88d8UQrbSKySstDnt1AlELrHZIWzzV3NO26X5+M/pIbCFLmL6pXLHlsTm1DPA
3zi3N0snZMQkV9typ0QPNYurUhegR1zOpxtAqaJx2+tfb9V19igP8ufcbrXAWEFfQg2M6JfMUE9A
QVl4PbsJMOMCfxB0Fn2zHsa0j3R7UWymbIenZMCRelMGqSIjcnvFtaK5aE108cQmLrOapuC94+Y3
C1YHG4PFLIEYA3yIuq4FO/kmh8wMHBBklLjSdIIWUnS1saNpZyaniImtJV05kpdZ34XthLFiKAlG
RUWQWo+qgjQKaHBl5LqFC/seYK/y5S8kHlZrEaKFVdprFsrOGqiBuIVJ9HCHKzcHPLQS9Gab1X5U
gpyLhkza8K8PIpyahSvD2fkzvQVc0z8jLK7UEzIUWt+CMNFou5EVzuqEg9uuUmQTNw5vWtEyExZH
KqEs+pNzrDsljdNiGBQlGW9NXMPG6fsgbFMGKXiCVO/xdYQ4gzSTDgXEm8WsEw6SCwMM9jMWTECX
2UwDeD6+vdIQq3LB3Jgxv7T55N5Dm/LPqZXSIaZcmo/VR0nUVqEkVbZWSWoOJS0O5oi//Epi72pc
vE6OdHoCpnNyQynFVriL5N951S84DE8w47g/BjCVfKyJWfXs9uzS9zpEyHftCoKRL2R+ZnEdiNjH
mnqBYQ+hv5+ccGExLgXg5bLAbTZ+KiUXtDXNPHyl7qLrfr4MLyzwRYRUX3DFIsf/BQi181ebKsVQ
FjwQ/k0lts1Ad4+pNuWe5HwVwivZ4K9d9XDaczzsqQV+aH919uy14p0Mp4vw3uNut0ApAxXVDQeA
URjnjKLTGaNE1yRw49RYQYSUPLQ8FJ+oUwgYNJsdKzMVx/d9iQYA65eC3NUfjscCBkpEPsFo3xbZ
0pUbC2EsWE3swwxQNGx5UQTq5sNJSXt2ddkLeBop8i7ewpNZeoYsgPYF224fT9tiHilg9sSLgXdC
UdTB02ugyWL3dkr7hI/YoZXjIVwJsdK2fHkmq/9RoFRFydH3iEdsAwKxHT/Ph5CCvhWF/P46TQlr
LVGAEeYcQEuVq/6cJ4023ihddj5bTub/lbZLC47dZ4YaUtOtbJ6yrZJO2L+VnCjOcNFXKm8vedFa
xWxVNK75c3MWPo7jvI/ffBr69EYXZUCMb8+jiCtGLKCdHJ4PRB/RI3UsXdazVpCRyLPmTqaE1+YT
WY2Y+oDjq7y6wCOR+U19lOnxxM87KKsLP84uq15yd2/bVX2R/mNRA8in2xgYlqVKXU40o/w6Gpid
h9pzmPaA1P8Ly/dtDyqkxsH+0xsJlkmOzHhnhcDzUwB/blblLQ/xLu6N4/V0Cec3Id+j1UXlR799
sReQECaX53HjfX0KoyoVW5FgtVqxonO4P66CwuVliD7SLX39U9p0egrix9Ama+9ekQatgIISYaKi
cimEeh2MUoI7Uaq0HmNTN7Jyv9b9PwWWXLZc8Gh5aYSiXYoQ4k/ZAvcNsG9TSA5b+ROYEbanv9Iw
buANrokxSvLINLMBYAh3x8NOjEfXNpq/7EIb1ldfqpMqIQO07neM0NqZOC8V6Xuhjmr/nAO0EVFD
hmZYzjskXY6yx55xCPYPcUkKg3cLa5TfYULR509yvOJv2fUaI31W5ox05xKRGXuJdmL7XENA29lA
6QlxXABOYjaHTq4dSZAahLqrXk060whKqH6Il3+oZMxoVY8PKYB3NNoAojGqsI1QXuniJ1rM2AJ/
MxJ5y6KlsJCWOsDXiDnStyrlKIViGNQi4I0uPepVBNu4hqJQS41vNN5HRgt/NCcKABKA2uGgLK74
EO2ubOuhBRAGlu1JBo7IWWSgmdGcQp3aOojkyN4eiLkDoh1iTIFK3v8DZEzt4i932TGzsNf6LZcj
B3ffyolDHyE1OvViPLN4w46nVm/jSDeYGc8r/Z11jVYysf5p/or/uF5FDY6X9YwS5SapwMPGz7B4
9I5k/kmHWGQJH7Z3ySbNHQRjoLUWK8DuGj+tpdr0foJJXpPc/csX7SgYC1rZh1Y7PDXq9zmU3keE
x9nHjNfkw3/rRXGeJXrLJqqw3krsj35K7wOUpCeNNoWFE45FVGAStmaz/+JdEa6wDqCXYOavmbji
RP27Oy5YAPItO7Wkxd8H2R9XTcon4Y/vuzNKGbEBSHiXNvvKw+9d0qYyKgMqFWhkxqy3apbryqFU
yprZp3iZ+T5D2tEZJ5sm13Ox0sKzLse/ugKogSWGP/o0dOC0x5XIZ2bO9qhdw4+0w1A45+TGiO+M
puBtG1kXnPbz4UEoJ5yhpwudm+Baj3k5PJDPjdJYP+RgrD1366oQfJUrbsstRYU6kiPD1Cgbo6Lv
G7NaxgFhbELYzFPaTPnCLXnOJXC6LVAjoCTrG2w0qE2uuOFevlijUjoXuY9Za40cHp80HUH3SAsG
MW/ApkYgsgupFiT9J81pg1DaAN18w0oXIY/jN0XcuzhWcR93ChRaWGR7sNZSFi+hGvPYfRVF6/9e
6x/iaVPiV677d40PKhu4AFNWVp9tDVkSz73S7wAexSaIRpIbET25CyXHGgx/03pkckXk4obYirRD
aF7OAHnOQbcuNqVpjpUFTWefkn+Io3gZEexxzOA8NNi5SvizBQ1+YixzV23bKsFIFjVvjLv6j2hs
bq/6ngNf3egsIOsJVy0Sx6dz+ZdE54DVndPzS3jY3EjMNwm1/7qIIpMBpvPtCxDNEHh1ehbyYiLJ
pia8H4OgSkVFr6/cs3va06BLJcgvyXcYyPmJeCQd1gnU1d9r0ktkBvqGHgNSIVqYQ0KBaym+E1KX
BSDoJChbhEEfJIkzexkqZIoX/zS94R6R3qIDk/lBlAAxMjSBZ2alaujNz5olH2QlEA9vWk2luqCC
pQMUHrFUjYiamO4alkF39sbC7MO+494hW1re4FECz5AwMDitsda24a6QIrugZjdtmQoEb7N49VBy
s5ja4N+RQhtOgLwqvD8u7gETswQzpa3vwAaGXGyCBl0oITT4vsIZ6tj1FlsOGieWb51be+LbqVRj
4rp5EcIxzmhSC39KtNkdAQjqUyarTbqtGhf5VdtKk/ld0pMImoS2YktJqDpaLv/URL7ub35W+8bA
BgMcw0ruiKWVKVIsLGuiRTWKh7QNKOhb9AuBMiRdJa9jbxoGSdzLyqPHbc080JhT/T7DsNN5g6qZ
nCMHvKX2LP07moBlKzPBZZ/KD5p9ZE4xwglGCtLymujgFSGKGlhFgDbB1b6ev1TfKj/couyYNKsz
KiCJYxCnTLwbpD6YZKeBxFmIpgKHnkExPTMSBpBWpk3vF6IkGxmLd3xJh7Ofxsi4MgIL9CQDrjhP
eJOhkkjupeQe68CWnoQaStr6njXKpCVVEtDNcHLMwCCgE8GZnoct6mEwdhlNoEx/w/Uu92lVKe5b
nktn9s+uoPYE+lljmIeqgMbl3LpKmS1cW4coIg518Kk1w926N2zifX9R8fXHEt1mdkJr3wtgQQKq
KvYgceHPdNkgdBxIEXbbdwD5GCCiA47Y8UgOe2BAlaKZWytk/T6lNXdRJ89jaEwE/4sjMps5oVa3
hvzYy2rrRL+iGVzwLAOqngW/6KdOryJ0omJ6C++Uyj1CXBKYaZVCxjW3M15pXFZsq8IZAOO+zBpu
73Vv82vNFdqDV8f7G1ZSuK0xFQ1BhDJIreW5t/4HR5w6SYYgQPKPBl/8GKqAtJIVCHpIzWUSVdnt
zOa+A2c8t49UXqJvzQWyU5xLNF/yu1SIf8R8+Xn7ATMYEy9hRNyVSXxiuYI5OBev9EGauA+8pD10
PAW+epOOfW8woJo1ZIMr9ez/c6PsNh5Jz6R7sDCdYkmB7lOUzwtfsb9R8n4HcA4lVvIwbS2JmKI9
ttEdEh3JPBb3nwlfhvMZ6uhGtNJCchK5nOyo8AMFBZcl9FIUxyCwIhGkifZHm+ihn2cTMbRqATp2
a+7tNlZEDcZ6uY/zD3bI+OS6tsn2nWQ+y1Z0zZQ90s1RZFle+uqCQeUP4ODsUcVLzjiGcWHxGv4R
3tAp/taCalzdcwL8s+8xpiHOJHXwTOxDHGautLoOw5Pfh6J5G9EQKWtrm9AXDEBO5dtUyytH1iFC
M6woP3p+I0u33JBFpwFDrLy/3vrVTo+i+e7NaAQhJ0YTOXySKAq9SKc3/XMt3EWYPffUM07WqSId
buzBST2cYQEXTCyr14GFX5Ukew7wXVIXTRLpQOu+by2MN/t0H2nYjL6GClSWNvDI4rfoHf+xX8tX
anIHHoRkHh4LaDkOFgsJwr+nGz4/uxyMpxy9meaeqIRn9TUK3sLsL9INDWu1ICZddPAWRlAKi8ta
TEKhatJdzvX/Qp3LkfgigxCreaxKcGEt1LTw5Rwe+8WgYhedBQUj1vYluemS+9b6pBxE71jTg897
WXteiFgehPVAoN5U65dqmdGMTUaDKTf/dR58FwX4jnKTCNa6FicW1PCtSBt3h4zd3bwPuF55z1EI
x7z+dtdue9d7VKJPZ8jZwq7uNtMZAa78q5rJ4f0OTc3kS1YpTZPQu2SQrmLgOXnun/ZAbhQsgntp
2SghWB8Q0uc5fGPDV0D1mhKxkRhS16bljcugnCOnOVA/j/vxpBU1Yq3fuMJmB1/ma3/i1AJezhr0
menx3LAkY4WM9ENyfusMbAl4V1KhJ/vgWsf+MRFwCOZ1yxjVdQ9zom0U5MntcHA8qwQEDKB8W+xH
QFbhWC7WDCS1fsGyjZhh/ypS4jFql+uciK7c1q9rBbyLMidprrmkue/ei6vFkrLD242C8w8NcPDW
ehl1mGia3sb8wZexX3kRtDicpwx1XHZ8C/4U+tBKHI480VBRxMUvaEcOhKdLcctTyZW4U3iEw8wx
81W29zLja+mSOQRyaFkhuBUVOzqeS8lLtQ44c6f0IY/Ucbs/gdH9dwYMCHyDJh/SkCGUnFsVDEqR
Th6NdoSWSoe+HaVEug8lHDzbY5PqLtg0ZdDXGz4YHbIB0Yzp7Iv3UpYeoajQN/QxRFm+r4Df+jrB
LroSao2NCZz2PabOpRQ1eO0IjLRp2qdCZbl0zIubD8ICcBeq0NTSDWkFyQGJae0pq/pdrebV2DZ/
uPjHTLmCD/5ezaRW5tMVp5Evz3SWr2Lbp4BMYOwrfGlu04oxf319KGYgPaAZCeCVx8bX3KMXbTDF
lZQe+JvEV5feAoNL2YYuoaqPaCxrm/uYXQG2lTkE2P9eW/6Rv4akTq6jXPqnMz3jJRWX2thXtBrI
Uc8tU9FyFKGw6LowxkWv3C56BOmN5RpUVwdPRY3CddIyxeKYy4sqpReJsHetxNS+FQT8j+J4PzUW
1R4ST2dR9AEqhKS+KhOYDSz1mHuVvWO9Q2jRepBpieTnVUhzp5v2BHhuHBmqV7HFg+dj6RfrRlC0
TWGk7lHoNPdj5dWEGk7To4lfCppJGey0V2qX1Ait7yBRVMwMszyDiEZqP78Xa5XZRkzn1lfxmHDs
30CrxPFPc4e3MFhOXFOQrMO0a44O/sHd9uvZlaC0y16XeRoyZNUpg06y3rtyEgz8bRdCqlbcb3xJ
N90zuT3AEeBnJudqPi3YxClt8GM325v+hV87SKMA3to0vxrq0J3gh7V4nbvZjl2qEWGikx9bLtA5
twEzCwp40E0eNa17SVmM+cRphBdLokdQKPs6xXd/CtwXNAy/1WD3olpe0HsLIE5EpJP2omlN6gYX
umJhV5rMRKzXsFQIGj/cXfUw9yMtJaFkTpGDIIvb2Ul/cQ1NCf93/y2tzfaeF5sHbsx46ny7KeJN
ivCxEyUBKHYc5GoL661Lhg3LDzjQ3u8VPbaSsDL2DEGe9mi3iVqoKhrjZdt/ld+5+po/S+vtKUp8
Kp8EFPY8fkPBBfmKIs8h2Z5z51pS4m0RHBldJY9whEbdWlb5S2FxMgO0lZ7ovEpgiGnJy5rSH5HZ
RUJvCwgM0hVoLTuNVqM4SN7NubLJBZ+ckycf1IfY+4ZJ2mopV+o46EEhahsQsyBAS6mvNWLpmCQU
OaWmWd8tjzGeGccyEgz339dfebnyRz5Uu8QMyGC5llrWBuZ1I1FBKAxsr329QkrT0bzWI/eiPVYc
ATUvTusNQS74A4zi/RwPjgrgcLsE6XgRoLUxu/1w5Q6U9XkHdLJ3T/W9TymV+ClbBxbUyel0sNr4
BU1Rn+Cgy+dT9fOiAKOhWvLbiT++zF5Gf+GhXaOIx7nDwAJxvpUCellg/9QmjA+Gy+TEAo91iC9i
ta/Ezed1lJUOQ/B0VKK8xwlqQt4hH5NwjCbBMf3lUbC3/OUH9nUXZpeBsvHaFjIyrZNhCnmhbtHw
OueP2at/6Iazzo5eu3rlCwk4GEP2NApnj7giVrC+G0qfkcfaCEyJuLgVkfY2szRos504S1Accwm0
ectoXU8d32ThWVV9af0WaqqMkCLnLvGbGgdP4POZEBwxH+/H5fN9NFABr9o8ojydtxHZfPNLg9Qt
gcP+PH4TOsI1OS9UEx2CqYRGN2QuU3Hf2hGp9d+M0gpMc5ChkxXz7MubffOSjzuf1hoX2dVJzXeM
hplkGgWgYHxcAUTktv3y1G34buR5z65nNhd6T+dk3KrxrsqICGS6P95kAD9VQIYHYjvAheXR/69W
SPe2IRu7VhAlXTUIpY0y8spB9ccLzOn6Hxg55grikDLJ7qk0yJKLbakKchuGacupC+Yji9JncOok
x5h/Fng8ed5q+ybnp5+EabLBEvODxSabGg081y23j8RYxC/5EbDuocUuTcF+U8NNyBJ64qtQqyBS
hhjLdZpAnOzZiHte7rVyagO/6jTteZ/bCZVWuac85APCk4EnDhC10psqbxuxx8jBu3LLXZTQ1IwH
gSc1gmeCQaR0gzYrzWE9SjbOT7k61vt4WzRp0KpE8o3/95KlCVTSNOWLCi8zJte4oryGiG6+57FD
Hi1BZUxjRtqYMlvslwAuCgDOoGv4VMIdGE4cCVJuEpcn6nke7b2hIWy1SYww0Q8oy0LDHvWyEBQI
Ukl653wk4IhoC6kkQ/gpyk55Br/tYCcEz7bL7Bj9XiHmPzeoyu4ApsJ8kPOOpe1Ld+dlkr2bCTBy
hq+YSq45LaEeQtyMVBCzDpw0gCq9fwyVFOpBQYXqkqjrQAqN64CX0hkkgxVAqdu0Druy7kremZQF
Yi90prsGf0wb7NJJw6+r55GqWYf0Dc0kLXs0ynku8Ir6ENgGowHt8Wk4NCDLsWKHdxmpEAZm+xpG
0mYOX7OxPSI41q88maErMa4SQ1Sx6jdJY2Zhkf9iy/nA/3tqhZ5LfGV92vgsha0TH3i7UwKoXsl1
PvhqqrIZud+BmxXt4HXZepzgUHJ93jFcc+oT5myKNb0e7EOnv2M1xVkR5Tobpat9U66FB+ljEWvI
ig88a5nCyE+gSSDQMu+hUQ3nf8kr1zYx9uo4TvLiWRbrAn1sAfCwYBVJ5M5wqAKbzZufKh0dvsXA
vXe6FIxCBPb2KEl8zxtIzBFDr2kKmbhE77/4RqcS7l9mw+aCYHZ9sg2BqqmvBIhAs9QDulbvdjXb
L/6k7w1BTTpUlbEAiaVDm4sbjbCr3RFJ5AjpW1kf6DKPAsdcmgA9D4xssEXLizFAPmkn2hJ902OH
YSpeocTL9UzYmYhtp6q71nMCkMlsbdH9IGxvBM3kVuYNRb6QMAVtSWu45CuAzLAHdeQEURq92TAf
8ezzhsBPsa6NCJHj7QPC/2H1X5Rat1VdRLhqmZZ0RKTxAnW97ZeyJXqcxUkeArk8PGaQvCAoU3NA
GqQ+6a/zyANEUDhMBXFJd7s+VmWXuv1bbS//3CISrUKO5r807iUoXZp5SDUnQLxFjbctrLPfnsFh
Z0RfayrV+qcwiiXoctVrt89wNur+t1LV3pDQOQXMKC0fjX6+2hzAW7ibT0b62UKFgHzOtu/2RzEK
Bk0Q9xqLYU8hxkw71XhNMaEq9Fkniu2iWltaNPHpYyuCTuiNrpcy+VKrvsBOjB4wliUaXaorh0E9
cfQbzumplfBRr98dS7Vg6NcYqYLQD8JpadOQ44+OhYs+mHeKdexSc2mJbpBp95kToJ4IDXkHkjsb
fhXPc4aeb6RgmFGiQmCScTgo8OOLgeE7z1s6RKO7XW3UAiDzrLodDVgaa3nwfR61xWmhOS0rXwco
j7M4CMgoXsrfvt2svbp+Uq/IE7/HPJWaXb9e9gjvSY3iNRXSLEdSZ4nerGYYymJhgMEYpdPXAUXR
TOATIQzptZqOjRsvuxibQQM+X1lpv5tIDcli5zjdgjxJCuB8+vbAOLuOa+sEqJA3jkiy9PAE/O5F
G4MyujZMeoLZBQD3Veg9Cia+gJ1trGRDnuCvn9ATsBYiwgsylmfHRwwO1mL2NBvHvfh3+/GUn/Ll
/rkpwXCnAGL8brr3najVujdqVU8B0iuyJGF/lFsQGXR3UFx5FxpXrLUO52/2GpXVSvXai1PAeEXK
cvLAb9w+n8F7uBKTo9d6zp58/ESTLyufUtmVN2AO3yFDzhlHpxC5OoxQBFqoGvNJm/F/ehGXdJNA
zS/Y40KW3x061X0FdtZnwRhE5G/TZvGQbtEdNBfZ5Jfcz6qN4xLOqJ2Sabdc0Bzt6LtsQ+uoexqI
qfjvWjWoU1J6Qx3nmTR5Ce/4gGwETJXaZlRdDQxNJwwOtQLDluX+JwPe7VHFKDpjMp2nE/xbVxsa
wrBpL466R0oezCU9gaLfsqlb0xgfQtFl7G4+pzCcahym9iOGDX7ybMXdarzRomRwgugqlmhzNYfs
wwgqmHwVHlqfrcdoy3NziIQ7MZORtM85aXnAL/1Zjw7j73d/NaCPrliYXsUxauYvj+WAFOHBl+A1
JjFAu3i3uYD3HczZ0xZ7sT/tRx3Ecd1fvvHdP9A2q6TGjqWG6uHUYnkQdxvH5Wf2liqSPNquyg0Q
7P46J4ngyEgFwi8YoB7KfmuCgOeN4ItYSahAgGPSr36ioY/DR+YcXbietZ86q3N3xXTJO8If+mfb
rrZoC1KfUNSiYn6PpEM+e76GF+1vP8fmopGBtu8+F9ZSOtfVJ2uHrlWIXEJwuf23lYp6Zd3FjL68
6tchFDF/NfFlWuFJCfhR0CDWUgThss0YCd/hZtXP2FAS1RZWf66ShQ1BYWpZndoua1nR/U//iR5A
oUz1W793pXuTEPKYpbuwbykM5564aTqYd7keq6yQcOKRsWNQg4MFbrTbss9rhjhPALy6V4/2t/QL
hlzvLHtPOtKKfAsIwKALqbqfk447WrOAq9I+R8grRN9662kx+w+fQ6Y6wI01c55y/26O1rq7oDCf
DvdcrdqFqHXAqxJK0HU/o+v4/pdx6f65n/Id2zEbWpVLi3Sl33LQpcXRA95PeVPelLoWQWhWEwrS
TTKRnyDHXabGXbzCA8hEgaDQ02dkV+4MShOU1X2vRowNrFHhaiqHXvOnD/KX03Bpo3DyhC7yTzKm
lfLY5G8eikmyeTS9qFXdRWQ4aD0Eb3FlZBMQk05RweEieNCdltKD7+rel91FX/eGhQ+DyGehwlkM
JdnxO3hBXj/hg0WtYVU1eQEYhTJyv2khPZTLgl9hgm1XYfCW5r3AYHtq2WPcB4vuLer/FCXvacBw
LMLhM5y4nTRkrYzlIByta//CRYKVdRozlXx0UtW7PsBYakfGkyo50cRHkpu6sgtAPVMP2vPA+iFV
ud5qsPQ5go5zGx00auNvTSTWMmd8eD3HaSD2CD0EKUtK9cEC4GlfPB4lO9Un6HmRchhXWraYF4bM
+gsJuN7FlfZcgbQtOndrvbLOtFjgJDUUb6QANlSkJyd1EFysd1VgAL3NPDTbmpToG6+LJ4/VQ91r
EDzB4mme6zVktIaNbKkkhcOAWZsJ46vd1tCbDfCKN3wXKqVAfvmdq4zwWaGe7b5/iWjSzFfUxCUs
Ijo6F7FvvgTZfOCxQZMOrmCAOWieT60vqSTvhEAQAuHUhMk8TrL8elrR2TL7Vko23owB8k3rq69+
IueNQ4AU6xYGBjY/sOGXPYxnP4dzSQkM95CRU0/EUj0XiEwUaOD5t1BH9xOf6BwinESqUEphmKX0
Z0gnUMVW0LMcmHezMhbfb7wfK7I9NFzJBOpGrPq7oyONxMnJD28RZXpDEdfk0vyYEYWZbcM+ypn3
xuxFd8VZnFVppMPydEhb5YzYA78VTTLC3egJCGSHleLN52RWqG7NkP2ISVa0DtuaxWPIN1VULfNc
taDZaqUFnkIabkc2IsrD/fuwR9xzsTyhqTEeF5FeHkie876j7HCjrZ6gSAveesopTR9GVVgvO7dS
L9sYLsPSxnwcAjfBycda5/SX1dSsz5XBEicBtX2/PRT06llY/km83ST/4youIjD77VJsGQSigfvS
35J3/ppd+bXnR1bwVcXHtqFnwF1/4CGrnttLmsHQTSxmNAy/njzCNxAEr36pzPWr1oTN/OWdtUfx
Epubvc2l4Flj34iilWJph4wTv0iiZeZk1PqGHMLAMgqCaUwUKdLcHPxmvnwKiTuYjMTOGNVgSmA+
TqEAX0TDLYW/s6RKxLYlmLEXnLdxHg6ZYUtl2hXVUGh+5sIgdPNt5mulA1CeLCgdqXV/K3/UWVNG
y3KpIh2umVhNGW2iRAtkQrJwyu2dAY+NcjfGjW3jrpFuP70RryQJNLMRXF7grpyYSLpaY+ciSDkz
yHDCYEQuJz2vBRTDOqOKGxD1buxDj0hDj+NMUvqQPfWZGLvKA2UnJCSoK/+ij4r8h/QNASD8WQh6
TI7+MZ/liWNn368qE56e19l/ztxSdi9hbG/lx5iGg81HBDM0+j/XQ7NUb0TsE1aPndSotM3Jp0Bm
4FOiVrUrWbiZb4CsiBG2cBVTiM3rkYGrfRdtED+I/i3vIZ0cDlBrqNGoGbGzIGfw7CRcwPfvkXNt
zUackxWLbID9ymwsZjzffHBT0df3BpFLjpfHvN/3tUoO5EAPk0rwOR1oJkZQ55HvcOetQXeClJa+
Y90xTmq3WwlEqsEuIcHWM9jOFgY40IIYTFukkiaTXzPt7pfrtbuO9nZ+4kzWg1DsKlPn1F7nitKp
lCeqO8TSGdfbiPv4lWtB4U0X+RhtBNi4Iz3jYH1Rs4Ilff+EmrYgOCx98uAI0QFOxvoCBI84jujy
SCChnJy0RiDpzVFqO8DPGs6ISj+eQsoIFnYfKdII34ocGEFsSgds/nWkMXZMnM+Hd9WLOCzVV/P1
OVPN1cKzGFwXe/YnKOhaOREPjSSh9D75pvuhUbnqCyHl8hAhUGRReRCCewcMQOAagF1fgXXL3RaJ
0pTR/TjfyiX+YDyDByDjBzHk9VrBvVi7c2Gmlb55zooj9DP5347rWbTFBHTbtDpqcITHtBCDfgvZ
9rTpkfhnmJszUz9nhgu/d3yCGkvRNlpqM2KLICzuems46H8u0gCrcA1m0QLfrf2to//7ImBXyGFz
tZI12DlGZsRW5wCI03uzPhCEt8dTe9lB74Ya/sbMit/myi7+qX1BauZGMu8YW/KLKrC2ro/REjg3
bOxOfu0zxai/Xw7Vzbnw/1o8dINND5Bo4oJTJmZMfj8jZUcz2cPKdilUXxRz8Foy2wmOlvSti+ZQ
v121fl3un/Bd7ztFlSOQNndBkXzMr0D0YEZD0xzCoEEBJ3Qbvh3oNiA0uH6jPPAwkYCcnGHVUMF4
NMUahPW1H0wxyNf5HlxCOd8fqIOxB7KqetI36hap6/kVZeugv6hGHFVmDY7BjNXCZbpzdVMdeps0
QGkwd4d1OKx8WIqRvWe5pYMjzjVGoUgCKYbPTyOc4DiU/ufZ8P3mG2F7Q7k073MLtAUlPEu18YLO
ayTlUZtGwXZJW7dsw5MmjMr3sRko8CHGFxCpTrPe8COfv92TBo3I3EKLkctPlKucf/fFQXbKlUQK
A0CRvjvxlX8Q8oszNVkAkNGMfuv6Znf908e+iRcdnvaw6Fy96JqAqK+9fNa8X6vfR3/3UaInlubS
bDx2bN34WaB2Z/PC9zk+tcVeDaX0ihT9sHEjkbFJ3n1prYrOVmzptldjLbPjt8584NN8qdd2x8O9
FR5wSRKDpcfR39McyDA6U7TYQ2YWT5bfJFIFba80pY+64Oo4M/j0+T35+UAn5ZTBYaTtpccdm1KW
eVCjJTKJGL4uXscaxZCMgp4/v1Rvd3fAP7xFN4wpo6Gc6u1FjJo9KpKsrCVmn6VKGYnYW7sWuJxJ
3qMXgF+k3h8Efuegh7FvX/8V5sYx8btPIPl//nwM/b6Qffl4uScQ1wkpOChE6Mmaag6WIPgqD1ld
rrUcMybwrXtIVTSo0l+5C0YzglGljYkJhvAUPYJUdvvwqfMrK1X6sg0w+4DVqOUZ8iAKmrk1j/vU
jETs9zi1PlKLSmKCyd1FteUSgxGy/owIIg8nZVW3ZWHcNShoxcEPEoTWZNmUZwfIN05ghmp8vSf1
IlQvnjZuQ5djEVNO2XcIGaUOarN+B1zSbxuw1tbVLJiOG5SQ1jL/ro5/t/Xg20T2jj/0gOzG4UQr
q4PIHAaFyBd/YeuHxWQHdmDX7w4wc+7FZvcUYjHDv8niOGT0XiyPRC5v9Tm7gjCrLceNeoRi7U3C
74Vfhl31L+2hB5L61zWZNf74b8G0rrNI5jL5MYD5YOY3v4nH16N4SqD/4TwIDiKjiU6Yv8M9bl8N
lC7k2gafbipwolUCprHUIriz0Gb4WXbB4bNAn9Mr3AZFCuA6uPpRgj3YaN1Hu9IRcCh5+4uIohGj
1oW04EsRfRxHo+uDfQNNiA75NB/yygLO9Wa8BliLnbmFJhJYIg6t7SWpH2Iwv/u3VNLanZgGuTr7
SefnBRp2ZiUWtg+xlDroIxAzBOuF8+v/tfnx+omxdf78Mhva31wGGgB94WEj9x+pqNlRl8OgSv5q
j0q0ej6dROV5oW2XVSJVl39iJo74bQ55gj0VIOKLEWQHGUeWh2Y70YafKc+FxLhfSmCQfhGoe9zn
uu3+AVF/uWebCDI4kOMoXItA/q6DUky/zOTWw0ETV+IeZfkirZf6BdpnH4HhtQbo3upFffoNlTK6
BsqzNrTCQdXLpLXvm89YYnHeYl8D47R98GS6p49HcJJrdDW0W161nZNqTdOZDar4mGudOaAt6Rzu
scdfP//S/7jki/eg7gpRRCs8vXPlOy9oeDN151PnDLr3oMNe3LwmeD+schUEdI7MqZWtpL1HdXm/
uEgYTjJHwgo/5PNobLJ+lqgtGUFeYOWppltYp0ujizd7Wb3FwWPPYTTSiHlmys19ILpO+2IE2KQT
/dlV9RzqRupekvfoMjcX5nmKqjTMfcXIDZ4pNAWagPWO8jty00/rPlmTmVnCn4LGojglT9zRUDJn
sZrFoLmCM2hZkUlX0KZpND0mPaUcqFSgtURh124uL78Bayn6EVQtXydFao+A1aNXKeuzJcIQ6Zzi
dBPNJowrXoTAGJ71EOnE4pe6q8p067omb4RCAwP9IvU0RVkQZNNAeLTsBq29wXNtRDe/uUeC5ViC
/GubcBIJw/I0ucEJfoo2QCysqjFPLpuXP4Z/nDGNrzFDIl9bnF3xxCOTazFS4Smr+iIRe9B9cjyO
dHrnGivXxPNTtBU5E/VP2xCkEZmN9eVHEUuIiCDcJL4I59QQZ+CWqxOHQ/5PJLvj6PSZUwsie7vB
qyD5CKJbj6OtG640ptlgDc5eRaQGUDg1R8U8XSYxl9L6G8cgF/Ll7hcFLU+ZQxfXIHzToizmU3Ol
KJ1zKSVxSqIm9V0kA+oUAkAK+gdKi2RV/2rQPsFHJc8Gfm8gVYd9w0HdlBawzDEDel1MNdBcB+Tx
UXT+dFCOCs7Lt8FIFC3CKultd3mLmXCe3md4p/uWVYTKM6sN32AUnbJsKcmrQcAwTNwwDAooWNKy
qwh0dysFQUIePWZP1JJm7aKpL1Dx8v4WJ9ZHnWicIbbl9o5gXq9CQhtbUhQLg3KP0cyrYPjKf6Xz
JV04Y/3vqvOMXpNANgAbvdTaoRSCnxZOJyo9bzD6gudRAT6Z+0jzKjJCMJaYl/TGtLxdhsyrqROF
SM5m9jFIAarE2v0A3oopvYiyJSJrz76laoUH0KCTbPFrNE8xEoqiikv/diKw6pTBgCLO5aOrURnd
qOTWNreJ4Dgu8d7sDgjA16n2sIwCPCGArueKLTqWHefJvEg39OIOD1HPdZjmt11shUbfjwbki32I
aUZ14pmQ1VjSZ7DJ6Cqhfx2/2HHj1FDiomlMpEbjihcg/WgulesIk95PMKpkQojXR4/CzsJp6QYg
giGTADL2C1A6Uu5RH4Aphd/g8BduJIWofhwsOfncQ+z/4BnIOMHfGaUIYuyrNeNBr3ZQaFFGE5xh
y+/gxuMZgxdmPL/EvUafa7ecgs23+pgFaSFOTBZvQIuFvw1uecQAyQFkbc6tYlsGmox3+jevoBIc
6AL+DHyyuvMigsZD6LQglPGIZErR0nm+HfDToyo0A7sekSgBwop75rc2b4ruK7U7zftWmZ4+4C1I
BZu0D5FYhWxib5hu7W1mHb0Gu/IASA3uQxl3BNcy+08tjzG+34WkrxJzFAt4iX+0xbfIOUs0DEpH
bLiaICSAqr7Ob+R1yyAWM0g+5qYSYF+TyAq+Alpmhf+Ni9374CvDeEUWNPERfEejhQqtfkLb5fPN
g+iJNzZLXLQTuLHBEi0nCh6dLl0zeNq8R1n/O883Rcr3ogwJ8nrJv+b5N69AbNGivMnGnYQhIIfI
xlxwozgA6CbPcOukD4xsphQJqQHOlUu3ZsiwQ+1E4lEA9pyHfGltEhsEMTgORNDdfsS44AicKihD
TBE2g6E/MQvbGhIZhFrxKu229TVhi3aq5vrN1H1seJFiB0W2/qu33AO9+kMupsrKZXVz7453Zgbo
bZHRm74wngntiZWyzHKiE3WSv2C9IkruXRTLdRgPqwtbeqYv5as2oxTvgRclMGpp9zRTpYJ3jLdT
mUSFCgwXa+gNpaDhxt2it9efLCsImx8ABbs1XTP4CS9hXyEj4eN0F0I5TcgA8n2a4MeYooBFK+lL
7MU5l8K2sHPi6lPthUGMkzmWHBxU/vt6MpkLvbf+3j1rCvqGUMVss344l2y+ima9yYwEEQlYHscD
QRY73IJVXb7jYe/jsGBY8X6UxLJfXiOmY8VKT1kyNkHguZFZMx+8MWX1oMVqn/wziOk47k6UOwe3
2Km2GRtdMb8fV3wE+bbKnHwGXIj43y0dw/GcJYCxw5rrokveHyH/Y+Bo/giELRBdtBadOrj5jpG3
fVYhvEAJqPruLj209Rz/81qynQ0MEHbuhVQkIIxl01kQuQHdvmDT/obQxGZ1zKpl3Qss8yDhWYvO
clRyDfnBN/ehVEtl5rdW2Yt5CZIpl3wiZoCqnG3UaCEX40CU3GUWTyeFmxkj8LUSVqUhnYz/iqNu
/GtM0PsUmDooI3u9+nU7brJm6gob7guVjucA85V4ALWV9o4oMoaICKVjRwX2zoAl191qqgQwH9cp
vGU8bEGhSiYPAtIDi0kulS5XRHg6ANsRw2qatglQ/aK/E2+vh3fmEMfjvJU+b2Z6YWyI3roqhGC2
yjJwlzNDFBAPiy0H5m30XZB7Hpqq/+lzEqvnhW+3BcTcrPOrzSTZOOk0l3BDb7ME7ldg0kDR24+E
y70969ARg5w9h1R1Zt8E1Uqx99SODmIRRR4bJc5r8BZ9m1LE1mxazxVA3FTZKOvcdXo/Lnw1VYJV
ZHUh5JJcvlO98pYc4Mij0LSe+Q/Q2o3rrQIKhMEhPkCCTMI1H6YlZ3Y8ih1MLGHYbkT4DwyW7b3z
LeLKc/0bPf4TPGNxhQhcyQOVbSgJHuhm/ExRzQTLkUNb025lFrceoUN2Aovl5xDE3BaC/KDxObZq
F5D40H6PXDfvvKIg6lv06GyaiRAJ0HLp/9Sc9TMKzHJgn7aOEnC/PhbhOIiwkRmFJ7Mw5TwZWfme
0f3FiSjHagmF4IjW3v8zrZTNWmykIrVb6rkfF7ICtBSlY6sIlJWRN4W+pbr0P6wFSaQKM5xg3LyT
vVhNAaOLnaK9U5aQGUZH4X6350YEn5Eh9cPaDqVTcDATVCB0oAdgx9dCUUocEDe/g07poCnckAq3
BLxIDxl+Q7dlKSr7qiQafyMmzo25Qr6Ntd80upGObPANl+hQr5DOnDsSNTi/LjUNjFa+yYpyTE3D
X4iqSbGmb6v8rRAqqrNUnkV2DSZnRnLc93D0O5aAtqswhR/KJlhOGGKybayKdWdw8sYGK+ELXrZF
pSmV56BpUy3UNnAvrum3UkuAXpEtq1Gt0BHYCEaF24liWcKH2oQL6kpjCf/bcgN44+q4aBm5kU9S
dY9Y00Lnr8AYKuTAEeUo6u7MwQdzxeEYWVMM7AgatJDQobK23uFTjdLUnVhesslKvcM7XqeymKAC
NUdJe/O8Ueg54fI0QR9cJzQfwoD4C8nBrSf1puzrc7D86YNlLqTwffb5T3c2Gg9mMd6G2IF1r1yg
acueskNPtTPF6CqxmoBwxyDcOb/0NLefzK3RNlkp1Mqcvm69dWSpJoOfdVSa86ANlYB7QjdCaui7
aryE7hCTahrrMkCg1pIDACSuK33FkRd3vRiS9qSx7zJr7gkgyAmj5RWORAc3gKYvtywNsPSZ/d0h
oSfPFmoHTXI1yrZ1L23etDbW5/lwNkcodDaVGxo0KRizExVG8bcUCw+RkMbuS2fd1g8yXTG7cmoT
iLN8NLeeswPfuwI9vhaNOP69FfgcVDgVq/6BlA1Yv46PTFfRYlLLqDddU5Xk0wY42vQZRAd0Njhq
sfcY2BeHqcmjDCEXPbbsNChJPa84luUxx2X13R7YTjVEqlbl21eeInrgdDgkK8o772xJDjwoaOSy
v88n15GfRi2jftnpMjQhMSV8heNfdTooblzq7BeO90ShkH1S5KZbSIPCsAL+CG/YQZ0rYFD395kd
R3CQPyUUHzyfGfv2tnApiDIIJap+DmDj4i/qmdFPplygV78FI/JYlmQ/7+O+sGIMtZZbLAzMg5BX
oKDZB/rP5kyf+ELR4gWY2kUKBefrYSZiLsxGULW+XY+Qp/Zt3xeDA0ynnPYad2RfXypaLptqwutm
cQJmI1O/YVm9VM2hTKOdXll3BjE/h0ekRBFk+GcheJ4Y7ajNnMXJl0U6GxqK2mbs5Q4rPkelMvpq
Brwyvhvb/2mE13Cw2gH6clwacMjttrIlkCb05xpzkmTa7c7fh0OAbZpHOdxiPpIcFGM1PDYEiukY
eMM0gGbr+tgMkZ+zmLw28OHmgy5jtJEipL3qjZIMd7S9/6Y8rSs8YCdstpSDp1g0WVxjcVFtcgp+
tuKZjukLp2NX8wEtOVESIPUPaX41+3peJryfjQJQZB95EC2hTdAt/T/HP5dvhj8FaEdsCPA8Di34
DoRWMDFqpRKPLcEDMH8DEGOLF2weLe7nRhXUgOjp2/DVSSh2PLPmNjDyiYkUhee3xUgP4bG+Iaz5
3ugagpjUNtiDwa9XEHTrQpOvbabC+AV6xi64av9J3gjvMkRqmV3LTJLs1z/X7PFI39tPGpV2/7LV
hVeJU5r4ilpljGGLmjybxSQAE5htY/TSztosPrIajOER1LaptgVzHn6QtN7DOVrD1sq3DsO0tbfi
z4uvzpm8/3K8uZkNr8DusJA+8tM1kpol0UwLA7z9BvwUIuuFzPhOciGBkT576RO0pqazCtHBhinw
ImlsxFlRLFMvWeUedkVFEeh21uDKgDj7OdO+xJiAoG4iOqPJ7wdBj7slNXr+G3jVO9icdFniVmok
jd+IKEv75weO0VTYZeGJdtd2YeLVr0zUf3MBUrEQJOG31RmZKG543tICCFMP1vh6Ww7QTidPZOIp
A4VTHXXfGVhVCK4oTTQlaC6vr1XHiV9cGxDDQh2/3KUItq/HkAEZ3Y8O7nisYlXga4YFZXAXdwXj
xPKibE5q4g9SbHAOsl7h1in2brldyeG1kvoeU94Zr08cNfHkSP67201VkMyMMguP7/h6MhgsXyUp
2Q+NBbMFrtqR+j5zH29SETVDtKOPrnZw82YsWT6BzsSCFFFS7gVWyWwnQO4EjzA10F6ddin8/IcT
y1+TMWxB0eDkbrgpTAAr7zbbtLBEbUJdGrn8cal7Nw+/pHerBidSV5tNAncwNpB2YwlXMw0fpnCS
Tyg3EvRJpuihRxR+9mNfGgD6B1ifzm+R6EvscJ23cjSejA/5T7Zk2zZnb0S6oB5IAX/9vHNcDbpe
K86R+KEcCrdMS9O4sY98KeCSMC5Yb3ArD8AU7DMx36yjCKcrb2HPjnrRJ5jvtxbTCNxKahnQfypT
9XycXAwxOW+E/18Ep8JSJNG4Hdur5AzLfz7Soe4uOudYbLprtDr2ZRUuJJSCgDrI9SdBbn9WNgVc
oXl5yfWcE5wYhqs895cuKJCFfTqxZ3910T9iGne3fdVEYyfiYt+5Fn4Od74iWIT3E3iCN4KPky2k
f2piG40P3dvOottkR2qv58AlEpCjCQFq7IPdbT2xVWB/tyyMHV7RwDmpO3FALpNxx/abr/N7LWzk
CVZzzfJc6Wf7400bCa1Ec8UTwlAjzJp/IBieLlWxGwtc+7mbG8CsOylYrsBzi5LfAa8U43wuzrKW
pS7ar6vHBgbOLnZV5IzeEXjuPDJgaMk3Ko6PHv1jj1b+xkD8t4L3ac4OqU/klICnQ8UM9pelp4DO
NEZowStXDlg8YjjEKOkk7GN/LxgmZQBt7Fj30Uwjhqs8N+KhsDlhbEr8lITU0r+ubpEv57YyEG40
NFXu02hsbGrCH/Kx5LXexog9XsMAbiMGAyZf4AlLsnOHxZ4YWTL/cTg4qBOm9hwdlECzbracCCUg
bhJRoTF0qix8KPQcEMRN5QgSsh7pmlmyXf/acGbkZynTAQa0xHsARU0gIl3pXCRrxm+7GJbzZLIE
xheF2RGUXamq7ZCjbaLQlvad1lkV9vbnqXdch/w7OPoAOjZJiOLw4L6GgwfHDg6nyKME+OVl3PAV
Lcj+RdQhFQxlNQXPFj4rdCg4iZsY1qj7+WNinQdzXwhIuShG2obs4yUV0XFb5luygfmyA1FV983n
XemOzLVe9BrriQUax8lMV8Jl98D3OACHoKu1EcH22sVhn+WMEVzyf2dzavsow7wyWkLDoe+B0NM/
hYZZTqvfJpeFqg7QLeu7c6j/Znoth6IHXcGzvEHJrQ9USy9zb9wISwFpYqt+lyCu+vNLzW4mtXHe
pSDUSUSiEpWc4VyfZTpis/zggkYHfvpnfSHZIt1GFdFYrnDcnNZcE/fowshQoyFkYqkGCcvVT94D
Oj1f/d9t3YMsRsbWg2CeD4ACYn+ppSESJoCR3rqr9NgHXdrScP41Joq6MgqRNHB6hBH2xYeFH9OV
l6BwW475sSsTKvktTsLpKmM/0XfuzjGNCgrNETwoLc4JQYITY5VYB8s1FLnC+AljpOP6/cQv0Xoo
ggo9ww0WAhuGlf92fWUt4Wjy6Of3G9SfG6mo7uF53DqmEVa/2M8kcWJA4/eQsmb4TkxL/KHsWUIL
sre2xI/FUKR0datjXKucDdIVgAzQDi1qhYaz+woaDVXY8j3xRRdmwN6nMOjJafFP4CoghyumBP1j
MkpEP9lnObp41IeHTmvpxPwibdmY8dF7qK0b3LkdHkMX9G8nvcoN4zRMIbZBMfSeL+lTt4bZlR8X
9RVB7ZZ6P3mJqkSpr83w3L2nng5yFndpw7IkLYcQqNOPP89knus7T+fpELEfHfcfJKFdwEK5dl4W
KK9xQxopPx1w08AQHi89bSV/WR5hvd7ojv3C/h50NQQejVgGu8xXsTdnIF/zroiRDxXX6j4MBZmq
PXmcu7rjk619D0LPI6pYzbjprN3IkocTaKkGjtUshnTY8pdr0aJmiMBwiN0UFIXaMJfPUrbKE8ab
9P2SSEW7ms3pG/lUBt9dJ0Rlw2pQoyhPizmzXkJZx/hvowlZYhgNs8Ogz1iXEiJ52hoSWr/LsVeV
qUonwldwP8tdwcUVF9Q7BXui5QCcTh0GUqykNB7ria+ZKK+aIYK1JztvLVBayoufARewzoDbxrX2
TWfIOAunivqM3aGcv3KnEwRggS/OZX6GoHrMG5xNLq4nhvKLnkb0UxOHQ+tSJrtfVjUoMS8rZ9H3
aH3qS2229XzK3oKXQXC+jtgdcDaA2/WqGPRmpgVDOxDYj0OhaNtAh8tVdNgnSuDLi1mYPkulaL0B
zw+c7bUJR6DPR+Rk1QCBuxOrcTHwi0BVPCkzCLao9TQDA0kTkVRliAXE9LYdIf9mRqlo9NEkRwSV
G14724JxlxsJq6+S2TJTsSxOLkOvDzVIYQ4elRutQ3W8Iz4BpsvcrkRFA0zA0wzXLccoDM0ycqj6
NcLuSKQvyM9ui0FfrDg3FRcbiLCX+K2Qf/arVHirjhj5Ckb7SwTNgEfFOJx4rBP8ZAL/DlKYbOfw
dr7D3rux+WqZyg8btsHGDEWbvVljFKBjtNc274tpYLCZ/H3IzQgMfLwtblwSNcnO2DHi5VQ5hvnu
yLTaexQhBlML7E/AsWPUZkMh0WDIEjDDt+Ntbr13UCSt5rW3yxhNqsyZDfsgUegSmW3rwIbNnvAV
zVnpbVF4uYK8T5siu7pku2aQtC7uNN5WgqkQEbc0KOwiZaFJMy+4YOuP1A0hmBtht4hfu1LW0LhO
9De3muZbupj1v5h2CFm9nokYVnQF2Qzzi9Qmcl8ZvQdOyB7+7mAk0cdTC7dqQXyRsPn6OPlfXZJ8
cCWpDz2IO0J9+CESr+UK9X7wRg2g/pZkA/YVjTCk3EuMOAiiPBlyS/TA+8ZQ4i0ujfsMxfixTShX
8OLxM/pyyQbuSzte84m5jUqjha7XthfYBPqYMnAIl7fgJBa4WaKIF0wCx/kBLcGty0FOYrQRxMnZ
PgkkSXzej5Hpt+hKNCzmgZJVYsQ7yO99bT4PRCS4PXDo2l78wQZs2S0A89tr8pVi3ivas+Q9AYwP
PTIclQSgyHpwqk4HCN3T0y5wi+gkxK8sHQytYiJu1XUEGwS0nJdNb2RLJFKx6BGjLzgDLpUEx7AJ
dqIFAcWContfM7jpctlHdOZdFpVPNmTfsSRKcyHzHHNJD+8Ny5N7PNzJea9byJy95ZZzFItOCAAH
aOaYDzeFPsSZmEexEP/IfMlL7M8I11eeYFjAbsnUWV13/PXqV/i18a/7G3ij1UalPTp7GPMymmd/
Y/Gzb51pv06JJbdl9T+ameR2qHpD/NutRHU+CetfSQ5MhvaIdYBI7vyn1cZs/ndc7gKxlZpdGiv1
JQ/IyoHWMrExksRHo2ym/ZMnij9jw0Wlyx96LbNwGP/ZOgILP5S6OqZxObVueTCk9oj+FT1y6JrW
Zdd4C6a43GJ7m0Z0N+25WDA+akk/RDE2caK8dc9eJ/1bmRtvknbg8SMUIlbxwJVQ6YU3CjrbRaz2
dKg2EOmvQs3+WGw9XavuwFuvk4ggfgN4QJ+Qko6mf0pVeg+JYf8eeyWwDmhOfb2cQYneNX0IOGWC
JxkgaMu36KdqT8DIpGNbik97efkXrpzsHLq9lADlVd2q1/ajUavOO0zFrNN8nks9lYpbRUTPC/D7
LGH1/CS4RSEBBoS/uNT7qaUj7XIzR24mdcyO7iiVa0f2TxAq/C71Qu+Y/M7A/swe0jb19ERDLy6a
yXERWlawuzl1YXJOWJB1kWiQtp21qUtKwvuVwL7fBDQWJXn5SBbhorzZNOtOuyEsyHTaR+8jxVaG
YwGkt8Pwoll/kXSQjMiYh2RoYO98/WI+mPGhGCPH/X84dd8jrNppT0f5KQkr+8/nNpteJ5L/NN72
e5C5C/0oEODewTbjzbdE4pXNQSV47J3I/9ZCGi4QGzMpvaVTlU0aCZonGLtAa8gfs7pSmn0TdYK/
MfxXtmJm/eWV1HdD40+dL3Bjsq0YgmAb42/44Z2JYpnzEPK46gROtAKUnZScD385HQ8PvSAu9O02
drpn6YCCKMRtnpu/IlFwkQkz/GzhZOoY7vsOjVqPwawg4ofdrTSBQyjNn3SWNeCKND6ZG/svY/Zk
2X42KdLA64CjVeOvxdKj/vKya+pBz0eJZ99Y/DdGWzOY+QC6pWPeXSqS03zSsulnBVqJMgfFqBZt
XL5tiv/8gKC/g9Ghwjvmtiuasfmd/VZ+eRT/Z5OCmsGYZc1Gi78Xd78r0rcrHr18LhMLmyOIm5MA
hVhRyXr7OI0Rpk6eCXUeppGol3MZA3iHl8SqGwInyJ7Nrb6vqSuBof7We56TsRuNRK3UaL+UpgOT
Gd+ECtsg2DFFlD3x8tn2s/60U0q7mbt9gPZLfIWsn28f/EHydjMN4a61qcBj03RK4nRYdyx4R2e+
EcU8y5UivgEwjoAVIp+3Unk9MeWHA4lH/EMHavR8UF4TGxyx9Kw+PduROIvCoHAxQP8ohUjndWAE
AzoRYYrRlt43AedtszfT2K2u9qjkI0sxYE39TS6Zqm1h4FWGHfZ9m4gtO8xwZ08fJGjp+eiplAZv
+gbLOBoq0rnLJzt8dx6MZ13gT8InU/6McV2bxio3LgOZNzWUvy6Vj6iDwTW336/XEn4FO32sVbdb
pXtth0XC0FPYlpOIRpZBeWuk3L0lglxZgWx+qqV+jH7ZYLIiQzzMUJlGK4wYb/PJ8ockrhGFtL+X
t6iYuw+R8Hb8eXhLMlb/Jk4jx3xlxRCFIlNkL5AykwiA8UYcY/F0msHR3iqRzWx9BgJMnY9+C0BX
kscIDK8s8UEIdEw0lmomdEWNIKfcsbHEiZWHexJOdvW0E8z2s3Vw8k6yrpCoOrbraK2FcW2h/olm
PbyusnfkSldPtGVo70XwOcmWlAgSN/oVc4uU0eqk3eGYLNqAS9CwKuM5jTVmia+dODMqBIkSBJbg
jepexIVoAaoPtmzY1MPZzqYaPcy0QhzQwe6c7NVahKGx6QtZqTuue7jN/FpJW5D0A4tUgnBtkXB4
MDDlDjx1EHt1YRbNVDacjqUvKYxedzW2uElEXb7ArxMauXKtsYO3C2m2wlS35i6DUPhxdrPb3SX9
hf4LNKMsc9a7mDBbvQMxWMoJzlMehA/vGFFZWGhawJ51BQKi3HEkGCpMzGPkBNk74z+i1VErOknh
FxcVdEIxOsWcK8XW20VcotCtrWfQb7IARyqdfq0P97lQmEKSjWt8w6mxrwU9ANuLzXjLFipwvUUP
PpPwZaerUBhtaZjVfxQ6CsALdRAKfW1/8QApyVGwhupFcCtrv6VX623MxIS/cYnYuaZBlwuoz36x
BlUL5OQKuv61PrCTwu1RaICntA6HfBJYBzmfPHmj3EtY7WOjBJXuBCB75teepNZ0+uhkyJl1IECS
JnP01W3BzIizHyjxZ+G1LW+NHl+0/H+ZCw+UVrqczZMcmuqFf6udNMFhRVp3k7iRTBB+gnyZiw4v
jRf3slTVOCoFL/Z65YvqBOQ7ssWMB2l/E33wAj8u71qc8f91xz1VCHnwwh36dxG8flpRjBQrNxEq
XTakIc3WmCZ9HdESpeRF11AW6t8MT6TPbMc8Us7gXM801rk5IP6oOCl5m+q4UjqLwZMo9qzGAT1W
hme5FGA5VeBqEqG4dASiFQDEA+JSZmHLtm9vXO28ZFj5PI6BU4/eAtgFoq1h0YBaKIvyRfghwgbX
btMQhWIftknuFuCJ4f0x1gkgqH+mZdEmvPtqAqxNLq8QF9k2TkdcSSF2PnS1cxObKLl4kT2ISWwo
pukXnXlMpvmKWGZJrPus1KiEisFgyszGo5367ePa3bc7tqlDy6dz2JiLQOsbGFJC5//ABWo9ZnC5
ddAIEi6feH9N6e1X5jxiaxmv0B/0qtYMBvcZk2ZFXH4u+LwyRRN5eqk2EUFddhpFAx6+p0L6S76z
hxZL5ia+W6GDstLXPwusSvRvblSr6xQu+6CnhpLAuQWOEwfO1neRX2RAGpsQNEfiJ4D873QgLpou
gjdBVzi23ulo1BdQ5LE0O2+qLhDqgACb07F7Z96MODzSWTYA/jLF1viS+3NXeZYo1ONhbt+ldVWi
pAPtq6aRvY6KHoeKc+m161XguicxqiZvDzISRY2ff9j7T9GL8UMVFBKdI8d+FTqzR/iUv72zD0s4
01iyq/QyL+uZXaocXesjBFrtPRHJ5DyTBjisMqNFDMtE6s/neAYl8bcr47zWwIcRuZlkaYez26CT
VvRya3grLIpMxz0tu3j1t5C+Xv6LoRnMAormtserDn87TV1XqDjXhAa8yoKZOjcFhIj1m9SYwGFo
tJOvoAtAkEa/crGSYxY5JHuMce5Wk0zDAVQl5nOkQGBI3oFdQv9ich4shxnnPQaWX49NWNGLhbVW
lVoxrm9AT7u82iOUvWNQLP1yAeEp9orC/eBpv6/E4Ah1LJhsQ+398/zIh/O33LbagTl7mZwZNtT4
hxBV/9/46tBW87sZBROd1y2dGhoEOJWZlrJXgJKovrsSE8q8nDENu+kEdG7Uqk7Nl8UDWb2sAkjx
mRyyJMGfvGJJn7zVfWM4X3qCwlG9mNV1yfEDaSfpKZlyTj23moP/q4N2IKwM24C6f0Gdo6xdhNmt
v6iHzANoveEh4WAag+wMUMEDmqqk7/tHCpotixHZxU5AI1WDwnXRNlEToaKgzhlBt9lntXXusvcx
e52/Zf4J2Vy4lR36Y2Mhzhyj/dx+CVDoHLF8HdlubP1ll7KpaLk4Tfklm9M9G/+LCRu4ATUJRQ3z
Bhy2ArGTPgOFzdbQ6QAZlRxFd1eC6EPByze525FJmtf4eoOoxkJ0Ml2pn0TXFo3aBHliuVpm27Vq
9ShjVIy0WcXsCK2uroWHhCbkXXjfxjBSwRCqvGSVHP4j3RwG+9/AiYjhBuySHIZ1FmgZYeC/Ed10
TNNfMDdv4ZkWbcJohTMQYltBZRZNkkhTUQzWJGuZDf6jV8qNVxLkEmqxM5iTjcZBiWKPdXwGYtJe
ui+Ec5/9rLNjeIhE8NLLt+OC8wRxytAl5cYAw1ua8goFspZPdNu5Mf+2S5oJreoqJDO489iHYm67
+n4jaKTkahNoJzLU2iaYgDo/Vv/cCXx/UhONvILLXqYIqIMjGpnYYNCrINUjIov1heGZYw3DuR0M
9O808q5Yr3fZcsEdWo3DskocWUED03gP/6Nqqic7fDrMobWihih/sGIhDdMoH+AomW9PuVxWAZxz
HRQoQU2UdirMUG3OndikTgwdwcFydJTdbB2gM+/1o/oTiYuvsx3r8q4BAV7smB/GZXx1E06pxVG+
4LRoTr+tu3lw59oIt+l42Uzg57NwgGzJNFKpVpkujVJw+kxW7pUg1KBjfFutrjJqEkgxnwnEVnw7
eobHqSU4lAjK14kWi3bGy6y4MABu3hXG0swSgKVU2Rh4x5nEqMLQ79pDgzGjCGK54tWlE3f10JSV
v1LsI9zx/8PAQylrCi6JBuXh/SmwEuVQv9D+ndfA2TRHJRIxQ/8eiJsAysQS1oayFCSUzzgPDmvu
zXJLsnEMkvMPMmKHZNcZJlmf7QvzdOPVJMfxx0RqJKHi1Xy3+t3pLjE2LvlJzRvi916E9Hg6Zr0p
GWcjcmzlRDwPQ7ZEtESqiXei1+3BJBSAYZXX19GHVIveF9JcaFVRAMa16zz6fi3gst8ZIYI9FLO6
dN3V/Ecv3suqImjn+vLGj+//oJ/OuHsLyj4oTxYFGgrmg6IMAEWCeDA0qIoXqyPnwOwjPYhm1FwR
ll8KefnaGotJSSmzvLTgfP83NW7jrXvBohU2FgcQ7L/UMwsp063Rw+Dk5Lu79cv1Og+aSR5z40eK
08NdCeu45lwovPfyjF8GjBxCPhQ7nuYzXYp4rKvyThuQEWmZu3U1/l09/J0UJa930LgY6xqHXazv
8FUaJIH0sKiddbYjq5GfiKgkTe6g+TumouSG8mFTjhEcWJy2/xHZacfVGabfauXa7Y3twxWUu+z1
rdxAdRCCb5/OWWZyjwchngcxu4j2arZESKwrJTLLUplk1FstxGL32m8M/raXpFn5p4XJ6VI7QMsG
g76R6Kit+bToX/isQLI7lGo1DTAStZ2ca4atyQDZ9bAYocE5uz82gW+HrpAV21qaBu4x8QCb4eCY
Dc/jmJq9go0eTIJmedwZfbzCSOmVd6O1UaQs21EXg36vtYFxl4RVrvE0F9o+zJ7N1oLpWIstC8rR
P6XfrlvikLVjnjlsN78oEkjA79r7zklSxUh45oY0DjU9k0cQd26TqjG9EIF8rOQ8B0lAngtITpZK
gW9SKfbyDSkuDqSUfZWjgWROEFlhMy5V27U6RtutJa52p5c0uXU3SyyL2fBCQQEeO82dyxMVFFLL
UG9AW33S4TvMZbEiTCKHxgnaaWEQ0mb1gnToVAc0jIgNWpn0SDM3GZQxDeJlV+x7N/5BChVM7ii7
4dkW9B/Q43JAx9otALxe2G5UViNcUFG12O7bDa1H8zD/WTlKkJk+oo6Dd7YR5MSZiLFDJojLTgD5
IdxTMFUr3xHguazEO76E6vPj/rCze/bWpFNqoh2cUyCpaTKIOqxhjSUj3IIScpIc1AGWjQsjyR1W
BI3mkJyG6P6y8mrvi4BJ3Rr+32C5wLvLzUeel7sN/UpC4SkwfKLiq71vjQhVZVIUJcDJvVw1KywQ
nm+tZ39r4Kk8pxXOk46/RrQV7Z4EKPu4SB+vBaZ+Pj1+VvUFqIUxg2A9uNKmvFJRIhM0DFTNZfI3
n3y5exQfmlXzgXP2scOnUf7LxxCZEr7HvZajJeVRLPHkv+Zh6Ithakb9DfD5SfdPet//P2i4GrpT
hFm23MgNyqJK3xkuHdwclOog2jwWfaM4SwL4MJ5Lc2dWhb9gnWqV0n+UGRbqhHTOtc6BLH2e+Pj4
euEoWxm4KcEhx4t9Smc9+hvQ1AIaQiMoZOaTLm6+1YPklvu+8eLnHif7Z+PqsxDtcxFF4OjEC+Ez
hOqircLXTKnUsMKqyldzOSRvXPQhI/yWgQTatCOs8bVxABAmTIHyNGDWUOybYZ3yXuc5AYDrB7KQ
0X7U+k72ai10BD0DhjqgKe9Kud4EljKHPelA750Pcs+ZSIb06nR2Utf9SrAXlg2LTtFR2zDwUa9m
n/ZXKABkLnPUGHUhRF1cfkpBH1QzSjy1Va16e0bkHQoyvc/clm7k8wLNgp+1yIgspn9dvItLhFJP
f+W/UA911fJgR3aPmE4tC0ul/r3LKgi+ofI5XfkKUeLjFoNNuRWSk8efOB+/VRQgPGNwDAXR3B9Y
VnAkPw/9AIgJ5ZcZEfyWx+kBJFQ21gnWoJF3rOPwVrZN8thygkur4l0c9e8g51zHJfq2v/wTCghf
0pxKErDiexyS0ktmip7PcntAseFDCVTkL0s2u176C3BnFL8OIYFeGej/qlIGd+a0VNNVLf76IB6D
ifOQQJMtmJtiVEPvmHGk4y4sV/7YsEU/gQjNaUx5Pd58iLekGZLtAwl1bA6WDYXO4OZKlNA2xHDw
p3YIhVJMWZ6ae3eVOsXNfVu3rtgYgsj9iOQU6yZMRUU1ZGyeGQ4Zf73touXZx7sq580T2LeU36C3
eCNC6d626OnJLKwkAbaOoBI13pe/IpeuUEvDJifF1bYdM6REHSxNvoJ2cjw7TxGrbIC/j8gSEPR8
70Le/DkL4ZAE+lY7cbl1Yy2/jEeM169cftzKmfMn6kg3gQFCtmXDhLLtFfd0ZzZUjOrdFSpK0GZu
QTzEdSyKeJm2Ph1+H4xTq/xmXC6bVJ+ypYFsnB5C0P6rVXxOffQhaYPFf3KGKwgVHjakY10TbZSX
0nl0GkEoYqGLZmMmfuOUcIZVYAyE/05Vf4RvmKj2CElBoKYU8ItMmsBvUAD0zBq1ziDT5ezwekZF
79ScBooM0EHjXuDqastf0VhiHpKlxyyGIEqTMCFatNbTpsLc5op/S20TDYPhCNNPXqD9+zYPIgem
t/dvBOOHsfo5FCaUJHq30CO52Hi1VxXTh7zgOh2SzaSlu6h5S3N9PPigmPuDDijyAm+W+zDb0/nG
/Uqle3Fpey/m6qf80boRYH+PT669oENFf5Av48T37QNyfySO14GvYI42eynJhRtvs8AGsnM2b26t
GwH7CvQcZo2YTW9RDVJRnEQZcsTjdczrcBcNIV+56dMtbxDPVcM84F/kHRlb0L+FRVBM4n0AmhXe
cULj1WjVJV/eHqVdqXvY3IUl7tDqz2zTrwHGxPB6p2bpnRRHGIIYrGIjl5O5e+9iCR4iU1y7OKQz
41CT7bSxZ+mLrm6p23+gNG3bqDF1EUWbROOfuDlq3YegAuNE0UwFpDWqwFggCgwOaHOyTrqEQPMo
N+oY2LclUO0htdDiyebz55im5DM8mqir1gT2GDKfRS2SwrhrXtSEAfTYuE90nz6ndC6idOUbEGEX
OTSjDhxILzmqbLBtfsBIhPxKA1cB8yXsyMv+y/IHploHnix/mCcB2BX7BQUwewJ2DUmtmC1VdjL+
ey5CneixDmpWjDF6+LCCMypsj0uYWjTmNngaAIfJEulgS1iscGvKKZS+rdFcvCVOwaM61a/JFjaU
X6BDOQIhs0/JiWJ3MGhWE4FlAKOGOffMXU5YWGaHAdt5G0PKh5DizeH4NUavS9o6+F3TgzgPcOug
c+Fc5lPdxw+nmWOGxhJPCoVj4fpFPGTk99dKWpUtA8PBFdDSuZq6SXFIRrgpreLK7Ws7etlClj7b
JyLrgt/UDctnfWYts7qoaNcuUJAWWcUQXmBYE8gNdbkCFN2cbGYqkvvj7fUd7wW0WpXHijGG5TA9
dBDeaKEyPYuXXce+5uj2Nb7WNm+ZWbfYQjENIvkX5NZoMgu0aDkoIjV5df9D6YzGUgfG2JuQxTqN
k+cj3n42Lc7U6++c7TGDeNGYLUhoy1nEV9OZrsMkM+18/EKVpOEg0v521HXOqf+TVTTgmxK9XFbk
/rGstOz0tRa+ljvMZDhaRHH8GDbfSGfj6+RPTs52eYinAAOU8aVTtmEilIvsJYMhEtOHi4pqBMHZ
IilEcFFX42qVmtewLhXeF1IOZ5T3NsLasITKWlZ3lRxvzqpp0gZKp4d92f08fdwCeIIEUKnFhApv
tyupfDvYj83dzGUUz/SBygYBgp38CKIcEiKhkZx/OGy++nG/UWYr/rgskJwy+9BAIIQDbxtcEVh7
bwnkwlWjNOGV9fTxFqXlaUgjzuIEa/U8wlgfpaM5RoB5OfMzfGRLdC0kxwOHwQPST3QJYlZe96Df
uG2eYQNxLd9aMnNWUFh0ITWxOKsnFNpm0Z5RqT/6yOxYLB+NU6SrhSMenMPbPa8ezzhwgMKQB3w7
F4QITu9zgeMYz/rAZo46pJwuz8ZWj5Ef9lC7BlmmXc7ExAoOH3fvoHYhbRbX5E6I/7SXiJmRLo3p
IPotkzceldva8y4vwWRtS/rqroAag0QuNtOUxbzUPNeP70yT52oOCgghSBD2slzXSmS228WjK7Bf
NVrN1GJFZJbeDejY6sZNSONSTYkwLfuc7XB2FhefI81eIBZpYYWce/+5/Ymn9+ltVLCxphAtGvgR
Ts9ovN/4ljxhgvg6qG5PBv+bjZNmxLb5j/FbqvDRUean9eFQGJyVHivSlaUsOwAeJD3fJKQrs9qT
Sbz7wWB9Lilk2dZpVVtS5AZZtMetcf8MvVrdftwEY3iGhlFjaC9o7e4bEFNCANzvHDbQXKo5ZpgA
Rt3JglpgQ8lb43Rh0RfRza1UKf8w6QEij6XQY6xahiGQMfRc5aLDThop4MwmYcqbxiEYsRa8qlaO
8gnzYO+T7Vl7/JReYDsMY9s2zb6Ydeh6igqzNYNeEik9x4q9TmhB5n0CfatQetRUXiYBIXeUKtZh
Zq11k+CNs9PJ654eBMdeAT4P3W/YlU9wi/3DiJ0BLSM8g98St95boVEoMMxUPecxBpnc9IPIUAXZ
G+k1an1JOY1jX6R1J3yJnvRGDmClo0w7l72xAOtopwBiwN4yYO9Vg+3h8Uz5VuiVD1jC4JG+zquO
mxH1+RJNROWsUoEQndlFgpe3ppXJ8SKerASgXRIUAlyi11vJxv+FHIOYcVTE9bVXT1rO526uevRH
z9FQGmMOJjrAwWijuBUcBo0SAbpvvK/vecpgwHu8IQhj1ayojEmYFHCEvS+RP7YKICFARc421914
LDkQ6KO7xWvmHJUnADtfS3vf9uToQ56Sgm12+p0AaGyP384SX26kL55iGe27AP51bzGvBeFjOxe9
k0BgyrW9PSFZaGyAUwQREyVaAqDXwrxmS+wTsEdlaLqB2x8Liyp/OFPMvSetQgDaZ5ujajJz3Nb7
/ecE4zvDqh5Kc8KNna6nLa59DI3ahKqVXEL2qIxUR3xhqf8xTsolO5i8PADP5yvFBkajJ33DEjcw
13+KGUm0i7Ll/Hj0uPmHMNd08+L/xxEvZRizXgq0rBOzkFmfR1TVkcvBmWguYIXu6IX3ojjfyvBi
UsLDq1wj/5I2FSJH/oa+iyOd3tqghNpQSBcQerpjX+cmlbnCjiKFeJPCH1DmY/OXIQ8LXk+e2rcu
sKtQPDMSxwebV5BCRNew1Z538aX/wCyZw2s+dRO9stuTZx650tuCLDJu6zr6R5isvVx7MRfpzwMd
IGNtL0N41NX8A1Vk4aMP0MC4BGUSBf+4twk8H6TCRY83wRQw+WDHZc4jqsQ1jmHuIP0UWm4PV/5i
AIPJ/GuC3kMsv13EQKXjkGrdkX03EhYUBdrqYnvGAWjiUkyPLe7J+fXQZ6TErtVVeGJI/MN9e3wO
CL7RUe4WoXIszRQaVmSga+hJDS58ZJ2eV9MItIqsP5C3rYi52Bc5MXv7B7+BSpFq8g3SZzs4SF0V
8bGxiT8rSAZvDkY7tlfCIPOpo8ujuNVgz9hACPbi8ro2e8oraJ1hg5nigZOstDKj9GmoDYuVv9yL
Osjg18MiAYbDp8UyDtcstDn7VuNPWIsZMQmvBcNMcCgJszGjy66/qXivZveO8xJGwChPEhfaypIp
obvPgIlztjEvgrbq70LAmxllWMWRumo2XEeeG3QOULl3nw0hBE2zXOphjntuO4RD6FZPiYMdYzvF
GmXRkBkHpNTWXBmnwG98+adaJ7GZkbsOfCnmxbHXZER8k+TdMt4EitZlxyP1jbUiFGJfCNBvHVdh
5RNDrzjwf7KFJwPF50xPYiyp133z5xmODO0tMSCD5KLfvmf/5X6XcL5S92n2tjc79GwH7kYXy/zG
+jW6E3+1pHG2ztlKTJuEnO43xOURwCgxtpEZlybsd/56026hiNETJtzwkyPxYeUleuJosbEN0osv
joSwyy6IX0emR6rme4tEm4gX6Zw4IgRk+pe8H34NxrBdCerTCA5vvGEs+uk4UWB0vtPmy+N6iZiy
qmWUDDvnfh2iKybWKv/OlbCZ8D5SGFjVQ5pzDhcc+LE6Eyp/kIJ3XAwvbf9Lq/Pjsc26k3DaI50W
4tbrJ+zBhwenTF9lrpYsc6AVpxLVUKSSe5HR5FT0EZwX2g+IwRRCfE86cXymtlIXyY/En7Tb0AAY
xT44V3cWbBTCeZr22l9YiFzGGc+t8bu4TnnBWUdGv07e6lJjctzq3jFYjJA7yAhYZbEjlmpRf+G/
CRpt+AwMjmGXPKBZkIver7nLrK3/t7YN0ptNablad1axx0iEP56vxGfOhtd/yc9M5ZfQHM5muiDU
WoO7c+GEpgekY+JjAFIc+DSn6uE2m+/LlMRxOksdeHoQwh0f9ctiWk9LmqKMlcuTOO6tcJKmDMvy
QXEG7FB6vT4FWoxac9+ah5VGIGQjAd6G1gUwiyB6lYPY3uiKmwtMN36slVfFKQZucNdJCAzVWqED
2dZ59g5Qa2lzKhPtXIypmkhGBphQJixlA79CJFwhQT8CNeJR9eHJiRBhJ47fP+sooCs557hj7OTC
L7j9612ERNWaILEGuEYZXvgR/Oifc4o1Ro+PlT2HwngEjWJqF5ZeVvrewhltlbaSkiGINvoI2gKT
vu+EE173pAnwHcBhqAs1avBUtKfYJ7J90860BfS/lqLI/DF64F7S3wgxmXV7p5ETRp5xS6FifqQN
MVvQ+iIzoU4uNCuZlBCghWz8r2qsDmNA1AdhuOfurzPD50pIYQsn2CKCm73nHA7LTbki0Axtazly
O89tiy5qYndAhXlfM9HiEr+29dQi1yBXLoftbA5mhnbbV1AJmIy6btdFIeL0mnZ9cEITDS9ByunE
di16lrhFBIERX4NBkXgWgBbqCw7kM7PD+CAQjjIUlXT2d6neljyTmBBI4wr1zxZ7d8hwxjZ9OFBl
D0R6kFKsg9W+73+SCKZtAe0laOxueHlCatw87H3fw/m8CWamA3m1xXVweSK2nm+GVSH2XAyM4pND
Ygoh8Qjgtj0W/diQqKC0bCE7HUW7jxIfKsB0MgNMAfeIDDAnLrTkd3G1NIwTI4PQ6hwAU+yfvDmW
cYSAQCHvVXYdnAz2uxV3VmVq/zUZyL9P/160t+1rkW5RTlycJI7HoxO0+Gg6iipheeSmFoal79c+
rM6j/hRNrf4glAueP/gWkNCjnq50Jfj833NUs33g4aqBehRVtqTneyObWs2rWA3Vi0RyV4JLdGkT
5oyxGRhpgetxQg+7BD7qApS8LPi3jcrEqs99V97Zy1JWswhm5YJri46Bf5s1UvsFpDxJNiJNyCUW
iBk4Qa41Ghs0s/urGIdc5e1SZJ9TJoBruVCINxB4ylBA4oiuSppmWI43rf37v0RGXWbYB2sA5qVp
kKLew95TV2slHGDbuACMYfbhbXay2K9HniAvgEum82zaiqv/ZmfjxCcDd6VIhQIdIoH7hlVL8yG3
wXQFXO0eMxhWjtoV+Ma+Cm8xxtwTkg1jP9OyvnGuvnKaIw7glYQDGsngM2a9bStGtd20VEoex3aT
A0sC+9/3omxVE8uQemSpETiRwXhlA3tcFS9/JKEyXJ1n2Rf/vznywOzXuifI9mEjr7rpP7E+2M6X
+gofBhwm5epOvQXbJnRGR8sMbrz/4rwFBy0/VYP+8sxyKyCg5V833UIg9nbzi0aFy8M4KRS1jVz9
4bfg4G0ki5ezg4iuSY96LAPs23wBMzP8wDRtA6WBcACAku2jwd6shIRvnG6Q888lj9QehRWiVUJi
xo57dudwNNN/AXVwKbb60XEHAnG8RSA5RV0tO1USXnRwyJEmzoso4ewQM+1hiNUSujbbHW+e37kp
zi3n0/Y5BrwP1sK376bLc3b2ElFtwn34PJIAH8cZIvnfUbO8CIpfz3i0fVfVijwgMkfozpXMsiFs
jrIFZSAUNOI2w6bqQ+UfBTrM8BFQtL/ooJfn9J8d/OFhh+lMLIzSKiBJulQpmtiODTlZFAgbYEME
iUB/oKhrBEKNRSBZJIQXfPyjd/lGBv7gFN9iYuNST1sO5VqwvaXWQIdq9JivHTVChzJsBsBsai2O
37GRmCGHf/QNJrVekbWxjXnVZO3pvsss+HrZwhYNyYB+K2F1278SJ594LSPHoG0zFor0bLDWAox9
RSCA6xp2g3KKWjrfaVn0iYFKgBz2ZnwyTKhvi+UgWowlHsbxDGM7Olfm80XsWdd/AyStO/aeIHdA
V//TOb8fRiIu97Fuds4pifwi33Z2P4agwLOJwK3rcPDlP22ynDRbypfcl8/3NOH0FRPSbESno/XH
A7P7Z61AEuPGB4a7cxHN8dwHuVJ4DAH+2AfUw2mEaWGl81zER6twKsVRmiaEH+neg59CRWZcOqwu
iBdKhynTlCmN8jaq14o0JC4D3j+CYB8yNpOJEqHKl/AIB1sEIb3s0DcVzfcolO7WNSuLBPuNe4Vy
j32TqTH+R6a95Ie484W+QlJR5RhbwT1Mi3n5/karuDt4VF4ErlvZqeDIDWjmbxfMQ9BmVLFOUQHD
882JXDXmHwo2GYQqhAr/ZBCcKA08xHRUOdrA2+vh6GQoCSnoevVZQ3B/DXUbsf2Py+VzFrF9M5EN
UT1T4SZLmBMrD7RkDMMmeBn7K+UYYReJ+O+GsSCf60/R2T/49bxJBzYFdNJE3H9lU/Mp+hZmEZY8
z7sx5+PCqQ8elZO8iJEDgUKuyFEFx2j4+c3e5iHxUOCxxN34P/UH05zPndo+AVvHtX5bte4fIVO3
jTwbQ7t+w/SD5ODMMjx1EE6P6hdzOqXghSZguFNofR9LPQmTQ3oa3PrBobpB7GEHqClNwHj2zvl5
ZsaWAPElZp0+bcwCnxqGtolk07B/9Hge0dDi5TOgqrkb3xwQaOepRieNK/OTtinMxjvZs2q3Crvg
Z2FkFY43rd/aAhzOd2pEGxIl+8AW+Z89rEFBEod5EBV+F8Q+VKTgxbkx6PG9OEehHTcJxyh/yXNJ
RAyrlluHD0/EWgqkYYH2cUw41UPW2vMIxz9mD6wkPUQyzFXM891/q3sVXPzR6pIhusHIUVzqFI0w
FGZoXQFU9IA8CP10s7J6hDMzohoA0vNAmJiEt0I9VpoTXHt+ZLzzBTHy/a95BMS1WiArU+i7Gykk
Z5HBVku6BdCPzChuCigzaCdhUxI/qLfLP90enU8HH+jhLmy/T9FcnugtjykG/Z5qzorUrYhHlRX7
5Jzu4vidZbwPOVUfp06GVVNBZWcyv1ragHEVWc5Sh3qCBWaKGjxhmKf6b462Xjx2r4fIbd49slEr
Av4fs5pLq2aaiIoP47o9OnWl8Srf/kwuxwLT5L9fG9b2ew/RDmrsyA1wNCvIWUZ0X3Rx7dm8Mt2M
rRDTp3NIKj5GKe5LKG/TIe4unJVCixCTbRZ6RVex0PUPW0Bs0QNz+iuifkywmMfZeHZMNawtZVlR
5ZvZse/JZ6hEDDhfxxji/Mic4Az87K86E5iwuLyBGLJQhwOmusaZ/+OE+kecZ6DLDoypsMRDA5ZV
bHFney3DuC0w5vYAzCaBXWGoLNZbJv4xoOSLe8bUuCa4UcOb9pedrFdKYfxonUP3Ye6zscYt+gOF
iPlH98z79hlCgse5k6S8Xnm+AjCRWslcg6qj9I1wHVUOmLgmnmGXysGH0+OL3WgTx7CVXI0kcRxu
dirCUrWDl1a38YedPuFy6TsqMGYUM1DWdnk2s8ZlHZwWWP7abqxbWKt3htYWwlhxyZQ8YQLt3+C3
84msXY5m3eXSL5jsoYQxneF4qdeqyDvQ6aqlCxfAFoAzqwmV/kSjv21hYrG0R872i+A/MnDiY76+
/A6E54tfxZuZlyYttJU4c4OQCamW5GIjUDTf1dA3MPVz5GTY3If7l4D793NcL0Rimb/ggiam9w1o
151y3xp7S9kfbOWaqbKHE4ESUhrUYI1wtApo0SVbuWWesm3r+mqib6lUaBlD0PRcBkE8+PCfMlFB
xFruE8P34aZbr53V4raA1v79lPHJ1yj1MVKkPjGaTNTh7AXrIVmph0pmuFMhp9Br3r+y12sQ4kIV
QIjZDO84Yd6GDUNG/Yd3hUwTyTWnQ7Y9HlYN3fio4p8wYCb5PEMBjucY+8G6WdLYUzlIuORCe9b9
vOACnYW4CmXuRNhOlFMRop8OdRFnOemUSYtMyopqRJkN8M65GLVL7Y8b0kKBUhuB+7PE2HaTOS3Y
yBvRxEPXqhB19IGrw2JV31lBbiidgQjTswrCNA6pn6CgFH/EksrE2hiu86A9zcgXfsWsTgkdgg8t
Y1sG5DTE+7zWg0wjbHDtcnnm3NFnP50op2b1zURc98k2Jm0RIrXNS+xT24yCuiAPfm6DK5htLGyd
t+IsSW+pPVGXxgyJVAbo+UZR74mvWiHcgIlNscQaRLVZLEt/97i9geUOIlychCJdirZVoX5yCnQR
muiLGiOV13pgTXYCMPrhVT50lUlyerv8peNqnD6asotRnshzvRjbGMIf6BIcJx63nRFWZkwHLcNR
/Nn56mSqHGVBW9RmOWJmtIngpw1/OZ/boZ5y3r53a+sjCerPcXZVaLJfN/2e2Z0ErGRQF1eJnizV
aXOe45B3149krzJ1rOLslomV96XevluqqsMwIlUVEN5fT0Jdw6zGmsbFu6V9OxnFGZS81IOcGDaK
b+u6rWAC1VeP5yKVCjJ/kqaEFZgHkecPBt+9HnEaIrsALmeVl7CWYJZTqV1nd9R3UpE6FRPw6poF
aSC3obO/Kyb/FHgQ2zK1b6mM9Uqg2upcDA8sp85MGZn1h4x++IoSpARiY1kX7CzovpZbJPs5+EGW
VDbTe2d8jCjjR3ma/28Nt8fcZKvmr2oDEkJMUPqe23LjpwMqKi0frU8AUdoEbe9/fN9EOL/lxM9c
7yDoRHgjZHk43q9deDIhzRop/8T9kwNOM588v8icPqKmmvVIWNU4kj5OLqRTrqFh+LFpLf0qK/JU
kNZAcvLkrVzDrkrWxN3xqBMNLlgtjMFjfp2PVoBWDEen7kUZG9cB9vpnW8u1OX+Khj1SrtpfDrIO
9jsvmY8dfzUabiRlZOtgpQOt6MP/bTatSD9tzi4nsnG0dbpLPGp9OqtoZ7wv/KdFFhM3KHHDCg7p
A9i2W6OYuV2XKdO83YAlIuJmuH9z+jfZgXQjS3rfOa5SwaMddv/D5sqEgZexbLTf4yb+qF7uDXzZ
km/ddWhZCOKzLK2EFpuBLJXItDTbE1kjYVMP8ftsdfsiZgrIoX1ZmG7PfCn+LDvwOWgTF1xCd56l
e/HwE78FISCDOgkpKlM4plrOBCxfqf9nVNEPMII1ksEDrnkZ3Fqxp5xWCM6zZ5xn8lTvinMaM33s
SrWO1ZLg5oNnupyRyjzAx3GGFY2qNsVchZdRhSRh8thL2Jz/jkIcC/lEo9Pwrg+Ogt/4uP0dhRjm
jba5PX8/y5vEqP01QTJmlr4CjKU9EcdxxYFBVagIIPPlT2vioJne8cMhDPga2Yr3/SYhvdqtl1bj
KwgXTavmlnuX1YyjlexKic1JIy5peJ7oSCiGsa25narTqjX67a/oD9UYw58ejOYVncrU6ot4YxFp
Km49TQSqgD+fmmctoRHJ+MLJifF5420ugti3OA5Y9gTMUOhKya8QJfheXSGFDPLmYzlZ7IMRcilE
t8kx0/k7CjA3w0luakV9HaVYc3nyznAfkq7N7lEdMiBE/TLWtOyp7ZFVGpmuE7or5/b9M1q7l9Oi
95zx8Lh1eMy70VoW11Toix/Bh61nNzJnqTUlltFYtd0cSNzC71m9VYgQGkILo+AZtdqL7qIlojBn
yv+mFZWRlCKLYNNpMTqAtNVwjsR3HPGDSqU6acbCDqToGvnY4wahkM2WLsc/hXhpGzCKqh2rFZLW
6kLE7p1Ma2RvIy0m3JvCkzN/FxlJfLaaMEUatN1QOq2NRYemnUUL1zQkSym78TcHoDyDTTvQdYVb
VcqurK5K6B/mDEV3Y/WcmjeNQsWbGeTEhJMerIKNtlqCrhPYhmkxZB6O+sAHz5dYpe0dSTKd55rm
I/Ki9lpfgkKArKHvnHOu3VklcGVdnxptp+xujUAAImji/CoJhL8AsPccnIUVEU8iVJYuNx3z7OOk
WgwW7bkrhG6zkLQlajGgTVS+6j19bIDkZm2wQXjvAWbn0JhyBPecWYF48xyFwl9M+t58owekE0GZ
IZ4LFV8H0wve6HSKLLQxB1rXDB9nebV0bR8U+EF4k6cv49EnIzF4JgMhOrFdbG/sssrZjaEZ82Zn
vO5A5ApQy9GBD4Y8/rUQ7Ab3Ck6FIEH9aWZz/9nfVjF7eZQYlVUPNouGQQRmZGY9LQHd1UeesDr4
JQP3jE8kRdbUCvLRaojeQvUo6LX7PmrQnFK53wHx5O/3lRD13Vc9G6q9Mw3+Lk1YINhFRhuqp1VQ
hP4LN/zcUGtsunrdKgqcfazJ64MgaP9J4LdrfaViAo/GYTCzGqfFYzaXPS3XBWCX5rFQdl5DN4iT
k9z/q2AsNT18ZvfImWVfxUUdUYwXcs6X8tDbAIOnKFbgYst7iAyytIzxgDoT996b8n2CDf3XJuoS
DVOuWb4P4aAZ0DW1GUpGpiFeG0cOI3GiQfC1VKZ7HOaFiXBKVByg+1vXlNMzf8QqHVAthFJ7sYpi
VzlmXqmV+FLs9lwfurvg/BrkihGJgW77QfF6M7j3rzBQXoPZDQIHnUhMftWmK4CEYXot6fUSgQo+
X285kbf3PhLG0OI//8WcjmLGENIsLp2IPetghcVUbYiWH19by77T9jFwmU9rCEImyAk2b0EAhZC0
V/65GOZJqKI6y0j+GuFqY6dkOgG09KKo7UxC9q7CJLP0ABkoAR+GtbogonVZl0OWIbC5jOMognxa
iLxMvX7IC6f0OD0x0aw3v70ZUwAAl537FNROr8tsuDjh5NtjIhaXxMvps431wdkZQOgF0DX3GdPX
nPG4BMPrxSPcK3jUrWn3v/B4bZjUE1YU3G8YQrPVIFf5wQKOESdzblAfGVZ0YkjDc3b4k7AMAH3l
l7BGyeBUk9Pjyc3Mc+hvfHxY2JsMiggmqEc6ruTOIXAnRu2IRPxrAaFrxh8/ZJtrJ0/eERku10dQ
w/JZdHPNtZhBLs/jvpqK6LX+I0AlhHhMpF7aQ5Fwj51ZpFOfwv6B1JCbEJzWduLmNDI86WNwc4sl
SCIeqT9HOiF++aIfjrMfNG/50MXLQz74C3X+BLKFdpUmndh9oexnSmKoNoOMFGxNIc0vAQhwJXBi
F0idIMPTua7zfoIWpuf2eMfwvk3YQsM7HdqRufqvZxPTIkzA4JcLYtxAJsVP/idgLE+NnYbRetA0
CgGO0T571QVeIdsFEOk/5vXvbvH9RXXYTNmkoaKL2gx78pfTmCLd2IWmrZmXM4BxDLVIoCdYPXpu
QPrtSxKiK4TS8CmHbAbVHnN+15wzvo5LUc7iXz0+vGF/D9PTGBasEAfx7CYhpC5SJFTVmJ+EsI7S
wRmvw7vwxljbX3+gOqv2IWPhfNRkUuE+tN2QJqhjZ7uwK34HEy4C7S30g1iVOq55lccrhQDsVF+s
TFj7g5VAfoAyZ4w8p+URtm3CwrlZmIPDenjkJ5sRZYZ8QHlMDRtXhgPXgUfXE9NnHx/1CS0V75+5
sl2PzZRPFAFaJEpI/9QB/mBo9dRXJnY9QZRlEFzLNKELHCekjUix2o22Z9udYmFaiCmZqyVkZDi/
ypGbvYgwPStdmqhvskVFulI2pcn+WUIHjAw28Okv9ekBgMr+zJ8XpvG7yPntyq746oKF/jk+2133
jvPgw/6NTLevzSumKznEis6yHo2IriXyN26Cv5LGutK0xmoWgRxH5NN4zlaNDbFxEKUgXriTGExC
NrxA2eObeb/d3uWdF76Wnnyf9hcGOtrv1hTzxY1Ucboy2ueSTrN7QHy+iUR0bwoYLcJaLHir9ota
aVSDznKVl7D+WxpRlhDg5oZHJBmbNxN43TFfPOssDMqEV/yGoWJ6bzLfATDOSy+MLKFcsc4bm5xc
XSAVU2iYLUG5Gg+I24M/Nqj2PAYj/8dB8ByAdaSZge+HwQQ45k3mhY8+D9Cn8juuiPikaN3KMl5P
jBgasghv6st9l31kLIL9bfqRf2EuXL45pZiA/mnPJW26RxI8GfjMrDJEpboOtPlUBcnQmN+YNI/Q
I2VakN7EnuIW6nwOwXKzdHH/fmf8ru4Hp99XvNNHlN5wKt7OTBgz5jTxUn/rcDw5XOGiwCTUUY0F
JzrC3COrCko/O48IwrupBwtz07VusaZMumd/xhZW9cDGR68OpegWf1SUYOSy5ojOhnabCxPbeqgk
x+rKNxrTh3SE2DPBzta7MQv0ctK7RjpCusMGzzT96elXYGQUhNG1h9DHLAiuiL+VguB08I9ai/wQ
yRgotQa/xeuDYoftetpQxHa1RiFBdwL2gkTvm67NLhtvCrAgb//UR7aj+gZkjM1tLNbDJ3D6yuEH
zRA8HWJlfctH6YywFfSuNvDK9NqNGvd7QCjAAcXKR5N1ZyU2Zb4pKlBS5U0C62+JUHv6v/58g2GT
k5BFJNOrNdU4fXzs44Ll+RipgRZLRykvaBkzu1y80lBGXlIBPfPTaVIh/zWam51NU58Jc028BkNG
nKJTF/1wq3C8bvPDOiQGDzD4BbubQ5zPd3uet/DTNAQsWcQhDSw7SMdilWyi2MWNGaAIvRAIkgKU
G4i10tAzJbbdX/v4FtBKZY1PsVcio+7k9ouXCwS7O13NWhWDpKHIAFE9g57n/Z6ML8a6IT8TKvju
tqn8m73dMeXTrXJgSy3XqbNfBrTnAWTx3dNEGW3sFS4oXsbIl1W4OXl1/LC1UmK/+fHgF3KOXlWT
R6bmY7qVsPCG03z3uY3Vd3DBMetS+xmYDoEaMsD3N/E5CajZb0vYA1Denf3ctuI1QPgzMlArn0J6
Kt1++mRgW0xdirhgJD569sCE1InHWPOi1/jyrE9Cds0YiVglyrQNmwcmoX7tHusZwNkA9/vgMDiY
D5mO2VPGx9LIbI8w8SQWbE1JXHdP8RdtVRk6aZ3zi07D7RuTZkFYoHESH/cz7kyfKKFuRtoQg3KG
jwhQH/AgoqiBBlRcKG0VT9JJh9En6q6wvViN9diAGiuA/m9IQeUfCYnYTwuTA8G9L30HjNh5H/aN
WEBM24ONVdsjTi48V3r6lkUoP7tECHbI3fyTQWAwfy+MN4L/iko/nNVbpUckbybKDNXaiUZx34m0
1NgPy3La3XLp9ez0mmO6lDEuL7l/+Kr+kjbqvPnP0sZQFvqIQFMk+et9WhTnDh7d/cOPNXXnBA/H
3kXesobqVaKTha1tdjrxgrjaxQraCQ7bGw//HtZGmDr0DVyGp3z3+XzHmkJv3BoC2hloYgjID5XS
P6e+DvMAv7jihJAcRloRaqK5jBQLw2Qhga02jnnYDwukMlPJ0rYcWfZJ8yHQtSnlArlBUoGOhxwp
ZDAWSUVZBWpgeLuzBV2sW1yI+GVW6J2XI1PY/B7zZIeXxlQdDuYu0t6r2pFyV3sfJyw5kRHZgb0D
x5xLxPX6p42bTekY7zJlIUWPpR0WV8ZDQGDU1mF6NxSicu8USBiaUj1VMKRTeTWpk2t26hPip1WZ
gxm1uxsTPHMIvAlQV3MmExnwkJTEUUCcc4634yb0xosOQOS+tt7DsltAwkjHTicdvguazIXpfLic
Dx6kXhTMpOYTiFUmWbXEBqOLvKzeILcLJB9PGR4lhR2pihHLcWxmO6Sxx58EFryLSkTo3LQ9LdAh
gmi3dAOGv3EViMACpqlwlqGWTLdDfzz15jHqhtW/hnUA/+CDcgyIUGP6/c+iM97qfnjiJA3f/oc+
C1JV/OubE5G0RCpmQoyM4lg/7THXTo28nCzfNN3Ewjukg1PPaGpbzYqfCNqLx/5sEq/BjzE/TWtW
afYWyQddLK0fGMCwkiKTfecpYsQ5NRCK/CWHWrUETcw5huSQIeSwNYJOGdMQLuo34HCSHh4yaa2j
i9LLI9k+IWRKoSthgG7w8jCoiZInan7Y3o3Hvt1PDz8EkKDsfBFoMG03E/DpPPxy20sHDHHjkvAY
DMvUYPxCR1M/q7q/UFfq8vWTwB2BXe17KVgLmSenAYGmPXq+Bqs37kZZN1xYpMwrkOdUaX4cy9rP
rObtjCqCo8eoJWLOCpLJESkklXf0T+uK6GpbodkkhKMISjIeeO+JeQEV8I3RDrAY5XKtuTc1xeB0
sJg+hTjln2oDNweIJfe9D8zHZYMZoaswfEowppReFPvYbO19iMoHr51DI2Sj7q1E3bIrAr+jELm1
Xfff77IGYR/nkwf0SdrQUwEvIGV5dWad6viodUYa2OcdQ+cQmpA67uy5XaYXp1U0igjtWM3L0N7s
0aMKoAamrQILpFzrRr7L/JUvxRRROBgeTveiKyMuiXP3tnbnP+lSMwY9ys7FbVpsY2sgLlWMNRhj
o5rv3vRq4EI5WLcquTCzvHxNPY04E+ob86nreeziHkaPmb+U6xZqDXp1n3FhyjoZALb00r2KWwmB
Cfc0yUguGdEmqjfH45pAyIEiVdHDudGKY/TjKeo+pg9gRcu82hljrTCPr+12YDDyx+JT9g1myWsq
Zs7Ux2dRPXk6b1B55orgqviORsfpUo5tWpm0MPjv6RlXXvhN8GfFDdarGIRfz9UPGRmhBgirdAxw
yeQJj6zTX4ANf/5/9hgfpy5fbABpQqrJx5l6bfXKC6NkZ2WSxRMKa873pRUfNLm/KFHcsj0RJ+ly
6Aiqu/RimOp8dFWD4URfh9LviOLTQh6RZJgjVe/yqWbKVrwPBNk5GBdJ/+/aum/qAWCcbGDgKsvC
H9u1Vn2OKPHV89bfgTzh25omrUOBzzpniDEl68rvWCttfgjpJGjKcu5RD7roSvcLs+UigJRRnMGJ
45Bh4wFvncWhBJ4pb2atNoRfZB75quc7Hnp67dKjrRrH3p251E8A+A41n9vwit1NkmNCQXM96TLP
wkqt+v9chM7QstCFWjIQXBcqFoLv4iDDjqDqvnFZLGrUb7GcocGAHd8p7FE1R2wu2sTUU0WWriKH
8I6aw7QLJVWJwJeJVBVOa8NTGi7MVbbfIIb3kMuDYnk112aj4ZVdFyL4X1QKKyCQpcZp2FAGeqFE
OfxWey+t+Qd04sCeG3uXNiagDKZ0D9bO/Qx7uWqKqAVYHc14ZYncCDuIvboeoCvnvpS9e356R9Ty
QIu3xlHKdDxSAnEuBCC4h9te3mwSXUbnnZqY2+I/gP4buYBkvnv95iBcaudt1xg02eEh1zE5lN1Y
gQOUrTegipJSq02BPSHIVStzO1VHtfyngBcyqAwJGSB/AkTIrNhkKNkjPh95Wk/NRAfkIuNtu81j
IVuDxpHDqoLnjtdsguA8GV9T0rLSd+pvQRr7ShJTNikDyab/XKrqa+KvSQm1CxZIxjbW2CU5+5j7
4mmRgEqgRG0GgsgBEtd/NvKgMsaYNcgNqkD2B1QSsuFvhZoZCRYmaHVW5+K4G1818z8TUeAlNRmj
CL9X5e46qramFsLRICVX4sH2Pttey6vnWYxK9QxiWtlLwcgk4mLHex2AQPA2HReUayBa/WejcIpS
D2Wt9Y2K+NvKUY3vDvzKvz9D6pdeeY+OOevLvjP285k/lUgzN0H2+jsCuBur9ttrz2LRCReUoqeN
nzkZuLJaJd6OgMxhelCruk9z5w8UYYkOqpWsqdFF+ogWLGjorDuhhVtx0n1RjWZGtuLy/A+sAT34
UzjxMEIn1DiyXaVVZskX1QVcigtueCktgElffr8oY0NzXkl3WViBc8LRgWbh2swSaWnZWLRDjv+/
yZPcYzneRZOHR97TXR0xZ5nuyJXOxfeaPQQZvv1NEmb/XXEsnTX1wZFI0gt56TsTdn+IHttPSSNh
sw+kQA73U+L6NfNqKSAb+Qrabtk3wfyNceKmy4a6alwcj+qiHX6VdkvHa64AKmRwDNs82n4zqqiT
K1ZaOQjrO5PsOeBD+bHGQ1BpzVIORKtFdNuNiSS8UoVGWh4m1V0jUjaAQ0EcKxCDxIAQy+uAaXF7
yI5/Ef/s7b6TR2qJmnOuFawYRIG5OdpTTRXbBuDYFJhhH2uUeehPciYvZFl64F3vsRiQPOtQsIws
EuABvwBFPrEM/segwBwq54Z2xeR77+/DxIkgrOdK5gJ+Z73V2IIEodBqhsjri7+YLowbUj1RAC2t
co8Ztkuov2TFGxOEdY5kpdk13IY7dWQXRMj/0I1df4vXaFASHn3BJ5l6bSfLQC5gSGleJnCtXp49
mp4CHamSWD50pFo4wADZcEHLQaeXvUc2H2KhfNF1Ftw+6AB4Ir72egF3tJQc5H4tVUmZ6Vp0uvMp
20LCMcX70B4/1Qc1ZwPVYhYkgxU/pSXSze+rQOCRz59i5ZL/eWrIw9J6VVt7WY9I3Gku3gH62vGW
VEyDZJ+dNU+kqW836IxhmtN8satlSeZiAcT3cos3F4BYmQ8fQPQPzoJLyQmFIPfpyJQWS44oLdfP
gPfS4n7/S+QNJ7FFID8wvm8RmY2QDIny6pi4tkK4Njs/aIlhZgnMHkCMK2r5Vw4AnLe9FGznfdAT
DvvQNkiiTHQfvOeLqcSlhsSe6jZE2NLHOCT2IlSSbWMZffz57NdClSxewgt8CkmEvtBS144ukc8X
R5XID2giJoSKHK9MMSn5vwa5iBUu14ex0MyXX+Wfiq2TzHVQSo04LZBuORpdoZdlYVtbp94yyqEA
4omg0evfQCGhCoZ+9niBdxLq7Tj1ee8IEDZ4fTa2ElLusesSUfO4DRlJm8nAlkKhv1J3H3jC0EqC
wYfI6stD0mmWDubC3ayOVyNuT9WQl6K8aPyV4H+WvZAnTNMhRmABAU8syRGFFEZx9IUIuMsgzO2V
glU9DBmdIt4BvWAP8nEm0oqWXXj6C5DB+thvnaQ/o10NDF83320b7DZD6cEK9RksYUggdvsHp3FG
P/RpmCQxw4TOuj4JhXCMyKJXSeIEPw/5YVWJzy+PzVyhew0UR09qEOH0K9BOinFEyzHz+taU1vz4
Hm4DT378HNsB9wIlMlToBkCC686Db1ZywTrBD3U1gDj5IOO52dVZSINby1eooGwwplD9vJHBrsBl
EKvWov4lgr6D/JxcjDZecmeKVW+kwbpLFjV2Hb6RaqZNRhcWXb7RP/FGvAJ2riLmGTGPRO48YFnj
4ZZEXCdBVqpxmM9XhWlOOxiEDV3Scqxaff8En35eV8oLAFLCOUuPh1ajEojce9B4HvHxQRlIuy2W
dAp0hJGwyDuD1bWvdCCTlTjQx77glpkM8pNJ8gcg/NUu+gQJvXInkPe7ceQQtMerg6UxcFIVXaJf
w9PX6Uk+8OwIja3mSSJ8NkNvuLan5v2cOwzBl26+9lcKLXDUNN2zNIn8iMEkHM7EDND5LZ8qdL5u
i+lwouttf4HKuJRuSRep8CK4BlihA3HJD727RvU+ahlEdv4BwpmZrRsbpogUox97k8grnYhaZwLg
Yq2bRHTTq05oD1XRUm2WIoqDFy/xMUE79RUwJozMXMaJzhmCzXmscX4WsbvQniyrG2TtVou8asmX
mDkEfEY3ipDxiOe7jqPUqgJ+7ZlYOBZSWxEaMnp9AU7QujKRefi68yu3FamxY2Lo3KD1QlX/y5cf
1t7Gev82njzisFRW8/z2zBtmSJukyfyoAezjmBjZItFBd3CyCCUkXrV/mUNtjS4BRydcEEe8v2lx
7Qm6HAAm/qmdovFSeBBWLUUVL5XvgJA+Oghq6cjVai81ZOmmOvBc5PCBgj7MwA8sdTI//vuPnECA
OFpgKfPHDK+cPeUEXjuykg80XDSi4RVsYz5f+YzTxXde+OlA/GBz7PyPO7sxljNmTbe6hvJvXRh7
xZ7n+EGwPy96awjrG+qlWQ0Jj5fVC5J+X+JSPzeE/XNVdWaUbbBdE5ph3aEauapIJYkqR6YBzyfE
hVIF2XcJa0CZMMMpcWn2FrEoY2SZ+wbT3zlMehR/0tF4T8BDQz/CSEaeFKq/Xdcb7z431V3uIj7L
RpNSw/9+VMgCnuVtbak4+JceNJrJ263Qc3qQTkKJMXDO6eSUE7b2D78P8lt8XzCF+oV8lQgwwCIn
Y7FGDJp/Gl74M/94NrwIiUOrB7s9VYQE5zznSYlSmWqEdKfIZ3BEf2iD3yuXYv8lYNbkf1uyXYXA
wLVL9Lup9aE52qypyizEc3rkdAYjq4IELca2N0etsuyra6ifkIkWL4wXu3Wcgk/4As79dS6HV/K7
LdJRypNVkeEuBtUy2XhsulGoSEwfgBKdymoLSIO9JvFa2sVFjz4WFENRQfbfoRuli3EkkRgB2eXo
oeaTwirG8KC3m6j45xrmL/oI88XjoOGfWy9yv9qy2t8K2OVWz+J9DV5GHblOxsct/Xa5pAfRh2NN
pN+n6wEL1A5FxT3Al9uMVIsrCKX+MV4MX8zxHeXw5Nn8roETKSWVVEtM2MirPkO0CIqjwXX3Z6Q8
lhZQvzmfDSsYjG2KvkXKkJuCAdlxDGzL65Jnu6052B74fmXPdB4YHmnSBQ8yyuMaBw39rIIPVvce
wODkid5aoLLnSrecuvaz/d7nwXXbsFPfjzKYDPD0VZdDIsYUqJz5+TZUImG536aj0P9G+qE3XdX0
W07GbJ69TLgp822HZL18yhx+vBG1N7aKJ0FdY5dE7wUZttdVYFjQfl9bmOOHKdWPl2BriRGGUmcR
DgRCKOjFoUtAryIlxYyv1vEvSqxqOsPuUWxrHjbihLSb3+nmbYQr3eIlGgjdeYjAxffHjIbwkfKS
P4rcYBEKsHWFO9e4bAPpBvQ+9SVbSmrYLOCasbTdTz/lNdlKvW/JK069BqwAOFGnjKVZN/zIbods
DgBAofi573IrS8+J2BNsOtX5c3uREuml/eLlrRvKxPcrfhSf+Nn1yo3neas/sx5FmndcIEsAngyT
k2FUz+wtf9JTQ4+Yp9AI9QUBbSRz4mm+ERXpDBBOBDUdYQP4rMCX0pSKUzVjhJKyZySYHLiKdSjr
Ofr5DrhdjJmyepJ4DZPN5nOBc7YmcGkzzZ2wUUGtJsadiPjGvz62nTQpA+WclCygmWfSHOYK5YbC
k2ukFeQ9ldDELemag8VHlNOOgfOwDV7kmR9ZQ2z9kReMXRZ/Lb9RgElw89++Vs6AsOt4MyUhWQzl
eWIXE8Ns+s0vVC0ySWZdnkmr8E9Qk44Q53Y9tHfU+4jWynBUnfKQoyOp54uhfSKXAbIi8dAbM42z
Mj633l9lG7+uEoNedahqcljjFhbSwgeQ9cGJoI+OVDXdMPM0Ron8jqxe5kOtZ2Q93q+fc/7tOzCD
1TcfHNP4SGqZ+urGp/PHdOBMx6MfFRrncIbgiBrbqMwUy4F2KORW1ws2+8NKyEAJPdsoUanvPeb0
WQZVuTwhNEczrRLIK2/bI+RYdm6iSteRcBzYzzUJIkURLG9rjlKAEvX7suhycXQD61DiX3OMsfZG
MCFkEbODPLKajxQuON/s5TigLKe0yE+ZGCV4PORD20qOAia4ctdXLGuthWVaK/YCBPjwafyH36GM
vUI1/rBzqq+lw9kql6myM/7oq9qKDubuEt7Vu+J3BIoTIbFC4QB7L4Zx7Mfa5v+gRRjjwK5vlByJ
Z//zxrHGdwiuHCYQ9f+K/KcWeBlANQLX+lSTYfCSYHmMP0XikYrlMUl39bEw+FvXVOGIPWLzl9Ak
A2GkLZZv2nzPnyd9ANN85I20OZILo913lQ6/Lqt6DM/lm4sToLHgaPB9iaX6934kbWxyLAjwVyKr
R6dJmUUAlZ4a01rAwcyQUBLkl6ic8KqEpsVLSUA/4u2VSSSsSGjCWuXWlrk8cpAWWgAuSfgshGzf
ll4R9C/yZnChA6gtSw6sMgwp8LzuZp+tdmU0RTIRpB06a7wBZvMMchY7TCyFeKaLKufmuIsHHHJI
NBDY3q1+TO5t9UwoY2VAkK78cAU3O6R0M3cJrjlHKlQFPlNIREXKpZK0DCd/+WZMUM4pInKxOTpo
3e9UDIe1cdlI1dnjzSu5cr3Ize4+bVnSsK4NYNp29Gp4nQprorSDHofi7Z8JkH3GcMQkTIiZxakI
airfPYPmh4qNSX1mP/rPEnxEKqUZa+ApUILW/s3nW0TorGYPXYPUIuwiqWRavQgAQT4BaF7gJ/Z2
WKMHV4YQZ9Z0o4wXJL1LZjjSK745jjnOGinKCzdCoEbfNBFXxxzx+opOHPY8zKf4dmBby/5wCeQ+
FxloJEnFIKBIJ07X3bD4qQBS0nW6bnj57nvGNg0Q7LTDxJsKSPwINHcnNK4+AkfB+ywIPSeAPa3S
w+vB6+9rG0sjHeO/IsjLLcOBNJAMXroHRsHl7pcV5gm3dUcJrfJAk5LCNYNwbI4aDpyLU4D0eKsQ
JNKsnqVoauDSeNSe8gln9q95yGyW4v//fx0ARXzmBXIH11H526XeDKljyjGFcz3U6m6UY5aFwQ1u
RpLnLu7qrHsf6jwP9HF+mSk/nqc73/FvcrXetLZVRQLgTX3nYKrQT5DMTYunmAknYZUo8o5iy4iu
jOQtto0ix3u48TfouOD1CXymUTmw9khra1d0Z/68tgeVarXUjtIWQrqA+JLvz6u0tl69Yae/fLt8
YFmzb1IlXiWZ6avJl8JRUIprH/+44nDl0rr0o99dHmgmXLn5ktK+IJTT+kZhzsnLsPEMhVHjsMe+
fkAgHlw+1I/pnB98IOamIuhywZnhS7pl7fBAnsQJUzDGI3CGVh//smHC9y7py5ioFi1IPp31lUs/
0LDbD/yatMS6mUhgONtLpM3CH/2cBwkdR5TPYQ5UQ5J3H4KNYTwCsnOgoWB2gtIIwVaMjQ4GcyC6
Nn4on/hBhX0EIOL57WcFHtf/tZ5Ct/0pwumXi+favwDAZKxoCccpDubval+20GfvJOsch8g+JxWz
FesoPjWBZD+pZSvihAMBrMFfA6uMChizHvQgv5V8FsUWkCCFoblh7kKgWRYckGyy/n23VJXxGrgu
7iz+JGUVFwrEP3JMLiJlnTv29ToM3lbzc3gquBn3jxCAMV2CBzGJMAqcZeFYB2TU3GBM/yg6rwi4
ogd/iQ9aqSS2OVS1VxOZdUY+THvEJS8ugea4cB7JpaDVo6N9tU35jqiiaB2GmrVKnLdu/obrlfjk
ORa99BZHv6qqBjXbY6SGpr4yAR1jnf77ua8BrzUeotjnKHAEH/EtyunNHCyc2ZXwISxsvrJsCC7V
ptAwICTDU1GgBy+KwQ3La2t6b3XaQ/m7qhaIOKgvY2fCGSCqGQKj4nfNQDGEuDjIEkDEbAol65EQ
QO2GH3NiC6hszZpFhjQvM5uIVmYjHcjKsb1CKKpn9KKMQmfaX4vDuEhMPyg0uPpvCAPn68dBwMaR
4EbPIanZRo6ez7ouc9qkOl0ipphjGwB/kSbtgUm8D4jM0Kw1TJpjLzdOUj1v9sxuZMrLrMRUk2h3
GzkeOjG6fVy0hDlih71JCSM8Pd7/085cvdE9n4jhPBdpRbNIxhAOs5zkWgz6B/c1toZNrrpSJsmX
HxVjlHuUiSu3VjLHLfqbPwik3s4+quQO+TwrCbFXVSmY/6pk6psw7XSCrznEJsTfmI9jJ0B50SwJ
ndEcvwvp/scwPThnJWUQesJim6gM8dpBAFW13ItxciEr0lg73kD5c39zbhq8CJpLazy4LzPtPws9
4wGjketj/8KGaQWRzDGofqgUkHQBM/tlzQmBziLi5hZYnrQiwNv4CBar9dpdNwfb+tAATF6HJVq2
GU3Gat4off2EfZi2bwYjWJ9kLlOmsP0PekK3xpv5ycOuIcmmX5pb7SRjDvkx8+VHUwk44CVcPpY0
1i4I47/VBD9e4DQeLuLj3tqs+6b6ZhMbcZhfS8kwj5Q0X4cK4x8AFzkQwUjwO+R7losKTnUqRDpx
Loe3ew+plbJKYMLMJq4YHZYb7jA0ZNY0ZDkrDs4ARi4Z25Dz0TDn0cjCYu+S22F646AwLndgmRjA
8WcMn15P12k0YzGCIAlhkf0mz43DRZ4+iQAi3gLpExj/dSJ3YQtupzWopGGMzaJMM7HT7/6wZIZQ
O83GEW/Q5hVeZiun2n2PNlOgkb2An6nWA9i7dlGMtyVDCufRGSINP2QXIaEwWMDnxKZ6okU6dTch
e3j3nSu7GteU/wfy+h60W3LLQcUgdD21uF9G5y0JJieXNO65RegsFl9b9fAW5G1gOEQAoFGFFkJA
eC9fT5LHiQeO4hp2X4tSHzF/S+2a7XDEhLR3nSPsDa5DDMs9FUsnxMYqZ0AIjJba4HNkC0wOwtDv
7IgBf1cwmVPOQ9vyF9xHlK/ZhPbZR9ozqRk1dbCghUPnhMJ+HGXlqIpeHO3Y/DDCR1VvZ92xsX9m
Q+o/pXjYQpnO5WAbZO+tEBqXq6FTiwGRBT70e3xeTlaxu54fLqOOE9I0kELqGsnLvGjzMXVrIQPB
tlJEztkJ5AUtAaEEgLH7L+VLD78SMLjutVYSX+oFjhiq6cqwJZB2ibUqwnFp8/imvC83kmqwUh/o
P9k13FOnOU684d80kZxvQlluqx6B6/uPoJoArfrhlbKR/8O0bTpGlIARqYII95xSm8Y4DYNyu1gL
KqRBTCFWJInR4ZG7hdjUff+IiVaQ1sucGPo1YUl7WeNSHrkNniw97ZNmgU9eWg6G37EvS4Y/KROw
4UXDqWGW9vB/eOXQ5zSoxu0X6rqobF9Hkiq0of8coDbAvDcrZUHn4LH6iaGVdgLKlJ9ZZz/gO49F
zr/mgQ4sK3fG0Lav8XvYEBqbLqlHJK0Lduk9NBrOGZW+IjZGqyp7xRfs8bhE5Y1WcnXprZ8JJOqt
NvxIw6UBWaagGV0eOAfOSI26fX1ajOpgXK9JIqyNhf9t8qtwdLFnlMj+xudRGleAuDx11PdysldK
Xmaxk3xEx0aaVsZuocdWbGif2ieww/CYFb5Tc5Hcf/elINvmYBH2cvLuaglbeP4TbH27BF5t1c1+
49nLpQyiAyKukyg6PhjJ/FnLWQ8vQhmLVbQYH5koYP/NIVMKig2zd+htUhiO5dG7TPb5/rRwDLrN
7ONj8qTIzMCorXoA84uH4NJVyCXcKOfpLNV8OR8718vPcDslYHk45V/EaoxRDlbASjH2JkrEpSnd
oW4QecujPQzqF8BqeoKfuNeKzy8K5XbaWBIpfW8WXgLohFi2DEfL2dDYUKL9e0Dj3GZBMigclRI1
fzse4yo8zYMnBbPk6eFCIMuBMQCwOYwcvzuSJPKBnMQiV35e75L0aHnR5DXs5W2qkKf/o8eCAKT0
z/c6BPsMUbTPnN9x0ki9JPTZsiezdRyi1nhiWyG6HWwCGgNTmsUZPUav9HCdmTZqEDeu2eKyv5VQ
3mFH/0zJTyzVFe3CsvFifk5A9GNDiwM5OUDKhjKBiIdVtW5Dzi3FFpdVnQcwq4dIBK0lKjbbjPzF
gCQJ2Tp0/UmgapUu7wQvU6cytf+PoKtKBWvSmNNr6ogvPnN4mfYu4G0sPp5RT7SwkPFosH7Uhwl7
3DgXfTuq4ChNCVlq1t1Ryxw+yOfEdSjxuW0sAoUt7/AsxniOdUw78uBBPia0aVIEjOe52ekbvPVI
CX9eGr4bgoFEg45kp5rv6mJd0wtsM/rTRdZ+MGwxgZ2/jfbom66HvHIbBFSfdBbMe3tp1t39wjOP
ZPyF/o6vyDWURcQCCPBYaXXzvOqDnZu84NAGQt+PApET0azAUotMWNSi9Ao09gdqei4gPFY302CJ
2ReVvSgEKFyznK01LquH2IOPbHrHCQvrQkfHFkldUd7xPeGDKG/lv6wGSwxUWDYDl+2q0LgMpkbF
sn0sdXz0exRH7l3950tUpaC+jBz88CNmrAwqTI3e9HxMGSJ7M8S7ZxqQkSpjD7jcOcP3IWxQ2Ipg
jtLVm6BuUM/1ZG9wVSf3FysSiLbMeDZCbPDB+IrMB/Xj6JTgXVMRdsMGJ7e3k+F1H7fTzqdQ8hFy
jYtPzHXWrxWfE1BwToVYZno3HZg3L8st0TjC/8CRGBotQ8REg9y0fLj70asMBKl+mgGsCge7P+tL
H6LR/oOyjVs+xbi9386w/YF4LnH5exwTWZFyaPeJo0QmU3Yno0f8JPh/mozvYtY2PPwcPoBDRphy
K782jH8MlGwdN84bB0pPjicuebj/XD61ZkKTyZ6duKWWLhSqMWos1vOMcymjb5QPuJV0+DROu856
q5sBX+gT0vMCEMLfnezIF1eJurc8p0mm4KWvmPupmpedTNVf0EXjDhM1WBIp2T4X7edeK9SJouhV
+35NXtxymvsZR7w11tK2F8c8lupEKVkG8jv0vClLYJn6SWfe1I4ZJ5nI2pDV4ZBmr/bzbhUJDhhS
lRbwKVFNC2q3lEp/ii06SRDZJHbmplnmD8cSVi8VKlSCpi5UkvQvUeWH55lVV8KIjF9nALZPTiIY
30u8jXHM6W74QRu5Bm9mLrUdTEcNwPaJbelJE+uCaD53DZBrPJkNA4WFKBiDV88fJ3ksk6i5r2Yz
OH4oikexVwT/v+r5PYZzAIXM6YVKQfVnzdY5lcStWjYzQ9bY36Ruyc1CeKZ9Os+ST2teoktTPv0C
I0Sh+VHwOXn+L+f/nrcM74T6119/LbI0oEFjjhkSN0sQH14At1b3IjOfpA7NN8VM83mpC0Hsj1hs
6D6Ycyn7l6fWtEa0qSdxUb5TOOl5oRlBHPAf6JWg8ryJe2S3U42pzd76nmSohxZxLc5bM4yjFzdm
cLramoUxRMJWA3N35vrstEm21awOITrc0g4z7qvFGtZdNjnGIvGGUevOeK4VGfoLW0PLlmvsZ0zT
nuMh5dxlwpDU4EbZKz0nTsFgB5hl8Mb+5aB6y1Yns9xIsx695HQEqQeyz2iEw400TjEw38BS57nr
TqlV0lvz6TBsT4rv4qIAkSj5s31c0iE8nwxavTO1skT3Q6XLXu7uWyScoxpvr+7814YqoqtkaPj+
M3UkosPIabgs53zRyoe2lYkQPggVAl9Eca6AEwYQuO3vT4p5goglUSIZdM0Ec0ZsL9VzS6RJSr6J
kWlQxV+U0EIrp1a2UtLm2QKV8MXj+IRT3Xc6pQ+UczMdSzswrrPx2XJeLPjeAcV9CurpfsSfDpux
u/SjPa3YFMuH0uUU/D0MDKvfzw2OZ5qzvsro2uZv6u2KUvklFzFeHL0vLlzRoWnBE2iGJyYuy/YV
oYGh8Gpg5XKUoQhvgwajpnA0yBoCjDfBwtvibSwNjvqLr6ZvktRctRighg8O1JPIS9yfW4FxS/ST
ghGNJA1E44FyZrkylwCRetn4K0YQ1KKpK/zfjEV2i/h4s9g4WO4xbnySvCcMmHq404W0n1XSbavi
uqc8iKA22sQMrLIxOoF4EqlQ4GFlzR4qyGGQ181jH7DsX8xTKV+ELO8RYy5vLaMxC0OJId/gS9E4
qnFzMEEb1xQu1aB7lBaKrDnJCg1q5cMbyizFKCt1d73RiO9uDr6YGc1ICJzT2aDeG2NEDU5wXamu
CTOPVbs8Cg2dXo06STGJ0ZEDIYBvRNlV+pq7NeiJo2uP/M6pZDWS+ZtY4zwUl5uALUXpFrcRzID7
5Icpy625O5a+k6mOrRJILWd3mmmE4ruuXzj9cF3g0DDQu6SdvdClz2zQw87XANjsRc7paVR5DPlC
P+EWKbrxVv9WHrSg8zr8dRaY8VIR2NJ5dvlPwMEkAaOhzLqgkiDR4gST1kgUiW8Zqasgc8ApQOtI
Ix3qkdrkP8WlfMJJ/K0RSzh2lQNQqKgK+JSBnnZgz6xegbbHHv63F8x1xTeUZ4IM6gBHzhWC4TNb
XKKtSKzk5LPWnH62cdqToG3wRa/lulZE3zop0Uot50I3pmgd3p6UtW8RZ21207yEiyuqV5QDLcug
WVLhLrUBBhh7NaTiUJ35l/2ZvXbd/ZsHGXKL76+xqg3GSNiOnyJW7Fo0OKyb0SZCDnrHG1dSoySO
PKB2qBylcVlDWt5/1H9gXvL9UJ7b5l0XU6vWS25lIiM4xgnQZOdosWAUAIYc7BSB3qidI94Bfm8h
Th9HbmuQXOnZs/nN6/V7NsGYdoLqnG58jO+sXALBqN/iJYVS/HBS//6w9su3Z6FA32jTn85rCQLr
yc55qtJ5DeGv0n55LpZN+r1XhSq+PAKh5UjLVsm2sFcFqJchboSSlbfSjp81691Rglbj2icHxTRB
esBgbWqTRGrn4h9Z/shIaVgDgnpf8shh1+Tb906gwuiswd8+m98Rd/B5opnckpROwlPkEntILp+o
9vSdFmVWKjicewqQNY4mKjbSKVtYniRL4uvWbvzvd44mL7PQkpXQj36TMN/TibBiK/FQUDF9qO3/
XQRiZFgCXkDHwoAr+wTOVl7PKySYSpTgvUXAss2dn636PJV00/EchgonGIuCIFxSCkEMAAamRljW
Uh5OgSA1TKw+qGS56a0FkWkIu9xNvHfpafibuoSP4Von1exD+eUqCfBTrDd+dzJ2R8wruiIJymUz
/y6hhsppiiN3xy1+mu0FhDTA9R1LanfnoJDTvFsvWbFP3RsQyJjxare7um2YAXcwUT9Jpxh53uJq
ZGIVD7s0BPbx5bF/gi/q9Cpiya2dGnsn04XyvvT86bbxSB8+3gRf43jmxKeYpBMa+8hCO5pRYgy7
/mSrcFW+j0ufggS1iLNpvpobdGI+jGmZ9k472JXLTVuSzntGZzwTcSIUc7LuDwKbvRUaMESW8FhE
SlEylvZ8FhRJIz1g7Y+kmAqNEE4aRAbWd9XgCNc9u5XlgOTvd1A6PL35ISLIwxQea3XTuPR7JnEl
X364lDG+NT9/iEq0lw2L0rvh+k96RoG05cwEu1mR6Yr2O1IPRO16ltzdXxkBOBxZ2uQXTNx2Nmwi
I0o8M09RYRaVeHVZxgbZif3nrveDWLtk3HV+358oKE3Q+PofMWHZbFtsi2mwRFXUWS+AqErr177h
Ma+HVgHnAKo886yB3gF3bbTn+zDAk3Ru41zgUHf0xEO0uN0fxBxWH0f04owjriJQPSjktwsuwtUG
CvrQEVyqMqCvnbNnZwLtICf7hOyaNqjZN4hRPMNNv5RP2kxoHkk2ifBDwfACGKMG+cQTo3d8CF6T
PTNw2Edwh8NIYyudgLNarYpnbtth+qy7J7HgV+LuUrBh0BXTWFY5sRwc31d1jkkn6ude9ai9PL6Q
A3/JKB97MSf4BUSfVbdvq0NiQkxYLQ6lUV1XrD4BDl8ZVEf/FZqziH5ZbGWWdjDzT97HbvG5JDqf
JDtsiXB6TKh9yBt+p6UyKfQvOj6f9bH9tPfgHKbw4IgClI8laBkikILt8Wb4Z3XcrP1xoXWI1z0X
m8zj0ULIgTqnVViRkEsWMjMk7Vmqrs1YzfKFBHnwoVBe4gvFzLEhv8MA01xJAWCwPX134OOu9+1Q
2b5B/lpdHZYHrdVUNQhs8EjhFCDSXAm5wUnsyu862i86TuwA6ZujHeiRM85GWwRY6XGg8SOciELm
P7F8ygLzKdn9Q3IoZ7XlH+wt6xVh9yBh/NEmKAJB7xSWlx9QkWh6JF9Ao82xVNt8TH6Pz4MdRWSs
IQh3pz/DQo+S6q19l40k4ETMtzMGr7QKTbA22QdxKtWVBIooPRl1PiXYSc4tkrzx1bn4pYCST1lX
NwPJdur48P5bBtKTqlzLShJzWudZ1K3c3+UA0PpM/eP2xoG5jJ1btdp/oqXEW/Uc2TgvDVS50KpL
SwugdGmBX1qe6Eqk3UVnPKUNm7M/whQ65S31tGxrd30vT87HI14MkWKIGSBMydyHSJz5W+/xnAkN
YMdIThsBHchvDEbB4D9HqXr6IO666W6Iu0w2f9YQEKRX/Ng8G+5QUC6fMfve4zIxgi4mvpqJeeXq
cjAjsOg6Q8AfDe1F26NNypct7IU6DQjuCerud47e8BtVIyk+7SbjvKQJ53lXbsPJQYRg8npWQ0YP
sECj8GmjUm4ZHGQhLcWLgWl/mJhlB1RYADmdiWxCc8T4v6dugEY7JPs2nV+3zz3vusxSwTNmDOMW
JpDA62uDe1ye8m/EcrkWzCTa0PJsLv0ICsf+uOZj7j/M+ODP5jrQC18u7iBQOw7gVjXIV0rZsHUg
QrYB99cZ7TlbLFKLmCY0r0AGkpjDsooQWCPcDM4ACzuoGwOTp9JqdAzpeFcsyo1IZ9aLPKAXWIVZ
or7dInKyjUrSnKkT121fBDxGRNgb6M2GFlc3iMriScZXD+J8RP6ygz3BjWrR6XJzF+rdA3KKQ8bn
K7VOB8MlSAIJWxjQyB2+33qOhknj7YB4lUdp911p4wpgJzuD9uRYmqjUflAbiYxtWDCF7IawyeBV
6EL3gXj52mImm257rp+k0/VXg50a/jO/BTtPs280h9lisiO5L/kXNThB1mSLKVP4fEaIsrHXh4yU
X2AkhCA1fCgVsXRrE7wtvVrsB1DZdMY7rIp+WwI3j+GnzhzpdxN++6ZofWwDQc+Q0GsILxhYz2tp
uJstxwsR679PJD4ZYQalw+t1RFODD0Q6K8enVjpyxY07rSfCrXyb+OE4iIbIVyuvYA4zhI83BP33
NwGPEh5wO852E1tAqsTbrEBAHIowBIQrgmMlXONUjaQbsMtApkxOaBnPDVutssRXEgy5OvHKn9kS
7g09DmwLLMBKTr4P67jUmjcryy4k2QBOIfxjE/M/XpR5Had38jLWrhBgfTTfthGQQrBLCkC9uVKq
h7hyd7rKjXChFppxcDXN5whsjHowO90M88/vHi9CVHvsqaXhJOh14VUm+aTr0TApksQSBbbVR+Ku
j7N9hnl3THbqxCjFm7rLg00G8b6c9rrgbsPNYJXy7yrwazw2170QtBJ2hCPakf61+P9LGhei4FOK
u2p00v9ZZk/XrvgEcEnaxnY5p1KljkHIwl60HGqUweCv92Ti86C6uS7WA6Tjn1+K8B0m7OXJXFHg
ZvaGbR3Bd8zSoINn/ummg4oIi5yxFYze/dhr/aRfF7DG7QzipAXHo8QqnINVVqoiKJzx+a9pXQC8
xwXmY2dqLcJ0Ud39lsmmX+S1DqUD3pWBFxsbXUt+ujuT4ox2Epdz+pCghaWXf2SgoKQfXQHO5LMI
52r314lfYl2lsHyI4y+OlREqq/Or2iNhmYDbzvJ0kPXovSic6DM9bIx1ebgOWhfDwJsc/SkAd8y2
d454FHeB4aAxJiQIohMq5RHvAE0gbFBwgdzQ5iP/14IsXhL6w23b9xHTrjS+TKVeCCWkYKO2ryrK
zHZtQowmL5LtWNUgFs4NzpXU1bqQ6ejbjEvd+PvYBD9C/51xHrhw4FC4olBtUBAgH2f/YgBigMHl
TxPF1I5wuntnwQ76HW8eymshQ0cZ+f4VXFhmoNBZp0TxvJ8qW0dx06XkcejeXACEaSwQsrtBzljV
fcE4vXS9L4fmeiwdmQo+hWtqqKnA7mXXu1ZMQdNBmUL6FMJy2B9Z+BeXpnsqYArM153yIKf4hXLf
KpchB6tRcvdalXlOt4LnKsjHEfKUEH53U5qqOraaoGXf1tjDMauO0GuWfA78W4VIYA9ig1U2Ti2U
Qgv1qiPNHOGKY86KW2Zq7MzHQqIYydVIoPHnTDsHOsGZHGmaFRIL9LDHxCiaEaBAK6XeIT2uDWXs
srEb/SO3beSzS4xFoYAlCX6Evn3DUaEH0AKj3e6mag9Zrkyw3iRfyzdMwXn1JNzo9R0m9gue2wsZ
fNA9ggbXRw/tnUdNtD3D0pP9NpbwyRyIltZoKrk+j4prCEyItIsmuWMlGxVa94/f7BYDGEXWeu7K
m2kCzSZjzcCeGe2cTZqV/avwacTDWICMxFRyXrY0u1PGvV3+rXvIzTMdgpmaot5W4YWUPbwyjqlR
lmsUORJEUsBTgzp6esHRQEdWygEuKX0GR1YviMVrqxDRxIMbzulTTuFlVLtBlnk6Gv2zfusQ7mvP
I6NC6a86cFcXs05I0YaF1ccBP9wPGusBAqy9wmhNOPUJf9OYUXlsEMzPQ+geCohV57ApzZwCPFFB
kPW9z9pxTQERsOBC1bYLPSeOC5BmxczGmkuCnYWFtnHobWk4jXG8iWFYknNV0wzgpQRqFhOArDHs
LEN5miYB9nLlK1WtdE8UNkG9cX9hjzFVugQOux4Nh3g3k8c5+zr4CuMJ4MWEvSi4KydgxjjLt8eE
DCcZqYHbQs260DWAaCY1JOREHmrubh0fCdnHWYlMMWuZUwCiZgkryacOGmYYQgYlkSYqg1RX3l/m
2G6rz217wN/SKBDPQZ1BRKZWVfu8tm5qSKMHcNW3mCmtGdJihsqp7Cb5DwIXsQOrCSNlybz0Wana
WX7M9TNDzKCpRT66oFVwIrQ9uUlNT06XOG2V3WNpPiaExHxaj7ZofzUmT7ehRWQM4iGIMxhLgJGK
mwofZyX8dNnasWE7duIka47K8dvTavGF2uxSlZAftV5Rom2trWTHYGF6vP8VQUy8Re6Bta2qmNcr
c6QyAYVjJRs4s2MiWTUFOQUtfq2tlpxerJpUITAUHvSFjLRTeNJ1hPR6GR06LXoJv8foPwZQsAuu
plKc3+kIK1A54PdKrP4FyK7FSUOWNeICGJ/4PsN6qZhP2+XBI5bV+N4WERHKkqhjGyo+CPg0OO6X
wYsU9l0tPp6HvDUG3v8ofq4vH8j0lmxVEhkECmk+ksmuvAPJrSkIk8e6Fz+NPxvD0nIocblRq12U
FERpxYAZtCiNLpVAbFjeD0jqh6P8pGg7Xn3HE+IkPijNDdEgGeJfEL+L61aQaED0N4ENehbY0FC9
9Ub7jXYCCe/8XneiTLmR7tWdMBmF2G1LXa8TPEQLtw65I2nD79yjweM/HPCCZTD8ROg1npLK725E
POPDjPEiIr3Ci6oHSX5Y2RSvCdQWS7oYx3Q1Ab+W3sGg5okRmzThjIVDuB3B9jixvbcQTbxlyV3t
5TB8Fp9d2l2Lo3JYxnL9F7CkKyd2nFi1eKaV4sRt6gUVE3Y+QGo4sFu84vAVv25Jjbq+POeMPhSL
O2I6fKE2V7L+aPGCzDE2NR010jPzHUvHkQ2CaE0iRsj2mzSxchi87lcYckGzI8ixeJyxUseN9OzZ
NIuddj3jH+J6VcB86j8q1XQr4sQg7YW+XNNeA/TEl9DN39ht7DbQXczbj5dPPaxGizL3aVLWtXCo
Fu3YgySI+VEnUMFRWViheRDK9QPANKccjwhZOa7Oy2BeHXy2YA2FF4DRPQnW2N9km1fjQGF30ODr
NvAoCQFFH1eKQhldlM+mqtlbv2ozTFv95ENIxlvwkxogi4/lG5gct2tjwucPndNoivImGJUQ9PCk
njr1jdiWPuHb1yzQ4IevOIgtxuGacZpEmzGI5Bt5ocr+0oJIxLsw4GMcDDOu+s5Yc3vauAnriqVZ
Juo6RbNI+KqUr2RXZJb2maT32sdkS6+NwFTAZtiJCz3sTKMra9T2IQqyDTn/YtcgAjFZl1q7fpYl
Wyhv5jX0y5uYbiLyf0RZ56kYDSHisgEEGyTqV6FwFCY+Zty8wYpJsP3CmL8AeBzEEI/bVE7AA9c7
fZ1j5JdpPjLVASwqB5Rf3jbtJ6+/9CEqEW/5o8S4vrep7FlGmkp0gwbeJlN8vl0+/PSs0D9fYUb5
Hk9012AUjXPK2U6sBXpBZQIdWXVR0Z6ympFVz4dyCUslOB9658MG53GUrDWDd/1V8blusXSGFGEi
gG+Y3nuLJcQSVug/Ho6p/JGlXvuTHiXobuZZN0P9LtZH6kT50MNJE4wEUgKx7WLzPlW4ikULK5bM
OUnMb2UeU2dQMnifEo3aZvzdPK7zNuBl0lgRKQ007CuSsi1vn10+aqD5BBa2ZU1mew48fNIaWX0/
0RMazYLuNdJaETOHtk38qdpFf4HqfqD8Ro+bvp2vzhVpHxC5FdSpXWtTeUg5unk5i3tUQqsNtOyD
FWdxyLH4SStfV6CE56kT/ZRwDWQVLEbSYkcW2UR8nyn3JhqY23tE4f2gH8EFz089wmW5S+dtre1k
jeKcyJ7z2kB9TgJiYmluzQhh0+oCtgmn9TFQUyJPScikqL/WhXsoeZaeMHUGfcqYF6infJYQsZGB
cNYSTveRgKsZC4zXFtb5ivTNJDdBJEjNmdQdZgIXvnE6aaK8N+6fwJS65/Nf2GvMuEhPQJV4lwbm
wVfBGAWyXdD9RFKRYqMLGa09jupyTerbZGjcPjej06TtnKhfBeOyorCyrcnfLrz82dsJEJkPJfpH
5QDp7TovYrZRhW3XaaqFwaMlAcWDZtQW1tHK5vIRqdlmvs+ieEFKwCeWrAiap6HKDVARYEj3rsFT
aNKpD+L/MxZtvpt7X3DPBfp0GJZqF5PkPjTnlC6MFWyr1HArMAa2j6OYZf4u3FIM16TEYge8GsvV
PCBBXDRctVlXARB4aY4SDYBNsP/wlzfO4zCyRUqt5i8KN/lH2S9lH98G/at6SobtIdXwKHHRXo9b
x6h5xst/rWq2q/zcQdIkjs6+Pt3pRmGn8UVQndrcF9hUesuojMmtZ8iBsgOVlpNaM0BELp0TbaRF
zOm1AlryVhmlnqS2TTB7raC+G5mXNiOP4tCVBhtP5Tfm6v/7VdpaJllymLQ7ve544swfi/9pG9Wl
6SG9AUK1YCBm7UhhXHSgqUfq4VOcPZ9e8RwwqZZ3ZOLNzgU65CL0yJDhEBUnH6FWObZSPTt8OCxP
cpiZiPq3rdFquFMp8k63AfJPJSTGYeQ7coV/tvr7dHmiz5vrttdVx510H2s6HO4ZwPlfkCA02Udh
xpG44d1gnokWjG1XNLucVkTqSujp0f9yCcDBV8/EUv5ArF+ApFyqsZ9ZusZfSDLOmA5ukVyBKHAs
18inygOU7DLMQk5BbFYDBtk0JI9JHNrLz8s2FINbjU2vZ0sQmFX8B3R1EXHx0DF39W8DrpNpVqxY
SmxtrkxD4EV29LFaarkA/GN2FMMBpG7S+ZSw51sdieAMnXRGqNKsATWLNTvGr+FUMpaElNLJosCs
2vmrRz77DQ5P3/V0Y7UKHJIQ6kw3CwJ70sf4uWJ98g3IeI8gSqmncNraYyxLIehMEjqhAr1Da7l4
SO8HkWQh+S36NFusBDJUanVRSv6CB3zQwjnzWG3a8VK7j0ZqkgB6PkJ5j8LRO+rA0KNyAte5kG7a
pPdyE7Xe6bu4vjIs//mMo8L64j3l3Oj+pKxWrbl607PI6RjKQa8RdkVyQV4VWY0vdOCaJlpPjtd5
UlAa63tfoD1YhuxdlbPHO5I0CkKOz8S8ZnBboMDLneTRBDTgDxxU31tsD8La47mXJMgS6qrh4hfM
sX8txRnrU96m/9E381HOo7TyMEVziVvNsTWyueqLhVseruY6iPvN0Baa3mzXzQvrWTzWEZ/GWaC0
luIiXsKJB264oN2FSrHRy3/aNxaSHIR8o4o1+n9ZkPpJfvZ2uRuhTwE9aIY7PpZMdv0K1j47+fxe
A15FxQh6dUIQ4cG1r0Ge7Nh7YcVCvLG3bkyjNAHdo782sHHyM5fT3Onu/KpX/iAnrJ+V7txR5Bi1
3uF6W3aqA6JlyQoX4bYqp8Y37APeJm3bfbUDBWWrsucs5WnVQNJnylJHHjKtFes9Ny1SBj2mD2Ey
bD5HOwDeiqQaxO6Au7B5IlUWCjvOJ55gS4J/7jW03q52tSXHEvJ1vvx4vJmP8IDnC3NFegdR9uO3
GHEIdOpt9etu/CZo1A1OWGAt7wR/bc7UmzMwo+jlMMYvhto1zf+cI3dXRRXy4a9dceS4FDyLE8he
eEnsrE8FbCIyOn2VVWGepwYL9QHj3dlD8w8lcuc7EQic2SQu/PMx7iSk81kIo64917e+mGA+7Dey
wJPVMSZsN9Hko8pBZtZ9wvTeolnXyHkMScg60UsER353ERpGk1sVi2HqYGF6Avwzp+fzSjDx14V6
EQp7bStZPXWPAwbAnu3rE2zqraU/RjVGHINM1vXWjTvVhzAvP2td3Q2mR5VN6iIYb/3rSHYwW+BS
f4AkutjM0cx8imA8cSnWxjNnfcHwTuu/tiA8G5Y9ockjYyoCac2FQ50TyyLrwCY3yoSeShF2YEmi
exXgoMtWTjHtWyckN9d3QkTUi4hdQD79ercc/TWuZr2TCUbC+OvHZp9oFyRRgzm9itpQSiRMkJm1
C9URMPdFYe3qq0eQJGYYVs95caCdrYvFxAa1smrGNDAuWYzkLqlo6fo6b6IbNKt5u+onqW7g7FAP
3BL/9eGGChR9i8byIqPr2FFfWMTuXwFNtDdLx7bH5wyG1mY6jg8AG8UlfdDRxxMPHNnjEdSqe7kn
PcDY16XtnTfnha5eFWtbQ52/X2LrQ5Zgc1acEH+D84Js6LxPQUMT3q1raL1WqSoBIEfHnZHILUez
wFaYVTNLo0AMRSvfjI/d+nBYgMVuTQjVjA5UcKR141QmDapWXxRM5re0czjvKZ9i06rgJEIJLKPL
54d+wPX9SVf8eWcOlFOOWZdXpyP40Q/pp86Ma301lZm+ZmaizoMtOPyuQYd5OUPYuxO9VGWZRBdZ
ISBWFo6btWuWcJ2UDcslM1ZAY50txgGE5CLr0a82au0Ik4AbVkCripnBrA9aSerzNXQAd5l+bNWm
TL9gxNEFfvs8dSVJ6I43hje9buzkWeGGrT0i3WHCnelWpblKGN98qdM2rEkA4neznoAqSS9Fv37s
KDPkMa6FmBGRmp/QhOpjRAXIkluSkxSwGpSAWEPZghOpcFvoq954aK74eHqID57sOmkdgyr7iVLh
o9QL5VSMuQQDCkmcAWtGV/A3bNoEoZgMddaseKBdIo8wKkqWp8medBL93pFuiYpC87XSVrTi9atE
RPaEK+gL+r8hcG7+YHqe7TV9UW6zdgrB6t0CLhswCLkg12iYoEDrdKtXxxinlhoGQDC9c9pbiMq5
raMfoOuEU0cVQRgclUcsU9DGWaQ/PjVINq0zYoadwfPZpa9SvdCvuhdxG+e8s76BJzGdPO7qUA0v
QkaDVmmrSs2lRNspR0pH0hcSG1LRFdbj8TNcV4t8GvOR3sYt6BfPXYU3KrUdUiwUdvRxJEarK7tQ
rGr+KcwZM/ktlRh+QbK8WUEoBG7p/vRDQyqMe4vCkYXncgQ6W+jC4s6jteyJU40HDjOLDlCpkvtk
hEmAOOKMYwOZKE0E1gURWiz7GWIHHEoCZ7Eihr/ujoclH7GZ5KdmMcB7NjSPy8oPSGfJbHxSP/VC
Kz0fajnQ8ayxvSZhwNaYcPrN5/p20tinW6mh/blNjvry1aGmR8yWMSmywayz+GrzMmixgQlilluY
FUW7QMhnhplpJMmXbGFlC0KikqNmWoHqbXArdziBXNeZAYp7juNL+SwcoUISEBn7sqPIQq/f6hmW
H6/iGRAJOvGzbczuWP33510JVvwE4VB16hSWLxUyQpWlyYHfdImFxru7v4kWfafvEwqdLwSpOSWw
LpGGLQ/9x3qJqRgV/tWg1kMCNhzsDq1cwBwAh7E3KQC+4ZOj/wgt7QiHlScDrzDMFm5VC1yRzDlS
RE6K0wXtZ7Wg7OBMX4sO/29zMLVkHFxzNDf8LHT7iWFfFlBImSBLLE2IaKjR9zeNmAI6KZJpZ4RT
Nno0dcMIdH7bMtMSot5KiSRPVU5GJLZ4wLa71jvJK+OZdFCw1ex0X3yLJgkShHIuz/gQrv0Dp1+G
di/FJluFJDDICWbGT4LcfVwB8bHB96SExWTOyZOf9dKjqu7YzuPkb7gUKixF/WBND6iK7VDnp362
ypp+LLH0mnNpP/kRjMBwXlOXj/HEAJoTebvKsxfTMATI7MQrcJMQ2s/1xUC9R7ZrAee49wpl54kF
Y9P7Kly9hTDqx2Sdf/aiunAA0T5yc1WcH/M1k3JC9BmqIZAkOV6vAaOnDE+BlzgoKUm6dFFtI6g7
kwGeMF5wE7pjf+QE17wTX9w3ZSftVuFBscX4KSR7CzCEgFWHJhKkPd180wZ7PrbHMpQKIvTJFwZ2
zwzJ54AMpmkAWubbgbir3CIuE5+kTo+7vQY9ng8qVQUiemR7ZLc7ZMNEKsQ83AViF0mzHwmX5MMl
9PIlYPrulNgDiL9Gwoy5On1MFSuSftcWVMH7uBovHqN/Y6IvdobXZxzFWQLTjFh4bxVKji+3KCNz
Zmj5TyxOo2djAoSjJAbblQHtXYlkaflD25GfMtMfha6amSMhoCrC1tAOhwa9h0d3L3d5qBMDMNxQ
LbEYpsxMiem1irHCXyHKXemhg0F4+CCIbK6k9jYIwy9mNH499hk0tAecwV7gG9hF/IljKCWa5oLc
krBMmyUEuuVHS7gFFhv9FbQGtXqlZLt7W4Z8mMBl9lfVqWAKL4i6Fy2krr1RxDnht4bRUhwFBYar
RaSkI9WzddIl/VZE2YE60P37SStKPSNlNHokXOZGXoglq9Wzk8sARP2z13Z//PHOP9LVlVFZiNBl
iZw51XIV0dTQk9UQPFt7vs+8KMj5feSjnglePlUvyyd4Sy5CVl5ScO+NFSKcxpC1FoCV84m0NkKj
CLNwUszKyheHbi1ZqL17hl96paLrDZ36KJgZ1CCkPkfuTXLcZZEtn/vnYcjVj820ItzN31kB4IpC
rLbChU2+u3zoJr19HBNpSOV9bb1ffkE+Zu7ZtjkMLs/Nmit0bKwX16s01BFXCX0NQwWFyQrB19pJ
K/xtTQ1SzciJthK+igjA2CbsHWKA+ebxk6liIlAh/xYBlpWK31FZiG+BLKdsLhEp/Lit6vI2HEMI
0hPoAz1G74vZ+WnsvNLuLzSLr0gj7cP9WAkbX9U+7f90dJIArH9fiJg3JWD/5DnYRSEQqHFoD63T
s3oo41hjoT9SdXtq4I/HG4p5l+YXajy6qvK11cNUXWSNQD3mFi3bx7AAyvHDVW4yCOHpcn9libT7
+JW7c2iAGT6jwsWT2+mj6H9KGPltWhpiWARbkLQhlePY7xNSYBWXpBXmGV95ROSm3K452J7wr6Hy
X0jvIRg/7psXJ+wwhBnd9SeLw5nbAmJSwcVCiszkb062y33H9ceOjPs1+Tg5xZFjexPjYUgTFiSE
6rD1q47Uahzy9QMRi9Fbv6Jl9DqLNVlcFPlxQUYZT/fuvjxCnKrJgTH/qqQjmkVTxj4vIMMsJaC4
V38MvpDV4m/O6IVeYFXe3bbNod5JvaSa22L6KT6ZWUNgWiJAWzFEuKG4aRGkdC1Bzx39YmOzmkXg
zufcw1joqD5D5r1m2MHACDiurMILD68HVLE16iSodBnvkrTzRzj0VmB7Esg0vOAcqKddSQpD690a
gWd1BL5TUFBMRm8Nv5t7erCjw7hcnYIUsVQOAyH3oZ8KKxHeX+7puSc6DJJBA7cevUM0cP22XaUF
1tjeNlivSTL9dgmz1F7GcYBXrsmmBpkMBBuCSIZvgguXOqxB4HwBhdOV5ty44k+ym97V+cNu9+sM
cTSBUcCi3Qykyj404RqQkvz0zTAVFULY4sTOdPZ3qW/g1v85Hkf+e9vhlPigzjta961HYUc6RaKw
0ScuGtKVAHiKYMAR2nHwQlY4LJk146uRjBWH/AdxJw3WNr/mj8dF3ai2fVbNBfcAw+71iP/6Dj0E
MsKIvxOiL5/H2W0MrFUQuL/nxbntbTWohCNXG6f9bUMpe4VfiNXr4dixzMxOERplXdiAUoizv+sW
reW+gIUF6M2zlZDBNUzwo0QrIKJH4xMohV/p5f5yGRTyH0bgoIxusmQ08Ja2BA4hCPvIYhFrRdTN
+zvYLrMxyLP6TAogBMZ/8lLIv859HiXVILp2QKIuwngRyOGnj47dGQXQ3u6dsPWbNfauzOMR2704
wIbPpwu8/xexhwO0ldEZGHFLnpL6TKkYDdLnvIkDqD4/J4t8Ix6Ct38HJsojhZK8eAseLlm5sNbR
vL0CJxyyTqJCH+SoE7Jlx3tXt+CwWoPponqQrombE1zz1SY6B18OzPl/paOezXhccRzPXqZICXVv
Rqg5TMt1okgiEBsrWXHdbHjJKi9iWgfvTXVYDlK07QzNq/JAwNcpvXyypZePkRVDuLmkWcsBc0L5
QCWnl5B/k35+yancE+eQZJUt0wyqcv8ZKqQDsozpvsPYqHq0L022ZEdvvNJjOPegf1DPXn4vm5lq
G4nu1eJ/2QHrWOEqq812eydDquUd5N9hcP70KEPIY1lbmLyrfc8ximnsp6QzJAdb4JBt+OSod0iz
8yWDprXFaXyZgmJKhBIRNR7AuzMF8fki98HkBjrYlAQFw/Wlh5z+s4d2QT75/5LQDoAv4aftRbbT
TGfKYql9RQtufDsvziRlcoWTvbTreoACt/uV7YSy1ulkLW70otbUqQqQPWfXhIt+91dPg15rRN9e
WwcBSu8DAf7l+4i5x9YaznYimIfooLTId+uWE9eMCwMMp+ToyfVO7BeRim4Tu8ESnkh1QDHl5M+K
kh2pknQud32l/J10TNWZq98uu0HbFw+TBQ1qQNFgnfEf/qcTzjLMRwPRXr4Lyg01QQXwN50r6HwK
vnLIdxmret9gJ+GeeafNqV1mymit86tsjpWsZAudf7mUgvM3K+2i/XvSsuoewLLQJn4xOsSdKXOW
G7V0v6qK514zSdMerTq1zKmGmq8rRdRNfq8Fu6yCJPjTrGOlcr8KvztLgJW83p6PNJKqTnJiT4Eh
Nu57HkIH/Kl/mGPE9fsIZxnE6XjVgno99y5l/hXBP51kfFpg2lH+uMSJ/xhZvTSThumJZ0+hS2TV
DdM6fx6o5INnUBaOShqdagyEf0Qzj6rzWx8EhbcQ/M9XPqnXnkr92ZcefXQ3mWyvVKXGePBEUACM
/g4DnNEJz9BYXtegvO+kd73JE7rCgGRIWVdl4aqIOW6ojB5jvOEf2DMQ1UuLVB5kXUG0VHvg2BoF
ljL5ReYqDLf7Cr65g/7AIAz+sLfQbbZXWQLVWbKws2fBi1LMinRvpYgK8sHoJ7RBG+WtiuTBSo/J
bU4xwnzwhkhX41yIiCyyMMmVAKMUzmLayxYIvq25XCFP/mIySPhUldkjifLY0W0IhvGROYmeGHDf
upDZR6i/ed2DjVUdwdx+XoftHh4qPxSv09qLE12/+XwS9wMAewKa1ObwrloUi/SEtU4KPyh8g8cl
ETkmVKRGt8w6VcBKKXhnjBXyUbTBKXbYKMvwKON7m+6KqJWcwZ07gAGiTkwkmDuYAw3ayed0qMYj
/yFzl1NFtnBGOTTMIDp151A+W8F560zTM1WjaAOD/q8Ewf4NHMyzOe7MU6e8l6q/6m53ExUMbrVo
4Vp7jS+wnTPXEa4PGHmXYoMHT9FZC+8Om/to4AfgwVSmvVpfNhokJSqMJClMYddPcPcpwfqObZVG
HKAX1y6Ab5dcszc8Jrt6a6kAIvNg58uP5UfhcicHLGj7Nx/kKgSISs/j+GbeovSmcn4TXmXrW1GA
OlsjxxYoqlkdPJIhr4vNdiKdbL8DrqRee70j6lKSDwFnFAlXu1R8ecUDf74T9oOc9pMU/ToIlfPt
IbMSMHsI4zXoopM+GsoT7dOHnQdCrmSDELTjIFsJTo7s1Qf/WSJJScQLsIZSHGiwFkvkxINprbD1
ThQ4d9U7DKM/CJzkrMOmetOpwqO+bI3pbYrTVDbF+qVkxARqK8cv3sG+vlUGbvhSF8dmWb5FDFlE
AGlGOfqzWmvs/VERBJdkm4ChDfQL0UCvdlIVzry8vu8WOLC+516sQvIWNZR5iOEJjTwNMWB9amn3
2HVMzxzTuqgRpp57VWQpabre/LzmvXm8zrPYthe84CPzhg1L9PylF0rtXk4WUqwwVVa4MOHYvagQ
gckOUVT7EfmWN6wMIiEKaFPvLsoVS5+Ozcu/bHHSfripsTSuRHTy3jjUjF6LYmBD7w+6hDZ9hbDA
aIQ402zJIlPPT/c4pUZnygCg/4784b987HBvFsOb4JfqFzLIbBG8KiS+hZ/BvuLgQJ6rstYEaq9N
U5X8fT7uW9mdlQ6Iso2auea0Z0N9mgrrUlfgQqCG1u8EPV77ivloqR7EgMkiv7x99qurDUkZk3/X
aFkrid4/nuzQEeH+05Um6mQwfd3pJ1gv4eS+Ilg1xqPQRFzFnyMcLU/Nv3/BiyJ6dAwxb0FZCdlQ
0okbXn5YvEzFNqeYKUf4Xg1CDPgknK5J+D+UYm3CzNGKnC1Xf3HqZHPYVHYHHntCH5ICrEp2PJX1
hkm7D8T3ZhQmA1ZdPKLRf2w7YJ01mt+CFaGUuVcURlg2OONBCHDWFz9+HZ235VNPARLhNWWGRaxn
6IVH5l+LMJ5pABsEBWtvi3SzwFC56057bu3U9SZtkMHh/JRh4rox86J7+4j5SIuMcw4m+p3TYj/y
8wxxjbrTEyoomRaefJFDgp8BvO1BbOAsn2oFHmEptXxiRu47wE/pZ9a3rfAVCTNjIOtglE6mBHL0
kRC8tP5ERsAeD+1Fjq/c++Eo+BjlZThbCjLcI1EqYk9dYyu2nRh19/KeL/6bUGBym5qyNGZNJsSS
B2gdOrZscDOufxT4HXrQducJSg1hYg1F6JzlKyIGtLTH3pcZaDUKGhxutt0ZK6OOgrZoaqt+fzWz
J5yc03GF9wZRE2YnCzYg9nAlZnwMKq2ezZcnM9ifxtfmbJhO4knzJSV0zp3zk4vgRd0OcGGbIUQW
yaGp3QOqPUmgJtacbhV2OMid2y51zhwkWgSn2p0rEGYFFTCwpH1GcRtuF+DZ+Gbcyy800MEI+a5D
HWYwNv188sbkd7iDxLcxCzGqTntOYvFP5sJ/YpSO+ISe6bIMTZ2TaW458OS7+RD+wlzJRmxaZHdq
zP40FcnDk2hkn4pvmV/HYPDthitIrTaK7tQ33MfoPwSRncFyf+nmh+rswVZmUB/mjoo6SFpvpl1e
RelCr5cH5SjPnaWEc70YaOzbZ2wa+7v24dKrji92iSe4Uu2wGSo7e3vV2Hjk0KRMHgYvwdMN+XXm
Om2xr2rcbvKr8SnPUlgBsh86tPU00KZglMmws+XSOPbqzbP7VZuqJbTplsE0EMgNuF6u69oSHtWL
Bm9OtsDYEgKJX8XzH2E3d3u4fBQOWZWkY3Gk8BFF+O3GChwMyTgolw3Rb3cAKi3kBnnwh8YKr7PK
tT4sNYvkDMof8jSkvcQCVO9SOZDvCdUsoQqKZBuJ5ORFByFgeyPCXTp5ttanK7sLlqA6fTm2emy/
cDrAF65fbIvPf0+E5HmFlfYJLtV8HXl051WsKGdN3S57434tAMHh7ss+t13gQzJE/XvyK275p4ol
aNvb1jNbLWjoXzfomsxCnNN1HJPTB+L3t/CztA33PxugA1T4UhN6XgqsyTLsajH0mzZmDnA5dJCi
hOuuvQ8/KMyO9aHkjwZy4NtpCpIbHJojY2esgToDTMqi/G8CbcdbKMvfWtCmFcHAh6aCi5UHz0dP
7GaIavfL533eWpQsyhy2uXocXIshF6wl4WqDJWL2IbR/PDr3rUhosb8i7AaDUvushxh8qQrkKkJy
8jTF9R3QAxaPeXE3hIRxsJlxiHk32TqZ5eqCFKx8O6DUpBKgEP7+lizVmf5Jl9yDeIbpH11rmEXQ
VbikC6l6mPo0+GiS5ZdeVQWeEgCiaA8GgTGbqsDrObUWstw0mNNRz0aLAtJ7lF92DrWBuhTLWryL
9O5rAfQJSj62seF7cZU4MQv2yEcB5LT/0SoJ5NnZs+FiVTUHnukk51VJCnQ89gcCqW+HeWo869Dl
dPuJmxh2bgnArOCug+QFpQgLSnFyba7rC1NT3VjgEYvefc34MIokCAOpxVXjElHBzX6L+RIitjQ0
MGin5yXfjhedOgM/xgHSrguj/ycosMQFRbBQo2fh0t50aJi8Hqm77/CIXaUEWshQf+m5o4HQJ8BG
+9ugfNyNH3tmiB84ikPAS09hJ5QOUZ6w2WNXCZLaGLYXABQ7dnFLjjGLbDB5VcTc0bsA5nYJacVf
wh3azk2vR1lAQWsRscMlRzlnRhDG/GX53AcB0IJD8ZjSTg0bv/XU23oF014TuRt1O03AtuOVe8o2
wxeVEJ4BKbkiSmFXtj00krUCf1EEqc/ZZGnMnfkzQYlVFihHQEfuIw7nw+uuKuPc7EydCBHWZKqm
qwvSYBv4ajNdKi+MKp1AGRu2UnehEGNXPVq6UFryuZTU0eeRbG+ZzweoXlVr4gwf8BuefXi4MK7L
lgxT8/B5Xv4VSTtNKf1UtaknYctV1W/cLe+gFbJtzX8uLZMpte0E0728eX0gWY/B2ah1FQ/k/mIV
jzqFUGcA9BsAmqwXxpMVb8fZEW6zQ78tU7o7rMFCKgctYwDIvmowESsiUK+YScg01vzi/S8Ateje
EomKBUiKsaiwBSnoBQcjIPeKFqGibt5iS7icSWYQYfFkozY1I/sHS1tfLfadwlTLT05y5+7VJZ4C
kMdszNlUSyVXwzmvML22/v1oTSqNM5v3hIQ2UkheixmahepNdG+HOVjJ+SyMfmnU5cI+l3thVC6T
4gU8xK9cPtAIIvhWxxOQXsXl1m9TIuXcpQpCVMsbOTkuxrqjx+d8ROIg1e418bhOZ8GywYSwkS6M
HNUWle37wn981aPiFUHfpTmS0jOKUesW16omaxLJ3P8bZ7wB46bvcQ9J/880vGz/N775K97kwKCn
GkatXzvcXrctvlz9xEVYiBIiCDE/2UMqld9ulZzyeXFdSoGsNhsQ+efzAiYUXxB+kDkijUdY+U51
hzvK1u/4P5Zw1aX5XqAJW02uJLzbuyuyy90NY951dbXy34CM5T+0jcvGL2crAbzhOl8FIMWxvi/E
vCBm9TwYciYjnPgg9k8JFqkEDtmMnXKAgz6b7LlwkrSUEG3k46J5uEp3tkvnertYBgedzWP9nFx1
PbN+vxHpS49ZCEOxnxL5lYXcqllHwEMJwfexHLdoNa3JazDlBG+tu72AwnYWWp09GFNnNqxxUApj
8M7w96Q4mkPz9AUonm5mzNw0aXiW77n9V2mDGiSdea5zkuhKJ47rlLxAJMCHPPPx+t71dGLfSL6G
yLRwKYEz5x5OsH/h5z7s0TUBl4zQueMbdF3Pt7OSXwdRoYUNXt1fB/wf5Svoy3+KiLFtcT9joAEL
uPgyp9dCUdv5nxIRU8tW05NwUGdks7WhiJS3agJ6UDVY80+k+XbOcL+LVrDvPJtolLG3FX5sFj4o
O7lnpM2Ah6Xnw8nsbciDVjundDx0n08PBZbBpCDDyjBeNddDWe9IY9a0/IhJ4kkSh8ngmuMlWkIq
0sYA3DrKd9saW1yRtubu41E3ihsoL2NLu/ct+wnRzZoXBxYC+ycqSiDuCnM4uQNI6Cho6E5NO9AZ
uxxJ8BV3Wa4ixdrMdH2qLpXdnb7JyB8GCMiNWd5KLS0fSIGOnwZ4wHRNK/pAIZmuLWQzw4U3Xa/J
d2rCce60AWv1TeZ14pp1uK6PotBHNRTEtMf3Ureaqv72fuZQnni0fypmOtUB0NhocFn3t4HYxeYm
DjFl0+TYCV1L9sMIF0KgbRfSihhkn4uvqNPVZFEfiFa8/WVR/+N1rT9knwiBxkf9bAoSH+35/Lgt
Zdc7BuRYz4UeAjSzHRtR4JmaeYaEynYHB4UCCx0bNNvuK5WFZgoH6OWNTNDp+lblDYI9a7k/O/WR
0UzIjDazGQ1WJqBbm3pwp9Lda1yQyGK0+w8hubmrdKPkswofj+tA64vyd+kU77eVR9lPTTFrDiTW
h4rOT9eeUim7as4CSybRBt7+b1rqxsPfvOGUbroEGPSstjiUahjwfOBZo2mx5g7Vq9PRgjF054aD
3fVwAWuFYZ9Vx3B0zfPnSc1xvKW5q7+Pi4l0M8zmYgxo6WhW2XmgY+CKcGVBhxAXoyQXjKGu4l3U
/oKXJyod1TckwwZOLdSx//zdGWFayCVVJfZBE3BJuwWwfRALXpq4NbWny5QOsExY/Xm4dmEk3hwf
4JnltfJAfiGQC8ZkhypaN0Jb96hhx6aZ8WgG0yx+zQ0+3tPSlnSkZ/rihgVdne90NmasB9y1OWtQ
cB2B/BjqPvy8flr0mMV77PuhQriuPobjCl+m7B58UPPXeP7p79JMrKuUaGSxaPTBR+e6xhaSe9TS
nGmi1NtXXMb1JIv+iELgSl0a8dW9Mlgbfh6UFDF/4kY1Gc20WHAUI6r18ndSHOZ84UtnUWLqyEKz
/543KBb6ieLT74Toe9MaekN/ZyjnpzrWxGpSBYetRBomyNMnAf6ydBmwWCU2tPzVQEHwqaCqmGAx
PQLUGX2jzfttYvCcqjIz1IuTx9gXE6dDuPFeGtMxXdVJ5uTmtK/yCnDGX0bfL83uDa4HFFv7VRS2
iVs2jKE826Au0j/rD06cT7VuhRBsfd3+7oxQBLDZXXOTajg72YsuHJvwZHJP5ANDWJelNSOz4oee
srQQ9UFtcbxTRAH9oxg8OL4ngsK9EOg0UPck/GaDGvMerezooXnTti+Bsozeiw+jQ+NPgDODbkFk
zgATqF1bF+wIdkjPz8Nfh7O/hYAB/VRyhoFsQ76RM4UZ+I8rW/rly5pHKU6mo/oLmCFZ+gHNYOv6
3CPxx9EqrcC6oXwMsC+86zvKfJpPjhLawUbbSV0CBbL0gkGx0lLTWddkWLHFGBNyjJVvCipCmlM6
7zRntlg/mQiViNGxd9xRjpPmE7fw5w4QlEKfboUes8LefVkYlbljwose8MUOBa3aZEv4QfZJfj91
+MenjmMfU6o5Adoc5pkz5KcVxhpYK/d7chDHWk/mFdWUSpXFHL/M0BOCJ9yyGU2vJDXnBPlcI/Et
XzU4+95XZil6Zdr1n26irhJq0g3/YvEpvsYD/0YRQqVHGhPgXKugHDO8jAAldEz86HaqmJYKTnwb
IUi10ZvWtHds5qrHemMw3GxxXqMwuN9r6H2yx7aTVr2sPO0jli/8Mm4i58qpDtXDaou076XgyGZ5
A1YwWhF+gt/oXPEFkUhXvH4nFiW9p1h/u8bhSvgQ2vpw5Ajhr/GoLgrPFP+yPBoIR5OrdoaBEfh+
0QaIRy1ESq1FrbytPs3ymXSM6+cJmpuizGbt7yHUMLHr+h2Dbnooi5VGV+TVVWl98psf7pzYAet1
tjZV5WFNUTxTmbuUbCfazeg4GkI/CUY6/Apzc4x27UtPNbrWKQTZoLY36oFK/iIRWPz2MOKVKs/A
3yjHsIkPGKvDcHDmuBWyx4uaWlGhOu/kZxcC2EQgQ+ZZhD5RxbLFVyKmC70ealuHU6uXBYOwVQ7d
TjCDFTqYKcu2+VHtFG8JUBFiCXDd8j/A7Lj1z1vqHwjjWqEPXKBLzavF9GdVGVtFLnVBHBeV/rHo
LNfATSvyvWFyaqzO2IiNwZz7jRgJGWCgP1dXSc/SDzgomUYcIREsWxl51oXiWDNYqVcF2/3KMVRK
nUqXQVh+JmEXgGx9pZsTrH8PabBovFVg/VcelFLQsRXgiyHD0bskve9AHddVKRtq7PDobd+yhEex
MNoAUwj6PDptpNXvJTop8ZqnSkDdbMj+ZwkS72IAmEHsVFFvbfRC4eF4rFC3h9MV8Coc/GW4ya+t
DfucO+0EQQvmEdhvIdBS7BAEiQOg2MEAFHge0Y7l0vTPmTbwIIxTYTBhrB5XeFzZCuSQ4821sVBw
J+tA1YCgJ8ujKfHd3qCsBafRMH/0KhMru659vLulBmJqMSFfO3S25Uhs24Eu+vX0GP4HSuyI9wUf
QnbqjHqQ1ox1fwWGSTz/WO7m1s1TA3h4XiSudvmaYR8yDLJ1HDcwVR6laF89q+MpmIyHJFwtcQY/
PaWDtKb820+N9DHRcBZ9iKsK6mlFy/rqUtandf7VJiBYvTUi/Y4lLE7FMulEbc8uYYa/Ozh8t8zl
a3fLXMIF2+9R9+c5zqsHXYgFihaN6JGrrHKYicw0Ol3TQ8KIXFxkdTi5/YeVYN93lloEbMupFcnM
b8sz3BWZu/cmQsqbiWkW13ltWQIYqFPpxxtY89vcM/dZHfipc/XgpuF4AN+KAWQ1jPDz+j0ddccq
lvj6mDKBIqS9HQerh+Gc1ZvRLv+Ptooy2C+BrGL9kNH0DPnVkJeXP3KrRvAyUcj7HfapakSxaopz
LLU0aVh9oQtnkPWz6Ay9EuFRQGjIXH2PctREwzi/V9hAcMc43aN/3fuN4igP1htQoJ555ejyWaF1
+xdrQeJa9BiqkeYBasFizqHuVUyepl4y5jhdVzcXqyDrjS+tpDZRn2+QTaDf6jgt8gfGX3ilTGQL
PoZsENjMPchGSNcDIkTYw2F7zihojuatuIT/wJJhOvG7zOxqLomWlet37lfvuhnxQjB11orl3n4i
gPzTxMYbtUZ52tQeadZrl0BXHbI4RFAX6FuzvdyM109OA6ZgQYdDRSNU2K/yaZtMJXc4iIA3uUyt
rOBHDP0pG4ywghfcHiI9m2no0Wp6qpS5whZrCFVm8hh2Smf4t+uqd1Ta5aN5Ngeu1H8hpJzftNVK
FNFMoMVhtalUBYqzJdcHE+bI2+s2Cu47lDsELUmru4WjeZHEkBHPTmF9Zc/+to2hU3EZ6WaNVbAh
+l14fQJXn2OAyle6YAOi7+XsRNpbmtN0TokU1d0yi8bYkvD+ijktvO3Lp88JgaYsSKqZPRjE6pLR
8MGK2sEDVtSmdWIRPJuEdw8csr2li/WySFwRV0C3+JjKIYpTadmqn4LVYnNaqFEomT5ngoZra0XQ
1IGyVekBg428UymIGlrG9gdijQtYqaC2VwiX0ypIBsTwWiBL/17MgLSQH/SLAjkfGi2fcPSBQHsw
+7KJdPUaj0pd5bPisqhizv6nLUg3ssbhAak9YzpAyhYiAwUv7H7pOFlpvBR3l0fmxLImLCI7HpT7
adLD3lWPUnv6s1muQfJWNNbzyQjH5Y0sz7fY/RN1HBH/Zx+kqRYqTF0h5t63ZSCxqn16o/p1Bh+6
eYaPRz0cAr7+sXh089w0SZVrDQLHFDLIYpkZw0leI/8nAwn9Dc/6Ct5m8G6bZbacLsUvOxPbeoAY
ErY0fLNd+OBZpON+Z2gguISGivE56OYGBVYFDPf18omvp/IZucEfBAC9DQC/brUQSiMYeex2b29m
khE7+3JbXjafIrU15sWwaB/iDyTcnZLZGws+S1SUTXhNtojYmnKV3mIalbcswnNzfVM+EXdRqH3j
/VIndgG0Vg4h5tPHlXW8AdC9VQNiOb8pA7Nnp1tA6hR835bvImxRc90kpbjIRaWW6kWXtTBs9P1i
2CzihEG4iMeWeAl7SEE87FREc7nSIEwBvYb61vDY2rgjtjEMpVfOMewamOrDGnngWn9j4DsZZdAA
pmAffgUkzzaVdNqJFDfEFUpLIHeKzmTgC0YB7xA9nSSDV6o8jeyjmwlZtmeSCNzsg3BQZ6N5JYYO
4WjFzO59zSxWs3myul6EjWSCjLnWcBHXgHSD8EvVagpucxLMtfjoFDOsvynTWAalE/5aNf+ZkpWA
TDLvJZtHSXqeeQKSgayYDTeHC+MEhjFd4rKRpiRTAQOj5SjhQoqGxiFn/5xPkpNhUyhpl7f5CyNE
sIJPJz9vleJBrXSYlUxdqpbJr/G6B3oYuc0f7zw2hVen81J88Hd+P1rw1F8jeCdAmOgmT1BHZCub
6STYBY7PP7pu3nBtgE8BqDCfgoeOD+vFe5lCOAckLCwBF34gnyuBbuctkvIuaUYn3gIR2vGwsFBg
fL8ndeBFD0JDc2Z6kPorXwEtteFePZBFMWfrK013a/gQbsS6bM3Cq79doBuMhHKBazIZ3LLget0A
im2YuapOpv2K46kpx2dOfHZq6/0xX1fIoizCQMZ2eyfnQoxU800y2/cZziOXafy6mkTULrhFZqSZ
WUpBqAi4iBrgEr53NrfoSsQOLO+26fpQpTHBB7DBHiRoTVAQD1j1s5uGsc4Kt9Ylld9VHCOwM7IN
3ZkJcWimqR6yi9KTW+vBTO8rmk+WAVYAaqS/KB5n6spJqmnTeGHcvRVXJx7XzlPebWndi3PBDKrn
BDbaQtt7iNluPv5UE2unEQMFTYLZZ8fSJ4fDvD7FIjKtxlQTAuZ2L0JKCrnSo7PBZoq/EFWoXiL0
pdC8o3/6QaMPf2xKxFIbExFWD1sBmYb3NwT5IZsajvaugFo1vQM8cvkRDmA8ukYHb4FpqWqNbj/D
sZntIvm2jrBjnpQ+MvEbB/q/e4VOfV+PN8QeqvdsRqntFbN/coHP3Tk9sESSBxpXzAV8fH0fvWAc
ipRW1MYHEUzPHaaQeTX7h1E5s1yUiOLs2Eke9mo9anxdIMU9orpZMtnrXLOFYLkK6GjqG+NoyD8S
1yvpBpS5M/gGDOLKDn1+D3MaoC9lYEVfGQnNUQlqx4PigsUrWhIOeXfZrlNyG1a0R4lIStKV82wW
Fls+3xvlgnTR8u2DhWIvIIfmmidnazCXi75VvMChZKisEpTiCnTt+tdkBdOMNvXlRAz3lmBT5PuO
iva/7M03jLKppxvmg3ItQtVdg6RmpVUZBX17464r62UFuzdZafTc4Y8Psf38Y1RetY05XiaHxUcq
6sue21Fz71DWqs6RvnvYPui/6TnMOVO2qAbz3os8Kd8YmSLN82uco6km+z6aBChJ8bcWzwcPOPmZ
wU7X5RE/rwjWYQQNZmltDYRdsLVR7qYEW9xb6/CL10oS5wW8M2jpCkCplPucsMoKS57Fc5MT671J
Ww3AEZBHbNwS9JOambWcReg48ywEPA+dXcgv1thyBXnAmBw5f3uwdIHT2+yGuusfG+ewgnVlYcM1
LkgL5Zu1GFrftZFun9W9oyVakQ8bIfe5+O79r9D9WlKaVRjKhIC+w9Y+q//mkAWIFMY7Vf78UuL8
gFTkNZV1O2IvbbAqM9iayJBxJpiwpMhRD5yvCfMzEfErtww+P9Ak2SuLhnVnhM4IZvCLv2BFp4xj
N+FuufJwmBZgshX8eQjwKKwiXEGdjWmGFTiM6CXUHlZCZJrnXjPcfmQ8GJTvPQHgW5BuUbg9FZCP
w8RNnPCXSKijvmgoCXVd6THCU2LCLxi/RFmDUrNCWd6YgAuK/Yza8D26xdE0idpECAjxrwoaQIyR
+jo7ZC5AkFEk/izBGQR6u6LyE6gcqeCVtaqlxWNY8gmQEFJyf8wvzAtVCrrJdVFk5yLbrIXdx2Lk
FyelLi+WvHsfAxgBY0esOjvJHnUnQhep43V1vuZaCbcyIV44d/W6+Nzg+9+34OdyXVQck0Ug1Rob
qEoM1R3uhqmSTyEHtv3hTT5Lz7WuYzeIQanPxaQ7f8iZ2hKzcv5+pKecRqSi9qfEWh0S/aTRh7/H
NdP4g1pO21KqJsBBhdNLH1J1R9yGSiuLPV5sMrXxx0es9QH23r5aMBig3IWK/OzEb5dVzhTQ2sRP
iDG1hsvGs3H1XbaXMCTPR61O48HBnWik3kSO45qeyYz1h7UHWP3CagC5BCYK5vkQ0Ywum+/918cY
gl8toLTcyAnJt3p4Kyz2tH6lop3LU93yAdEeg+l75S576ksbWhY08y7Wqik1g9C1yzuMMpmoOi4a
pKce1peMHjaWGECKE3nPnstpaFQR3P6BsM18MWxr20zJ6ni2UopVeNShctRWUgzyipWhgzH2h3Aa
l1CN8vpGm3+Fvbj20F480QEq+yZtfvwWxRug57we2hk/TdCztbuux8xudN5AO8/W8OkHaInSW9zQ
7ydqy8NqHZ7gyzoHTqjcYGSe4XkCKbzfNXihNHx3FZbFwQ8uOHn2b5WfVZ+pgA23bcouhh+o/++g
uiXRWJZS8dRTg6T6lCXll7k+E8JM0PngmacB58MinW2nuHGe2hv4oOYA8rzyHbNvTrp5wQy8wJEZ
1UajQOEcsvsnaNZv1Edo3n893ZZw+BqsvLBB0tVFPQRvIsNbVhXTBKVpf1tQCFcnsvSNcgr0+QrD
Vq3gUn997G6BwTMFrDxPYnOvpdd7Xsw3GjyPHeGUxeOULWyHEY3GGm0Io0Rfd2l/QGkKKsV3VuGE
q4CaEXRKdUCV7gfd+/+8/so3lwyfQUaKXFlg0NEjS1HW9v11EGn2pxB79nZPSuI38sBK9OtPQXAV
2NvrILz74CwmxbzPgask7YPv8qCxLUh9OF4Lnfk+nqM+TJW6El8YfRVxmJtRn6yVqCoQbsdMGf6h
jKh0bJ5e5udJucUxBNEFwyjZIOfkaSrdIzVHsAQsaSXakEN5bi3DD+KBRJUAsNrUXreXpb5G5dBe
tr7rbmMqvXNUYFe5pV2BR5+iCWp0WuVz3CZ2z2BJIJE3mEf+ObDeYv/pDeM2z8/tBFfGa3IcQTsF
3+2E2DxHRTHcM4gUOfD9SSB1iHvivQu+TSHHP+wAdCSZjxdnTh/eybxzIYpWr2moT3foBfiaKuD7
rLUwnkNWe/v597rj1hhLqmx6EKXK60CgXJclQVllw8b4nGd2UKyJL3x9XcmfWifP6lO8ngy8F+Xe
0t4D7HdnrOl1Z8MkxK3GRH5FQlY7jFBpeAXVmbOxkm1SFfCBp9DxkkxPaX7uNamZOJYgMAl8JMK0
EKfzenQO0l+Yf+4dVOAviHVuoNzKDEsWYcQ7aPfk7HCUreEV1W/aeYwkihFT94CqtP011z+Bmo/f
ScBKyZznTj6o2s3hPmLNolO0kdPUaISYUDjuP9DT/9ffcqBNjc9zvyc59RyIqpuyu2e9x19cSuAo
2Zn7vYSV4MYXKwBd7Zlbp22WCe1vWSMOZYxl17VbzCSqYyxIK6tB0dTuTtm3IMTRQyr39Tmnmnw2
6h39D1GT0QSfHYI3V1PLRwFw/V0wjuqgwffDNfGGH6pgWLzRZbU6+Tt18ws3AtizLToyIdtzCk1Q
t3jO/Gp7sxVzo96x9cUNoaN8F1AL4qo4/lIaHDwA71jsTzDbWvxV58F5/F6sRu4fezP28ef0bLqD
m5JmFRKtmBWjK6hsG0rH7kh709zLgW9hqfSQenAVjhOUqY8hyHqZjoBVpTttrDOEdGE0rxr7N5gV
PYl0xrYVaFZCi7dwP9veAxzRwVotzoHNe60cxjRNlAPQ1hpETqhJyxUyEUmfdZtS2CQampCAir4n
xqUah9eSm3GGJ7FB0RxB7hz+jxwAMcbGlVL/mIxZcuck8rmCLhjOiWVkzSCEn4I3Q9jcIRKQpf94
MBhCP470z+qc+q9keUK/gxxEP+JQsbp0qNj7oTu1LukYNj+JI9JbYxF+pLFmKnuX0WyqaKZ30xvZ
ByuIvT7dWxDjwqtMgqUkVoWRkFCmJgxWwNXTZoo63B7z19C1iuCdgyx3e7a41KkvUMCytSDjsals
a6sFgSUL+OS2I2nmx7IV3ZOtDReawezF9qRBczMAWaPXfuBH/W4HrwQA+70aEn/38topqaHQQRc6
nVQvqcFR51VcANoXaA5lRdH9kSyJedAEhUHWMaUGvKRkN+grLjq1sUCgxTVoyhHLI0Rdah9NKzM9
HpC5A7nnPnV/oUg/2DwpZTZbVnyrxrnfSPesML3zq78aT5cJaWwwykdD99WeWMaJvr54lK5YARO1
8C3NVF6Ih9KUUYZhbaJDb0nEXCkKCfeAlxw/hIArVuImx8Z4OUmM1Cjs1wGeKEVmLDpJVc/xYtC0
fSpWhAvy4lH7uYN0FEofNQhrBxtSOfea/Z/yEJglTTy1ZqhQH76WSETLedqf6LA/HJyk+h0+Onum
cm614fQ3PWB4WZUW2wDvyjGZXm/A5ePd+exqoqnxU0Pw69FXuuiCMsT1z/Uwlp4yJS2Hoz4sLzQl
YXRrRX8uuPkSOlI4tD/427DIe1ov5aVeXhLS91graGnHgI2K2GzQ/UJjAX3UWt4UgnAMhBPYDA6b
Fn+PjhyCCQt43ST/edfckz8RocbVmfmyygQ+m2Xwq1cVDg478fqwjsCuZaCztZajUvj/k7GLlRgW
eDJkmEFNcJgEeO3B9lFAJlt35QRMEL+SIG8ovzsrtwMpGW0NoBI2pelJFZu/LkD+auM5K3a8OJ/N
B7vOB7mPOg6xr8N83TeT5kNCH4tHsGETALFQCKw1A3BS96xEy2GyKL8t3H5QlGEVhifO14jgWQzC
LhuXb3JFXOQghHgFvBZlz77qACadzWHSb0eeNQCUmbB06NrWnfgtsc+W0Q4tnxvJVrknKQB2SlAi
P9Q5ZOS4PLSO+MmTyKtoEF1HY1dKpN4x1EMEWa4GvpKwdUqLIp+rLww416hDuT3kRK+DWF12Iwis
gpZwSq74foqgvdbaw2+1P+1oVG606tSeS7Qhq6trEUXXkigpVbkaK8EQLTrv6NiGDK6Fp4UYtJJP
hjpL5bUSLp5wvigHowg/jBtUqgF/Y98Gk6V6XOlxNM37w7APl4NXhh4/JAk6r6Nt/YSmt8594qQp
BbvsC2S1aq1Tz5ZXZSVz7PYGtOzV3bnpj5/nlcgqI62hBWBIZbzciMwvfgVhPAbtJNnUBmK4ttjZ
JOJvNdFnPhUasA46Gnbg3YYpCuMNCw8ullNDeHCy+bG3WPW44IuFeSKuR+WZsy9ARdzSJcGHdmd9
h57lXLbtONa5d4FMOQVZXtxTjj/ID9YINZHnn9xlHy+4Gxp4iwI8r7aDSxO0ifNhZSLm2UNxwcgR
SVMU9ThPjP7bAHl2ppeCuCf8HnlEcGrXqEjqBqxyH7DMspg0MYFS3/n1x5tNXlV8xUhhi6oCjM/y
eDc6hz834hy9i1ivOwQLG76jekyvfj3Q5D8CgyZfDof6Rucb5z+ifnvURp191PCbFIFTr0wZzZus
2JSFHTjufrpUF7ND7aiQSskSsfm1lcckzCnWGL6lf6bNjQ0VwV3xREsNsZQDBQao8FRC4BPm6y/g
gcXTo1fXISu8rw4jnsYvg47UGzJ0hKlePKG65z7LO6F4CigjTLD1KiGO735yFt2bcsGT0E4A83U3
TaYnNBlAwSO2XNsbIcDmCBTZqgHGuWp5PiKgp6D03I5PZ9e/cthrSdU02QxW/MGMVQbvYd9vWbhp
BSz2l9D/SwswFLJnS2k4L9FtYyFgAcfzuHaxtrf3NYXoq2hj+PMTiDVsvloK5K0M20B1V40Ol7Wy
c8Sm/Sim3uHeX1FxiKQADfDXia0NFzi2c8x+/HStukyHQoJ5BkcvUoa3RKN/fmNeR+Fnfy3ZpxkM
yXg6ZzXMGLuI+bKRTdElmTlQVZ2RjF+leACsCDR8LdjkiD2hnTDfB/tlTKq34dJB7/G3aIdcIIFP
P8yDeFPeBMh8LcfeQWXF60UhwShhPoArNQWWFNpQxSDDA6upVowkeMjZw+ts+JA1/NWZ4snrPuP1
swBBg+qvOlFqymznwJVN/kj+WlTM+9xhokRmAwgRzgMAxymjzD8eipING1KMVnt62Dc2/7ke3yUm
ftT9df5RwKFsMxcWlZWm4J7rYlcl0Xh4b4EIrJvPQx/tEPriZETKgkIKLXmOYKaISlWdRhua+PGM
l+E+rEZsY6X/KYb31VPBOlqjndF3aauaVfKT/PzaCMhIhjfPQf9c5+GB4OqrY4I7iVVCfqRK/IGy
z7vcbP+ZLrQr4CqwxnoXSJsslES4ON79zDKVI214EdYC0Q9+tRmoEgnTtRPMlhEY1W7yxVmB22HI
cZ0Fj1zSov7r91D56Hk4668D2snTJs6JtlTx1Aw5tHArdXL3XplFhK29PEuYRVNtHwWTHtWcXcLY
fcGarA+T8xZ4aITUXADmgbzSvnkA1dLzaRkrNwSCpiH1mrmbzBHan3gcCsem2YpaA/01CbjBL/B7
9TxXr4fo4ZC3B5RS9QgIUzH7LrWePpuD5gbLrnsab4tbMQKsC5iUCsri82rOx/mOwYSKglYlbw94
/X03LQQ7Yi6dg02XuR8bt6G9ll+JC031t3DISOJOWNFY3J5GiSFnqBIxDmUXddCSF4k2WJl2kpWJ
G9Jjg6I1E+00AsvYtYLFupy53Xu2SOszJC+0aYQ0QEZSmZnryfPjS80uecHeXNZw3BmzKAqzVWKl
icrEU/ExtCg4C6q48iHGkEiudPr1j0h/iLdN0l2DFMCaJ3dHAggXcFydsUf9DcsfrtWRsNzwFvT7
upB71u/G59wYdmwak5GxI8h9I6s+60nwNkr2TYAKiffzJTcY4s1lIfbzTyIpmssKHzF1oNwZ7J6Y
sduDGZaH0WL9PFV3TXItsGVRQRmXtIAONuNRJsoV5R3sK532rH1hm/oDN2+mH/IHdEX5Au0Cb0wn
SzP4QV+eNxEyaoVT678ZpAlX2WuimS0CJQphXZuTWk1UycyZqZ9I65JpFDjMex22W273ACAh8ZHD
SlAd6LkzdVeKNv2UvtdJNZHs5ybtnvPZJTT3vjoSQj8Rqjthu8e4TPnf4KyMjLEcQ1HdfxcC9LoH
hdofqzHyfKxHAykJLU6TUd2NfWV+t0nU1iGY7yQkB7iIWzADMGkbMCCx6+vWBCtqL/syWleM7bMF
gNADNN9tfqEBqvZAYQLmXCDQhE8+6juqdLVdEy7s+6e5MDgcYoArAZ2vo/Pm6zK3Sl6aoobwxeve
YWeSxTGucTKGFCh1B5+njkYqAL++NaRRcG36F6cKDmB5QqC3qQLGPFS0Kzqp5O5zZGXwQiFP4H4E
sUAGtCtnL0sNeflQ+QgE6QVSSq/1Jc3W+0mn9v4jR8gWtEw4PxyPZqcxT9Daug/BaVuwIXRd5oU2
IkQqaQsme3ZtWPLBOwzTKMIY3vKfCEoeSOvPeQ2geVVGdBFxUV7gwhSxHAAE+3bbfeAUlzaI3Ehw
ZanXaS6mHbqKx/JNlpZyG78ONKuke/Yt2RkN8nPADsTnZILBpBcSJ8+VPwioXA0nzPq1oMr04vXk
J5Kruo2w/4g8cT/sZ3J9RayVYxHHt2hwQzcCOZ4UmlZwZRCmpL/ol3SG3EjsN+JojjBPIZyFy9fr
Uu5vV5vemz7/pB39Tb8wsiR1878PmnVmBUMqBDms9dPQAwizgPDV/ylRO4STeQQ28qPwcq4ub/oZ
BeqwIQhc9mRYfY1MwQlvT15ri4NPuDVi4pX8qutpykfCZOgIIgxTNp5jTeDKu7gGom0ZAXJesXeL
RWwUpY9MITLfMR/q4hlEeeTRNXwDMo1/Aosy4HXG0x1B2Xj3C2PQx3dXEBa/KbvT4nwLhPJ+ed+e
HO496M9vElbHO/xM2lXiJGoEmYBi+JpChrh4VVDh6AXR+iwRbAAqNaHBMVon9dAENNcqMHQLZr3w
0bQ2mLuypZLEMGK9YBzwo8p9DPlH2HWWJxfY/363fc71vDLXi3FBFECDwrw70rCVlQE/9JWGFOtR
zK5H28y6SIUZrDlwlnlvdlzcGGK8VWZAt89sds+yiFjKQEMCDDIMVdG/QAI7Jh+Owt+1pAluNCTR
6QFKqktHL+Lb/fdMdL5EJr1NqSJlJLNa1/w3THhamQiNGX5N9N7xGOkwY5ZfdfJddNHND/Tlezju
k373j3xS5qFLML9sw+Xz409/LAT7D7ZIhVefWnHWPtYBP8AJZwNlyv0eMRlKIP6JThqvCOJUzWVa
3lUNAtyzDpcH+9RnMtdxM5eQG0OOerXHclqSR62pjmS8bnNRkvQmU1ve/i3u0DAMPse9tVZsENLp
2Uuz+w4SBiJpIHcp7A7zvdmWOh15i4oQMFyIRgVXXiDZ5vV8QekoDS2W5foOPLVyGbqQVqcVNOAI
jIhhBfCVL1vOXcmZtVtWgCxmzwE97fUnoV1BqjDeh7QjJaDIaNj8j6+KkZAkn7D41ZDSu5/9kGjb
L4zk257enXjde8j6IK67lMn22d32jqrW7LxSwDJkvlRghfu8happh2bXnof/fLxAzATyHXEStP2B
ntJBP92WAx8BpG567b0wqCqaAucsU6CPVEdwRdZXn0dVbjvfSFJIj5PNWj58AzTGi/0wKrk+kXJQ
5ALuNWyhG6Ic3kZYNqpUmh3ALAWvq0aYThc7WrB5xGiNGS4OQKUyyLcUaoAQslOlbu3fllXo8gQN
ArjIm5/aX6kmWgpQpaH+hdPqZEl+ud4aoqTbYq5Q+Gl4cQ4AeadVzIfEb8UpIohLQJjPPLuKkSEp
B+1y+IcVkGn7xJaaDdNgMvCB18mHTVQak8vMumz4ZYKzHsVtdZBgCQk+zSWAvacpNTKGGxisH12a
ehdq8yACpGrtj5+KQSGdHKZejYYpqqid0l1U7azyTD6w30uythSldIEz7deAeGaRiWcbTv6jEXGX
ls9YW5gNWngdYPRLW9CmFlSuJonHvELLepAe+iqvjvBEvxG3kaspf1B0DOSwJzAUOJfvNGylX0GN
gKz2JxhH6TN4SESkh9Imymk5NMv3oLp1ogUB6xbdGN2aE6zsge/7M2ZIMu5zsRnqUoY1qtOqzw5b
0Exwsa2OK9J1pmBmTevX6GeCWS7uZ1rPhl8lhm8YnMN9R0PA/iAxVQPL4pFOYgaGDTXOzJ8KYNwB
nPB6PkRK3z4qVfUiYRqJICp0Zoap33vQXXvIpjy9aBcnezMYfwwuMezZ56i1RM/HJA30rt4XYbAn
o3QYWxrRQGvKDIbKqznijJXWsxPbdFkWtHEXcvb46SUwZ3lzp/kf0aBM8jW2YRuFIKtPKSWoE61E
/wlxuPCRgPyfTIS9LtVEIPysH+2IeiIdEEDt1XeuCCa7YzR1d2lN9zEVn0FBdaiTRpea/bWrsz3+
QoBUOgagz1kISDbGo/lLHvOdDrYfFZvoEjOPMcZPb4S8C35T5glhoj+lNBUAPikA3LbMPddTAuLI
/7lZ5wTPRyYIJWUHSiFG1jyj6QyehDtU/91vqbif6cO1arBdd+npoaj6qw8GVLfzDN7ggiH9pifL
c4kkZaHU2iT6bIP214pr+1f2jH4CmJIyEOhDgg6DL2HhwbCBhagxDa8qf1cleM/QnzbPHIOv3HB8
vdvjJA2+qY0OJhDgbMqDQ7K0viQlIznk6K3sQqArWUGqSbmVYU/U1QPbL9tawGQzVfwNY2N1wl79
IkjG3aNPplnqUWLqvbVlgPJ5lnNRHxwJG7BS3dFGZwd8HtqybO4ikd2ZjpHXyS52fHaVbYFgB/QI
x16mmcivwp76PGpUzK+LSNS0WE7xh4EuhJDebdm1ltDkwUnP4VBmHfHK+gOMn7r5UfXBWKB3wXgA
38maLbhT6Y/FgfDtp/ri3kUTZNG5HkmFKCQ6if1l4X2Tq+fODIXx9dnaLS5dHdCAJzw3joYAbcsb
tWeEwqBjr7p0V9iYL0DWLkA0Bf9R+37RcJHVVARJOeLN3WJCC2RliRxWY3HldgXcQt6hjoPpCBTL
VLN6Y3IcH4xXINhqFQOUEv4Aovl1UrWDCy4cNQXeRVtfkslP6WYwXiuTsf8cRoDM1hX0zaGa9up6
tmIldOm4pFlCRI3Lq463MGKBPnGDBksqLGRBrFkYTdhZ+VbwMwB6X4BEIUv4KxIJfvay5ui8Om5e
smsbEWlkRt2r6HyDWz+vjGGOZGploZMRiEeSey4uj9QeLUmRh5CJGa1xKRAcpFKyqbAjXpLzcF+E
UiidrPBWaCmTLShPLJ4yWiCtLlUZyT/4fT4+TX9sKQEtrFXu8uyQsrIqF5NKHDFQeiousNDqOaae
/PfApwVOsrG9+wZxQTAg4GE2uI2ybujEpiS5G/dgQ0BLD/ptD1LMDbn0Ea0wiCy9RMbArQJUl/sN
l3RCSTlL82ODNTlH4H2MFQz/ulgm5SzSrMzkL8Y16twIAVvSIweBmbiEaxxEuGGwnAm6xK74xW/h
T8h0FJVFahFr/vGCLUrtyvejoaClIiGOKHFgo31QEyd+NRHbTcJGbaE2Mbgr1iITjBi5K4KyiwwI
2Khlohw5FPW7r87YIjnU8vd73v2koBdRgqBdtokNqGvtVvD3RpmbVqZvU0zGaGTcsisB4i93Spn6
6nhgS0kdGcNuk/2B7sftM7ZurlakKOb3Ntd2T+8XmDM0dyAu0Kek35w/akNnBQm9PzMSqAESn0wX
GitwIW6z+chXBXZzPxtv4mtCIxJ6zSKiqStEOQsZdKRBq8JmY8zZ4Nk4yB1peZ0/2s7NUoDnS+yi
jaYxGAYVngHRdqASP4xb3WS4OhNaRcNl0DgZANoQ5xfBJ10LEGjxPBfoy2Bnw0xjS4AjmafbxgUK
YGochW3K3r3XtFc/cN6sEWhMJKNO9gGI8Qe6Pw092kbCGsT5Qnvuz/V54KbDoxg/lUWDo0DYXIUO
ffPBCHMo42xJApWeJxGrsr0CwCY14RsER4W78d8KsP5/XhGodrHjIijpvJuO2HZEIsch5SNSRlOl
Zty3fc5/BKuE5F6tAu4s4HFYCeOGMJyqIJpe0dZ14Y2sUtI4I86cCAGvINAzbzjiMr/CDJIDHRwZ
AC7DfaS4Y05j82EhnuijBh3vl1TOEAL3x6/Zd3j6/L584QujyZROvAyL8PAllaoC9mrNutDsjl2T
6PFHHO1PeijfXJwyK1zgNFFuVRR9C9blIYTVuT+ZtqxzGA4rLdb0lLCG9+7Y/DV84oW7/J6zcCm9
n2A2dfyeOEcG7dCYAbrKkRGTqSJrUAjzds3MfZRS2tT4c3t2FvZ82uFXar4TlSZ38PaUvkR637Nb
1T+z3zB5JIp/mi3VScQRHhseD9ri1mb8ZGP1BpDPWT4ZGR23viNKiuRs+lCtoRoBr5M2hbiR4J/i
/LJMaFmzW11dgz/8TH401LnkhfK1F0JmyQg82gZq+5rFYoyOu6G22a28gg7Igt2SPMXJFZSy2bMg
hHUBXn3VxZR5V2ifwgFdQCSrNfgqEwFQ4+QWsAkW1+xKg4cuUfZQNFJW82yJgZx/RR3ejMX+yZ0b
z7jUcbkmPcEf55D3Lgf377ZKkdtKI5Lo6HZVdWlzBGJ0N7qRR6YcTZQvW/LLAcT9EyrD1RtGdR9Z
rONDASf4Lw4u+OEKofB/u3ktwZQgqFDDPB03rU9iz0g0QqCdVaspst4pus/hDyjlexJfdDd/xm67
aYef3MxvIUkMlpWmVOKbPnw0FsUyAXiJ/7v8uB+E71AEYIs+kfn3k5JlHp0mME43j58gQg13ew7u
Jtcc7om7ufXsth0/XHPno942E3JYZeaXQjRMhyD1bp5MMrp57HPSJ1V8t9zY6cfT0VR9eqS6UIO+
jRdb476Awub65iNcC1Bf5tuXtq/+g80P3uNXIt2xtule8g0kfNPcAJRYSwl7GmO867V2YWJ8lp7O
LoVnMflVQIp5C+venVrNW3350470f1/b3GSMb1QRYsiyRWqXT7YcaygVrJzM791EqDx5PP76fxdx
nTxetFOqf7Qc/swWh8USLChafLmX3m3VD9z6+/gNMc72g61xiHqBYTY7kCJ2TZoM58/wzWY6NBR3
Rq0M7j+1Y4fTX98xnBuczR76aZUAW/392C4FzP8rqKQxxVKK1amfNAYcWK2ygDr4Hh+R2jvrr3G+
6HzW7pEK0dK6ati5Az69YTRaDD0N7lww99890guB/4JGdsc0oEsdP3IxkVueq5FTd8wW1cCzmjoj
HzrhIho2z7GL7F84VJ0oSS/6etjx4ao86gpwGpn+2qhsCZ9YPX+s2YBWnpwEtW36xdU9jOIKjZ+S
eBn2vOz5lXs9g+7XVSgzxHLEXHe8Y62jZvG9ImK8lRPaK8P5yQWlHKEmLBKuQMpNrpDNCtmnobr2
O+eJvQIyr50jVrZAwogJQfV6MgYcd97mrL9ExDLUK2pZ7ghwtcsbxzdlJ9M047kMjs/lvolyHvdH
YsDRj+IHxCkPePly4TXorCJ7tH+xPk8sOba9pAjEXpLhMnMsnQ+hTjZteyVUCL4K6GO80Ta/fXq8
mjLX4QTRTTD8N25PUriSj6Lz7QAToijB++H/DvJWXFObnq+cXF9cyzcvwMCpLr4IGvczQGsqQC9z
ECFrKQbMUT85BIUvA9amoa5KdX4po9cH5zk/i/mgTTZjjijr2d3+7MZW8SVmkKytvSRJLKD+/REm
SBE7exwLBWeD0lF7oU/7FRSSK4c78zXpZJa/fRHNidSj74hkMHvfcLKc5TKav3Y8KPI4qI57NaHB
DTWqOMpKs9BNNYbi1gc5HiQL8WKyoCdwdSoY6N5rUH/tZUNqHQeNMIfxl1V9/tEcEVc8TluMLP0H
oNBlDuvXLFUN9aKdq8CKWCXEucI7HoN27JypToK/7MNE8M7dd6PcSh+K5PpefwFm0sPf9hTUX1s7
nCFaG7Ev2RGI34pLgUtj1eGEgdHLlXedykuNJWtPBbQQZNHNpBbAjeYWnvzgDzvXaUARBNbN6I+Y
GnTPpV7EQQfC4lCq78kXUTtlSAloo53EhVlefYnZuCmalY0xCLuDSM4bldxU8cMKoLE+xrs4hGQn
+Q3s4FXNvqnn6amawLni/n+Oj9m2FjxUnyuyCybUBCh/PJuT7iPXKyXnBiDgl7fNeBN2FNl8K04o
W+roBYGL8usGeVY1WEiA1GVYo6E8d+ftujKaYhrqWbkA5W0wnJH/mK9ShDzzsYbfm8t45531OuG7
gfhUsPfnGvDTpyic954+EIinoHW+4kkzbl6FT8r8V7sKukxxyHsnVndICuiZPIyBItk5yVoPoKbN
Icy5npD4LcAIUV+f4Utq0tJ3hXQTSELBWgs6j8XEDwHCto5YepSLuxBF4txi9R3mx1XIzhaQ0zsY
j4VtmaYX7fqHXwEBi6rGjifyi9II9ja0qso3iZWyd6dDWHp07YuNAMq9Uipx3n2T4LCGQdNrurap
i+xmd1t6/xFK/JjlkQKbi+I86sAPcFFPcvIbGyGbgj45RhJbYRTCPvldC5/toqcO3Oq3lTlTp10Q
/47E7tHUzJ7FFpCTob8kd7wFSTo5zsPmPV5zbXIm8c405m0DYHalftACZzV5uapQSouCcZ8pVBLp
i8iDHhXOqbcozUHHkt19YLUPbXsRQ7lFBPtQRM2uojkQx36gtaoSkKo5oJ3lwQJQ6XR7FOCmJEBo
PM7R27NFwe0yAAzRSLKZI6Nwviom7AnlXocQSbeqe9eoWo8qX69Qsmt2i/unAYCihWKIUnFwZ3R9
hcLBaSq/ZtV5xH8xJ7GEJYvbxQpdZxEXsqUdWr6XPoOfStm+AIZ+Y/QxqxIHugNC2K3I7+j1HhXz
+gq4b+jzphAAwIrvFRctuLIa4y7FZDTTpIifZMEELCB0jNKEAx3Sr07hIylEFhlqqK0vYJqIbxmg
f3HC0iefJatCcUSmFkwDKzkTP7oYlBs5Xns8Ux1xRyk/9+b2syWAC/SJHhnJvtS0eoZqMw3LQuB0
npiaynGeebSafhMz4ab9yeUfVKbNw/qm6TYDR8HAe/tL0b6tAnhzoiUijl84qdpRHZ6p+86QaZ7O
7c5tT8eOk32sFwWJJXLsFgy2cV3XqGChwjZ8u4SFh0uZSSGnmaiFaGRwnQeXf0MaNwL+fE235vEs
IoNKOZK58rf/IOBrDz2R6+3tECPrnE7B2Zb2Q9dsr+mDqG+cLjM8B812ejQK/W//yqUY4QE3SAzN
lTUhGW0vSW68s/Uk7TOhOk/QsupadduAHmCrtq+KTEWFsARf94JodPOwFp3+awfx7EAGLAj4oSZh
FUy7VghpcERyFiKqUlI6MXCMDrUamA3OSgN1bxy8TSDumavTnGIl3HbYUX7vX1LovD7FRR+mMjk4
CcM7YCW0VT2ywbgCtUKcdGLJ5tTXek3ql8WVbXAYiAQZ2qqwmRS7RCthQ6J8vytG2l2MfdfZKD3A
PBPWJn+srJa/kmZcHCwj0vd3b4pPgVzUH7qT74cPR3feI4DRI/H0wV/npK1nFdcNMlI9wWtq72Sh
+uOSAOXIZ2w/rg5DYY3faledWrzEa9bI6x5YG67z25MQaXQF6sihs2UjQlGO/l4i8GI3z5FRexn6
kHTJ8pUltLR2bnMB4yHb9mi7L5YaE3boso0PI8eMtrQIyejR1+A3rnjhoIz4JeGQFKGHySe8XsQj
jWyPhqTczUYPxoNklinQSoV71PgtP9vWWCG/nGyskgIy4VSh0zmpV4x8amcN7To2F/LdyMk9km2J
gh2gA38V+QN6hKPSYQ4Ren1wf+KpljMZtHN0z4WJ+LT1ep4GGlOEV0avXaZZ/o5phnEeSRGpiPUF
Es+HLiCh3QYiEbGhCwO2YZk5szxVoYk8CjxwGm4juoTNPUpBwsZjoD3GiXjBYSswC6canNKZeR1s
/vldundhKS8+7TNkr/gF2AAPnuFralIKv7rVnn/nWKiGJI3grG79oi0CD4urHFOMdo04GZ3tWukP
Ncm8OB36O0RtPtpZ97PNjb5JXnARJ6sCKCFnJcGkedhWwvD6D67qqsfdeHuLKRrx1U39iHR6rs34
ifbZ/ozBRKNvqeM3i9b4c+WgWMTYuKh1M2pZna3bwTr7mpYsqpYvybOUy28as5E9p0UlsZLCDepF
xLTmqTO65bSusJVjMBjjwlMRgAg2oJW2/dpdbVtUTi+cF6ODvpoKNZJhYm1gqCwysN9Eik+5AS+/
63KK7VeV6cOcWD8ZsvuBpFhJANEvDHPnENK+utrfgBzzYysiRIUPTsqDGWpvhbNrphb0ho1XVPzu
Mqgm/+PkmHFg/4pOxU5KeUDjn0JV+txtLR8DRTuitCQL3wLuUxbtPxijpaJSN5SV4/Mig+dkdg52
invOTYScP7Zxog9Q5UJRQVfm/Nm2cwnaXtXKPvUIJ20+l9yq4YWCM/s2R60HGGmys3Yx6y4oKxJT
N2sMzo4EZemZeNCe/4UvJonr40VJi0X/JczdSjEwDmAwstPmNzbti/tShqjXpfFSMjYxiog1I6uV
x9zRWC3BC8MVxOAmFIsrms0jdp+CYqWbuSAJuQc7qbnu2UJA2qBCeMg2MOCkTeqzCQmhNYvsMWtU
2qi1vNaNcXnXh/12vpAgGGFII2nK29rfR2yRy78KnqyHbXzMLf04e6RgsDX7A4AbOvHYrywDhjfo
Cw1DoJs0Dl3nu6qlnj5WSpIUpOf06gNRZAvlDrFa9xNn2/y4yR9xwWL1gy9Ht+0n1Hqtg1J0/xyW
I7oVWQsKfyW8EEeWF4Ohk7yE677vPhR7MaHn5up5JcyzoG2z+JH6FrmFCZ1mAJRsBNt9gkm20XNR
iQmaxiQ92OMwZeXz+4tMg4AUGCpNms6gyERvhyoZIKSLVHxsw2F6uj+ViKfJtL1wBvmU1N8ktmfE
X+eAFd/licEAh9/x9hjDg883WzRGkhtLHTQl/LB3/pJk5V7bmbQLmUC+c00h8XNhlI1RITrc/nCf
9znWLBY0dhz8sJJFoMYOrJ7ZxUsBVrdBA3NGorxgxk94zVqHATbM3WCTlQHFAxlUSxI6aohZOtNl
PLplg05cdx8YRisDVsNwdJJD6PG381vuZ1OsKYMprKqx/EP5ngYEcwYDsY+YDyGGzJcVzhiKG+1Z
b/hjnh0fymvBxxWyfY2i86djzPy1hYE0V2qxG8PIsdPlR2cUHKwBOsuQ7/K3/OR0plH0QDOm88Me
6+I6uqpbuCozCV7yPTwTU39dSgb6fOLm7So81Mc5p88ZSYeNVGxV/HWxAd1qhKxkdHJYYoME/1yi
0ojimZhqKKQSZQE4DUfaRiVAy6XO3WSI0qVqVnu2WvVGBGkpNEB0wYEuDvnxSLyjpGhXvgEfG/kk
kI0+CZ+suDFmYIdofhPgwDe3M6bXy5y06IX63+tDP7hhoM2DXsQ36xQlEVsxVgew+SIsbXAvyfgL
S1Bf+hQDh/tbQHuC1K2USJ0LO6W72mSDxFFzzo2yLag6tIzogfrHHgOFvTWKn3ZuhbN4m346MU3p
lJPE/Qf8cnibcutbDnZ8LsPLLgsCkUUH1vaDQ9yMgOXbRyb5cp1Bc3AFQD8/px3AhMN7hB7HxMCc
V2cO/0nr+Uvmit4goix585Lz3GqfltxvL9H3B8mJhVkiRcP+CO70l/BSh0mq/Gdm7oUNrSQNLb5s
uAfHcgp8JbS67Q1GWY/BiC9Nmvg0l1tJFg7E2KPNaE4O7dbes4Lx88/yY9AifZxnGrHTxQo/j/8x
u+fvDiHfVXLF4fgrj0GQ/gOt/rDjjF9bzIu7NOX+xfblJ5S9xOnxuw8EPGnb8DgPIdAEmRfXOJQf
4YGR6EZdat95cizxMSKLdjf9MJmhjIma8EJMk+Ie5fesHaONcqU68rqYovt0PXBMkWjMjIYomUOo
56U4+T3wbqvH2zxieTQYw1AqqojSqHjFg5YpsB5kOTcC5OlH3od+6fM2GmduIUhb9ID/abw7W7uj
GHsayaD4sWobbymtma1OdrjUJp3eCf1D9Qp9O1aVPqJfHy9XM5jZEn/1OH6lc7vbajEQf0nsPwM1
4uEQmkXI/awhxn1o6bDDqszuhel3GRv5fSXtHgtr+5H8UvCOGbBTnH16S050/BhMBGIUIX/FcykH
eQNtNa4kJORZ9gA4J6k/AITOpXJsMRPm1ZYJxRRArl2vphtJ0ncxhIwq+7E2r1t3Ob1ib+tkGXMF
FN56e1Pk6c0CgLf8nm/eUjo1e2YTqbdw7j7CMmyopiWFO/n28cHjm6xloIIHpUukFvz/lvNngeZG
dgXYS7SGOvye9/eqW5sHxwqC55r2WA+idkLXjd3aPe3ki1f+DpzAV1q1BoK0YYi4otMso9pCOeV8
ZEW/wA9DP0jQzFtPEAlDfH36WXKsipEFZKc18WP7QAOV8MGaOHgp4EqOOdVBPpeBaHEJozFso5JN
PBWzCPrUq4RVATb9fH7nQHzrkq/9py8DwieDZXSY0UJWBDo/uC5sXe6RK0QMM1menxqk5vP4uonj
grvCllMBdHJqYqJf5jeoGRnL+WMQY/rJKKHptH91oyqYBXMNsxdkXVslCanVYdjWLYuudVg4C0Eg
WJzn9hY12fegjA2+r0YxQhSfEIxz8Tbod5K1Qv0Na2c/cFUn8Nls162x+LygD/Gs7mf8qowPu8C1
lBG0FJ0QBS3JpY/To2U0CzuO9ThUgMishZ7pVPh11QIxlDcx1jGl4k4XriGsdmMkPSczsU4i0ot4
kJ8xCG8Junk5I/AriIiRaZieBilE1d26DDu8EPOcZDnQv2heiQsmABuW9l0CSc3PD5ZvOP1kc8rt
509NwycQMkHvD6UVmdDRaCpcV4GRDgNPQgpJjx6TtPCQ/7+XUDHN68svORAFW6RRuQbAOTbN83pU
6ux3+3XgeQVVW6mtgUEfkT+MdKPs4IMq95AzNIQ3WplOhYxe9nsfmDtGTWNhLrxXv+/+PJ41tj85
S6RkdPxkaZ57ia/+HkbxBXUEm2iKXuh918cLeyd2zy1wfHBL8N68KuQPrOe3gypjNoO30GCCA0sQ
uAbXIwuGN+HxP8SyPBM+8IAguKOA/+7A+t7NrjwHmtMqUUov8PjL2FmcyBiGKQFnbUiquPUkvMM0
xBnM3aSeJwe6urCmMrMGP2ft2ti+2drNkFTAztyaaepYuBsz7JSWf/6/CI0TDPSKwhuSbvv3TAnv
0XRVImaC6McIHNIIzNrGVXlvSs0HKlwR7EmWvKbLQHMkZZaUiJWt0Mp4sLcDTslxGP+j/IAdUpZC
vyv2QjH5ZzC/eYnFs+0d6zn7C+L3sFuj2Q7n6R3d+wguIGIM+j043G4JAb8EAgZSRuWOAaT09yRb
4+9Lv349vuMoFAJYQS8BjW1ULFVvGRaztG3/jSLkXVRdx9k8NJ+EJtJnIvjNVGMSYmeXFBtDhTCt
aIOmbtj12SCGs9+qE+GEy1N16vY7W0zIZ/vI4VDfHo3RASHIFf8suCr6r9R83nm46D/u/u/dzUqe
IxPBjYrVrB2YdYyBov/SizDbwst+h+aLk3pJdTxSGNIM8K88G2x6g0AYldYjsISraBmbQLPF2nDd
2zI/oOnLM347ROF3r8pJDJpRKgs+vggyBixa2EeJUseT/j4WsmHF/aF5HKZb/kQs83za3m5nxamn
0r6R3QZGEnO4oSuqiShKdJDZV9mYJqrmNAfO3P5ZFLqLQQ89VJWTXtSYjniqlg1eOt3wiObzRRUg
FxPduSzl/+oDSAdRwKEZCpm0o4UHfQoVwjRQ0CY1S3IFiH6t6m/sprAO2MEJprYTELzpoBwebrM3
aT2FIMyWN0lfGXZB6y/u8kOzWNHNFRLwtBmxQP1gie6zcpGLIWyO24xeYjkYoNgmiuep7UVNKZ2t
vbIeAbwLNp8pxiNx2kzHy7CKaQaZgEWNVrl6/Q8wH1o+zGFSS6ou9hdSmhk+rOFLoNrHPuog60Br
3AsZfulHdWf8SLqR03plcjZpCeFdKnwru97WRqMoUKR4Ic8jdRESwzNJuoeREDBVVbqnENwNikPD
rSETVkfj6ufBR29eQPQZeA8q6MQglRWkRJSYRBRFJRMj25eZX3rl4XTb0S5fWfWCSspyTmbRKOT5
7sqBwDYXn96bDfelvkjIN9Vov16DDo2jPpMdO3gpFqzmYCsc43laWslIhgMz/QEeR+T3+J+Mfjwr
//EOEf03yLC4T1YyYcqXWs6dft1l9v4wFQZDWFvPBib6M4M/PxDKjbLdF285Gabe+me/dmmzBXHZ
tHlxWpn25998OUeD9Ae7JDCoe2eidfPI6Rz9nyC396bBeC/yxXOg7VX5J+w6m5D/aPzVNI3pDH97
xdY5ShPTM6lf2huRuJ+xSApDMb4a41LQTNo5oE6D1nSc8buxj7O7MeM0Zm16APzv8k5mA8P/uRgb
1iAwHamvVPC5wOfstlk3iJ+xikRb6jPAIBsWHlB6KG+uDGYO9vU8wSfQ156FCqJDcWNZdiGTORCK
Eye8Bx1BvsRoGwSYb5dpWCZ8RecAocWF3s6AewF4UXU5xxGkyr2VgJRtE75g//xZyUbFZlj/3L5Q
j2pr/8p3GZnTIJ4Mftl/RUH01sIrotSoMI9TJuj5QCdUGdpKFCeO3DehVkF2jDXs5SBObnui+kAG
yvz+ZS46MJoOZYKSsNfV06rs572DtFHR8Ydajxo/mA3tS+giQU71B8MI6nwsu6czjx/lLMY8AUHQ
c1tUuhYwi0JoBty59zmniDUxTVAel51V7ef+8D+sHgQ7JsepLBAz1aT823bhwXbo+8AHEwojYmkr
LmR/MQrxP4CdPtoozJzNllRnCvD6F7hxunb1uIyboDqwBr4w4whdmKALlCGWpWg+3mp3G82wIWQ5
OpORYmPaC35fku+y4hPtPPx6SYA7BEJA0IJKuS7/zwpBVs5VKcVV9Kxlmralt7sxGM9Q3LwHHvKm
etwdL6ER8fnKaqCsyDYEiQwRyMkY/tAvuO9n3TnUN8OJuXhf7mtqFsxf+wTccTLTOnEafn11XOTY
TCW3Q1Wzx0j5KPWlE8smxlWQ+ic4MeGK8MmM5E8TSaKV/2qrHiStHnLNcaUTF26ruxmCjXInUNSB
4vLBeg1YZEbvG3LRO+iz8bHT0M5nF5iexjrT2aO+h6eMsCXaiJ26rQgwI35ZlfnK5qlOoE1oA+9l
sej4ynTvG+Ts+KBI5sXWL4x0yyh+5tC7oX3mM3HjHpj7EzxO349cVx37xTqTR10qySO1OlH+ACLc
Yh+XEA/oPs0xRwAIHh+81yF3J0n+mGMTw11TR0Itjj6KPN8XOyuxEH27nK/gbBSvr5drDyF/s8j7
FHh5hun2RnlMMeahHigHXR9NFBxSzTsjIrat5WLKsnm4hJjzFO5iWBLfkicpUtvr1dV5TQW2dEgI
ajOw+G3knSxd03ARD7O3y2/9Fm+AvvMFYAo7CmApNvi7QY5Sui31CqZ1VsFUU/32uWuYKr9M0rWi
VY6LAIsM/r+hkq9z4SuggaaTFhL7WJOuq83otwOxbMqY/yOWnPHQ6TYVRvijakX7bD0cUtYBTVsC
1mx+v9w3V3GkfEa7jFyYYgcVWyedGXpKkozWb+tDIPhMbuBO1a1dNnmHI9oPORCHNEiPo0vZh4GL
elY525g23ttaBNrpUB2mUcZLQccaROr0dKDR1iga0uH7NXw9o1g/CvfpnDiEo7p1kMjG9wvqhTZM
t1Uk8G5Ihi0KNoGaLPFxQDru24YiGF2v2U8S4UZUkHxFYEVnbvSxOOf0oGZwfxUf1aEA8F1SOHSk
WglzC81t9Ml2yXM5Y4tJPh7R1Kdculb48J8URx/ap0vwrgQg+1ZFECx381yA9M3g+XzN7dh70k6Z
Ig2SdlxsPU3fdr4Dfc7m/3qurtbblAWtc/6Cr3Qt9rojEuJZxaXJDES8F4eS2VJeQ3D4y+iegJD9
IgASoB37byk/cOVKW2MSy3Ri20CwE1b8+QJxfPIUEvrquca+NV458PIX7xtE7/oNu/DumZjpDVBf
8l2YoZ9pLGdCfh6qWFP2pt0ZYpbPWeegQN47socYyTblanK9uR63lYpHKspya3xqsAniCiwyTLMS
+qrlphILWVa2w9f2zgi5XGWfe3ofvHGcIP1U5AZxLh8PrBH9tG2K7l12wcPTWBQrY8g4gvDAa90o
4KmAKO9XGsPwu6sO+/PfwqehCBpWGzIw5ZbA4R+qJ2zLhrqzoRF7zvCs1xILYMC4CsHNwAOhNYJm
VMLBpXb+Qg7JlFy0GyCaNABTcvLMZzugiqz/Ayd3Ycynhp3i6vnfDg3E4K8qvrx1eqk5GRFlHFXH
eTZgTGkNsMPqtp5pnFFAaQiillCFO7G34F9wKpx5JAddyKT5eoJjqtahE+WN+VQjxubMuWD73ge0
C0DPU7A4OO++iBpm7AxERZrLJ/6zEkeOUvUMU1bOz3S3EchwxsRTn3ykjKmriUDLl/8BK5l9AwIc
T7A8p+9eXehMqOnmiv9AvxsNQLd7Vykuej5ru7i4pqWY7LLJY5BVZikInqUl2OXcJPQwhs/1AGK1
xqQqSTcu4dxkv/b8+1iUgNthPeCzD9uvovAgDLhldInqyrFTm2rMz9zCKd9qEh8mA9n+5MtIEuul
IIpZ78XtblU2oKamj/asDBnfnuQ0kZ5gxxiN5PiidbGqj5V53lm0+gjUuToxaiDvV9VIcLd6KmE9
dbzLLG5yuLBHJN01k1bSU9tETp/JxKQxHGbg9u/wSaDiccJBG6lSpojAHQcktPcksPlqlYN4rPm3
GotVaycYkztsgDouGu6I+k6qP3sQjBRAWsn0u9tV4hiNXQqmysfJBaV/JRtvI3Pii/qMA2QYht51
FmSrXN377stND+PekL3ZqetmC0egd0Bu1eKG/qes5MNOTKBCttFnW3swNdYHPv7YWJ5vaWalQ6NT
qOspp8QqX/fVHms5yUt1t3B9368ASS585iCmSN+S+8BDlJHj1stI7MP3iq3yBPOC0wQlUY4eawJs
0l2/mqULBlbwE4hj6Qqk4cqJ2ptVqrnVkdDEXl3n0Z8smXGIJgpu+Xm/Zn/v4Hs4tJBHN4q90f3O
BHvy15MGV8BSA+2lucy6ky8/yKJvfcUt68kcMkSSv/FrbrE4F5IQVfvXUBSEj4DqNrr+Qdxz1R49
7Ig0t/Vlmb3X5wTAN+KnsQAZgOj/cblWK6QWQclfJnCtkBR/hksmmjswSDgstp64p7Px/tT1EGUj
8sgPdVNTGu2c/qK8SoyJMzH3jMGd/8KSHoyjfVWjXJdD2ZtHR4WkDB9TKVb+g/2YzDRXXSVgz86i
D19Sq/Md40/w/OcyXReO92BRKNJYEiE8myy/TdiXrJNeEVavNNbB0D+GHINlLGo0a8u5fttY/Cl7
dJ/D70LBwrRvDUZk4Cuds259M2lV+oUwMzVQNzAXmTrqidTBYZKnbPLbAwPBgBQqlL8Ko5NAlEt1
MeENtqatyiE6eHqMTpFUqsC66gCqp69N8cP8OQjsuiDoyIWfjIX7v10l3sznwNlqkxQa8FO6pA7t
7yltWJOaR+/nVMXmO3l/88Rq1ifzsKgsX6kB+EAOuU2AdUv1PsSuvjpS1zDGxwigZyX+o+rQv58+
6fKZJShG9ll7t5Hgtfkie8442LJKwkahad+a+HjpWOSlh+ZWlnNd5cc/PZiZVYAYI/DVT8321vqz
6lneAkPgZdokOXWJ/1WX4VneNsu+mJPpWXsi3hR1aW7rj5x6QUiQ+h3uMUCtMKi2JBkb9fyyVpAI
btSjt2VA0pl8gt5loGqcMxUZai236QL2rr5cRF+BZflYfwOBUF/fkrHeE1AvkMSuQq4d0mLNEoKX
fs0yWMjCXZvoHAGKD4TZ5jDCJowE+Hcvu36zyRedpmRWa7YQBRJ/JDgcB2WGPuyAhjCjLbJeBhL6
xTN6C/20U2kWH6GMU8VzeNtJg8Ad39102bG18YEvS44ECazvCT7rlUnTqWpb3p4R/YZf/fVoDzK4
IfyGD2RlbBnVZTvCtxKuqUs1hink00xVHjBTJr3J2jZ86wvZvyyZ5NPEWsZ9YSYNFutAi3Ltwyh+
YW7pt1fygGPSsIFTLX2y0XeFCwTvzobgF5nS4f/dsD1UhdhPYZBKpzR2xDceXKtqvCFbsSdWcHZs
RNDFE69hF8rx86OwpsAZRmg3aab+EnEARy5MxoZMGV7l+I638bviNA9pJd1DBt5RJcVwLHcKDhtn
DkMOM2TxuLKF4/X7C8cCpDPcJOk7sO66BdqN8GOtbIqWXH4DUncTvDRAzrYrcKOmn+1FeLV8oo3n
+pu8RgaQ8sc5Wy3Chzj8vb//ya+khZnrHJJo1QwfMU4peNE1pGBrl4YL3qgGG2LRTMIV8vgavFSb
pCo3ucucLi8YGIPtbMyqQeWgq1n2m3wKJ5nCJFnX3sBYxNu8VFkq+6XbDrLk65mLB9DZm8mz3u3q
q5cRjBMOwMyTdOOZhReUHKhKWcIn2ySs28tfFn2hqG1lj5SIMN4UTXJTWuPNZmsx3AmjvZKtneHF
0sIwEUxo1UezTh+HkETLiK3LyyxBF7rPWNEkOjC81yrhPT3EYTxpCN7gxBytkiKE5lWllv2lIwCo
JtffSbWRUoQXjoYOY1ozQzTb7iEa50p7di4vqlTBIUIeuaP65j4gCKy0dPLdgxl9h1RFRUqpubJW
Vz/C6X/MZReEiNCWN4Q5+VgeJyF2R3u8NTL/dgkRZCrmZ6S3K8tRDj5zI96LG6MVXO2Ufdb47f7f
GCoLoNbpL+PwjZY7NGOUKl0iwIyd0pQ/iLJhosQTRKJNlUv9TjklodQwTzAy2T1jNZ9gz8CZ7LTR
IzIDOI7CS3cYsjO3LA7kF2OUfmotQp4KJ/BEsGPig1kE1qapMN9ag/xd+t3AE50MOiVbY5IO66ls
W5i5/Tu4HQKd0cb4JhRwNpP/Wua7VEJbJDTws3Eq/QTBFiIsjfr66Nta3kcLnaJXqYkIkogcHlxZ
9pwacNimqndeuCRi/titxzriWUZzUSVZxhk8/9n3um2kd3shuRnFWkRdIy+WfKwwsmoOQr0mTyIc
g9iaHOFp4dRW4+SDEWNZwXlyLmvRdyyfIyl7sjO3r6OVEJYgodZJw28EiLXp78fW5coDABy/wRUy
cXkN8vwMUaI4L7dv9OxaV57yMNuBv/cURq5kng3DN954Rb/vgef1alsnY/Su9ZkVvWVJrAOywHXY
28qALL3SBG1dYOVFUn3cBr7Dppsk9El4KYlNRkhtQQjqP9QwcW6P1ph15AuRvE2V7qkUVffQBHVs
PEvScfcGnXqEgJ9Fsen6I77Zk4EVxykx5Ll5rOnw6sQdQ1aw0KbfxiXo3QoGXBjvn15Enk48g5G2
JFhDlLJ1mMOniGR2hyC0s3mKKH4cSQaP6DnEZvNOkgIB6hoDbJriewcKuKWTbGwgnCYtdiUn48PS
SoVXy0pdxTrfthbem3Jpwv+NXEZaJodJRb7a3q+gZ3RHgiDlFcJpsgLzRusdXts5Pxwl8NKF4aRh
fMkBN8orNUdNW0GamrTEU2T3gSnb6SBbgYXe5vQuAXRViMIajhXDbfj5pIAQDUuqrFHAS44BvOyu
ValwftLSnP89vrHtQ/aD139eiqHYHW26TLAC4eYFjCJt3IM2L298zMpoIZKXAyu+jVty8orhpBN6
krGRUI+9QPVDAwJnrXGUtLWMoEnXGgQr5CHk/58Z1TMtjo9L4+QimP0uaNRJHjmqAwxf3N8HnTyg
5LbTqruLJxz7pPmPISxviE9n8vRkYUmLZDWtHDXlTJeqF/ixuOcc06/tCQJbi33H57qEceL3HA4+
mVEpx4FZ5wLLAx3u4KaDRvA5lC7d/1Bs3Ao81E2gjb6FoKMlh2zRLjLqgDhHzYm8NqHXokB1MLYx
EE5UuOTOU9utRYVTYtcaHoF5KTPc0ZiyXUf5bcfnah5fFzjCLewlKoZjC91w1NqOHdWriDrCznUo
fZa+vBT1qDRMkSZgX76ytwtbKV68EZ8cB98FyHGkKkuUevuoSgI5M2t5id28ze499RtXMBjd7gXM
b8WIAXFj5gF3FsORYfJesqM0R3LxZDk+SOjmkiy+MsA+W5jbhgtuSNASlLNL4dIMHbrLt/x8cX0g
CMhsOhhI0/7ppq/3C/H3eoZ69VjL49WxarVA8nG/GRpuDzznIYehib00ilffnx68wArpj/KLV1Zt
I7YFTfdCpFYTXDgrD6hPWiCiErV/jSzdPfu/OFe2LtPUpCMJjOTenIqNcUlQOssNDjKtexEkSQfd
kupbkbSpnBhAHBzdX3ZBZY/wSPsqutnWrqsZQqEIfKw074vOhjvY6UsmznmjE7uCv1aoslT0GnY3
/p01m66oBzac7f+qD4uJkIGy69XfU//s+pHwbPF2R3Rg4GHF7/qYvCsrVlBN1G5DvVZowLtVZtFe
l6fsVcObRajXrdiUa7HXCVm9OoUYw7/fAP7oarlhqA239FpEhRHXOuj4y4UCV4TwgASdIKZhxlcw
NQ9B/GGGhnkCVLTXxsothabPj0X8Cr3oFh8utWBFpPofRbbc8v5xB6ZghchHstzPDcp9kvHi/M1+
5U++LA6QiNJ3Y/XH2HEdyJ/1YRC4znxZc4tSuNww6Wyu4pabjkGmDgjDTWeJSlfGttPfopUTXd2N
iTnnfE0EA6e1xpYGLM/rYPjEaMh+gULDSSh9/nkIf0fx8lGb6SX7Kl9nIpC3T1GYDZ5ZWfUJL99F
Djk+99Rk+n4wOoUxhUbhJ/4gQ3JM417CswC488l/+qVkI/xJzp+2nk86CXt5IBZuaFKDTF8T/chw
w/dNA0+fD5m5HkxBieNkZsyW8EOLKiV1db9XYEzyFeVlzNKPa46yfLO9oqLrg8nmlKq3S0ghsKR8
TGM1hXXriC8/+pvVr/C+u6v13DpzLSTZQqG5DrcvGH2R+966oINUXh94KtmMbCzho65ntx7SpEFx
53iNN6XV/jr76Fg7qKklBcMVJySHcgJuwF/M7sryV7H84p8LNyLjeBVpQbEsTu3cOnLu0QLUjg0M
xX1SXQwTbXFkM94X7b/D09lkaI74oOWiemVqDfem5/RsJP/swQ5DxXK3963IxYGBMca2eBpe09eA
mQB9JoRwU0DpxfVZeWa360jP9SREJVvaaRt709Io291tEpu25d+ccOEHSY9XlgtrU7ErVPcpCskU
/KIzTn0TZlRNALGFzKZecTpYlRSa1xoZl/SVe8DMu9JNHzaGmD4AeVYA3Nf7EKZz/D+JNGjs6WiE
rS9FzDaci119857slp1PZ9omUYPi+u8MMtM1DU4vWV5hGlAQ3bZeIESm57hnZAMlHahlqx7QYzWT
ZPeJbB4W1A9IAeI0rtW9Nbii5hYAExllf6aT9x2fw6VgpodFflXz3F1hMFPTTGBDDMKVBhSVeJIA
Jim/1NnaUAlExoSrRt+Iap+fFz3k9wy7cG9P9gSel0CzsvQAtQUIlTzeO4HYXtDIqDXMa4KMMpeW
gSzYsmCt1l+WnrP67081IxzVzOPwX2bYXqtcq0aDwtIcnPM0n98nxc/3Jb16Y3F2qk80/eLls0xX
VwW97B76od5PVazSqRClUINCSiyZMa0ObJOXkpkv2NtHrtpGoJhRYbXoX+a+lpKf0hn/J91oU6oC
24X3jUnRhN09U4JFO/au1dUi+z96fqP6FtFA6IQTI+agJB4gtorwWd8V8KJMcbrzJoHMa90ecJQm
75VssT6AwxeiREz2kBR3jFNkPTYGMWcvMmu7Hlwir0lObQq2GeudE+fE8tWyJtdgT8p0H5AiyWSo
BWr8rjTNkg00UyMhdcez8wk+ZxOeHDUXcVGFzmeJHosVJeaNhtTnGLMPZNiquI4YQe+Xn6wtNcXh
M86fqRQWbnl8qiepUR7w2dV3+8APrrK8gnWLffYFB+uDNWVOowYOgFVKFOmtfgP5IHYEt3XI6WxG
NfKI8y7zAkm/yBn306CRQtJ1DR8iDZ+zeKXDYgWgySY2Ld37nswl25BcfmybeHi+K/d6FqKd3dlg
mEAjo/jYaVEBYjoMa2gtPg+W79zMC+scSD7atDI0ZyrdFgDLSn+Fy6xymtCinwL4imajITm0dUdJ
ztrex6pIOhDa7hUkwrFlgQPgVfCFXBgCzKBhFg+AQcaELBqIyYUYhgine0E3pTUTny/LYvdgcdw6
+sM86qVXvjRr7FSAM2UcI9MafFshE+NdX6LfoUul0Eifb9jZmjIXpptPG/XztDAbVhraL8ks/WCa
DdQImmL/IXKi4yMtQvRnH9+3MmGqBQjR6jyWhITwDQTXJpXRnOQUr8jXk+kvheIefCR7rpevtu7d
GcoQBXA63jJ/tp5FWbgB9F55KLFcI/bAFFQ2hgrsGgktBevaxje4GBjSlNSNJqJqeLZ3nXUOtFOl
u6IZohpxVeoBSyymIFIfRlhE1bLCleS2QCO6xdcgl0yHy9MbHQ2wGkap2yzqR4uw58pOGBMy4J0F
jcKMW2Dk00CQy7ivesA5FXY1DKXZFFsRNYsLv9zoaOGBSUO72LBfvgldoqCvRfK/a/wgzaGNkX9g
oTNjVemIkuYif3481Enqr5Bvyek1o2dNW1xfkcNXZRYlkGx+F4hvL644FvLjN/xckwtFzuPp7tQt
lDi0iB4XaIyLLPf/0kQfk/CiRoUPz5l7GUhixKNGGCXSOqM2RGNHqVNUjkfSvSofn78xSG9ucepI
w9qkmKK+pKEtQIetp0/Ma/INs9Q+ksps8FfzcCv91tyQyPm8ZaQKvt/3OKDIP22oBxIIKurC+uM9
Ce7zYkXL8eBOjOm7Cj64v/xTcsYb0eRegR/MJKXS2VrkfnBN1DZkhykjTYl8GgmMjfjVT9GpnKkL
+Q/qyIKEI1p4/mRESJgYvusQp8I7zyRI+j7CUb1pTeuw4YUrZYO+6O2cUiVkxDv0z3OfcmVOBH4R
uqRnNVPBgUhxiZ0hg07a3AkwRZ5vnLO7NF+gmijkOuzHqnqWl8Ellsgl2mGg7NY2TBOTF/kj25i/
VaWcMc8Ma8apl6P/FsuewJtyTzi1jVO4ERByB+emSf9hw2YoGxiaon2usevsdvQvaSYOrGvJ4Gg6
VpoAWM/8bKGpDL5T3DvyMJD+ZEmmxAyk6Ggd/Jrjm6PeWlZ1StF/fK7i4m7SqmAIPBYn/G+g1Ldf
Mkn6HLCdvPHWkITn8iWuHEIV5dWMC3r7VLy4pDWvF70n6wGVo6KMAKlqv+7zlESiarssxw5NyNut
CZohkw9Sj3w3X7wEAnbA0ctchL6nfhc/b0aS4QDqsje9TL4T1uaJrVRLFwRfMC8KyGzlP3nOkVN0
DcAb7f9anUNhzRZlb0+Fvp7Y2rGZoHM+qlYXoW+FzePUYtRV3YYXKAwYmqf5wNvv10MikJ026DFz
uMYUMPb9IGH8poJ5jhYP0RXWmpMs+ydYdZz4KO10reHeh/NtXxSB6/30F76XETzmb3XkA0CF+YfF
JAl0pIxJEutqv9XBrYv9NiqswfbjgZY7aL2xyxQ6SUOKqmUy36QANjW7BUGLzSQDxTIs9EH4CJPx
05BGSBUccIgZ2eBoRZWd+HzS2Za8s+bxl8ELtUbxmgkAmlWwYduDbR4CjnGG6INmUluj98XZAloV
ABxO4U/0K59Cv6sn9xMzjA9jkS55TfViiI+/Y02RklzwkoYIiTcaNV+QS4+r2TcZVYOB8fOrQLgf
TTiO4zd/Se+YDsbRIncPDONL0nU/jmuv5lgHVW8Si1GWHvg/QrfPc3D31eSwX9oQzod+axpzjxD5
+yTo4wpz5eBmQTVlJxusAznDew6FGnsudhp2zhwFkQRdD3eC0MHhFKHPiWPnRt0Lt1OYVQ1K9IFv
30AnB9WT1+LrgZT5hkUDHbNfM2Vo/Ge2P/37UIrX8MB9l0TPCbQVd3Pc5lpPCQrVG5zb189Hm45o
3A8gYmnCSrls5uWlnhsW/ENOugxTq8r3/pQgCS6cYmG1XV0Md0lzG9JjDvifZURFiOpZHMQnZlNb
NNrKN2+rKMPNRAGWErgCxmq99M5vO0ylS9svf3PTeCib9HRq3jXZl3/z9nRL0DUuYJr4HeCa7Y4F
NFZV6zthQ9j6UtU4wSzhEi7J7MED1kf6X84TASjVsMMJadyroMJi3aq94x2B0dVbAoQfJ7372t63
+oGIoYCs94eTT9xe89mR/X9cNncKHQCXos9jdzAGqwuUGxzf3eKtuWaIwKntwK3mnIS/TIW42VJ0
YwzNh0mjqDN+hsiBRSLX3LDrPdR9hCw88yMOXm/sMJ0oAr/yArbN7vJml0IVBAHgmU1B2eXjZgIS
OoFuJ716LPfWIq30X45jQPEqFzqrROSG7EkxQA+dqP7yFZdGGHlwHoo4vKsQWoDd+zrNE2cKjmca
zrjXlPQiQmGFmpt8RnxPZZhDDxXB9jeRgn57zUTatw0OJ0xZfVODa4L6B+iF3ni2SlIN05AjnvsT
W8Uc6yAu/0F4UVpsy6MXy9CVGQBaIHhEQN/JF1/xAsrm8g9mZjkz+W22R+d+yHBzjgqdlsKywVSr
YRDEUsN4qiCqziOILZVE81Z7jPlGhB89zLVzSz2TGzSSxH+xHLRDn3XSiijwg7V6RW97I98iH+rx
hxxuSkLOAdmz0ItiEGHG125z6KD6nHfG7rxKpRiaSZqTG4xHa1ZaLhk4nxXvl/U7phXNE2VGtMFR
OlrSRgG00udMHtnp1fXJqn0lrcbsiABFiKUl24yfB6UXizxEzPm5kmD80trTzeDeLqovTXkhjXnu
EI8tvTlzOsIUxBwg5i1MudK54oWhkNAEH0rENzzMNW0Bbd6/qHqsaGfMEEDwjBoNR6A3G3GCb6JE
9XzI+ti2lAGCKOLWzszPEgrzMYsxqV0kiN2FvnGuJJFEDV80AHoOm1SSNz0YMbh69oXMijet29mZ
87q5RzfZhWKaVvKPLaKnAIaJ6Y3yGdV3xzzIztTdGBLsxOrmu51S4Yi+Dk0HmBHiy5yVFhbnWww0
geIctyklsWszrL5LlVzA33sZ8gU6p1gzzAn9BiKa9FezvIyV7zNYYkB+BRT8jWMHMTSJ1fEfXhN0
LT3H2Eko14dva6nezTFFCb9etTAqNVS4SWx5OjqLwHSMHUd2mY+S6X+R/mjdfs1siH0ILdtOiGQN
VEQe0sIyu9ZmWvE8pXb97NwGxldIXoaNbqGuJVn+Q/Sm4wt7gyHmxEPEKsJ1Ddfl9A5fj3sDQUKr
N4Xr1bXC2Zb5qJDWE+q1//ygLWnQ3grGzBmsbVOuoJVonmkb2U44gqdbm88RUHxO1hCnDtLCiI5C
o1mgQ1BkgTCM79OQtDKQCu1BljldNUkzYYihgcgSF06EVGZgSGu5hNEe7xom0ZGGwPfzjyqnkGk9
5EHp+fNOuukZNR4y/03hchUnGZzyqbMg1aMHtDhWKA25lqGH1jDTJHOAvHIQPPgzwyJ9Bl2aB8cA
hZcOQO1IviEfapRzKvHfHDeYzwseZeUvBaKq26ANX418gC/Me/kdKm6dDyE4bbNbnHDlBxQI0UO4
SGb4gROs4ki0v04TM1NvkhaIwWhFIIZ8LGOp5o9TX1W22+5E+Aj/sxyAQTrD21qVW0bOnviybWAx
r5SgbBjHEDv0M20azRfAJZD7tCVCS64RHGsxLV1T00D3m+EGkgGRY72OR7N4gfC5kn9Ay3+oL8nL
9XEshPGBwWjBJtQ9aaxUPiA3/X1e4umQST4vpNNb2AfThvA55gmIt/nQoLofo4B3mzmF6yRzRSCK
BIsRqzj0pjfTqpw/gGyRfIMjoTvJwIBqK9tZDKxWhjRjL7xiR3f559FUyQ3Ep4pR9Y2tZS/QNrAQ
RB+khcxyEYQMn0YvtKKZ0VdRYJyMl28GoYzjZ3upkxmAXapg7qTUQJqnQbYhWLt9QZ4ON0AO5KQ9
xhMXDIKHHtqM819HMQCZkOU6XlhcIykuFuuQhS2Xa4D9jegu9KrfMZ7tiX45wYb5nKHkZcKwq60o
pjj3u0tKw4C8UrBtOP20X2PIe20MxsLeFs6kB0LH5R8LTq5LD2AjbXb6gd8m8pL9AvzCWpU0iqQt
7g0U0sXcQ6W6M4XLxX1o9AaNGwKuswNzWBqFJH2dWi9ul1JPfvLOSCpifOJ75ZORazlsQIAHdFpj
em+w/H5anMxn5n3tYhQjJTc3uo0pHtoqadmI3/cTcSqr2y+bQp5BOX8czIM9QU99DrGJ4yUvBZ7B
M/T0VhUsOPuXm5YyuhU2PxrlqBbZ23lc7NrI7+2TH0fPVSMcHhsDEoU4ZBSraMFP93lWQSHtjt22
72jR44xwDspdTLGBotVk6tUeBnyu3MCAg+RSNnrZoa9C0MZtaiyDz34Xb2enuuaDyNibt7BZxWsU
2Jkaq/PrNJI0+IjBCFIvVfSV1M04sImlJELtBRjBrYdwyvWVVQSrCSQhU1Cb6oAZ6Z5NJE/pNbZS
Jv9nX3n3qXpK5DyIMPUKjkuNZnabAdWsGqVy7xBLXBGYARiQH11iXN45HxAndLv2d5BLhUJxiqSv
WyOTolCKXp0O3Bu8DLrKEb+CMNZRddy3F2qoYn0+zw+6K/cyvv3Bdc2D47J+BfCc8Km/KglPSICo
80v9W0c9fy0XekzZ4MVoMLyEJ5P6Oz7SrLB7/kCtTjsN+/EtUB6S3gffMzkQ/vzuP2aEPLGDG2vn
IiPooeRREj9ItCDJYJlceq2WhYaqT+QlAp6FquyKicb889joxcWWZSatTcgayo53+B/guT5ZRRaU
MWPO1b6PQSZySTE/++HxPZpy69Br0lGCcGOBHLU1sinZ6x8FhowaT28m2PA+8N5aEaSo6ikrlevS
VSwe+m0LVJEvk4xtDLTAHfcbA09S3jB/3vB4BgT5X+o8jlE5ODdLiamRzxH6XuXYmMstrg8QBWiE
k6olYtT7wnz6PgKAENb3qzLIzlGrNC6sXnThNW8/z1Os9OygjCP+jYzpi1H8Y3O28O+VrwbzQrGb
ruZaEy13FlI9J0Zxgp2mO2PkVyjZ0PzqfcXL7Z5gJrRkkrsSyuUtshZb3Nuj1xzfE0bNYaKbGa7L
i2z3X7JnBSkhwJuI0/MwxkclIRdM5k5FxaUZzN/osM+/qLuHqaNe0h1CNtSZ/Z+OU+vE2cFxNGqw
l+jeEv9mMHXOcJc2e6meGrT4Zhq6yPPOCWg70+swLb2BKiX4QBFZglfq6Em62hWtMrnbgZSFUU3+
fpsPYzTFq/yLfX7DdWYnMY23HJuWMFqbL6wdZ9PqZHCM2sa+GDi1+jY2HO5Ru592u6Bk2a8YFvRV
xE+RshYElAPukM1Y1LQPWISV8yDnQIabsx6SWjVy8Njus6sQNBexlPFKk6SiV8lz8zCoKs2QfKUT
sFjP48wGl69mBWrJc/gqOX7YcMsq5QeANZPnO/MZpCVuh8KGL6KlTZXe9oYKRtWFUXsT6x9tbvOr
W6SXsICu1BvhoZ4hnC7iFZ2u6hGVWHbcWSlPZn7RMCYquBBHv89plbNtV6c99yXdsxF1HO13K/jj
aHvRlIlqn6ZuoUC4ayUihPzBTTbnbLjW1j8jC4VWqEHGaW9gh7agXFk/wcgfra27PaBmuqbbGybz
qzVdDn5rvPrwNZ+A27rxVK/fteRWHbJYUiH2ViMy2QyKpboKMKBoY9HCUSlj0VvRo5ouYDgz/MuX
cmFPmQuCO9PkPlejdmerhwAg1/a0IlE6+a4LE0qn1WZzAzNq8oO8TDWd9no7q+yYzCs7uwQmdjhO
JnprMaOHf2ZP7f7ECOjIGdG2eNiapLS7a335NyRlpA1HR2USVk6Dbpt/7qDnwWWnurjxPRiGB5DN
aLx6NLUcYu2KdBZVNBRlqzUCUGCO3AbTZ1z4IwuZ6MrDRQj5INxYtbu5tmVeAk62upmUzDuWKwXd
Th0pVn7ZTmxx0F1ejpn47Ykm/SZ/LWzt5ql5ZgPgZV7ECeeGbWwEZpclW3wq03PayXKigXTZk8lz
DIpu1B+pu31i34fQILsVgh2xFrxwQXbLoi8qJOSqTZOAelGytnDDl0SqXQ+AV88sg7lU4JJuAH4D
xFnll/N1gtiCSk26KYPezRfcclameJWYBBw9NOyUf13MwGok6JSP8P9X8QvJ5+k9VNWSsxtXv4Mu
nljBHz+/BkxkbYevtkoYWfQwWTqORAXOJ8Pz/mrORPclvVSpWXGCXNkDhD4qmvVDN5dSHg/qsDHY
Cy01F8EFZqJLF7YFiecHpznECNuyROp15VNnRidvl8Q+jNiOOGDU5Euu4ESUvF7doSD9zlfgS4QC
YO1ov3v1b6s7+J8ob3zdposaEsXoDQwqNsM0rq95Pliz+KkSLxEGC0kuc4pzEW9TneEdcKc+UEVU
iSKuyfEQvLnFBtp30JgyrLZF5MzGtQBSKg8xu1wbDks4BkBwxy51aVrdlieLyUxQULb/Q98rP7UI
H/IrMb7oqpmdxpt0nU9X8xL2NoQ+ZUH57zQGuQog7Ja+J10pnouj9FU8rr5J9Cm3/e0RL9D9nm4O
gnMnwEF9zGwPv4nMx+mJuLQxkJl2t7QNy6bXAlkP9Y4oOcKaMx/C9iBVjk8Aen0+y2CxxjPNPkN4
nXqEPCOPEtXsNuPn6R98illVNJI/og/78xXFcKD0FYGRqa4O3JiaXg/onOARqHXWUqTItANqkFaO
WsuNd316n64ZJ5OaEwQRyIBiWSNzz35Cn5YvCRKyTpG9o3MkchYj5DlBOka22S+RCFVlUuUkX/B8
Ppdp9qjxcD1pZhzDopoA+UVpItm3kEqwT96iNas1AcRCY3puQlj6wiH2Q6J6CZ/GJZN0E2WUY8pC
5V0kpFmw3vVH6ciRato7PXCybQhoNvYcb1GR2BhYoDlcDczT3mO4kUNpT49cG9y38lRVVvbjCxiE
8WChn3FJ+4sK5Q4WzPqBKyNKv67zdoYBdbAmWqUic2i/xrVruWcxT+SZgzwZa6J/y04TUpHYSM5L
bydcI25cuUQUlL47e8fapBHt5LnGrZuDHyGtxl2sDdyi/1E257S409YuVcItvF50YushOfxJPBwt
kwteTI+Xh6TctFjELnTOwealD9fsQVtFxmNKbGAtazU54/PqooKGULGoAKzIlTTGuT6ut/5u8Gkq
OhRaJXJlKv52IikvQcJFxjkkszLvpaQ7aWlrv2MQaOpIl4hOE7R1fcnZSV3XwU8UFxucpFS5FFWw
6wTOF6Hy/yPfQatZSr8xDtpcUnMkZ44x7nWTT/Xah9B3hU8GrmolpQZp9fKReGo/kLjn4ObCbl4M
hRUX01OVUhwpHuiIoLQNc47NugpbnDoGFm75XvyjwaYFJLcEf0G7T+BiQRj9mnW4REeYQZKirnRo
atlUg8JGUhuXdnZZyYkSWCaNnpDG3KGRq1o1lwtBwpvaT4MDE3UfMvUJk/8JDO0QEOlodPrGWc4t
EIWW8G6eR0VMZzDXzk9yeQlVYv5Vf/nAWS5ReD0HRoJLW3ihS7vFF5oTA8u13catpFc9cQFDrCEF
hqo02oUVR/mGsc82yaqg1Kb0+m2eriO304Oh49WDiNrgKg1AB1Sta598ZnDTc8aTHgJPk4gPveQe
98pzbe0cyQn98lHjNe7jvIfQjH60TJo2MWkCzfPt4jqAA0vD4pL74IVyETtvExBK+hT49tNxOwHC
x7g6klcRBs8XEmox0SlUvXwbFQA9pZyk1zTH2QjaN3xGngM0sg5TDzUTYC+514SdM2Zp/g6rWBP+
vIgKYAac8QZ4h2F4ICSjJuuDp3Z71/7+Q5m4oSLhm+KSDi4abAsMLhR/Lxd5N1tv/kxMM4pMwwKw
5fl1qvEaDQAR0HXBjcgXlE9t/jsf8amvbotGV6LFm/9cyESv6NibL+Nos7fkD31MP0j8CNqnOEzq
AKikEIpZuOJHpLiS74Znwlj94MG4a0vwQ94aERdcg1rDCWk2gGeVrTemI2htUdvPhHqH4z+lrEFp
nTj2GfAfa5EA/2ChYcz/6+X1kwlXk1VtO5k+l4hN1PoyWA7flgdZhtr7MBb3EcnCGshTRpr3zGuK
kqO67J/OVHf5aeabZv88DUaGcYdAb8h4/Ytyf5ldAMCkUpm7EZc654uWUqff6cKlaB2VdK+Tkce8
FAgEjkku1Kd/FmUMvnf2nL+xCzoKIxPrl1C+paCTHxPwSDYw7KO4qeQkdmSPgVDjwFZRGd3Igy7z
4sITPbSUvI5JvnjoYQIzdEbTqyt25C51QglXsC3DRzXm/zuqfo9XGDt4LP80eCiYrWZQPLi7cyMq
y4crYnlPtl2J8Vct2YXBcV6cdjOASBNjwSIuvGSaxGUK/3KWdG8okL/Iu1ICyxb9LJu/oZ74WpdQ
RB0AaOQfZDEWDTJHfO/MBueZiizIHGxEQlMPy1tjgDDIlpZPhiCD8A2RB2Wn0H0j3ZiShiDF3FMZ
2xnoS0p9Rcq5XB9jZb//QOFCU9UFMjSqDhH33HTh3Nu0ZptRxIbZWKeSXzW5PkWzzWX//faPMSVr
SOMoNeUYdeNZ4EE5+YVfZcUb7C5R+PqnOvxZ6SiAwMJVTVc7nPoQ2okibeYZRGiMXU0nL7iwKmnY
B3w/oeSIuiNF8L3NZD79HZuS+WC8B0TSHI4ZI44r6fAksjdGvQpF0wyUdCjNmAUG+4ciakUHrkCa
LKCDByBYYdATnKyGFalpp5/cCFUyTglSTw95rHHAb1vJsCl0Q8X9Z8tHT8QpeZVNhgZZGHhmgjxe
zVxiIRaL4K41P0aJ1b8dWtlsQhrVHFYcPndQmJ3WxKAZbJLWk65DPrxwKyJj/U2tyUMpp516GRSN
ocrljiI8/7si4UA4Mup3X2IJv9HUaa3zQ35OeWK6rQ7VvqwEiZitK9Pl1BSX1Www8kPCGqsdj8/f
v3Pv+1uZ+rKKkkI5ffzrSgniP0oKo0xeG+FS/S1U1PLg/VgniMbXd9Jl2WDAE4wUypQrdEHxJC4M
BPL8pcjTyKaUVzS0re9luyeD9WVYk88gi0GYD7Pj2iDeIaTxRiSyN2eBdF6L6QgOorELQDBkjKXG
f/sOm3DZwyPyUFsMbeSY5GdsHq5zrTJPbbfa9auU1ws9BryBZ+NjeGru9EdR5H0coNQDW+FWVAih
QRl8rvLn30XUAKHbIE8W42t80acAlgMrrwtPGxhIGkQ17RPs2NNvSjUTG8mGomyt7WcnbS4n034q
i44AijiBffnOkAWxiBeiYwmmPyZCW6Q6VLMZXutx6R2S3SwS8sRK2Q06g34OepkAJdtnbweANB9N
V/LiXFR057BHX4XfW3nwO/Bkij88cOU4NUt8docyS6nYcdTMfwm+/VZmR+p/YDfc02T2I0291SFu
JN3a5YB9TTX0gwpmSUMtaMMlYmxEn9evEK+6Bpsc28LelIA8Ans1BvWYCrMG2KR7SWEIxSR6TvA/
ZxFqEt6mZxgV5KA7zI9lxvaEf662Nuy+H9qpyvgBopnoshzIcPzz/oneuN3AMx0u9Fl4ww4/BNJQ
WhQAYP6y27hRDK3Xo6+lYbbWfPDRV6W6Q5qMr2kA8mMcvTTUmRv9LzDvdAjRfWtiN54JYCdhiy59
ZNa4K/98g1naf1JqwBriIabk2tIx5Rn5bZZLt9LIbMCXZaU0vIxAdQqsophamYcG3JCjDM1SLQxL
+kqqs57BLuasKxN0cWIcGuMpY6ptAsPDmjrLsx7qo/A12dIjAlmUUIz9XrRAnnpoZEb90S+8Dc66
IZHfdJlUnHXxu+mwr+PmLaIYeaAfTlxYGEIO3T5VmrvWm/6mW7t/JKalvQOAtLqFywvfAi3t2dfh
+6lPI3dwzLNK7AHsfZBQVFqE4wgHFLAN7tCFK20eWTQdib0HMnWr38EkVAPNu8/fPF3Yo2lksCEf
2uoNrdmZKNmPNPEX8nSWFat4ApgNVP7eZNkuh3mIZYISFWQxc9ELlJ0xU95S/it5H7WHNZb9dU1k
xFjrx9e0HfTnc5BIUas4pjY4MyeAZPqUkp9VQnbT1WQc6s9niz2p/WBKNapTXSXvxeY/MaqVi9xY
sjgqak18JWlKRYj+ae0b8ZPoWCZOc+XXqGQ5Nek3877ya4yOb9H17xPeV1v6WsyQCBZUesE+VYm1
kJcYJDSQL1FR5Ht9D0Fiu9FVB2g4M0gE7aQXvLf7bulRNzyUSiqpK7vsRCPJowttZ8gfv91RevWH
1XWBNYALiKUemACXaLeMKkg3FPtzQb2hpnEeNjJeKZCtxdlqx/mPSfCkW+LZRH+yEx8EDMvlO8El
VMSffoOrXfgShGHngfIMQlRc1pc7i7WFa+qbVgNffVbFfNP/39yUEGMN0+wrN8tiR9AkySJxjRcY
1uw1mpN6bBtkth4qOY9S/9uZAlGLymEM3YEws/Te6Wyo/kTaOXOFQtDyk3v8JAZ4/9PUWCI7u196
glOIVnmfdZp6rDZP/xhg59GZLswLHC9WLulhyI4azGVfdBis5oVPLO2mB1yqD6JvPuOzAogObAH/
YmK6CxaHotSq+lUpDk26ht0yf+I9pZ6usONDEL7zJv+M3mqlcwgWDVEvOTF5dgO9Vsxx04GIHcyx
HStkQxNbyTUMv+kKtwCDnoNzXvFnySeKB1y6yBtX7OlqC7wi0hDRubZiq92vBAfnPSQ2Tq7STSZu
1e3qKNAZphR12Gz9ak+/so4SFETSvQ3QtXANcNYxRwAlX1Dlxb79UZISjNLifB6ftHq9fI3w/QCP
undexbaUTTAJF2vwETDz7q3hLAnZPflJaw7us7rugEOpJwRW1RH6eTmvRdEkT/IT1ccmYUOPb4xd
nnU11tJ+vkOGtzuu+EZOx5MlxXNG3mePUA9AdL9cOdhBiqG9Bo4Lfgac8lr+qCjFP9FtGrdS7M+V
tHiEmeCMP9dwWrHJ1RXT6Brk5leINnmVktuiRhisRvCl403kMH7i+4GGDPZMkZLPze0K6kAK8TVb
BVvy0FlOPew/AXZ+tVXpti/CdQYb/ILxT/bfT7mcdvyEDsLyi2fyYLsZkw6SWiY+nYXNswynm+uU
AxGJdEPorG0UBzX+mEtsSEY+pJ47B7Ysgs2vfNIh6zYONc7cN3OMvo0zW/R69fSFKBRiunhEfojb
B+NHmS1oveUtrGcsY+qU2YYFsAzK7dccMF3Kj45M5yZie43tskg0/g9yXD+NpscgFa2tD6XVlBUH
i0oUTC0ER1jCARqpfh62IXZCeoEKF2VALqWglhmg5ebQL5HH2teCwz3S1p9Qot5UjYSWEsraRtOu
nEtF57aNUNsjFaPFQlGCXXvTt24k2LGCOLKmL9sqq85F+xWCuuZWHK4qd+unByq2r6nclPOitCEz
osPw0Pqrtv2smH9dXiGxB5NlgwpzzZAQPKEg435Zo9XwNGL45gPg8llAo98CnRaAF0O+qErp7EfA
H6Bw9uW5VJ7cey+wG1XpHap0Ngv9+i/44wwJdBnch6BQX81uk210dqGl9Xui0A5iITxNAgtX0aOw
xWYpyBz2nWVVgu9DA1ZdgOyCc0x6NVd3V6sP8n73HoJgLh/gh4eZbL/T6xC08TveGTokkhwl8fmO
jZPUDBJLIOXaNHyz9Vccw8weNpwmWZ8GFxNii8SsUTwQCvP9Q7U9IoC7SLopWn7UXDiGlDrhiKFy
aANwFaejPkEtZuhcv1oy71dV9JHc3XIBKNT0aAwrt3CR2jbhIR1k71aD60dMq1myOim8WB4MrDH8
yH2bi5rBoM8Cs+Hnm4uv8vsZFdQglA5Cd8HGuOiXZBscrwY9rv9LGXRHFAcSnut4WDJ1tZdYJLd2
FUF5DWTC3tk4+t5dnt+asBwRANC1aTQ/SZwy1ekFpAWE/gJEPusfqTRSYSuOkuSOPDUMvujEpM95
pGqsvhiiC3/hrybIqcTwAiZVSR1Wo0tzgFpa8LPFxb93aOPtTomqYlOCYM5VeDPIpr0pyGdidLWI
O3EJyW02P9X9cNrq4yuykVYFIo8XHSsLvZCSjIDxNSO0FkCUw2/rbyA6Ledq4c9J3LcBM64BAeSZ
dP7zvrfjpoJvDkgRD0KEUxHOQ3i+qJgtt/Q6CvX67nHbujKoSk3ziJdoBVZOn22IZozhsXtjepf+
ZdLP7MaIetoCLer1GH1Id5SSEcrLDBh7Hh5hb5prQYuWyF+cw4mdX5KjcznsfnxJRHS6Sh8ZCSco
0NOjExhQLSxjhvt89UA1RqyWPkB0m6rX4S/MZufcX4Y+H4lATNh3Bd8KS+3repLI+x3B8u+hkduP
ffFmO9LweCP39jgAcdLu5yIMehS93V5+nX7Xy8Ar2F+Hei/Y+zQvISy4YVCc6jTdmUf7t2kXNhhd
kKsXBGtebiMmxUCcL5y65psJ9CoauymXg+52LkJl4bqaVrozK/o0wXckdGJpyYAcLRj3Esx7h3IG
Z4oSwXLsNA175LLhzbrCrB2yRirdJ23eK+1dZSy9XUKfpS6r8bFth71PMNXlshW6gIAne6B6ABIB
aD1sYNj6RFUL1RpmFAXvmrETPy4DurfCZeOSb+r4Ouag95Jn0xHCzziakVWzQQahxwSZBTRnvIzh
51y0Fp8H53JH8/JfkxCj+J0yeDHxjHMrnOW3C5SVbtOO7mTWwSUeqg6C7jIAlbFlQCmdQN7zadvY
tCZiYb61k+cZlhUxkMFBgZxVuR1qXvLkh+zoEu6u8QxGj9Yeh0ydwQ+qpw4mTAzigVkvunHtds0g
tVex2dwh3qL2mP9+3QWrvTXfJ6VMROPoy3G3dY44wLBwk5yV8ZMLreg0MXq/k5lYi1hfojKM2n3c
DPHSyT7h8WH8DIsv2sF+oVIJKnu3AwcZtp28g4VDo2O2Uew9an9pFR8p+DRSvuj98wYcwe5lt5dg
upNlm7E8qDaJcJKXOBapNvwBPjH9KoadzoxHnhD/OPL+cv5ZXutlUJtoBZ9EVOEBm+a6g1Kc7tNY
qpywB20cYRVWAl9izlUTrhSzx0Gp2381tYWrRepN/0cvbRdwdOUiJln68/Oba6Iwo4lVD4h+VqdV
Mzhsw+i9sly3VqLcmmT7+2Gq4ZWr2mBATMrffxyDdNp4F1bk+rmLcsoBkw2PKL2CTuQ9G1QdPs4a
YtfSmHx5PRr8G4cAyfCQt68z5SfUCrdGavypVah4AlIs2XHQL759xLm1l55kt/1kNmmHHZzgeqov
qhe/vIPIArv+sHETvJ+YCy77zacPjmC38tS13BdGeW+TIix4JZxR6Zp2KZgoxCUoCCqfQGzSo2jG
lWQ3aZnjNBTJPMCJ2uL9rYXZBvcN73bsheMFVWePUxI8YBW1WpCm3xi/ZnostMrAEhn3bRGKjnW6
H86+FlbWuZA2g68YxHnQUbjDRUHN0GAuavSPX/bZJd8bcsEuHAWtBDU4cj6AsdXRzbshx+o5nvAJ
TBP3rNa7JhElLzbQqgNqV0x1a9KjigHiqUX3Yu44ZeBgYdIXps7JP+w+IynELxxQePAEW3Si5bJy
MQM1xAn7gpxDHpBDznvo+72lqjWJC0q8JVg0yB/hbH1g1FSmnBR+KopkIO9SB/7FvoWti3nV+fSa
6XIuQiK/+juLutymYa/Qr+5JETu5FqYITwisyVsFxuDSyQmvsRAWMzNRxrkj/dg+AMewyaCc+uAR
SxTzc8mva1GRwXjehSKNL1kaFaUnHvZFcVkIN1DcI1JfYaMq4HJmEOxC4WpA+rw0PnNcypNGZCuO
PWCZkRf5C91kwjx+7TkO1lVIT4YD+6Cb5nIBQCqcRw1lLKBOQCBDMYkJdnEjogFDaX3fXYzTEyVz
6NUoVCNe/O0yvrQ0INIFC18d0571v4RnaCKh82O/YgZIRpwxtg8zXlRzovZKnIL4fUbomJ9IEmn9
Bm25kk8muUo9TBedks/xhIRJ/mKrzzW3ErHdWw/ak9Yx2Bapbx4l+AgF3zWpNgQvwR0ica0jwLBZ
t+DmUFIuqlDzqe70590V6NysSWdzK/l9izYjKLn9WwB572vYk5qvaJ4p/3wXJadWEoRHTnP6NP4e
hti8PRs8NIcO0y2TsQX3d7GqeqUabjmVt6ND4jWf5m5SpWM09CkdMxVsmb/9eituxX5Ea3h+m09C
/Thd8clMveXrvHTXIPPFKXIp3Xtxt4a8LIdTw4AAoYksBeszAJUdxfpr1N8+nZTBt83bhSYq0W5N
+AmgA2agRuWPe7QlN0R953H5w2bD5rwH2qWrnaKD2RHN5BomQrpcHwjyeraFiPnT8atHqq77te1T
P5Jj7A/LUttN+L+IEplfJFvSQMrxQqZhoyiURaJzGlagyMaNVNl+ph9lUImm3mFmTaewkQ5AIAsQ
JMgFD4bkdtKDgc50Olq5tSETXlvUtzB6vYBpgOLlPeYGaLSAVCloYG2RFrBt2FYYcCwmqlezGe9z
6f8bp55UYFH5NZox4BGoNQ+8imD7j6w0ZsEfbW9qV0HOmm5NpAy3gEuIEV8dytWDGFpfKSxHGJlB
R3W+V1+7Wx4wSj67BFL3kRgePp/bAMoByrQNplNSNYV/WZqDWdebQEX0hpo3P8MgNYJXextK+Kgy
l7d8bLWRryRoGS62y6Wn0WrmNSbvxMEqy0Y8GJ1RB+GeGHifRo8C7W4onW2+az+qEX8SVnhhH0bc
xTM7W+otzK+ExI7oGmW0HQ2WCa+CzUrfqhdbu7Npj8+8pn2mu/0XYFkEBVrTmAq2KIvuvnyH27M2
J5Rmp897jvOynOFeP1GOMH53GOScaqL5OB3ppl4Vapq+jwYKecTOK0Xz7uXXaqxZ1t3Bdk0SBBo7
pgw97pywMk2JDyji+8dXC9GlK1Os3KntA03IhQblXrwa7qCCz08pssr5lifLpx+bGHj2tbAnjXjS
FKG0+CkoxtjtnTC2G/6Gc7vUoMiFXVwZQiEwtgd6Ss0kRbjg1wnqY88sRQO9NVuHl2Jrcw1sVyXE
lWUFBDnZRTGeIM3YVb6WVsFOE9CIaH/PMaDLPZkYZuexkLtVwnQ6uUpqeHHgmRLYqI1CYTN3K/Gn
TeMJbzCT3Hi+XoKooUl0aP/ASoIWx28mjQkVOJnSkKS8g28L05L+dsi7H27mWBFy5mJU0z6+Qn5k
+Tj52uB5sujNeTW5yEVu3/QYqFo5HTSEdp5iFBMs6ILUtkm4KOvgnwF3zBshqYse/gJ5Xj27dEt8
5/sQ1khZQRD8ZPugnj+oVOKSiZhFx4ktONhAMsp/nZNvil1nFtKfyWahliU4eaF/602A+Nshj6HN
guMDHbInQycUuQTXd+MfjGHL0k96349gqvu2vFLcN1n1VYXfkoEixOjAecCROjwsLOz/Z9j+zxFF
I9GVuQ1qnrKp45TAIfwhC7swzaD2owt5kADR0BRnsZSY+V4f72UoE6yrqwboC5tPMCqDyN+f0nhE
tFZToetx/iDLF8yBJ8KLgGxy+6Dnbb3z9Jc7pMrZh4KW5Xg1Cz+8r0ae/UzCcOLbGm4kFf6IxJFv
u02Conh1iRJgmahUtoKpQEHV72Rsnc3T2K1dL/IImFbDsos/HIZlcEzm/xJ9Ixpuct6KOwOLp4Yh
cdTBJk96thIk9vlgg5ZiOfk2j/8p2HYPWUtSREkLLw+XALC53NWihS0RmJenb/CV+n+UlvlUH/KX
PScBgBu4Oa8Ljjpt/y1BaLFcXRcJSDHfAMMDwg4RypvMEKX247y7il/uCH5inPDzbWe/JZu7+RIF
7JLyqirIvGuNb1uAvqeGWqK9g/r59Js+uP9coS+19HLhkxli0R3aewiKxqXtagNC/Q9qL33gZDKa
1QCN+YDodnX3ULgVlSsp2YHts7nkbP/BE21jClxFdiUHlR2ymMqhtcz59BntL+oa2MEhQngotRGb
9aTKk7ZDeOY1ZTt64dSDdOXVg2rzBw77C/qHNdC6a28l7qMYcPgP61LX/ePhcN/INn0oldkz277/
rtql/vyi114kLrA1jl+mhyyx5OAHaTZeLkYaGshEDzXwtrc4v94W1gqt+OBbE9liMj/X49h2GX6z
ep5sx9LA0J4xeVAL77pyXgSH5nNepuubdOpILsf7gwNxsjq2YyYnL3ZK0iohaJBJ5jpa4Dy+k2Yf
o/G7GnDeXyzRvUMJwvNHxN4fUE6JwCC0g92jTUIijehCw2BKapChAvs2PQ/q8sYMyqayagR2zV84
wz6aWquOo0wrIWGPvbGRay22OrJl3N5GKcr8YLTtV32oZG3KhYMXSTp/YUKAGrMHXv2TJW8SwNn+
6JNjGgfQlkQ8R08OLLsyxm2IqkC4v46+8qhtVje9aSuQQagR3peNpVWupD6GdxNzTEEe7t+p0l6B
DbrjLW2n0snHnptwsOKchm4bqKVv4jSlVWHaX4wBANA/iPC+kCEkgkv6Ovr8UvhdlST+CCmHRDSj
vhMbjFkKrql1CHnc5hyHadYYpCZzaHljO4oIilkfGsVoP8kuwQgCmg5+OjSoJqHmLWOKupOWKqmn
4PCWoF9Gl8D3lZcbaINbiaq1TxIJmEfq50SKyX2cFNN919hXKfowIkWm8yJC7FPLDiCEgFWmKwZx
onxL0GMS8VtSmqp86llVVBgr5nCMzh66kwDq8Lc0SdZNMX/91jHtpzgCRGfyju4XE082LFXBFM3l
yghywn7ctTVJ8JalbyRaqPMDpM12Ig8iU31NPlbvozUkd/1xl5blkbfqjoGQMBMwVsyolGDrVdt1
l+Crw+0sBak4s06HzabVGvUFzZm76dDcMimmTK0Q8Oh0Tc/8snxscfl0vy0197XnlhI/JBHPgZIE
SEP4+zTARyLFBds/0W45CQx5jxgwRSjMbOeVx7gdyjfWUEcKxHB7b0LZSwRpqQR0qBvD48ccu9k1
qXCt4RTpFHwY/eytPb6rWonK6Wi/QX1YaDjWx33uXmQVvM2feUXd35UePJkSSEku7O3tCmXYJuAD
h0rf136QOEjVZYo+Bmu2dfxFu2VwUZyfZBcHKRuTk8B2XcBafaork6/6CL7fe/mPdVewhIh0amKu
oB1bEiJvxRwxJh8wJRgGAR2VQY5Ev+NvZ4huOhNyfvDYPI8lNxMok85qIlh9eOlogNc5+TZ8ZoMw
p6+hTe/7xZMLaV5QP3khiSZ20S0uH8ApD8H0mixN53oV6pDd+xrtYiRWLhnKMU0rgUzCSCxKMlTX
pYVF7st0I9kMp5RpANorgfrVsl6bBUiYTP4CxEaTkQTszYeau0spCpKN1QANB40iKaivZmEqXvkb
pr0Mhmjkt6VhAuYr7erlgb+W/ARLIjh2XLleV+ItPuKdeoAUVf8aK4hIEqvfpAEw9DJyfjxsye/k
Is3Z5aOlqnOM2ImCuqkQbHX+NrI7qhJr69i2rM+7j1ADJsUWE7C7HX4EsWlQcmqFFswmcPXGcEiu
YZF+TkvdHSQ+ArNh7W10H7NuTao1CCAbHUFe6tXGpqr8Q6p8Znn8rRqggSi5yFldocKLtgF8K8Sf
UNbaEeUWZN90SH7IlBaXZvVH7NHHblAE3kHfQeG0iwh3737op0HhFWkYisFJS4EbUOjc/8E+MfRo
n+1wfyXQljzaY6DCtq7aQKTsIx5NWtaP1CY7z8x1oq/7aKH7qL8iU/xyCaT6C1t8llCWd4dyuoJ+
9W4LA0oyoTu0tBHhWgKoaEMcDJx+bIuxJmGzL7tFyCibGCGI/eSUgY9gSFQZwsOQvofdoRL7zTRt
TtLaf5j81ezngpN+x/6snoIsOs3zskl6nemx78E0M5r3/5llf0kccT53HGiKDFrN1IQ12P+PZubl
X7AGhsbd6W41DQZmtLEMk5vAosJRaO2RH1L1AU0lNgzzrUbM+R9idjdbWbfYj70joblP/JIpXUIi
8tsssgWQvww8CPNWkygrUx/awP9Cl3mraX1JmBL5ry2scE0L8BcSQhjVYgZ/TOT2YrgDy4L5ZIRc
jHZt/rxrDj9Oz1UrFvBxiipLXYz5dyguw5TzD8ZSDPYlbzPVws+La/3J4F2RZLi0WP/ZERWpJ7Qp
SiUZSuOeqz6B13DOcIr2np16/XJzO9T+8egg60WR/mSCIw10cTDEb4V7RMG6iHfeMgW5tv5ILaXb
tIxVme6Zjm2ajNXV3wUnW2JKGH75L6cu5FfHcuADiiaMVB4GHXTTbEXStaVWeHRATyDUY0vHbsvZ
JO5YtwEYNK9x/ezI2y44LAur/mAmuq5+c9BfufJAknVP3TI8yeoGaqdUZTYGhHYLEixRWZKMC8Li
fmY3sEW+nYd5ygzV8Sevd+o4Pt7LMIOsqLtTZ/yCYVyAkHifVXigTt3S3yqo1a/XFuZOdTNSWNC7
xachWxiLssvSk9/TL9f+UGxW8WXlS/UtUCVIeZlnu9Lu6Ta/IrS2rmNuBa9ft4vx4ZyjNX8ZXe9V
DvI8INuqTgGa9YwpYkchw6tRyzvT9q1RbSlraq7mn24V1EBMXrel73kMULsOHMwsUY5NFQee58Oh
dDl+ueNEHoDj4Vfgy9ndvdTf+R4cnEkYW0a5ttbrf9L7Vsn67QludkqLEDd8y53r5fIV6wNGr7GL
F6sMLeaJEvCqEnU1SVMySF+mlAy6ldpnfDAYOERUSsOFZotI1e9euEF3hIvFqg/5fzhBt1mftqfd
dgD4mPAE+w0M/1ppHyxKb2CoYvCYrbzc9OmnYx8zfAL6NwjWEQft8lGMwvHMkHtShhkJTKt7cOwt
7LKYz/ZlB6SKw/ZLPCEuErQkWkX3dgWaXbCJ6Uqa41sdOMZgByK12/E/uzNh3Tp8MYsvDHbVacS3
H2ewnw7Kmbpy+O0b4O5L/2tGLMR8vz5T1B4tFiNf3TeP1FDlqqeGZHqo3DBOLi0OJ9LXr//3dSEp
jltlWdlBwv1DRXPIDJcsx+jBehPGltJufWhgV29Oh56n3nkesNM9BEB6RQOlvoLzGMRpIVvGjl9q
EADCSInFy0V9mixp6CfZHJP1oabhjDU8sELudeAMa52dkjbo07gSo0T3vOi1MCktEbev473eO0bK
lIXmzlZ/YV5v1PRayxqUcMPLunEJlb//sUgRkpk9ZqWRgwkMP27NKyC2m5Xt66VK3CzjkVYHVQGD
dijVumIAgytRRQxY0cfdJVDX4P0W1GBTpcO4vF0HmG4VtHyrDCXp7koywdhJM8W0v4K7dfZKvaYy
0F59t+tO9C9sDzsPJOBhQPIRRwqavp9+Npo/KpJVlgKXXbR+cBszWi7JHqo6d0JV1Q4LtcC8fg9P
8eXcRo63tBePtB2IAX/kqPdckFL/lHiv0ADzC4ZrpeIIOntC4WkucGgpmi5TF9HhoA/lC0vO1wvz
tZHRz5kzsiRMIzjgqgcv5hEwaG1C/PZ1xK2rHQtqEn6d/dnJpMzDY4xkUA8LYgUDkvSXlIoBXarM
0jwr/CyOMUdGJFdqTF555UVe76HiS0yZ9HJKFtMfqgcdKfuMT8PaqJoRg5iWUm7x/OlKXGusUnL0
G89qm3uTcPjilqTOd3MIdxWo1rgTDQ+YojgfBLACoQ/Dv1Wh9Ao+YLyF75o9D6JAW1RfdTTH7ROj
zZz57fw6Di+cRKbBSFVWeJTo1T+NYj8Z4i+eTAfFpJ8LwsJk4WcgO2DNwTedBJBdAcz9XS95B6/T
EKZUjbFisL1yT6cWza2YqKy8jlDq41ziyKn2ZNm6MfC/VgkTPNfhKdSVfOM5TPxYGAo6tDU/Vwaq
inDkDvYtvgD+D8HokzgzP9NRheooadFFVhkcYxj6guYc7TghI5LWDUP7OF6CEZ0KG2OOYc54ZN8o
hPrzX/NQnRL36xLCEHqGGSoN7wCFIMZrHnF+DekOUb6pEXb/L9bjxES0z23FHiKpzKSdRnSJ/eiM
q5kjwbU9RqouTxojlMPftP3Ak/Azme1VIbjjvsoVNPO5pZMu0wf0o49OeFewEfCtFGxMvdv+T/Rw
UKnDouRnF1ceetxRd1tC/H+DEmW6sJMayb4wmHF/mZO05woaObZmnZjb5+9JTKPqGF5jlEQ2glQV
IGVUNLLb/oyuqOFoSYzJ/Idr/jX/Ju58jbV3T6C9Yn3Kcto9W0Ms4+rvJ9fYsCAKW5OEsTmaRN8y
HPQHh5DM12bZnYhtVByrpYaoq/rltysx1awIxICnspkaOVHQ0Lxn7TltaKiF8sR2synepXV60mV0
G2noZTvB46UVbbl2cYkghuYuNZsabAuCqU7nbQIJVKdw51FXGIOJBac9Yc+HeBnbDXRH2IHrZEZP
WDhqf2juZNo3DA2dtf3HJlkgO6nivftmxm4y6XVqFuIkg1XWBnHDFh13GivzROgrYtvirtNvEE0k
jkkpT9VPqMI+QIlUa0NEeb/RERVT2R4fELNrlNT4ODyLwwe9WVFeKQEYxxUA/WWkpFDOswzpHr1r
5aZPGIoq9SG2lICGKWpQ2d5bPFhIhyHwlVaHzHWSEQoZwaG+66wnUWjUwst7UgPkCCb9Hx2vH5Om
jqtMb1XJFFD5m3PAdzj7NT57H//7vlj11o4eMC8tMJBJjCyrbMCBVd2PNPnGibLSP1k7MM5JGrZB
/1Q2TlxE6LY3XUdQvTHhTkvF70zXaHuQb2v2ua6RIOWmHcHjiXpqSth17dH2xi9rFlGw1S2fT1I0
KjIS2uNUUtwmAj/Vv477avbQg3ENDc2PjpR/8zR0nchsh7B2lOKP6W3PJ2/PJRpWp4cQ9m4D3xpb
fwJgtsaBWKwhbvgrhkVRhygY/6xC2MTduPrGinOL8eztcs6hDtIgY83HGd1ifneEGTIobM6yjPb6
5WS3nAGnjLHr9hexaNMBMFEi+GQB6QTA5Zw4PQX01F/3vGDnYVKykkX7Zpq7qvgqoMJZCbjLL+sw
4gsSq6Jwk9/k4IeqcTdKgQ1VDeWcVsijI7iqnb8AKwI1JxewyG1HK6VHlXwALhFl+eJIGD5AE87U
B1iTd1cxCMg0ZhADxCqp10rYPcAed+K6GVqsVI+VZWx+1piC9Exmw1NUAdPNmHGZPB/J2J61IqJA
0AzmuweTc4bDOi6o7Ya+BOuK9AJh9ll4LP7Zo57J23dTWXW7X2Oy7Hg0gk0+5g6SEqVAk49BXbC3
7AT0aboqxQ3Ii1+PzPEWO7+wkp7JM6hGCwhwoGLKCz/BdEGqcMYahtgdCQuFgOMX6kRZo0jCKR0f
rizR09ee8lwPFHERYEyx2pbCwxE5VeXmu4/G9w14gtu7gbq8ZoAYQHtLL1JUO0eLd26iFwBWrbFP
ieNsFMHglMz0ZC6NlbR/icG6x9fw4qKIgRV+f3S7UZkP+HofSyH0xrxker4m5NHrtmjiyMAIs30e
W6MtFuAjj1gJHKtgUwXtmCgnl74jHYhLj6ZKVtXZ93AAMw/v1YSFPB5i++b58yrbodjwVEgB4IUY
3G1Dh1owZPl/Hrr+vVXjvgPLHO2CdUM4D0y0Mm+B2cFEhScoJwqGgrJiNINHUDijEeH8BG8OAwRG
s9BIzj1D8cTuAUd/H5iN3FFV+BJQ9CvqWG8UmQM+8wZMN8gHgO0we8w1qn546r5LPr5igX1LCGWK
yqx77b9BT5bpKLdZ0Il4udvqFmLib9/ZfE/MR2IRx3AKz6pjHz9H8yjSy/1K1bXauNtCY0EZ7Y7O
8hfD3FYLqG04nijzrichkOMRU37Jhvs1qL6MgGqORDZ/RWYa/2IlAVcKLQhkRkosDRFg+6ELDoH6
iI11Dtv39owotoSkGSymtVSwS0RrRJ4yS39ll0gjZCHXJhMnJOdstyPwFTZEHpFxFQlVMDzmI8HQ
ifXX7jIUViE3Vsjr3mz68qaMAgETTNahrcAyNVfPMuGFPJxa6PFzgwGHsGiAV5UkAd5CBtkjx/80
SC6zrk5kt2bhg4I3ArjRu3Pvn6o4pFgMrL0mk9Ufw7BA5h/hOplkSuAvq5eWnpaqdB1T6NI5hWs+
NXBC3e+DYqCOqETEBEqhogX5utSLtsJPNvXBik/u2B2l9nEs3UYhYI9HGyW4nr98M9yGomIRCkgs
1NojZ5bv5Cf+0D6St7s59xgwws0PYi59iDHpwAXJCBu9whH34R+NFT/hXoT77TUgKPGToB4uuQr2
KqeGg2n1U1nFWgm2h2Ego+5O77vkKnDEgjvh7OpDga1KD8269Fd1CK+UeOdwp4pioZra2fdlpDaK
97fXfKPQx2pMT4sbcIcrWDXhdFSufiEe+NGLOyyIXDP+ms4FsEJzAsZnaEfypYLrRe1VMvK7rkHu
DHqnP/GZ4wWlAV2kwx1Le0WS0FcxQLZvd/WNHKg1LD8P+ylWbZBiCslrCU2oBovUWXyF9GPdHFhz
vRuhCS2H4Mkn8GQaRmIC01ik5epn5ChFFw/rtaO3Anwf3gJKU0DVV9siZYU/CGXYTKuZcSF/ygc6
ERpaEv+dovIxDCFE4ONHijrlvNfs3jmQ6wdMQxrAcgXUdovQOyiAQF6L8tWYGDE4VILN83MT44+d
/tslV/pN166peHQiRyGNsmfwBigxixnlEbUEUiR8r2yWT16kDkHwQZmaz4iVKok59GSImza4Gr1a
xCei7FPvCRWGuFal+ListW52t8CcRdfIiEw+i/fcxDOlMADzykBhnfSfpQxpFmVIvDGt54ux8HNm
fZUoMzbyg4LjBjBBBed00uWTtQhYRLxEwxepDeuUSxlVSAql2STOjtU8awCqdKbav/VAnDGRa/+q
24Nza0z+EU3nSMFUnH82SEHxibxy/8aCe9k2N6kwrkYgJIyvYiBz9vfdrxcNXBdk7kG3rouTcTXO
3WNTIM4iD84Fc5Siypyu8BUMcyjziFEgV4XrzasDM0IlnDh2yRGjrVxDC8/CLegq0KIM4npPZ2z9
D5T2PxRMZjPUZqmSP5Z5KFqbT80n2A5Sz4ww48j4ilO34pVwtIxJ0pe+NMujGHdFD+9/thKlUUsL
wFjXENkUncu0PuEeTHBJD49hzsHgibpnZk50zBhnnytbyqEE+1a2m5+kzchvn51qDC9BGfiLSJ4o
3FYI61deu7HzRD8RdkuA1hSkd31+kOp7ij8AOJ6fU3s5JGSPzkVe2RFSTj0mdhKunXRORECYEACz
ZSowq0ikN21kTy/knnB8GLcObLSBUyWo1L2hDLucwDohzEF+p7pOXO9lSiU/KCA6ZVfV2d+ITYfi
OTp9al7c5vojcFKTsxojEjA2hwfn/G/qKkrOnm3VHLWuEZIVKKO9MATLYL0Vvs2t8apvgpAKZfKl
fxFfDbKIFRR/Dl2NmzEVQM9xoD6cVi0Aw8szHLvcLRFWWAlmK58ZIXDVl2jZOWb6eSiQ4kWPQctt
2LH9aprOw8ui5iQYiCUpYDsK7rZITJo9rsXijni9oKLLwp41bOuM4Pn7tNi7HeModZP9fjRrRY+q
TW2xrfOfFryfKXe2XJqPeX82SHD1Mhw2B2coAqaqYDQzHoZ97qwj45+yw0dHLCp4ug0UW/wEt9Sy
4OC6uKt7eWzEis5s9W70BHW9uzwPpOFvSDDgvTSmMU/1pV1a+apKAStucWjYuqEp+PN92LpQiZTi
tYA6bESXfwBskpOw5Ysc0PC1dGborLfNFvOKdgbG7kZv6aep8Q4cZ3YlOJ6X2WTiLeKwS7v7K6oT
H51Mo3T39cZkDh7mt5hRRtItbOvrZjIR/QHig8rHAFbdPmGBdfuUgB241EO4IFYL6Oe0rKiT7/w2
SP4rHAeo0cWr5QDlxW0quloScO6OGkZnmx1JgY3QH4GpAjGkEjkN0sX1qmKS0xogIdUCswc6lpe8
MZrvGrf08kB2Xnk7/sBMEoHBr1PWHkNb0EIx8N9KV6SilAYAbzavwGEFBhDWrkuJywyM9ajN+l5T
exGDmFlwa0+cxtj8iPjgw9b61tm72o+AudGoJWCSBfDDHemOZRd1yWVtz4+EYIqKyrcKKg3X0oKx
oV0iXxJ2XMpcw2q4ShaMRJZIlMWJrkAAU5YjtYm7b/GPuvUkyQKcY88cLndRdknUnLZF0/1D7/ma
PPVdTudMTyCAaXoPWv56isW51I2H0+ULPAnPnfnvYVx/ZTZ5Mi0IX9i5uE4PdXwjkXUQcN7W0D0Q
clIJlzJAJ4BCq4vZ6fM9eo6R9I13i+LoJrMZPT9jH3hbM8sEIER9482CtCSaqGB3Hjht45h2+tl6
AzCS2DowgQQQd+EjH6B0j7DUgDNWJViocG3b1yHsrg96FIf3fB3a8n/i5L2ytXym8EvHhCVBp4X4
W6MU3XyFv4K2ltLFxkgKzb+4ZDsOaYCUxwysap6OAfsEj5qO+2/AjrhGfw3IG53mzIB9izL25Dmb
ZP+YE/YqW4R97dEzhpMiyhvmMkCANOVt96rYXlv2NG2eQrQIkN81ZyKH2zypfzu+gSmcLw4U3B0k
bypiCGBBLALD7wBwE7TcR9ZhXaJUon1YLzMoXSDVQlFeb8FCWRAPa2cwr9fpR8Oe+x3wuAzAeL24
13yQGokQ+ijYeMKoSbCDRUVG3u5+cZK5IE0rtDvWiiGS3XGZvyOPqRxFxY+FqM1eFP7y8KDlRefQ
9MsE4j8KFns80nJvp7mDAKfgiWBa+WMRb1KOekQoCJQ6XsQxCp36w67rEnQh8lfY5A8cicOX4O9m
jpDudG/638yfWkraCcC3xGo8P8TNdkbqpX+bf4FCOydJr6Pr6bcMPtDY21NfywGk9/uIFWPIEIO5
TJPlb1SKcLWSY7cDSgz+Qi27Hz6IkscNrJ6uotBkK8GGdfQZyavgy3i7znbhCKepN6BfNYQc947M
XDgcZqEKdXE+KJhJ07Dm1I0tGilmS9uthUtXLV5DjPXWBoihoJ3y2LSAtEcKKn87kRXxr1jdVFcj
9iFE8GYItgT1ebnIj9rbkyLIKVR1vZPbqq/0tFfUl/m7w8X0Y+Qv0Vz9N+GTZzYzm/VAIG8ulRzh
Fv55ARW6EV8YFbL04S6Oanjx+xQoci2ho5c/F5WMsZ6zWydd02N5zHOJVy+OFXRXr/jesoPEZr1d
Yh5FMYLG1O4omlsQnSorWkVVNN1rCR9QGpO/3cCXaTIyiUaZcv/NQsf3jzI97OtgB3bcZ4mekdTK
8DEvU9gQdd99sXW1A2KxOVU2osKVKlKiBfd/jFfz1vXSKMBkaX+NGMPha6QRyH+c34pACM2GwBTK
pGHMgDvSaoanY27cID4i8/9ZYqGDrzN1bLtymXK4u6JRwhwuNJywLyHzYaKLQyYHpyMKna2cQyvl
hACzC/KG029/TVCmz45KQTNcerzsBWRHKjdso6aLto0o8HSdT1HzhCkWHQKGSLD8doRGuaIfFG+n
x4DJ38FCQ+LZdcofHgr2Xs+Je2qWFlU7mjePSNcjjYZRGbRjr4J8tTzR0Ixerm2dr7in/yuBs+zP
kijbu1vqds0gJkalWbDn83f+1VpJ6/IUTkIrQDZ38ZH6ZCbv3SYDQSksVee47qQdGh2mlzJrDY1n
JyAtIvdZcbquAXZCyz3RT2c3Ki4vecqDnudgadGDOl5jLEqtFRbNPYGcesrs7Li/aTyhk7XgrFUI
T6kmnM9IyzrYgisqQiKU5tixgfEmv7UkAtM8fxKPl+QNGQ81mSuzYDA3nNbLmKgpU+G50CZNTCUn
I1MoKFBA4vtgPi3eCXWPqaKXyPTx9mSpR1dnUYmMDvDGLr2sqBwWDNQnnr0vrDwMzjh75iPQyotc
oio9Wwb1Kx/ullLCcgZL82AI4AB+QAh64xaIT+nhLxKMUq9uio6Sx4hiTO26h8X2hCSiv90VRK2A
x6fv0SSHw10lbMAgq6tu//ysdN6QqnWngPm2KRC9rJTdooSuS8C0debWOI1XVCc4toG/+Ohf0BFU
jOBR72aAXgtwRcRSL/dM1HEEmGuVDwQWQMD4pdxCxa0D1rC7nrL/nBr5eHcRKqzWpFLPB563wJhM
bzYoiFkZjpz8Gn7inimI2EYQjsIP/+54lEOSgEEzfLcAUcPyy5cEiqxjNJnk5R5pNmQVoNX2Yw5u
sKIPr/ltv5f21IJnGPbSC+ggyBZaeJMENEpYs7uIstnra1RM5EC/BDVXXYS9hcSN4j2S2bB0uL3K
mIIhcey5j18sgSbQ5kVkvWYSdvYTqewrYwx/okQrtByM3K3OPEPP1YhqON3LwC6lKvkhTM8ruDb2
/bK4maRu2cxT7eYcsHBnqcJ9U7Wjk7yMRFEp7MrK3Ef2g0K/Wb1V2GIzvTSLpRdlpFLWMAelGDTG
z6Slzuigyf2HY8I/kBCVft8+izp+lqD9PPQng57Bol/CoZbzHK8Nwhujh4qEKx67lSXa0SuaQz1P
8OOOdF8jy6JxCGp2/qb+oJCG9Cyj7FBDQgForiJTx2jghUjLi90PV1wgAPLsKW/cFH+JxwqiE2OF
r7tqz2TIHy6/Sq3RLXlvttEUvpE8MGnI7o8BYM5+EqoPov8TuN/6gj7FknGOYPZkY9g92ny+gEYV
iCdBnGF0JDfOWRMBnH7xw4ISHFk7ZBhsNlb0U/sfBB+LfL65a4OnT/PITgtW3D2LbAS/z8seuqmc
zIAwZhqfibY1vh+i2ORT5cym8UHVpWQeNd+Z7/pKEL5/1B9Urdr3loX3aHEwz6nZT2kMnpN1FPp/
fVZASEWloY4khASB/h+0ACw3h4aAv4cdYYk1rpLzEGCmCo6D0K1DQ8H+KaE7+E7ASMuv11C9HHx9
881vsons/J1sqE1B6CNeooHHcN4aNqk53edm0lOjwQMeRuwSnz6NuHrsnn4u7G4rQfFfBr38TxMd
AmdKus9FrHU7t8GNXAo6EtrMm2cOmDGOXJWWVldIWY8bQrTlB1VFrkeG9cHJNz29ppWrU2xX17SZ
w/UIhrdGJaz28wNerklpAIZJm5YyZ4RUoloQUGrHeaMkn1fwR405IiBokUo+8A+Dx/1gH2VunvDm
Bj4q78nY75JIq/bcaJRt1DnlGdDzwMjLOsxS2T7YH1PWqrraViklswMYVgka7PEVjx7TeZmUUF1f
neXlfBVDl7TGOgoXEgwaAUxEKm0kKqtRpIu8kb6BRSNvtDPBZGaxw3QvP4khNrX25LslMmxpQuf2
sCa9WqKItX93DD8cJL4wvmfRZMaafakN7LNyTMyjpJ5sijjFVeuzKYHBXmW/Nf3I6Kf48aCb/JoU
oaUMa4uqfoU1uXJUqYuGCglC+HMnR7M6ylanBikSK7AyTfpimUBKLMPh1zo9HtltJnqXk1oGQBvn
uu6zMOxVzJRMq3+XzhXIhNyV8HfAVCMHvTjDl5bUk16BJoezVYtMH7dlFUcoR8zP4N8G8gktapHY
KW0dtzXwW6h5PL1x2DpVOEngTOp9+d99hc4F+QXUQCRI+XGbYJyOop3ZecofjR8wUB1HbxoiVr8d
kRkz7xdsXm29RxgY/QRbEQ6A7HX3JovByXWnaxOprnFTpt4abSX5pYXc0dgsayHY8pwoYkxLGL/C
+v6zFdgynT1mVzbbhTtE+xM1/jYZhw3S1qfDAI67zakU+D/KFTSX5nNQ3mZyyhdOXxLGIhRxv7oi
XdAguDREiniLecbfy+e8rKnc9pDEMkgl06AUE3aQzdb/CfF3sudZY7leRoIrY64Zl0HeABSuT+WR
is2x8TQWEOJyXebRDkHygFYbdJaZHzoHMZ0n5SBsp/tfird52l19Lr42oS/GTXeqKFdNXGMdtmfJ
Lnwo2GfVL7WnyzVmSi4q/qK+DKsu3fJZ5uFclHXGTn+0mJZ1kekydUp7UfvCxOCEOSVo/fbOX898
bFcYRgFukyWe0zeBDHp0imuTGydGYl4ENqt3kWHEEmuPLSZuZwnVZQbhiSAjF5pdkyFaMAqWp+j7
nHoj+20QDt11jqUhGqqU5aaIW1pkzZ1VW5AfqJE2lYitzRKq5vTDRan2s1+/t239+qHXxIya/qmt
KmgZfjVmYbxj/GzH4Am7YsMuvON4eSzT1WdTxGMK8i/Qwn1BUDR3u4evc6uyqK+txfr3UD++ZC9N
SRFF3ORngDgH8ubqyomH3bODLrzx+/nTKiYAuAqJ4GUqa2t14bLW4n/ZeRaqcye6FeLyVr9BT8bD
ZSvpbcgO1BlZvu1yPWy+E705hxhClot4nZMcj8LXCwW+S5Gw+TcGcC97R8bYw1ZLY5lfPL2IGnJK
IiIbrd9TEy/iuIKCdf2LtAlP5gPEm9Y5giJ//1nF0aDABO7oPpk6I6DrsfgwBpYY+NbDMWzDUTiN
jhT5229dyb1JHOicHNsoqzBLb08tHh1B75lq2AxoUFTp/T6o1Cekj8o2Dimcu1U3cgyns2PuZa7M
zudFsH5xsX/rell+OsEykOJ4A0Bd8Zu78tHpZs8K1/6Z6udrxXcmpJO1l/4LLbL5dQnjlBzNXphg
l2tfuUsrJOjSXHm+Cl4VYQTs3dZ+Twj1PrEX+hRX4RhO8BvGsnPIuACE3IKFoMfwZZKari1EyJet
SmrCBpPD3OiJthNVzpDHMERmQgEM1fJShhYywLYBYzYV25bukg0VzF0L5P44cPD5w1iumY1Xy36b
zLAzMuIC2IJebCAvhQPlbH6W/OZF2Ht9sYqA9XjA5NtwaS0bE/GjXLafgEejRW7pnzfP4kwfIk6x
JNlP30xN6eVg5YMdxiL+AvqEt9Ljq1nkJkTyAcTvbWqHg+NXoL9GeRTtuPphKfVVoaHX0qIkGH9O
DUuIX0YNFe7pJtfNG6ElEoAnyS14by8RVhvTBvDpYta0i8McIbBfcjexQV4kOuqFKhQJfHKH5Ibf
r1s9stujS2+wr2dMCBW3Kwu6A5UdyqKoGt8wzUbqXbjTxLU1nQ9iL/WaShByh0suXjZX456Kio4w
97a1Z4zhqJhdMuI1sQztG3nGptFqUU2EPTsnFySw2aZ6WweMB5/qM5QLL0M2qjJV3cJ9g/1UQnBi
Y7jPe+roGnaFeW9RDT09iIEsGYB2ZS6WVkpdRovTLdqYRLJvwuz3ZocMWAvq0+Tf7SMiCzfXob0B
lnxETxqYNjGLy4W5yGqBNjKw6m3wYV1ov5dtmsHF4gB32YzK9qRRVl0LDFoSPX58FvrAXO62qc+W
Oqe88cyXr4dsS5JoNsTiRmfiX/3DTyBjA8mkF2Wt99GRsUf4fYn1/eY6dezXqHvAzqCcH+O8CGo0
bB0c/NQWX9CScNCsK1IBg73Aby+hzVgy92YdkkAa2o7/IeIvI18kkSoX8T4MFNey1mTh+Ce47lgV
N67ksAk9RbGcUd7mdZE/KGOrEOio5j6jPc3OufEuGb6hauEdLlC/G7Bk84GyVvtv1M4+yXIzaH65
ktRbIDI4amYDg81AjaVRxctXoem6AxTN/ErH+LAirUfaNe5bEm7Kld9ydkxxe1vWuhEhFolEdw5Y
rPmABSjqSOtlPsgOumeUL5TLbo0gy7lfE1V+eISAVnOvzdKnRvD+etsu6ktVxPbj9ZqnhzEsyJwU
yK/FGuYSQxHxU+Nbha/yGszwgJVHniOJqVgC9Ez6o4nvL+3VWwv+xljflWl0n8u59M7ClOm2Y44N
8QYcv2Xw8oi9o3ZYeTx57iptRcwbxdidfzvtok0T1mRI/yqDnkXj91hrqFZNo7OBF6P2kz5On0ue
u9eSP3oycGinKNJFWCAMGYfKWPbiMFqpG9dZNElwm5Wl1WW4RiSNout7DU/2bM7gPLrguhGH2GDI
atVD82NYMWp7NxuJRmoFWtHIfrWG8G9YkdyjlylpbN8p+voWYGgfQPbUbPg3o79UwSeuNPNMQRAC
jZqKBU3mW941qOMmpw9hGQzC4YwOIfVKPRxaS63e+a4sxMNuHXVjfvrIIHFHlEmKEhheapHrQzu5
vL0Xj8HuPGsGDz5vKHQdo/FOloM/A+ZyoHm6ZDlnuKn580HUKii6NVLUoTy5qTLq+iedIg7jRyT4
7Pg3avQN86Iu1ZvzjyuRAzDDl6l3UpaCgiu5phgCnPT7yxc9FrSL5u1P+glEfzNNk/+8Mu/1a/G7
qO4rQc+HoOR9cRTQosgyWTHgs8zQRrp9uRRj6wgjMrhhKfR83KIW4Z7UQa27RCjPFFqha31Ldk5v
v+6tjF0fP+QKJBmeCIRHUvkNaKZsTOmXaHfxz162v21ZjhvodFPCbgvQjIiSK/K/94xSYMbFcivv
mbDrr/syCrpLax3ojzDfp7hwsL66SfHFG9wmajuLjq4WauLAxq/GOW6T4KywK1ybpL79Rng8PfQ2
UOFpi85x5YZf+a8D/SMOYviijMRvGWV7i/yYYAUcbyjXHY5OlGO1m0baipNYTLcsWlsrVq5v4MIG
C4yJfsVpDqiPf67YtIiOv6fWrmx12EyMw4vvYl3dwH9tKXRM+boTAJ+x+AFSACsoObVMhUhfKVi6
X09suHkB+ebqXAEkVPJA7ufSTD36u1iWhNhzxXLvvp1gjNty+ZiQ8p7eed9sF0SEEi7vkEgaG5W8
16ndmxyKBGJp89mWLPeUIYV87Po3HXdQII5KgWS2T/kWj2S9Jn30u0bYtTU4zlw9HkaMpPRkJEko
MdAkPBwNjjI/lUB5b3NCANh1wbfzmqco0Vu6XTnM3bZMrpeY/WZ1kC/+8tZcaxl/ZBqlaZ9DySH/
1kPypVRGH8rjuBHTKhimODydVFQbmTE4Gh0JDhAa5ztp1b9HSR8wEUnl1W4EK+EuIUszvOYPE8Nn
cNZSLMdxwUeZKXV2Myv+Ra7T6+iKgm6wyfVyk7tVQqSAm7U9rsYuUY8lmwYJ9xuKvmd254Fd51bp
UPzLrU7vTuDAGHkgx/tKC0yzcbmFIUoCUKoFeacnB1bUHNi0j5DeCSxnNHscBAcyHN3khM10AEMT
RTS8G+45j9N9+EoORID+c/9mCbpvHCxQlXZBPyE4cSBh4rEnHs+mampZKWW9gk+z9eIr55M2JMlo
oraOlDyWQOl6bc1fZSWaCP7bwWO0CgK48yHhu8UQvyODywUNXDr4tFFxXiPxjZAXAeNBfGm+DjDp
TqilLOMMae296bWV7q4XFSnmMRHppQWUFxU5NtLYljFzL+8Cq8sBtdU4u44/8ATX2rlIk09CqrKz
d4wRmWjHFSfagY2m4PY3AEWFwYRytbnHO8Pm8NynlbmgMKoyXDGoM1LAP9ieYQ9WdMcRAJVFctE+
EkDRXb9ysS9QSarJ8GzRcnGaw8PQ5c8l9OBPn7Gv7r0dUHEZFHCJIEr0oN448lilSnwqMOjFwby/
7vV6DlX5fA4M6zq8r1/wIihW0M3Q++7ynjob6gpcUeG0/FDfI5GRZyUGLH+jtYf0a3bUhColnDPk
o9/pt9Ysj2YlfX64VKi7S2Tz7dodbnUaz8MX/IfuQt4JenurDqoKmqdUFVJxyc8FAJNUjKWq7l+5
RsBJ8pLBkvi0I7EuiWZhcrDN0b5heRzlJ6GihzHqiP7fo7XGTcqd8gimNzGw4NO0glCfqiFQiZE9
IuRge04qfh7EUA/3fWdMXjp1SumgKPU+yvF1VVVqzGIr+enwdq4f4jA+Ok8GrzE9Z/Ur0KdrLRuv
rUkDDSChtFS1jFZP90PoszcYRvHfGA7PEYNXfYLuNrkwz8k1LmO6VqM+YOkGn4HjXvtVCyZYpZ1W
98LOUk1RETuF2pD858t8IjmocXzpJeUKbExHh64Rhl//GnLqbG7nrnBmMbudbagt1xxn4aXQkgpL
LQ9pp/RqzuUlUJWKQDHdIc7mGtFKrSThj8SWpZLdiBED+tQvavulZU6K7x1rmPovnWrD8DWoJM/a
oMTonOCYXpkCGDi84/uTs95GnHwc6PyOlW89hOCXH0fZHECP+CupfLT1QwbIQT3YeObre3JoFu2R
3gK7Teu5t8s6CbQ7NHuqygneo4hH3WxDiS23xbl6ja6aFucfj4AkgbxDvwqGMwVwZHFOlqh4s1ZQ
18lDFdmwfFctkDb2TdaP68yVIAn/QeHhOPXHjR1L96eKxcnWsPQJefAcZ5/PI1R+DY0brM6ULznV
1HPUH3ePw2HYqTcVUxni1puVhaOmlzoQaZFvaklq/oUyqsEO6aXBuugk7LdGnr+bnM4lVj15t/vG
gjtWhM2RVf9bfXxtTLYbQW0WA7yqB/x1kk9d9Oyr3M/uNuY8GX2gFWyAirIdBDlBRUMJ8kmsu+no
0kXmYKJ5Zkq11r2gul/aneTzN80FevUMAuA9FOP/bvw3F0oUln04nBsMRgGOmMoTh2tzs4bJe9cq
He2CEXBoFZ6HquqC1tqOQ4wqLD6HJDRhkk/5o1yb2UMrw6vaQ5Zhdk7hhd+XlaLesAZhGI90uOIg
PgEcI8hBZAAQskR/Kif4IQwhBfGRaCZkWBkX7EaMsDVjUkOMzFJtQstDcoSA03WvFjOXoicdur1W
qc5BpWPlYkDqMKdeegz9pWBU+TiKzFJV+GNpGSG2hPROMhhaJgC8tANEp/7pNWJEfGSXTxG4HUDu
M0fx8ZsXoXZ3p8v1dlBOj8a8LioBa3q+f4r2cZEHW6g5S4++3L1p5g4oUvJ6ncdguvyMlAk6THSH
5TR8Gt3VZRx4gBPGitmGmBprSqKY2DQXn9Xyu4E0WRZ2N5Pc3sfcRwiLYw75u5uKu6tDiV4VuyFB
ViC79HN+SrMK511P03euf9Ee6LFZDm3U7if/sHIb0V+Yhtf7/XcsW0dZ6qa4Eszbwtk8BiNfy0C+
xkH8PV4D2a73R7KEzLOTBY8rh9w6QO/BFydz34YkyNnylzp8LznAT3yte5ftpCUt9Trg4FVCKZug
9NC0LtZZLa83FtZeSaWW2wQJYGVVXVr5+kfHiUpB215RBttK9iPFxUd6yD5EY+lexWYOQ/sjYgXk
htlCeIvfTOl9wmZICUjnm6/9OAhKZi3Fswy++vbsPV8Hi1wONAkoxq64PKzEXyVMQD0gciN7pXcO
zh+pkJrr98nVzyXkbn7xzmZCLVlczvmgpEQIMKy05VNLzwQg1kKi3W9L2oPXTInfs5a+YpK1Ig83
QFufbTSOQUwATSLPgL+9p4a54m1Qy9KsHe84HmzsNfOXHwgbbAAwlF/8CkNK2q+cmDy6SMkaPyIb
dFu5w2JzHKKT4Tt4zLuGXFS4TUIwAJuzzB59z9s2qS3KjFPCw1OuXa+dLcSPM0PDFrzcqc8w2aoF
QxPJk5uN347OGNEhSXls3QFPRN+Vn80MzhOOHp4daUUFVRaoMfkXCCg6P+KuiDVOA9PBUckMP5ZE
8bUgcI+/r5Fai65VVBsQg7CW4BeimGYa1ywgX/y/PUXIcVaVX5eYQQAese+pOIATfraXtjP5A4Ef
6WxPDncV67EUa24pHBYXlTiJBAHFvSUS/pwzJfZ6jb2LYXvLnc5+x3gV7WJo21wLEC5ydmaJzLIO
w9Svou5cRqnnKdwbTRww0u4jzG4G7+mOd4uATnGLnxbVpCYLbVd0BIHd5XB8ehxN78yZQGDS7Tnl
XYBQHBPgTj7w0VohaWynIKfQXProuTr0D7v7ijS2GQGS546mI5+gm7ZMtzgUJ7tZaovL4VifcHWs
k25EAe4z6vB0swyS3iBdUa7W8pnwXmyj9uvDqxyU1+uYhOfnU+DdhPNXLZ2nEw/PIm0Q49tHaLB8
Xl3IvJbycGUATBpEaOL/hmankgTnxtrKcglykZDWlHUo/0UFDMt+KAyxiorefs8TMGLL3q0EGbn7
Ccozh1mTKhhR5Vm/rllGrqBISIGVsw3+DoXabRHR1NpQsGt7Xq39Zyz8nIu39SCXZSyvrRDck0Zq
Na49mBUsDzb8qkupjk1ouetunJohhQN2/OhAFagvofx1CnoVTcmTnFJ8zgycltXT0dGBMh7a9Plh
tqGjPKSvaL5xBqGS8SAzC10N0ZttERtedCv0BdFyM5jGYgIc1ksrb3g2Dy5719zIIBfwAgYyN0Mz
odVQGub3CYZ0K908qFJZKlHUJEc/k8ErhJnrhTgF+aBIV/DbwPg2U8y2adusNA2oSuGFb5ZC9t9O
V9hkanRXPG7DMl2N1ZUZuxscRugBsAvKV9QuZN9f9NqaKEMdql+ke4jxtqa23gYCU0qqZzC7kZM7
kJBpyUmpunt2ZHxOIexJ7uYgVoncSnk0PdWAYSQOqgv/v35TadhrCu3q7Jwy8CknsFB6M/wv4uob
pso7A2ruCeuAlXaIMQcm0PpSDpszugchqRlJewnezQkyfeZcMmQfNqEuc1dYhsqWRCb+jku9D15v
rUad6nuzvpu2tzwSG+xWiL94m4npOecrYCdU2e6U52EMagXUI7HhZlnrLkDuzcH/adUZHxQgH7dg
GCQ3s4I7yc8SYaGNP3k2dg9Ma9AsRjEQmyasukUmxmkTVxQVDmliGBQTuPDjZdc1aL16N2Py7ZWu
pA2/ci7gSW7yfMZmWwuRPq+UkjIcuoIgWEeJB7b8mAD+EB9tfGat4NUIuj+cZzvbqgkod/DKcX73
WVxvRjpc1AyNlkz705MX7IdNIHWLXD8P8XNqetesNo32Mbk1tIZJJfi95Ja9zjBUthC9Llh13/Xr
0IgzDaAh58ghxx2kOuQRu4AuFGn4/aojYElvyxCtfd6zeeDzdcPVnVHT8fuEm4kZUYdbcgqV8EDW
7iBXR2Mp94kjDV5VRGahr3FRAgLbAvij4Tw7KlC23DceH8isJuylnrUFvRpbmxpuPwZZOF7E9Joh
K0+ePbrapHzDOQig3OhTdnKeOqzcoAc8PeZDM7GajuanXdcylS2kHXuR5i9875R/4U+3H+BHonYT
r/6s8kYOADNx5fspTX9J7Rjg63N9bZAJIgqBvqI9uREO45PienoiDLGnBuwcJ5STmRGP99JSiXhC
EETePXiY3eUe0OcUUvKGfou9VEws9dX7dwr5mSyrS/JMSqJc4XWSgs6JQ1Ek93szqrxAqnmib38M
FdH1i1F2uZtEBB1+n8ggj6CKgtKxmX0kGEAl+evWEpko5zW707eP0meaRSKJlNVhBiZzeqmo4S2z
dPJXkwW1VBZ1Xyqq1CIIOFJpM2HXwpuGZPDvkFwQgyKZF/bUtGbmvoeNPJ8ZZ2lT0qu87OfkPXA4
ISYHTScIKkka8QYMwFY3BSFqgDlfOVgXuCaU14rbBWkamQ7FLWAyR+7TKOKeKU4B9s5g646Ua0AV
4b5K8GH9ZvaL0IvYrypd9kFoTKBp0rp0rK2sZCXL/q8pFy60kuHB2UeQ/qhwWYdSF/1FhnB3+S0G
VSQlgh7142VFLP+0c8qE/vU1vuRr8h52kK4OJ9dzY1USTPx0Nmabrycr5H5aNuFGvgl3XPsumbJu
GPRmZ0VKPiFiLhpMcHZ9jPgRqwl8l2b2Jhh4dMYKLjOoRQaIGmSyEgLNzxTogOaqBxo4/Nk1VUst
lgHCL/G9pjnb0k9Rsa7vWcn6JnKIi5oziKuFPeBTvwO+g+XY6r8UFtNuJufWsFnRW3IkgDQhwits
HAPS4+Xo6Rh+agXAXxnftWtUXK0z70/G2vdDM6cmdmxjxq4/Ixvj5VcaWCw9hxV1EpC/QzeaF78l
TgE3bfkMznsxu/zthkq8CsyaRiMEasf3xOesy4vjrn1uw5RB5RIb6sNhebYOp3zdasF0dvS2TFAS
d1ViPGPAxYbYMOh3mwwDkljktHN85LNK9pMmT3c4k84SkGkCxCGkFiAwmnSo55mrq2zPOLV9pUIg
/Yywj1D5ax76XbPUSjT766hJCJw/JPWUn4d3V0863h2hvSidBt5vPCPjLe+QlMcLWlnX8VCVqjaH
Zt/sk7ttTjNwifNApG1C35wgDkFGoQ1c/3P1PrBvTXB37xPF3ITikviRAicsmkhyvvNqlq/OqUuH
7f2v2gZBfRiAzQGvzx2VLPnpnqdZ/764GVOQfqlbkNKCn9Mm+scHFhGQNOZpFaZkhZlW2RB6AHSz
4uTge+0m0HZpqEPZeURQbBkqHQC2TU/PB9UbNrz71Sx3tjTgJfX4b/tV0uGPftv+TYFpjBeeK/HM
dfmHf4RqCUI1QvJrOTedwjxyGWGzRuiko0kBiQ1rj1zLmmlLKUVITX0TBeNOEWI7pzoEzkcRR3m1
TSemGbfGjSlDJX2Utdq8HUVlJGjRP1zeF70GQRm5hhv9CdHkjqJQtgC8/KCi9tAtPPVwM8MTUF2E
TgxtaHI1Yo8CEUN+cW4UMGNQ+MQdQqkVsLFHpqn7Kv5WRZ5Z9RzWRLX8xVfOINLQe/1sY71BsBbJ
kKzTzW3t9OyCG8xEiqHFQiLMwA6+di/OzwcIe/CUiEENllsyc+h19cgDaYo0PJh/0OTaVTe/0Kw1
ORRC4RFV6jOQB4VAmaJ3exR07zQE+yv9fP5z0foiDaEauOtHw9JK8KWkOn9sRGqkYSluMUBKsEyb
/UfFBBnGYhi6iSZGFrx5YWZNVe+h19LLkUY1ns8/VCpGIUPdf6WXD6ZVH88Jx0Nch7q27nuwIR0i
YfYu5+3sbHS14bNQ8NBbXMjWYpzdBrf+0dpMo2C6pjU3C4lQ/llZDzk2KjkmyoQ1McOgwof4qxUD
Ph2txOgEz16WkiyXJnaetwUUNzmmJfUpI+MEuJiMY+cqHuPwXYoG76xCH6qgCcDw20tECzkYI+16
XsuSf3PYviihHSia0ZKP0MiRFzsKBkLo/QOpVOU+J3WpOfNyMtBBu1nnOuQS/16x9jqK4+4SMU0q
uwq0nDQbJz9R80g7WZga35P26XqhphZqMEGclPGTxky1E1ynh3a1FLDgLvzyTnLUy/M05y7ozVc/
mifswIBWeDMEBZ6Vs9WxUu64f84NBPo8aB5oWfWFVkIKblyz/bq6FcsHerDk9ykLE56CbdwMiumQ
dAF5L+Ul0DadFVFnusBF0gEVeLh4SqHCU00yjSwJ6qJi73BLjob+VQ8xjjTxkagVwJDU2ivhIkQC
6w5NOKqYLI9pHnM2kmspJ9EMI+praaC2WG8Wt/8rTZAzjZpG0HJMYpmhbhdpSdEA57TupMJKZtah
i/Fn4snvfpwxXI0gAOLx9/w0n3empnWi7YMdAvNSN4Bt8BM5eNNRLEkkB7HPRY059Kf94zf7HVrh
UUaMqOTCEhbZQdKviFQgJED24vuG6yYOuwUL0tJ/yrT9Wo8HsfVoSk263K/hMN9lTlwdwVmecx8E
wbuHRAflcOMOaRJ6n2jhTyAOH8IXgm1AzdAqUjpJTOycAd+2nuKqbEqXuMpBEDzaJNAaNNBooDJA
NWDb4gN0HU9b6EuVaV3SVVfJwPVbDbYy/3cfxXzwBp+NAJ00TnzKt+mvtj8BrqmcoCR3ncuHn2zm
B6gWfFQie62wILVKMLlZBh0ZrBUDewtNeQ3LmFb+QeMFkBFLHUWNCCQEchoBKsrAP8nMgnSxeHTf
+ZXlJ4N2bin9IlhApS8f6+mf0bt3R8pzQGaZwau5rIntVMsV118Lc4ebZOXuuaqMQs76nQCxLVr2
jGgq9NNGuUzvGH6UT//XAin5sGHNw1lJ+1rjPwwXecerLxNzptzW+EB8nq9cLsoo4PAf2T2E28RF
hwV4ibJK0I/B9jaI1tGVaiKMZX984TQ8JJIlIrnevakF71ZsoyT/n80brxlG2O78nTmLwVRd4NjY
LsIswdhiQaQzfAvSS3YAct8Uy/zU2EhzS5wSPQ/V2ZOoBLOtbtvu/S6qPA5/cMp2n0jyV1I1enXP
o0cryMJ0L+lCsHRDMAr/qQfPXlVTHcdZqzV0P6tEaDJC04Ew/cvd/b3+jGkkuBAC0Qh349q8o5cN
ARO/0lp62/lqx3VDVjuFUkP18meKGJxCwbdURXQtncHKK1R3S7J2G2XEuOTefnQVGPhD3txNZ+FX
9JVhln2J64HfN1qCsMkWdH9Vpsdc3MLhaieDKSlCwFWHRzefouOJc+GOAN6kSiNP4kCkbhJHjCIq
YAI7UtXUA+c5CSlgJwecFDX+biKL0n7NpjWYmUzMyVIeU+xTGc9mY/gN59e/9dzY7hSTDKHitd1R
oJxuFgRn8Lv/Bjfe00D7hv4SSQ53pSaeIEoNnMjsYATr/VaWyntItP7BSp3M/kEOsIsKhQ4qVNCT
c68XYfKH10DPqrqjtUdFJGuEkCvOuoMjRjS3wISmyGtgR6x27Ff/if3t4QIj77G5oGCrG+Xcd+eJ
k4Vifsr/bX8vwnI0SW0NmJur19o6aDbgR2FpomJukBdiKxD7cTvG0IbmpAINSNSq0YozrSbDKw4c
ZYNEW6W+UfZo/sD5yW7jtDn0DYxRQDW4vQYQXGQVedL4VA+ObDseaH24q+kSEs46uMXG0zfDFJmK
C8QFLdeR+IivEXu/HLCSibZs8ezJBS3OjeWs5+lXmyWswxXztQJtFELyvAi3Pkph9kITPhgWnBxY
A0sGlUipdEjn0iDr3Hqm/VMI9ygbHatWC6HgoSFp55v3ARtu5fuckGig78OrYW1Bt5yfWnQvY7ZD
er1p4Uj+VVWxg0BtLjN7ihcNNgkyK2akmVTIogSuJcNkGRFopiD2fNQ4CQAub/bMX3xcCLrGCqlY
rGXJj0mKTH9qYgHELGYHZKcDqZlgUb3BIPZaDVAwZOE9+7QIKMgjIxMUtec/A4vvFzLgWODG0RyY
2hlcgk+7bChSsg7JRAAQOnbnOaREE2HKx5SQbxEnPYDQZ6x9SgmJ5X0vdHjd0aY2lHBsIZ6hDq23
BCKijrbAGpgbdEDy3ClelNcMYqu5Va246KUKRrBjD0+HKTvk70RpmujxLshDQsEWCYV+MiGbXWnp
/ebY0nLtK2RxAimYKKZO0QZrB+I17G9sBrVOpY4DNwN4blUpYDJAFrrKR2Y1K5tPNmlcr2qV+MRQ
EJgk37wq6IUGg6cA6RNVUlBFw/Ja3e5jYA6pZiEJa+nCyvfvcMTkNobmI8nDhabAqdaqymCCvyxP
Dl7e+G5MofxD+N8c5D/S0e5jXvSFu6dMO1NnPyxZjJbIhualuv3LZCR+4YQdJLaNLaIqsPfkB4nO
3NwKj69oj6qO+ykIDcw66LxQjd5J3NyizjMVbB1YyNpanvPOMBbJM1SrjTU+pzXiSTW02v+o8Heb
l1X/jXUPEVUAqPNkTlTWXo6fJTYzGiAJdOGsV23v+IGMKeB+79NpEoAta8Uwj5UrK1n0Wi5j1qTv
L/j+TW64oqb1W02nkXZZsNeh/ml+wQntytg4LiegRGaLeuUAXS8rtgTOkZvOV/DPlEkjMrMvsRAv
eW1GpDM8+u0+5Nd/T3XzfjDPonFD1ippxM/Ebkg+q1w/kc+TEHZmpAV/Y1ECMDDIkufahFIBygFB
3+FYncR0j5Jgp4MSRzx/TMYW6fo0027i9KF1gtEpmtqWtitjoKeJXky1D2FUsL9o8Chzjk0VMTsl
pe/Vg3AJ+bxbL/KhpyqvnTAtukzbI0XPhMgZtJNXl4y45zLx526jUAcgc+JFFrS1aSkAqioM+gJi
F/ikMl7Dw3+ksytDhmAYtURU8hawJK5yxYBS/O2XIIrhLPajliTgV4T22E9t9x5Ken5jFgxDn1T2
IQkvE+VgMlRLeR3KP8dzHWCQnwIKe50YqE6Gia9HFH5mtbX20zGsLTimCg8iUiHv3POwocpA3ggc
dMiTH3l4gj/fm3S594ZBaIG94Um9EI8sAmgciw8OF3aSkSFQbYPUqE5M5kkCV4CQTWSljl9kfCZW
HhdCcMViKVNEW5/YxWWaF6wN0ygCoHun7oIgA0xBb+3zuna7ff9tqO2i7fgiyBVdLtgu4aWfIktS
lNeN5BxW6GnWNgdxCFV5S+wSOFbd6f5uaH8sXddxERbkOEjnHfURVSzaF2XUHKl1LnQ6HsdOA8Ji
qswzD6M53wMiPSWjTkUnUYzjE0VzyJkdxYnnDSPUnG9NjXQREUVdIV8u3MAjmIcM4er/QHGsn/nQ
pJ711PX9PKg2WWh7rLGn1rAUoUNyxDqEMeUU0cksXdSKdjt3CvJYEZytqNjoC5yZwwzSni7nN/f+
FI/tZJP7DNJfrUv3FufQ2zW/grTjcE7TVvmdnDiFTYpbG/UA0dWzzc4liDZ9ArtUbOjU0kkylvID
BIbhVO4Xy8QRwCjSfP6A3uaVoGZSGodCJp0VzKpYORxvzr7Snn3mmY2iQbbDUxtmq06dYHCRU983
ZLT3dLaE6ILsOIn+TUKzpJhZmyJ3qx420g9DSMn97hzhUAr1PGkS2tpgWvP4V2b6dR39CQYPUvL6
RdXayMJLMoKS++q51skMWc1wDa8coo49RvDA5S2EbNYTjfEwR9xQfjZjLC4232saoAwZ+Oe1Ifwn
dJL+V15ctN/jr0zr66SveWxeTQkLTwhUr8bRNJuY+AEBlOAgB8DfbbfgO+fD6pfXzVQ/YJMl2E30
cJ+xt8UAW7jQGAPnKv52fROGbVFMnnRNBtoaRJHZQkSCXqWbiiBJG+pJiEPMSFl4EbFacmfTPIZ3
tcCB+uUPNFA9eTn8QdfLNz4BWs+tBglfWJedrcyiqMZeJU6RI9zgwinRbzmtDMV4pD1LZIxQtfxT
WJcpnhwtTGd5b1u25BpauderJsmwVFuU1bILOXTqJMe5S9Nww0fZNvjBpqr3vmolsHI1h8XgFj6H
5fh5ob3jl2AIL6eRk9/UBOw/Sss/zlCeaQ2EcM99izdNmODZM031P23teCcvWmfInJNSl6rl3H0x
sTGfD3Z9LPOYgF6AmJAuqEra5qacymGRH5wcXx4zD9gWgRF136J8s6E4B3fvr2/ImB+QIkwOsWnS
dInYCvsHysldBdjjHzB8Pw1O8IyaBUyss7JQ4snllpws74sefHG2kgxM/fH8Cg/hDXSziCEyWY5d
GNepX6dBQpJIMZfMDWrHDq5JldyqvzzlW6tn3hU8JcoXRfpDJ2ypPeUaFpkNM8z5nattbiqa5YTb
79ybNqfw2a/zIA9BqwE9pA9W2SkSLqJTFifcSDqYMYQXjdbteoiGecUDPsvSANz32JMAjCOKpa7g
K84ICH/oB1k6QHdNLBbsuUkanjz1AoQrXziJTnh/uzWGfGuz5KLdnmAWahfX9liJAIa4Ko01kAhi
MVFz0qrIpKzRy/Wranr8OjunngA7BLQjfUhlpEyYwAIjUgMqWBYzRrfk2Bjb/xWen8YpHeVbWMe/
WnWFHPKn5z0mA3+nwNyvktsepdM0USffPaO+3UUB1A4gzIPmVzIYRNBOewThEIrVzZsHznkO8inW
vWpsKY/4svbGBzKZLI5aXVCNYnNHnH7w92zL/c22BQ4rVYNKzf6ZIhlYIAETBj6e5+Om7z9JBk4J
U90NSLC5VpnJYrKFfJDILpezkriFrbg86yZ9rTA6ESvOzAEfh41tRAy+2GrxACxYkOaMbe+TQQRK
VN7rGrHnxIwRlzmIy+zAOzH7J6htymf+Oq+3F8g8VPx8i6S84cUP8hYQX9Ol1vFG2/LpjmMlUImn
yrOpKiSC5EgPubZiY+XLhEj8/0rcMmkHKGguRpc7OtYvJ3CGq0Wyi4ds5BBQrybsXNg/JYrYpupC
qULGxNr15NqYEeRazYxrFdWpGDWCmAWee0CyPjUz0hBSokgYd5YLm4QDa9jJ5iXndS71TxRhJGMS
Al8wwlcp0hMKmzY10+IgTTE3IBmxLq0qSFGgD/1lpDrEftwlafFfdzA8pz3cfIi4pkOqZo7k3NDb
XIAHoOYMSlaJHwIuBS+DMVtm4hN7FdeZE+E9EHb5n9CQbqXeaCz6vBuQEfmI+P9pgdbv0czO/Uz9
TVdy3CKgOo5zlRBdPdEbuA9R9RKPLprOSkXXgu377/Q3Oy0yG7qUhEJ6T7DMYme3fzhEkD2NOB2r
RihZ3ptUjWpNT0qxYqlgxv6oXSrxF87PvnYoolkkn7xDAcDfB1XL9L9I+f7yjjMz7qGNPqtgYHpQ
fCq6ttOQsRgBdCXs4TSE2ZwvQnVZWQ4Mwwk28AI5Y9/FCp2seCAjdBM6dMU2sRpvaXEyKU+c758t
0cP9I5A0LVWE4Y7evjDgD+uDEsyP0ivh7jW12Icue7gdbXPb5jKKTbSg7mVPYMAGRdbnRJh6fLey
yk/lzNuHVzSoAALQjpq+uQhm6aqCOwAXOkcJtPfXjRjBEzD/Xo4id9I43t6ErOVjxh9gOlUoVJcG
UvTpevXRjcgiGjpZyYYjfsOS3iFnbrgAZ4uflmxlwgHI3jesr5a3HthOimIvDS/mi4Z+39POOLgD
BpEEoxNXjXcjDRCrJy1IY8Ub9KXnif9ycbvg9EgyWAPda0crmEbd8QHfIck0NiYirxOrqReld7Nf
qnGQAe72t4bgHC6qpY9RSIT8vZMLfU/w+iJMlw1E/uJ7KJh7IeKuhDLsyihPrM8hLvZs+ujDDs4i
KWBiPl9K49ayswvcXEw29mo1D294bk/Uz9M/D7/Wsu9d8gsggx+gNidmoeJs4KkzjjkTfDzpL6Xf
wC7wXp3Ky8mveyWEJLKHMzo1Ih9HOaoe9sUZFG1mzNuVSivBVvdzq9+i4KPo/ocjId0iBtBOWif1
ZBH+Z9NGzRdN4TYIH87wXdJs11wb72lKB0lLtQss3yK5JANnDrv+f1JKRSXexBQ6VYl8CUmSkBab
/9JCBRYEyJm566C7m/J+pGyiiw+HeiQk1t5WjnDp9SaE1kyQWqbP01jw01CwfpKSGKAu/ocS20vG
z54rZoVEIlnJi/Aa9WD3m1FXan4tZIr7piI5lAXVD8B4yC/NvfiBg8vl1UzJt88r0TCrjZBYsm1N
8CJdOkjz6zYtVQxi+ZuwxUoyNoA7yOXa6013q3L/1NPOnJeklbw/DmC+hmTCgiBD3yHGOpm8KBao
HAL3Lc/DsnGKAZqadTfuu85+CCeUeVOxyX6Ct7U6AB5wPaD2VmvIwhrU0NA45/zE23GUcaJ3jJkL
yQn/is8z1BKrlcnPcXRZayZemq1gxMX+ZIBhs3Xh29oLRiR9LjhxvSzL+lBn5iWN15HVkujCLgk0
A6rlbcZeTKh/+i3cGqF3u9MjKAkZG4Hf1LlVvNk7ifrq11KuZN9bo8wPGZZ8EWJkWAcskSa6aIfe
J1/Bl7m9KIJEvyGKtlIXmOnLKd40Bqa8W9oKz1kdbiwBCa9Gz47gbvToUlCZ0qIOToxZqPW+IvEy
0NDeZ/MxbDDbFJkIejEFrOLvVZFVAcWdzxopjJX6d97CEi+FS1ZM7D14r0D2no1xqXJ3UFFF34on
+zyggfKF7buDKKYusznMypemRXqsU7yKLnndbz9Ib9qr4U7N8/Y6HRUTljckRFudPVpAEbOBIovR
6Fswc6wgJhezzYYbCn9T5yvHab+w++kSM4J58x+w2hOzqatWDrE0KRyv5RmRVYOoVnEwGommpN4G
XuH+ilrHxQNafdn0bFrVkoL0sPESvjwmQNI+UxPRDlL2dcR0z7kcmfwtincSrQQLrTOOyTSJEC5k
+uWiEOSn3uV8P1oBi1r7LPZ5peG/SDKA7fkOkXGzSYeoKEU3psv7N4K9J534hnmySW+2JPkQGpLH
htoyXhvaIyxhjk8kTPHqxext5B9RJ8rCPrEQL91WWNIsbJSF9Bw9Lp3sRxdtidauuCMWBLizDWoE
wEFmIUEgnENaOBb4nbJOoSO1lX19e7/QH6UOsxeqiPpQmt0MUNAWxLI2ZRv9WinHmFO5kD19BujY
hNbW6BkZXdCzVQ7Vzf4n5E5u4M3qRwO0rjaNhoP9RBW4xzZ1ZqVbdXRr4ZnoKmtwIwbvja5wh0HK
2IGIqBbuJSAh6W7ju08xRV4S1+C+4VnOS69rj5NqBtIsIoURCrAjPOMGli1V6e1AyBvBJl7vlMeO
+ngTPj3qaDVvjWVs+lDd/RyLxARZOVD9OotgxzACiSu8Njoh4niuqKUd6NCb7c4uAI1Vpor7M9hU
knaezA9WwiTack/ubhwKzJEKuXPsZ7WZNOZ4DBdohYXF7AW/4+uUM21NlHN2VN3m94RNs5RyQqEv
06eIMlSH49hkiKfevfjRjpbmXNg1zPeSg6xL7DWiJyV3Zq81pNmEMRb63fl4E70RI3nozTe3G4nd
j1P+pPBIfReg9KwMIDR4aNW+fwQV6d7D7woKFhGRUDBKnaviswHgsYt7KL+WePeYdC+/vxuOylTy
foKzAPdnaizkLgIlZR0xRWFAy1peYX2rEVA/lN6Hwdh9IZPPxsEWENN2x5phmt8KC2/Npnin+8XY
qBjtmdk59xtDFghqmtEpIddAvMjvda6frfV4vj70YEIQ0lvJEgHflSRB2qtRcNCYXF68ZYOx9t7e
3hgdO7w7vPEZEF/PT9nIYh/0r1KMEn5trWlo6HQivKiBZuc0RRZM8fhfAv/SfeXTuJ+jMnssj8zs
MRFQeuvpFn6WG33zcRkH/aH8KJEx5+4MM7zoWvJLI4jCcoTwXY82zFaoSdZtwvqaq8L/jUNeZxxb
OBfMto1kBcH6VyjFum890bHq+2JzUZL8+x5BA9laGNhWkqNOlzlMmK4kOVODsrhIScPxtOu+mknE
/WHu+ldw8EEjp0DOjLzV52pXhvjstU4ncEkSH2XkTb3EtoqHMcOxCJfkiVPTmkeqn4OpqtWfRk/c
dKRzONZR1hXzAgkd+OVuoZBJM1Po2s06naYxrDyUXhlPRfk6CwPWtDGfYSvU44x6wJdySLylN2IH
XccfxVFmDbP8ZNBL7UOeuH0mRtBTM0U4O5TF5jL+LeIp9bi+gOQGSm5s3r6Uu5CGedvFu6bb8dnr
W4Q3/DOAUDzLxPf7OSAPGzCrTLCk2r8AFpVUmAauv3DxFZcXQh68Y3kKkqjsa+q7TLbZ/x7m8wb2
c6gXYYDN38ViEDTo10bChoN11otMK3fpw+XiOhaVxnqoU82Q4FYQYPew5KktUh07PjCgsZeVK3aH
wpzYi4PLOyEhsHjSqaJvpGG4daFn2sHWIAPVNKvgLUYCYIm2xwlEXO6MRqFnCxtIhfsFTFa319NI
5q5vL3IZb7bsLd084k3SLv7gRAu7JIqGw/kkivScUIdmTfF+TT7sOts3hiwAo5rxXM4iiLHziaSS
qm57XhlXHIR58S0t3farU3toycjr1CEqr8Fxe7cKYxqVMlqvNXF7rz4mxgnDaYR+Sg06DxU1KWsD
yfiDQqbc3SEOnuV0+cIe7R6XVHuCAJx1jvyy1l9mPC440bcdNOV/3gvNB5Q93wd27RUUW5EMZpO2
g7NBQQHzAl+qBoz+yKsyJm9cXteHAHQjHbIGvNavQWqkTAhpiEapRQ7PtjAQBe1xgMEk8cRHz3ti
QDlEfry1v9CpcUpA2LPrd6L2YzOwh1Tpz5H0RY4kV+RxvPzeOYlwEPfXweJfCIDnbB7vAXQWKFw1
6v7zZ7zwzWNYbdiuCI7SP951mmYL5GDEGXfL+/jf8WlpZd1ox3dPoCOhtxxoCxfXYDeUFcgIzz2z
61h3/Y5BeBBTTA/nCAw+hK5OYUZHmZwaLVKUXWNcLImOOFfwqIHTCwBBDcLVo5Dy+2/hplS06EQ1
1b5Wtu36GnMHeoplAwIVZ9uiYnYcC6xMyywFjdUb6IvmxYCsqHUeqLbUsV/9dne+o4kzJsYSukNl
EThFrSvDU2ee1WMCr+JTQHxqBzO3R1lIvqHZxPfmVgWNE1KXsg1KiQlrSJ7hZsl+ghcmZPLBybmD
iWf1klPEvfzfc4SqcFLBclWo5GdwDG06SLM53vYXAqBKYT1R+z+eq+1usxEZOkTDSN91Dw5JwX8x
jrEmEO0OsK+dfvnN0Vruk77r/MUfXzxQB4yKERB+UlvTSlfh8O4AJ7r0TvcX2gHVManh4+agmPZ5
aSY09FGbJ7eoumkuozoFA/dLkMxHEbV9eTVjM+rzXijeX/UeZ9PPaHLCPbls5LcSEyj4wVBumdAL
qJGeHs7qjUl2LZl9iW7YtONQZZiSpt0fvdjkF57MS16GfjVYIL5Gii5Iywz8dzGM0bxif76bA+xh
jG0TKbCHh/ciIhRsZaZFAnt9WJFWtU7DSkpYA9My2+7wyCtcBzroLAsQL9sHNuOEAxuL7WEpVI6F
3WSNDn+imglzTWCC2trNIKB2Z9cYLas7ry1KEs/EY02YOq9G9yL94Oas88WBTZaDTCS5A2uMJXuc
9xhHxAHUdslbO8baqVn284O89bKfFMX2Z2R4NcBCuZwiyOzuo/OfHA4doia5L5I8ENvZe4FD7HCx
qhNq74Ogl3X1Et7g20XfT1A+HzpRiZxtCJzbvnC70c8opAZKPOyX4cJMrEjrOsIpMnOgjRyqcKyV
8WEUu+xZS39B3QnN5h4uBXK3C9K8ZL0ngbIaTRGhoavSTNR41c5BsXZR6sroN2Mg2SwbetTnrWMg
Gtc6bkt33uGjnaBFLNoA0sDVkHWQXfCYepMiEUuhe5clEyWq0DrI3JCr8XoEvnZWcnN/kFou5+hs
fiJiTqkPBN8qPGwd99myxC2N0bBuLt7tziEvA1uoRraillT4gtQlSTKRpgXbsHVT1+Ph5SWM7AsW
3tM0+pE8AnhEKXlfpZwyRZUVDiALhybSIiT+r4wGMTdkwga0T/V1ws2TYyoj8FzfXwDH4KdvYAMW
yiAGK6ciEmXIDzaN3Wd33LxM/tNm/VLptgaq5X0L3CqsjPN2aqLnaB7zs6tPuxeVM7hOkfGD2xqW
wqi2P1PAF/WPoKrIDoGfU+VXC1JSU/t10FIGqNRvttK+SbnDACEyPc9nT9QfurIbbsCmZZIyGWPu
YBVGpoiA2zd6OghU21CxEya9vS/2JNKFLYcg5mRhxsMBdwdfJVC8bvl4XdmsLssAziYsrjC0lPcF
cdOrSCBN+oS8T08Ly/PNJqc3AJw4kuA6jpX1Ac78r+SLpetj7p6hkNsqlt6jzyE6R7ASVhADfChI
9ldBm/RHDtFg757pldQW3xgqgN7i/j/HYaUvTuOSQE6ZKI2z9GPLhwOaYjMS0eEO8fCtaVLyP5Ff
NCLheg77kQOur5as4q7OFvvJBzS6rNDnq0QfUFwXtmEj+dk1BNzwyptXWSjt+BeqFD7KQ2Ayarq6
czeNd+mefRritxeyFqxEe+LmREfS/7ZBcJfjq8WPEOssOdd13Jvj7B9SNk3/iaHeDzktfGA/NP9z
OCPgsRy2TYc/j4d8CxjDQlYWvtXWl4A+LhDKKqFf2gplmuwV81F/FW9KfOYLCzodbaWB2opRrthJ
gRmEO/0s/iSRxgis19VFCagyjZ3/NaH6Pz/Ny7O93yeJrslv8TLKLPQRMnnCQ0gxq+o7ir3HjmCo
mmxD6ut2G2aQ7bvLDOCtJWU30oWRGVJgmstyg4LXpPugHoW8g8wBeNH6n8Lrl5FCDFqz+egjUMTf
i2rlhsDu5mtBMLvXZQ5f/4jYr80PvNb/31Jd4l3dRAkb8ynVI/63r8Jc5k3ZpEjzTmS7uIvY1LC2
oY+Q9baJs/LP6+bgZUKube6752zMFRl5fOmRSqyz0XrMw8UJ9WH01C8F/C1BpOct2LdTsXbv43pm
rxw9ystVQeAbf4A72hAhB2SXHmKcbsPPaqfR5xsT7S383aEhBbyhfFsZYpwzJCmHFDZpqnKnTwGt
U9wUNGEOAaye9YZQGFYCcLwmOxuNaJLCT8KyrRNdn29RDxu5Ec5fsoxidfCT/CRVXkq7l+HxtucV
PZyM9Oy5q5KRtXoW0Gx7KvUjTxNYMQABN4j4KHaSn2mW46ldgSUu+FCVvRACiYpMGThlBW5oO7ok
YfLeFN1CoyNZiWcbUh1dkHwrM71uMF4oCzaBHb+Igs79wjRkKxDbD3uv8HpnyF7wkwTMQJ/jT6wW
8nCfVyciCCRYJ+a4kLXuCDjX66yzesePF8DyyWgX/fLUxTgSujKqKuayE1agxaA5f23bb2wlhb7F
m1IXpBwlFjQVnCZuydwMaVLEoqtEMxIBQpE3MGNZP/qYOIKUSIAJrqejCGf0M/ZNEr4koouJMjq3
+GoyFcUiegZ+TkTaFGBcaYOExczgYM6ZjL37/TLeNeypvcZfI+QzRLdnIGetOT0j4Wm0tTsIkt9D
m9Zw7O0DW7fH5r7pQaAFkAvfv6Ueqv0drAKCxGaz9MUCj/K2MAhAGkjex+XzdPAVE9hiXfyOMyx7
urXlMTG8ip6GZ6T/V2grGf/SmZg3gCkUWA+EC2+6xgHCZ08CmPuj0/bvaQiQsMrm+pHapD95nKr/
EyZoXpPZEO6AZM0bmkjHqdGb/otSqr4nIN1iHfLd7YEBc5s0CqOyMCbT9Xh1Og4Sw6GmFnH0yNiE
vxk7dqGb0ZGvkAJ9bY0j+Cae3WKOlwQpabfeKUZcAK1lttsKfKZSxrpREiO+Me6x5CpQ6WFiFmpN
O6p7+g3c4gfuV4VRAlIAqor5NQDFDBkUOGKF8uCLU8k25tMjxq6z7i51cAd+6zvq217nOT3Zi72F
TP9whR3jqf+1r9rr+JIc/SBOlZyGrnwsgxPFrGPf+v+6xNqA5ExGQvIWfs8nuFPBR/fiXfk9dvhI
YsIqjErNdx/xKliHGoLoMgsLsuTyWyqB4oo+bjVZG8gnKiIHBPUg08afSEOTDyhLwBPZ0VW29pPi
xQB7GKlam/0KgyYVRwvizfqB2rVJZpG1LsFFKooGoJhvrAdiEeLTHQbH35AUzq6qpWXpFCU2BRS5
FZ9xjGUHVlaR3rVJELqXB7Jga06GB58jh84LqkbO9XG+jGJlFRhBGoGpFe04Egclw+v0y0uVjUtp
7GQDEDGoaVfGVIzbKmQQTlxqUeaM0glZwJJ9BWxHGHKPG3OqW/jZvu/f5LGL2zG50zKKsRyrJaaB
k3+o+b7xQbKU8h7zG2VsgRfz7irc7UZSgT57hG9gbbQF/4hcUUSG3B5oxH2hEwp7FUFd+tA951WB
LKwBKHMzGx0woHh5LBtX9YOAlfI6O6RGTRjK7Izt8rZKaXlul4maFZf2ebhKpVn2QkJSf0Y9oNzo
4YwIdn6OUuSXfwB6FwLFd4j+8Fi6WT5n2KRU1CEUdGEOGzwwmZZwFvWGwM525MPWH6Ka/+luAFY8
uTrTCIsjiMoj2tuTAG8VyqSm8py7l1Vd+BVdhHJ00VRBZuRqqK/PObtxsk+TTHu4hXeDQELmCxDw
MrU1hLmkJG5FZdxtzLOSCoJxeMWRZ0qy7hgvmFOEEqizWQSIX0xA7LIyDQ4iex9vWkTFh8+ZbaPz
/cN3k42o56BtAHBpuSqyNgCs7GVXAbf3Jrl5CRg/OVhfK7XCCrm68ppG0Qq1cJCMHU7d4Uut9Bqd
MNjDRWcb5kau9vNReIzznwJHOsLdMaHe3+KJEXOMJSy3CvvXFddv1DlY2RBCWhJ4/IHAruKU5MNu
fOzP17P8nDRU7BzoEmPsnc0fNAkzLHPJW6G2/r0vyXd+I/GachL/EYmEbr4W1pH+YvH35JsKAP/S
obiwxbv6tAqnVQKKW8if8avBQOCFimJhFf0lO60qe7Q6NF/rMwjItDw3y+E5LGbinwRPcMvuG4HY
rLWyLp3y9+nkiTsEdE+vIkSnS2pMDZGs2VQw+jyhayfRBffLz0Wk9NSUh7ok2Pe5qpc1NRnuSl8i
hTpu8M2HYD/vj05n2QdJwW58Ealnm0iHkDZoGH6iko8fuxu8lsD9xZ3wkaOMVKkMr9t6kuA2dWA7
uvHs0BZBAi2gM+mG7GMcConLU5BK91sy3sBdrFk4S1JZbz/lJva4+Ei4LpP8KPm79TptyxdJsnL+
XfLmtciDur0eGYm2q30tfDQZmpcF1gSLyDxWgitPxF5LIhCNIBudtjHD+all7C3N/YrZnOheRz/w
GEzxm5suTuE3Z27pULTYuytBkBKWWQTqQzuN+p1RaltUH6goJR6vNVZq0FB3X/0yb9cYGBzRtE2K
rz8ujG5DUrTLzPynIHuZatW0L8+GiNf1EdKjLik71AwDrFWwUsyRLUt5wuLgaDOD9rMlwaraCLUj
EpIHyQ1Ahy+Nd+AI1eziLsJYD09eXBKNT5NX8V260vUBs4TsD1CJ9xEzrP70TsQ9og/NgasfhcZH
BSL8w4kX8EWo/4jdQhv3/O2+bfeCZQHgtgya2M/joWFvq4unEfGC/8i3YjB7rLhg/IqOUkcOqZd7
H0tRPORzCAuf68APOyl/MiY6X4eSHzYn/8r1WTv7GGYtOJXYZiz3601zNBi7K5zyXijFD3IAza0Q
75Uz4dFvsPxSxdIEPtppPUoO5JqNacz4CcNozgCotBajBhcVxglCqeMl0Sbk/mMvqDWB0LoxEI9v
/ueEeIQRC/I8/PKToXbr2tjrd2T+3FjeBNIuUJiTQYnJW6fXH0nOnOu0oafRKgXU2IMzaNcqGMLl
G/IZ3wTr1UB1TUIA/WQchbQlLKsRt+2mEKU91Manct7xPBpUheikpMT2uxsjlpt1Irl9Iu4Lep/Q
GVNF31yBg/gO+GJcU1Cw18Y0Veejt/eiOebEU4pm7Z+qmMyEZSpiGgfVhMqkj+JzFlBqn/Uxq4nx
ORUMbQHPt/bhx1S8+OPA5/ziUQNQspsN8rE/DTIXRYZEDQgftVnEefyFbrxt0Wd51oE3d40RZ+Qe
o1bhm/GyP4R5Yya6vNrB+MpWHY5h0vzLRhWAufGCU8aofI8B6s79rfaxJ2KY4io8zT9WMpJIF4ze
5J3eKF11XwQXGNPCCfBepv8nZ36Py9hNCr1kS8HNukTd4k1beL6BQy2LIuBw7Z/GevyENHZCz6M2
Ef0fwYJ4d2XXrHHAswNcVHGzqqOJnXc/vxPEL1+JTXXbf/5mJUBnS9J1HvaKLgNsliJvW++DGuXg
eEOSOUekdLqhh59DMtpt9jI2PtuI+RM6iP8UQoXW5XfbDPwfN4KOPjCg3TtVkJIM1R+25sKcIW2I
8YAoDS+PEC3n5FtSWnjatWALjBgFC9rphkmWOEh7y2LXyTxeD7tz4CjhCOvAvy5u7yYegTkrBfBm
UA/5GYMBWuCA7ssbwIAzKlOActfFxhQgPwrqbir3KhESTZ/ScqlVeuLEg3oeED4W/3IVuDcI0X5q
RBsXvRM+UsgHiEyFW9iyb4KMd/GFLqhOE1+UvUrSShZDLtSnQPBz0GVsY9P2TxGUTVPHBF8+31qK
XBRmGWZ9tP2dW42Fifa7JXE8dnJJoNms1PNaEgg880flB/dKKa7wqjGcKYva9lWVunMjYJX6lCw5
XqNY3hdXVP1luDLL8jEc3KgWka+aeSAUe85JalDDXZOALaFn2rR/YwAff4TxUd2HYbi14zKZ+PTz
WvzTh8u3Byv+tRiZiVdnzPz7XYh8z0uC5sPiOy2IXa5nNw9OZwkVfog3BhU/mHbb+okCVDf0cmhQ
OU2iRYyUgdmZjg/8TM/LjswN+qJ8Lz65WnuMify9d8UnYL764ukh0/HN3wPBSgKwVjzs40Fqa+4F
laTnq5lhdQV1lQb4ua7SW6k/4aCLNgHNrnHYeOREJmnR1qUUumJu72bu9AO/9vdZGjLtCvOdBC8v
Ery049VTUBdrBSEwk6gyblWnhEq1wmZl75erzzNd4UaykUcqFC18zw14ii1yniEm4eGj2z/BwZUD
VquYZzIb0h6oCbkVx7alfQDbErRwhEQr335+T0SxJhgIN0BUPGnX3fNqGoqKgwDSG3XTKexHea8d
/J74zFMmhANB82Mj64DAvsLY+x7ro6J1R2xMO3Q/tRvwPvvotguDdjnMyIuEjid4JImHuRkMZPEK
nK9F1LTn6DFbjcb19A1doB5rBV+6Ha1ywYUbQP3N5CA7o0tqfAJ24ckbOhO29CwvEdojV2VkOI0f
d1T/leHt9n41y8tFFTNT7UPSgo/jxvwlRigTvLhjL4W1nw223fu4D4lfxQp9v7C4IN+ihFoLg6Q0
gfOfZl24cAUPz8U7QapLcXwzPROC9S6n/B28RtwDypOquhxzq+1DLoHRitsbM9Edl0hOGwDdeZ6H
E//5gd9UFjBlJhftmGf7sCqCu4hMdb0MkmqAFJK5kLJRLmAWbmxFJC8ibe22qzUM8lFoTUESqFx6
qm/9vxhJl/pkjAarrpBwL4xXLycW6U2rPWKThzH4QUXiGbrBhc66Sgfp+ctEHCAhZSSqjoJQG2Bm
lXjVSpBC+bpfNOvOXR8yUJS1ICDoFCyUY38JZ23G/x5aS2FaUPrEfNIHPSFWlcV9Z92GTgK/kRXQ
+G2FhGlfm+kl1W+2Pqq1MSMpJAvD/6naiMERhr1GrdNJR36NJxtFDNKqRevqZ7d0gqQcCxjIfPgb
zOnyvz930dgd8jL21+n2sJbZYxp2/uS+a5wOZWS2hozV3Es8vrVgSkprfyFeCe33aXEC7cys8j3X
VqWFJkDY2JigD8/v5KKdevmn2/yuHphfLn3goUgz1WLbIVDgAbAdpxmUP//t4a+zdHf1zlqagiit
KsJDeX2XRQc1RfN0uWnHR3kT2z1gwdxVVAkjq2gZliqmy7f+QSlKX2ufb+zYS+4N4kXmmFWNZw+n
jOvQ0/b3LOgyCKc5ZXw+QZ6lZRti2SjS1QyWqLkw6NZv5SeRord5sKGCD8xvs92Z6lSzZcA7iM3R
VyHxaClTkLFF3e3wIsJe0Cy7maYX6cv6fg9OM0ad+mHMiUxsQnQbdq9jlj0nFj++JYBuTkHaeimp
4osYYe8PFNyBI9HerVPLejmPVk3548aTmtOLNbSk49vRcX0+ERzJ1pP/qoSSfK5r8tWHxryX32JL
FLl8LeY/ro77PvO8uenPTftFpTjzvioRyYNSYEso/IYcavgu71T1pskvSimlRBio0sPtBE8MVKI9
zCjgzUmAj5kRcyms4iwqGXIiM+eET+lNGv/zDLJ4ETPCqaMXAV6nOcixLFKayDwFUVWTEX6j3Ir7
uKWnERDBd6qcrtvoeDiXkA7wCmnUzpkXVo4NL1dJlHs/gt+rYPhr952TRTdEy6emhHTUZq3iYI1U
zv/EJSXvhnvkbi8RSEJOTDNYTQj2OgmsQnpo4rj/tm/NXaj7UgzHT/PPRNnScGCXVUtwa8zZ2WjB
epU7gtjm00YkFX2nyMGf7ssr2jC37eB/SjupHkRNqHwgIClofCl9nEjOoKPDYOnlewuOfWAa5NjY
ilcOpP4/6zPWajSSUe49G2JR6HiXB3A7+1EPxfGwnlbrnSxE2LS109d6df1+vXQTMVOZjUrhT2Wd
snhq9TZIgHQ2nz7sPYx1xemF+I7m1HdCtvI1vhjf475OX6MB+g/bJu1PyxMdqp9B+xwzEFr7PsuN
v/74rzEXT0UMyLqj6T4uzbZ+6BYglbclfoNzvPZ4GzeOxczoV+Qm7bkUqaU5OfSaAptKGS1WHXJy
otBEtuR242nkXXqDEXA4GsSR6ptNquiwSSCFIzrNoIbVUrtjxVBkgVUeYl74+DlnnOQx91WmJqpS
nmTevy44kSZs0G+5ad6QeZmWDiHOqBOIR7+oOJ3oyERlQm7JOWL0znGBeF3k6+TaTVsBChe9mfO6
/JmsgM3Q06PyXn2bITuXjzH9dSxAkZjEyMsDIA9xfowl58/rnRLlHKW+YSFsHJvKeNWz+O7WYvc1
Rt2hqbPeRH1a1BIwv0yxKqzdUI7KHUprXWLf2Xjg1uE+3r16iScBqHouGGxEJBBIygw+Fx8S6/TC
3yElu1nUarQUBcuHsF2VsYOzE94WcHd9+ZpXDy+KHx26ZJTmWowjdJLwMo145/aieIPfrJLHb7/2
ZgOrBH39oAK0qYwBSgxRpzgGiRmv1y/bYcTs1pl7f9e+rE9axWiVn90OzSd3HCiqo6YmBy8mKvS+
dr+kBnGR0umUqJZhgnl8fXKu422e3k96mwmqt1ANSB3LUQvzXOT+OOxAbnRSQD98U7IrBeGs/i6E
AQlbHk2A/ojvCxBszkJOeT0pWIZVgZ5KW189ZK56JGPBKQDYfafnYeroq9fbcyYy+xnI0iN/QSor
Yl1AeVu5w9febWQiayw6csY2bqA0OB8Li5FfeIIO9AynlWPqpPLN/s0FKpQFPUW04TWk4Re+J+wl
BV4JCfb96vY6LUlJliUOfoKRJJBSgEfk0gq4CvubDWKDFVPiEvxqShYT6eBmnpYSNrb4dBhzaJHA
OGdlkHt1tQ7U20EFjXL4jiiT98D1T3jTS/in+h4CUwW0uEyBNcXbfbt4SPnDbaG6Pnw69DcXZLFp
80prXn2WG7kFPM57lNZLpi/IbOTOskwja0AMEuiR2McJIRgtKOZQv43gMzzAmWsoGFYnus8tMC/p
fcJRuJZIrp+5UJ/2QMIwPDwbPbmzouXaJanZ8Q2huyTOJULDk2huxgr2G9TtmBJOmPZ0K+/yf1rP
r1AiVb9DbQMUX7oicPKFnRHU99l2AAeoZyLlnUp4eCXPcvySdGskTfDM9vJMDs3Co/bRf3Y4Po9J
KplVRxdqPU7DkSCZpUriDD8piwZD/tfJR5vMOWVFtAEM33+Q4sG9+HTGkxwpOjU9wXFIItAAHWlY
PiEghj7Ahr5DXORztAInQFAxNINfGD+EZQZ38tNL3G2Y3UDWO09/WCEoQDJg27sIoW5WpBUalN0e
8zGXkWcMNneWkpQOGYlBBDwoT5UFBeVCYdsAAKslEfBgkvPFqeBrmaJTAWBE4OdIws5Fc01dOgaN
poNoGabCTAyHCQJbr5EK9m5OvnO2XcasVzEf9gr+HJqh3Pdylz/Ur8si/b8/UrBcfrBRfuCh2HW9
rCUV0bka2h5vHydDFdih+OLXZUdPOggdDmcfyzZi5Q83wDLnnHdlwP5leGYU+bl3pAzsFRymMaFg
8glOBYT44zv6+e2+nBk2gAqASuz5ybn5UENERcAUCm9ps+S53dbS7IueKeedUN372R8PNM30/MBO
7wX8LqppO9xslAQG87pp7NzNqKgrBjUhuTi2MLDFZGJLavLgPFfsJtWJr6taQg87DnT2HUkyw8rf
urrjM90rRBAzPfJFWsimFREcfRJq90xiFVP7m46OX1+DhyLtzLSH2DrjxYwp6Hzvzyy/orZAobhx
Z15lnyFa3DM+Xzy02cVHS+F9f+TInYBpNjJ865b5pVsAqiQSl56eq7OMYtxvnj3Wrn1j3NEzoTNd
XgetYzrOCKHMub2xxhDFRIyNVPmszXYbzAImIt3g8tQgnZtBujN70d+SNc4QcStvdBLFwpmNA3cH
uDuXTIqfvBlWmr5wPBoJxDvhOLroA9j+jexKgEff7ch0yzU0bWRk+xlObb6bm3lVgSt04ikZQ4H3
q8ocperX7ALytF2DK5Js1NbINdi/Lyr3tCgeJDuD8Fqze6RyeOgBMCZafylJniG3km0qv2t2/olN
tls55ewJwNqvC61iJS9cgN6ola3AZJz37WvKwFh1NZVqWiIj+QqYX0KBfSgTQlq8ukME8rA0txEO
RbwB/H1SQyEb/K98MeVCYzQ2tQm+SphnHDsLXr0/g9bna90F1+j7A2SYRBv2zbpALMaFUnCuoMjL
g/V99cR4LGIKu9KnjLD994Q9exSbepky0BfiJqVLrTZ1ui4hcEpjClzHtT6BFCV2d1Iw+EP1NAhK
OlRa/GG7/NKUVTy2sZ3KHex0CsM8ydujabKkBrM4+oA9j2a0fHOfwP24hi3J4VYtaqyoEcY5vo9f
SuSXKJa7ks+SEyhKG58Cw5deoc8JnYWimRfS9b8p7j+A4U59jiV9NBLBolkc3Culj5a1H847nR7Q
5IxtrypaYYONH/SicrnMhQu8R1JjG/15BY7/oECf3NDi8Q9equuIGdgN11OJ2eDXUX/idaUADQM2
b9MQMCq1vvxS/Y+C5mkCscQtjIHGxq7h2Whz+PHNDAMjeJFlCfBW/cMGGpozmx24p7IeQNqgz6Sj
HQmOk9Wd3X8WpMbkd/cPfzQkMkJISLFQNPTe4+iLOmR9PKj+qRTYnmwvV3/ve0rU9uV6Mbpk8lqy
wL9z/gv24Djqc+l28oAwrNbQlh5ZpTFKqijZxoi5mrfepja9T/+AOxi9XhkV+71N7hvKaENmcpZT
gI4K53aPOhQtwjUyMLgIMuvJP4Uuyfz2x9QBjCe8fhqO6dSvXPv+VEYsrI5XRZliG/aOqxBp29Mw
0CcY+gWtlYj7aioKP236YQ5jgyDxl389sM8xBs2IyFIfS+wdMQvYB1IFJTYwRmw9T8uQYxwxhLma
vZHVB8iixlW6kBdWH+kbwaRN/gen+FgAsVy2MqHzdZBEWNucHVuipNKNAFaljrmY6gD9la51jgWD
AGNNaQEfTVR7SzRP5OZYzZ/8k2+DHWxlPdg6LgCZYQmWj3h65XQ6uynAJRE8Vef/FVr5ZpzIG8yJ
iUbbAotB+1GGmmAkElc1nYgYOFrz8DEXYRtKDHTt9m0SHsxWO9J2kDD5XDmOfisIxL1Pyh5MRKfI
4X1lZsOBlwakWe9qaqOjQD59stBd0CfM5OJxqcR2OY8+7MPO8PSbVzUmUcy6SG+XOen7kZf4fPxY
yeinj6gMPf8/CzE3hkSy3ZVrS1aSqVtZCHySXaAzVQGBscXxa4h+hjij6fN+lLa43iMoxeDl+co6
OFnLh6A3HTtJFN+qeECGcwDhqOF1Y1rrb1dFMf1vTVj/OdmkUgDONE41qSd2ejAYSTxod7AwzIxQ
ymdf93RTbqSkSC9dYaxTf10+QqccMAYFOWEGzVinDNWTe9cIrltH/68E0Z0QiqcMannnBqnzFTfP
ol+D/rETrsUZX+p3IR4P3dp4mSVzuGb9xvldcjXTENV4CjcFz8zRHVx/czh84Ps6N1YhbQR47T/1
vuPgzz/Uy0/Q3JIiB4QFoxuAEDcCrk/mfx5P0rrVE7oGBegDRE/LaeLTPz9i64fNUP13thtmkM7m
V8l/fOJ7MLaz/q8XXmIn8TTTGSbcrAlJAFJfTnMpw8eV/P7S/8AZOiwiDnJ5r4b2Sw/rfGiuKMH3
thhXfrb0963VekvR4iNUI8bRxn+GPZycIdW9IwPtSNq5T3sjChNsYDkGGoN97rn86ccwF0KIn3ux
jLbBBaR7iC9dyE1fS9VdBuTU7Ju6lJuNyVdFQgi8d5++kED5j7CQVUHdkFj2ezG0gkk93ES6Ek5S
bX2kqePoG0QBSTzC2HcmcaBRew7T5pgB2c8drWmbVWtFxRb5dOHn1qA57Avp5wobfbMWN/IYmjLV
CqEyRxtDV3YnOXZYMApng8IoOYxnqrfxQiqIMimvtgfJL17NSNZDnNNQys5IXJ3oDdkfFXi4K4WZ
bjt+ZnjE+Tjsq/Ns7b2okNsreWWWf4/DnV72j6/qlNVvc10XygWDaVCEDZ+3+vapwxbRnKArwkPd
a3bYmcx/9pF/BdJiIRi+gBiNiCw5rRGuQiSVjNEpPHjxSsMS8EWcn0n6ahP8pTIFsh/UpodgVYos
L3YNLIT8f3uXyXW4JgRP6ud3fp9rsQ2u/IzMqNYcD3J3xJuXK4JczidfnAKWBjcOQnh8rpqtacPJ
77rSLTASeUal31wsGfKQw7SxS6LodoY/glCMoMfudjOu+yehCwrfAtkCz/B/o1Jd0cmOT6oe2Rc9
JXK/5Uu3cHZTYgeXfZcZ6wHTPGWqteqEkt5/tB/nR7ZzPV7hpgMsiF1FaFTdrqv1Jiy2iwMo88q8
wPYV0keciTkuBKNwoYLKpXq/ZG/eoUj17Ti5KQqudlCEL2HmMIDu4fy1VFcv63EStpOATbM2Hs0t
wbvgMxlw6e1HLZ/UMD7Odl2qqFfpX1KU60vPnAZy1bJIOu3jbNhM/XBLydqszsswLcmAprXeTMsw
0T7hqEjsrwIqmCF9DPdtFW+PK6BUjde6WrhFaos91y863C9XGZ8/Dr7SwYIFIMCyKK5hq5k2+VIU
hE/ch78iztlLBxSmVa6Qq8oj3yQgk486vJ5p4bF/oQez4NfiJsyA6kQgh0CyWres1mF69tm7UTXC
qT1hbp9W8lYuyTJjTS/S+cEllXUES3OSnpheVD/YkYJnLJ1NkHQEgdwFZOONVyF7JHHCi0Xn1jBp
vPTETWnuPg8B4/Pq7/eJpFj6Jdnr71Xuz6zibyAc+4nFl1u4+/qkvr/4G1C7LNZWaXyS8InfGlOn
Ur7dUgtqgEwynS7jxrMvxo/i2xp0nJl8OgqPO/9UP/KfhxyrnNpgaSKMCpHWUJYN03hVRRkpbU83
scu01cgllXztkvIbZXc/Gge5W4NdvnQBaYHy0VM7YGFju0N0TrDMx21nSlOJmobcxNF+ETmkU3N7
fYxLEbQ7Ymc77EMWc+9XqQAGme0uayvp0FlI0x9akfA3683dpOfUL9v953X2FRzrNBepNrrWpKCi
kZdWl+ZD8boYWS/4RSSM+dPyXbKMMOIs7En+/TiSf719hkwI/bmmG14s75DK+opXmeS9GW+5meRc
3aZmkgVUQLitN7VjED1VvyakY9HYKRD0rrrWInBwXJdYKWjUQY7Frcae7TtS89sk5NiNDGdcA44U
cGiiy0dTJWAetAHIHKdFXjMmZQDlK/T+ZMO/w7DEqDzizKZPnQk3Vpqb6OwdsXeuOkEXK54C+EW9
j7a0YLrEHkzMsawyDiXueiU007CSWbXguO1tvKvgcRKnuWvZL5MZtbjmBr0/zrmE8gZkMha71Dgx
ouSYF6f2PxIw0046Xdb13I6vVBAbV/RPxy4oJmPnV5lk5T/ilQfGnOMGZLfnD+Nt5VSXwT/UQGCb
y0RXSGSG2TuLqaSc3r3XyIZO8hAEsyvi7IuN+37F2ioNac3nMHup+39/ui8ooaOOyvWlonN3MA2V
CvyHEdttp2CkOvyjny9bntpVHN+h0u8PEtWnE8volmcLVszZ6a73659uCLI/To4UCJasp9TDihKX
K18sHhknOdEjZJLKj5ebSHV08JxTm9uh1NELtfHbCZeliErYC7CQraRyF86z/7TDL4L7fmwlw/dC
D+jJVZmLmZX8GK58AWe4Lxpcer7vknCfdpuXVgmuIdVN5MySBJcYThgbUItv1WYMBDpS4+wOahWm
aV+zO9GjdoGWDhtlakWwxXQ0sbb2pUFg1J1zTjp3QgQgLx6e+QInXM9R29Vr8pWI8H1crcWyn323
y0PtsqR4QOwSYCMo666kgWtmW+MC9wpuNWoVldGS09yUVRP9V438l01ttX2Bjkb+b5fzW+eb1Yg5
NVk18Gqo6jFo5c4vQiQF/QWL94xaLmLkV5Pod6U9PAN+H1imuKltVYADnQNp58uIz8movS15bPRC
86VQvthgm8Ba6qYWt6come8t08dEBevtcAE+PXgtBBvru0vgyftjZXUYXrrXCBrNj2SwYnc8Nvy+
toYrK+dLE8gfdeJ7xm3uICJNRYK4RMQlYx5WC1dR+eaYLOHgrs0SEdY4b5/+PUDnfhwKbLFkaWsC
Ic76hZTpT200OlY8C7V0t6h/l7IoPn+YVpRVh6HBKZX8WdvudwdYHZhxKljfzsOYo1kHPvpKsNKY
A3Y9rKVdRq2V2IHOcV4dLKHj1fuG5SIFIbBqoMqWO8gsYR+epliGwHoOM8FYYLEfLWd+1RrR5ifd
BdWvBHeiJfn6fHnZLbEC6fmn4j/AjaTuLeEFnnLT/GaHegIUJox42WnjkBP2fBRAqNDeYd6APr3G
SpNXQ96idxw893w7YetAklqx7GKcRERTH/oHSlicXTA5gh+jxA+OdVln3bhGLfTVJVqvrnSspcoY
gIy/0War34dHuUyrjan5Xbw0jVUi+tGKZlQ2ZKs7SQnDyfQBEQe3dKLKUrZhhvzgPsGV/2UOay1V
eY1DsdfHHu37pvzRL3MJKq+OzkvmUQYCj1Q8gPKajr78f3DiiIGIgeHbTESxDP+d//dTtHAiOOuo
AE8C9QzMl5zym6BecabLxFNC6//zPICGngd48KjwZ4gx6dnZVhKLs+KNRu6SV5qBZCMcwUN7llQ2
CV7simjmCzZeJy+ADoiWWneWcwPP8Lsc73RLyC+kbf1HAJxcna3Z2zdyi8clGOujnVOztX95IJpv
+//t9TPknyvvbhFjhskdAhDpXzNQyonUxCGa2LCvLA05xmDfGORqqcdeOAUS/wAt7AwSwbv1X1As
NAM8rluJR2X95Kt3JsAo5LeO0n1TnJkzqsBEZFJGM3hFxFkp+VTp2fUu5mul+87JzdeixHAn+0Gp
z+qOHeJRolVTZhKBrHTyBgsGeWZKbSw7pfZ3IuOoPi1xg9etZ1S8GiCupnBHv1AAdum6TOZ1j3ep
vp3xneeUmjEWnzHAiRjDNRJ1sRMkm1O7+SrCu2AzqHSlEhy81VibAusciMK0q9RlcW1fy/gc7v8A
VkHsIFky5AkoQqUGbkGfN4fWkfACrrLp6LwPHuUeCgBE8cg0ck6lRW/BkCvAqy/v2Vh1vclpLWzi
MsUMR/CCpjtooTNXJccYTJ6V0t3enWZrTPFsV31kcfTwQz+3M75HyN0NFYuwmSvBJFOyAphIDdhN
Ji8+Sl+n/4wZa6RmBMUgaWOXYWNo2PjslRj/2h1oyBtJOKC9GnUlNuX5H/qEyRAE4m7mJfAbdOea
ziHp4PuLZyX9ZNsrxeI1CRYK+/ArG83JhdHV8m9IdvAZuFddM1/6U5dvPSoo9TGPMSaDUL/Gy35H
QD4CRH7sxjHzzOUViHKCbarGysdQp2PnKh6aqzU40kAxRd1ecWb/+N8XY7Zjc8Sy3ekI/rwhRvCC
7aVho40IeYeH/dYeozjlTLKx/WzVxdSVSh5FYUIK4oyM4VnehdaIbZd6GSk+zsfOdc1x8Ktygnz+
hmiUWBuU4Pc6dnFqgRovZoWgA1dtb10FcHWtiAe7TuV9NvmQaPfj+TT0jcPPTqu5WCPnDzBNMWia
AdiW+2nm0iC2Cqybx7c80yOflc2qNttCp1mKS3gYYnT1bahV8cs8wzGFvxCXKzGyj9mMg3C9rKdn
hGuot2QezC5L79W2jNInzdA0lHDb1ALybo0bsF5TMsR3G27GYpzZdBBUgKuVLN9PArfIq/lrtwSl
F2M0HTahZWufxrzEjehGoW94JiJgtB2ipGfkritqv2EeUK/P4+GjhsujWNWyZxSccNkS77z6PzEz
sVQtjVOMNb0VKUFS56r1yyTHUNDfAJQjDK9utvM55hA23NbDYZkLo3naa9JRgUL025QEh5UhBC5R
DGVGIxUplp4gWHNlCGChVQSUQ5ux5aWsdSksRzFgQQCu0Ak4+P5h5MpgtViSnkG28XWeVv0hF+iY
3bJgdBhyrJoP3RUQHjd723973aFSqMp+ZBYCwljlBpBlqr8XpCnWIh2JieRmnmNWHiY0hJoyRrNj
NiJDbnXSREn8BtQOT440KPk35E3E50vXWag376+VtJK5yVpb6HD3JaSEgBw8sObVA4SfwqX28NWx
8X/8Sr+M0hdoCJRJz3XEF19Lmm3AwwJ8hAQWrKWN2iTJG4ZRfiHrkl4RGgXeBoeP+Y9UGCZG19St
xBJ26Qet5nr16Xyo82aMHVnnY/oUHXJpIAJa7txcOGAnwy7AdpPjkO1OhIrIZgosHR6T7m4gdfRc
gspesQrReiSyhdIXbVSAucmS0l1W/HXYAgMnqEN1m/X+IL1trX0J96Xv861+Zw57EsAk5U3RXP9L
3ttppykWIUK9JmJqHJBduhKDZJIG19/KStGAWwte3BQZfXPBx7W8Ufl5dghG/B3ll0eUkTIjvdC1
VIoNVrQnJ5cCPyLx4C/fr9jH/VA/Hw2N2kJ7Ty/pYttv1Qg2c45rla7qlweSHOFC30/ny7SvWmHX
zFcI2sChNzrxsueHGY+1r1iLfF4iZvN3F8c0acqNUHjaJOyWPVQf9E7r4RnnIolczIZBI3AOMlnH
q0HPxwbTsBwrNqazrHlx7l0RNw7m5FYEA/55Nk+THgfHGd6ge4fABRjT5/WwzQ7nYKbpi/0sb/1f
4FtiHz5l6oEltCvNVnDeegAKu4EN7f55/CCprZ/8qf//avEcAJcCEuIBNmGzXlHKQZttmNPDN3yj
8ZwKtgUlBaKKW+kDz1MhURoOW47o+8j7un0hLdu9lWHWBDrdyNDJuD11ItMM6FKFm1/883iQ7Qor
YwzjNEDcy10gViK7igUXETTKcbolC/Ogr9sgzGI1gOGQpfNrTU8h2VoCIZJMsKifrmw7JeOcdPUx
07oIl2WKj8AyC0dC76p1AOxlAegitMR63AQl8i7Fchux4f9YYZpJtxgr5QV5jWZeC5d9rM63/dbh
e8paxmbWYhB3aIvf8tnQz6Wf+nSnc1vbuEYjja3Fn3KccBH5RzmSmE3rYtASPNRT4EqaaMeU0K1P
H1QFHilOMuCi25k2FHH0h+UYeKK4NLy+r95Dx9ciGxWV5uUxmo1inqHNE04wXbzHeInrLogHNIxG
HwlCB4cnOKf1U58/yKGIUmUhHB+1Jds5/kwX3MZLVbeUTDLvVr8cKoMiG8tpbXIMKZFlZhH9g8rM
nMgdNJzqsQqIQGsS8Cbtq9pR9QIuRxQblsQ0btr5B5Vwd8hmwl4S5td66uwKUEjJW5krAnp+kem5
MFk085KVlkPlnUBum2xRQrMcR+T2n7c94AiGQZ8AjlX4dmY8D5OyIicN9K/LMRJlSiU7C8EY5vlH
RgdJD3viHPm2fhIBcqdz1++EAztUQlaP6nyzb14vsNW+RAFY4yIvyZqamcxXp9etuxcxNiqtM0K5
tnINacoxXw981cUtYN2huAMJwHgiooJ3Jan3WV3oZj/yqqIqrWSnXhkCxFopHg7xZkl5Ggb53DxO
ylvTTY9QduEMb/a6MhxoeITVPp2xHPLfOvqjbQr9gZ5/g4qONIBK9OYA9fiBMwNdpSQgc/kgZO3Z
XKgaZVr6K/AZ1zHFa8lR9g/ryegkUJhwYtsipAaqenrqf/G5FrW4TS88CDF7Yvdm0Ux4M+2rFeXF
GnlkUVrXidXvXoojxW6XBrDIRGYovNIVJEXpWwZHp5dsG7htq8ezGyytfGtL4/13PoLK4R5mpjqf
mm6XTGtYhTJCZuOSgv+NajHfk/b9QA96wx230OWagoOJIbgw8VgZ0Koyc4+RqNbU0JXDq1qV3ovh
opXWl4bRnSWyD3/JjprqKAdySvD5ClpqyjwUm48uuFk5YbdQNCFmzY3rhkU151oRJDAwR39kwa+m
rQivzPIhKdB0kKO1gLvmNd16gi0sk78VvUzZkcCz6KzveODAGkPZhrI0Q0N4fc7qk7Gl9Cp5ZEtT
cig/AtmScP+lfNJilRBdsbu9CHaGfSQNM78XWWFmTgdUG7ixIvdtNFqRJkk68B/Lb44afgTdaDua
egLW5z9+LWK6oP0iDBKKERnhsn4FeBlNOvWSOu6/pHFtQoZ5XGB2gneqFr30defwzJLLn8BA1xel
SpwvjP+q9uYn9HXLHnY2NC4Ms5++LIEt+XpqKoF6jIm27IK1/zFne0OUcgVxGXug/qeuBGmUeNbU
mMnTn8Dww13aP7AgHEdnc0Ra4A/YoMCFiXRsdPl6YT1k8PXkGbsFK6IaMSEIiOhtWImDUVD0BZEB
c0Ced5g/IzZgZmKJT2xZmY+JG5ansgNUWIyIbUE8rBj/QDOazv4St1ha0eiWIGId8uS9kS3ray2o
kNLeHtieUQ2ojMWf7mECeKkn5RjWRF7ZPH9UcwTMXWxqGoFbq9bS36/5J9SrWexYxDn5BDzfm6np
GkGpaRUSm0LsNZf9pDBjFRQSyRx1wCD+l/vuTCOxOcwRffcZRImk2HCtDO69ETYs9XyNwnHi5wxm
FBmQDSeLOkFwBh534qkxL0UlMhLGg63l3APC+Dalksn2e3Eshad1NRzZnCYW3u0dre/CrON9VGW5
JoTTt730tN09wRp40TYnvTaN2pccyTQJf+X8tsJ75iaxcgiiqhI6hNf2wa8RwZVZqAGI7C3QMcV/
D8VOt1+pLzTokt1jCQkvKco0zeKJ4yKx162Feycc/+Q4EGBIjA+JdX3kjqY1Y9Dvvz8lmjcKcGFH
qO/XBtNy5nTltpN8rfa+AUYhyJRLPCYI6u9AUpi4jIFIwJvbfA3tnYZJ3bTk9X9qTRexIJCagCFj
eKgkEulf924YsyHWDddV3XpgVNIKfrVWAKqu7h8hXUT2KM7Ki2CjlKE6I7OK13fJer5sC1VM4cYk
2e1dO7HRDR33YR3dJmYE2OKLnnAhj8tA3A6QlcM5vEw9I0d6/55S7IpkdNp7cr3qLdN0UnVjEBda
DYQ7/YghkinJZ6SYr/UlZUDvkcuu/wIJ134Kfwp7icu7W7eZak00OoZ2bCxc1coHcjj8r015JzNA
gwYW44AKmg/76x6ahMf9uHIUpVzexHSJT6LPnpeC+DDO0nSgberJgfJJ0vo8B9HjdmkUPTuBZGyG
LPD2GlrYNV64594OdW+m9ibGiH2J1Nf+xlHcSGo0EbklN5RIPjTBAQCI3SzhIZ7x+shq792tiwos
TCmja/MiJx8q3tZh9LVUoLeZRUH8+tsoVpf1RppFo7M+PRr4ZYFkvmHmrpGwNSJSI1TpvyheH6XO
3NmoGnIpmNDT4SPPn+HMMPYII1hN12vK0VdOcNTL5xKlGlxn++GLSdXhwyD08cscb+ZaEoGU/r8Y
Bgl5oWTxojdAGqtBAXRmIq8mwfpUNX/qyi+RSqsGzi5GPD3ArDoMWJ0eVTrAPL4ppkkSwy82ERKC
uF1wvwT0957/PbTbuays0soyTWSLFhM5pfL2xtl+oXVmAcc5y1SSRqZXrOQUAakl8FmOA2O697cA
3H3GAieMt3AYEYiDJbbXWvvl82M5nPzHWvzFw4HK/2E+scYO5JfurQhax7S3fgFBV4MsKvHtUMNu
kzZqXgpaBhIYRKeioZMLh6olxl6p2MaDjUjyiVPEb1mq2q/4JEpSZVRNfzjnyLFJ8w4mVZGr+LnU
d0qs8IXlUFHKa/eA6/NLiQos0LJ7T0UawP9sXudvdC8mBrNttUHPoSHscKGqSEVwDe7Di2Fz8/U4
5T3J5Vkgw3ZUyUEc1N2WNv0oH7LQQ291+oGWoa83S/GfkYiOGgmaNyuNCI3yxelXHRNbBicwyDl4
xMenUbbw/TIRHMwXwWKFKgANonmQu6YOvwXpBa8Q8tIZPK4U1iwuxapqTMZecNWLVC+i1bNCYw/j
T2kPtT/2KsHlYvqh7ZPGfZgDQsGPnLiSMKCQe0g8ZZfquRskCC34imSCVOKJIfpQynKBnmaE6rS5
1tcJkmn7766pU53d+mpK6MRDQZGsJR9rl3z1NHqOg940PE2DewAbdm0+ar+k3y3O+P23sbq2pFXc
DZ7koyMxAHhzC179Wsbu4jbZ4gPWo+MZoLqVyyRVZPWht0IhUMmEaemgMqvDa/mnAiiIVZrVf/b+
umsVaXeZo06a06e0OWmFY5kG3UzmACGhBTVNTaUKSjKW0a3+HYlKcCrfROc8O7am4Vl1ZFhld31Q
BttbYAMC5WAnPuZs7NAEeVtp7J7YPU07nHj3NOXbOqEcDDsctMCpyvRotTZ3z3WyFB+NJm7r+NJM
posHNbmyzd9zhNY+92u2VAGHipVOntf9Pgtz7EI5o5H90f11lVJmXVWX1A9qpLCu6jzk2lFRzlPI
b8QfLAvM5cVL+HKe5J7xG3Dmxn16P3gAwamoyzCKRvTdxK3rDlwcB6WSLM0xPszDvkrrG1drhzBl
kfV28pxFr/+2uX4P5cbbx0/4mOOiMw+WwyJuELSvIB0S2RxHC5d9NusfTtjXEqJk8rHI37vGUCW2
h3vU8bgVq6aMc0s576Exwq3Yf6UAo0vZTq9kw/C5aLNTtOvPRaEnhSY+dIB2U/Qr1wyXssLmNRAF
yg7W27djEpwPdaunGbShs/foQINbSZiFwCrLci+gj0a8CiRTP82k/OyJQ/iWvPiq5ZwO//Wp2cz/
Ofw1xON7sWon7mRqwHDd9rJw5WMxr2NhmenPmhhGsjxDFx3aThAfSgmJZ73zQDlWBh1JeI12Q+n1
TcZEmDKT97uYupl+H6u+eEwh1ou6EJIdP9A4FljJhjm4y3GbXMFDm3t+9F1sxOY1wSA9/OZQf00g
Xqey91/o68TdKMJFm58wFWOm9Vef45NcQK5Jvb6AUK73M4MleZfsACaM25DJXXbTap5/ZSLxbxSD
xv68/PhqDJQPlowl+1iWaefoq9eW41cYCOjcxNi5GZSLbRwq4ouAnM1tI7xHt17IyhIOGHRGHSIJ
WEdiOpdao+cV2hNlFHdDTkTrXNqPTNxiufP6oE2Ew3HJ/DRex6bEk4jBZHjYNvld9oAI8+NIDlE5
jIpj47Wgjk594vEvjVStMBMcFL/Ya0lvn5SWKWr7D7tPoqJVpxVSYTq7XUgwEqvcE5NPEYENtfN4
/Vu8wihZjSFyz3otFEH/r6ces8Q7VzpLhIMSY46p6/yyKR8qH+eoa84xd5JSpn7sbCz4FOCCdZoc
6HEdcTa4ITl6wVXQJ925SK1zji9BqN/wwbsLImGnmPywUB/F8s1Z6cxpT3fkfo9XFXZKTvJkynas
pyqe68FtZTWef9tSzhLEjd6uQTZXbMibgr54lP+C6iZ/gUxDqjTpMLwLBDjf6pJwrE1s1F5eIWkM
ACw/AlBnCtau2gkWed1c+/EK8+jQBLYaKi8HLPSOppHVqrihwKQRpvG2LvRmgRQaaHo8eoGZGqnA
IB/llXyKUtQD9R8E22THbCiDY4fLn9OtEA86iuLxNTqbScL+Ol5TfBiia2wE+PocsdPwCTxmTTj8
PkSjlw42LRJWM+iWa4LPB/D94mF0SxubHYBC/QoGPoG+VebNUb+OlO1A1lPJ0Swpmt1wBihhXD4E
wJNoz5plMbC+oZ+tt0Pa103eVo2SH00a3SEXEY8xsgaPlExU3S9Umj917TENUu3rEgOb8DifzSH2
vZXPHFKh2sRi3rjvb1pbOuES8AbEm6WSoe2vhFOpBkHQo4AwXXh38UaC4J7lxQOLhS9Y5Ugx+XH1
wZeDn8gvB0ZFDZ+XRE+oE9rlrSKxX+StPvRGZ+oXd13TPGMblvaQFIhUD3rWA6UP7vSVqndn2o3V
gsKO9bSpMeex/V54WwMHmf52aHy0ijgHZ8necoYiQcNPlecYpidQFVfSbhOHwkDoKkiax6NjYPnk
QuP88VKMCbZTJAdnqQyCZyQC2564CmI36mu/8CAnxf+m67qsT3SJ+JY1jjM20/7Y+cTKqA7dtKfk
9Fn1bqoWE3uW65qkYgZ72r8Ao/GnHVAmXPc97VOEFb7cBuJcWP6A5AjhVb+Sg+6/paJseoVYh7ud
bJNMYoAshizkzH92r1dCPc3s/GapJ1B1fW+mibSSjOhQ68W0qKDT24st2wrbygGQj303DTys+eMs
dt571mtTjnWjTFd19wKrL2z1Nqm8RB5fPxPCATQMxVBvDe5ZI9Yn76rlQwseS40KjpcYuw0UCRZi
XSgJ9B0vYdRq8fyfdmBS4US4huMTCuknWjZeuLs/iLYWSBC4JJcQk2ntuN+ZUqIjBT06YOQ5yFl4
N6O2rqCA6t35OicwujLJj7Vw/ip4yjRZts/ieG+cwEJq5X+s3eROBjs3kbcmLjkkBkCNCFWWnGhi
1HVIYLuMzKFHuj7ExouzU82gVeWvGSN6qLgZ5JNuERmKZYW5tcsS66csK9Fz8ldYDqIffjDEjgam
rAJBJ397hqRV5ratIg6HnWeJsWLJwHkn6cFKlCM/R6HAz5C/vBUfXuJwJbeu/WdPek681HF0TAqO
M2wjiZNU1VEZQWhhKTCAcb6FTOSRkXiqFNvf7qwasjYDVBwD/0k7mzCr5c4BFAHpH2PI/Le03eTG
IlOnOdMAizOqFv5Lma7DqSomXChhNyF8ZFg0ept2Hl9jXzlbB5NqdPWactf3LfZMP4VETbbbQ1fy
rOJqkHQZyRe6EAyX10PZOtcqiIbyf8uCG5pcy0DDtKsXQpNUIwkWEZ2zhgVRQbiL+cxqT5ctGo4T
lK0VynCfOLF2lm+zt6d2W1M/WGaj/+MNpvXfl6EoF/qNFj2XiEPauyix/+YEk7yIRq15/0ncYdo8
eWIhcvVJhoVO/PIIEqbH2F1/fnKsxB58TmKnpOIxV7iR4dFmaMhPm3KhUjd2+6VJUQvmQMQSFCnT
BLQ7zdt7I3tqP31EenXdwBQWuki2zlTqAMcbsolm+6w1NLZsM89NxT5ndKbolpcB89yYJgmforin
cLCZLxndORth3+GbM/u/hTAWxZmL2ELKxDbRkMlhrk/LoesoKnMVdb28/f2ryltBC2UPUwm2judB
P3odQ3OHN8RkE/qSjBaV0p3AY79eulARct7Wev/ouZpEoZEKkT+G8yH3lebbCGIQo9bzTGIn/J14
9NOHZvaYaprjhkKx7Jv5pxkAj9bGfo5jKnQ+XLi7xP8kKXFPVDfSGblt1WwWyrtaFO6RhILgb9gW
lhQmzQoe38aiDi3rnLErZmusM5KM1c6UKGT0WLw+8UhdKi+8/Dhc5I+fqkrHJDiXhl0zrpqnZC25
v4c671loGT4q3UsaOkb6jfuQoYBm8IYddMR4//VxkZE/0gDHqRa5kjoYo/cinq5yYYKzz88CZT0y
DeJpoFUbpHtlOZ+M0M8pHBtOsJyDUrH+XxvhqG5Xy59srgMoDf6XC3GMj7JemyV+BQhim7Ym01yG
zYPoK2FrXDQcoRgyJMKWt65AL+COcycJVc5iM0PJabYZH26cMoOWwYMNSFNixfZDgIIcsc4mM+St
i9eA9ZYW7Sgl25KiM0T3yldf/sKue6lKxAndILBwQ+FGmkqHsSaxtbyHkhpMURES7ScJYWsQVEtO
SEGgUmMwIFW60VZwFAGNDU+lR8pgtkO3b85LBplB4rr7457Q0tc9jHZMAxbhkoHT0nQyOnzXw82A
rzzdBTY9+GKdtyAEdNhcnsK9+NPs4bhRWU8Mg8s9PvEUCRvxC9Es4XDgS7FOXuxtfdY/coil2SGD
PBQeFq8fHOKQLSe/jpL0QhWY973J/ukR1eTKmeOrAIGUKo2vx55I56bsA3ZeBfxDzFM+fz+OiC4j
mJq4QWDF/gCBcu+YuXp9zLNXcrT5JhfOQM6ID214u47ltPiKd09aOtkU4IU8hl+jJouNyVo4Uavq
tE5BquWASghHawk5piMrncLZ1hmUu2igyKVwsxaPD3MG9iVRKvajO4/sJ+YRRHW8T4/FzGty4Lwp
q8A+2HRs3FbYRq8xae9hENv6khY4rg++xHbSME2zFzn/49ge64VtsHXmcCxlC9z2M+fqKkzbDlTj
b/VHyEZepwMDIBC8pJRBt7BkIDGrIabt5cOaQhWn07lyKTtFs//75vF0fHK1ysW8iJa4JoiU+Sf+
IWuwcCrlisiU9lFqyOBFcVFzKcka9WTC2363taz/FeedxUOP6frxPL/4MS5d/hLf04/lBftgpHQO
OnnnZC6K/s1hihBVe3Sqw4MHJ4S4DXkB0corwnRGH7WRq24mh7MpKJWtQxOyI+gIWtgGHn2+D4d2
Omgf4M8VElmmtzFb9xG/+E5X/maVXGC1OqoKQklsVQQI3kcWakOmZXMdrc6TrGRUf+StmHLKqANq
WlrTmcwHWpLexu8bqaG4ZYSeP9dYy+w5y2S0FT2mQ5OARoyOLXfrI/bOSC3oISy82e6+AV1fE5dk
dS7fMBQPESuCSY01c52ZbQOETkeYY+IY3DxHTZFXWiF7pgYxLCdveb02A1Sni3M4oLpqhJYCn0gM
JekvIrgOfo2ao4tF1d0SbuKTSNVBsVObAdc0Rta4QPxtP+hkXjseExvD/OhcGNxFr0dKK3LEV8L4
LnrqMrBY8Ua4SmXK41Ra3zhDD88qhKoAy/tE24NxUnK3u/XI6GQZcOhZK2WRGN9CUrTSYGz2mCuL
zBVdpXzSKkiilgkTTqpEF4ArqfiQUDB/xWKBlt2gLC5RwBIzrce7XlV2mJYRxZXnYfunmwFgWjKf
/OZJRutYuG/seKD1PuJz34k4lGFbrScEsUXm6VSpR5hSfKVNeWx59DSLYkPCzhr/tXcOW03pgfRz
pVMx4yY6CPM8EvJlrj7ZXUenuM4WWvo7TMsWWYMd8y4dnwn1gxzTFMnzuY6jmej87IYX6wXUPxFy
DdUpxkinebTHSClcTJ6CwoeOXsc5MAQXWZS9ezY9QTcZlSN4OTjUH4fF8N/wJNScys2roo36R6Gx
9hODNg4wjAY/rUcdXB3SCCjXXs7P9zqkyYboCEFaXYmtd0joVxyIkgd/KY7M1QqqpR9YNXI423j2
dteo4pcZNbOpwv21buBS3KQ6f6ehAcvvNzKml582hGSR/A9IL8lGt0sSM+J+dEr8qrZ+dlKuZUkC
9UfhXuml5N//gnFiwpnplBJjNhneztmO8ME18qzhlpohz4gIdJ5cmr1NBIyC+2Epi4E0XWfXv/Ne
RtrUMgfgyxdPf99nkiJLSBx8zjRCUNgPdsSabvHbX5s9NeAgi+GoKXsU6EhXX8nk2+DMTrVg5jR5
zL6D0ZECHBmCLHnhlPbBh1upH+PdAXAATAc1xgJUDT3veKtyduLclMwlgc0/kq4/bo2ngc0KINUq
wuwzjfHiSIbfVDb7GRVfbMh2mDHaNKUFJMXvTaO1kv/7QWskZ69Sgas1hllZXaCWY/cOYwhFqJcO
B03GUuJhR4412yFY6dWZ3WR1KBoy4pQTvEiqJQI7kt4RIgtxWvywP2but9D6oEAQzfXVUPN4XWYg
ikt2pTK5/HfwGKRgg7QsZq/n2mkabOfaHzCRPc60lAo2G+N3QKR8cAFKD6a1aO7ZRSQ6GwjD4Efr
AAFJLSbUGZZ2GGJSJ1Hj5IVxEgp0OE/3KlhC1FHTTVtkf7444JGvnptnR3iPnfpEAXZ2AtlIZadF
OISjzoAjdrWwC1oyRnsT31wn6LOXSU2vaY9xEEcI2GzgT+hZm/q/Qt8nh/4oYZgA+D/K6iSYPJQ2
J+/r7VNdFPbbQkwwMNR1GGW1mukhVRLGbjE93Tp8rva86gLuq3UqEgUbak30yJUOVNaqijohtrLa
fsaGhgKuVEqajb0KwmRUteXltUFjW2C7L3OZ75K3xqMkIgsENBJGduaFS63TzaYzKQ5qqkTfPpA2
oRQxKt8QbshzFR4Ggxs4BBYFQxd1II5wqsNUItDnlmD9NQ0Tdszz61rjIL126EBGCl394yi8DWAa
l37ZxUWedIf7K1/wXF1OxH1UuHHD3jO2H0U2ieKqyWX7Xtf2ZbCjIuEVrYUltTemTtLAJV7zL9Yp
V+Fn2aXxugEdTuGjcfnCkKMufRZOaqQxQ7UI8O8LgtiVW7xsPXRhJeI7S1liyYy7OdEJpeYn011m
FUIJ2gd0cQN73+j+D96URNTQENOHkJPA/uWFTAOh45HbVS/9pl7R3vBmPOX63wpMS77+AbGvjsLJ
35tMQ7QOpyXIlgCH7KqSkNBlXruTSdiJDQ08Yn2oGQ8WPycNTR+l4FXdMTjoJOLv1bU2vImzs24m
O2PcF6U4WghC4/iedRRe7DOi6czfohnGjRrKBPTmgqe8hemUTS4RmLXbOeI5MrxM1KhXAmHDLdAx
ywBD+a9wyrsOCqT02dSUf0I8LzzU4Df9VtSvvV79TJFZ58TORaYI15Zi6qfP30FA+1s1aaH/b0A2
OID2T5kJASMj/ycg2GmxAc+rQXSlNhwT+b9fz+RJcPBtbKXUfnObo6XXh3rPY+/qV6J9DiBRhHi/
yAQfSiU/Pv3pmGa7SUyv2n9Ngt5l2YBjlpc6SOGQY4ApzCYJ9yUC6BeBguOrkIvnqFKPr624NSrF
efmO8NlsbwBoMwx3GBK5B/E1jYRQR8fGAguMNpm0nGS5JaTf/cWzdC3YW5OlzstNe0AiF+og9Ftu
dg2DClpZsywdSIflfH2LBPOBsYXkVXZ1CNcQZHeXQnwxB8ay9uOus7h5lBfdg/1OEXh9bSFZRqwG
PE7bVbXQd4nhPeKieNbmmmopUFIbYPzmURNXLUrqxuL0UV/Ch3lTO1SRUrq+xFp/FDZkNqKy8MyL
ZgSglz21X91MeVHOVV2+MxpW4VuicbHG21q1yVTIOU5Z6Q/FDbaLk82XTRDrRrBV4um10BaSspSd
9MYHuwFzqXOyRba0l2sLPoUMPUXrr2RPimHXcObgx6icO6h1kEmBHCAQhxY2IRDziI3rfbbjDWHW
cnrIbyQc312wSwgJf71RFiTjakwlf1dA6auaFe1nzsPbLBwoAfNOfPk6OnTGRW2l5VDu/tGbq11l
szurNbaVzRrf1JpL7Zq0NVfm0B6O5epjVaT6Wuc/qLqAoWau1Wt4Qh0ZKG8azmWNP8T/EIixNH6N
jw1cpd3utLd/dIsS7Xt5niCeqk+8sUp7D1OODJAtgt3NkXoz62DoJaqSOKMl7ZEB8oFBvHK6uw+0
v4wnZ0VujARkRZhRjsdbJJwygomlcttK8SVU10csY8ZVL9He/9JRAdc2TQG55U4h5Nulbsvm51GJ
IuurIlte6rSBg0aGNozbSE3G3FwBA2NJEnvi8d3vZAOKMGXO+xn43Z/G/7xU2yvAvHgQca/h7RzU
iL7X+eIBbED0txveoVr3Sf8mNDLrwYlGMeq6VZEJWv3ETlRgoA+D7gbisqLxeikmQXar7xtG+IFZ
q55LUwyVSCmraYf49t9f/wQPlFgbhS2G9+vs7/r7zY+I+sAW5h6cjn48YDSYKoJuVNhetw2VF6cC
OM1UU3JtEKOI0Yyjc5XiB0FZIq6FyO+6atk5BPH9mRWVj9xY/9OvQbgHcA3JhSOE7pjjTmlqcxPb
fxtst1SQ35Kppz3EflCr2z58W75LO/kZNs1lyogjgWsCrGBPaQzHqYg3QdwKp5C690fcpNeSZpVM
VgIljjVYXZ1k5uF+mmW1VJJT6ZV9sPwZWAuVXYMj9+J5b51RsJC6Zm5Xg+T8nSskgYZfI4Wnmxd3
aAWXePSulCOr21h0Y4IE3k5/f4SmD897MDHWLE8BAvzhDDWbee2Irz9dxad2U7gC26Plkc0gXMM2
hUggTyY9DtWLOeDiz3UOi0IhPtvEgxXuRod/NlL+iF9TxCfIFpoKnYt9lJLuIExCW9OiXPxauYQ7
TMGQbH3I1m3JG9QxJX4bG2qTaX9wMMlBcy87zqLAI0qEP6V8ZSB+q59ZWb4APeFRdnt58q7wSX3K
RUjmRH30yLiwIBpyq5cHUC+dC93r7ZS/0PFxaFpr44PF2tP+0uhfi2uLkq3CqvJ38N1rR7nWSoTo
X7gmoZ36rNJ5ATojDQ8dg/wmzJBuIt89SjMzJGcy1vBdy1ItC2NhOwE1iwAPPIjdF2D3rQLR9N0n
TH3qejCQD9s2TjRcYxkPWJB2vY5YTY12Vy1CxBZSV/Vopq8HMd5j30qZk91hEvfDFbbKDkLqYH8v
wk85ZGoZy1FIlozDxoMdupofJbLmwpQqcoYYtK/mhjZC9OltwtWLiv9kIqDx7bAl2IygEZsiuII3
YmEGmNACSzSmbsQNrUAYyaei+lpErXEoGaw7oSJgNjLlxsZXe/BdIEsxC4Mp6DqTeh/ynW0r4K6Z
FOT6J9faL3ZX6W9xpR27l8mruR5o6MIH1Odq8ZblJ9OAiWDWywOF3ujniGUbXthjP1vhct8z8mTY
4S9x8D6uPLnd4WKYKxeDxHnExgWlJo2+xhIqX0pF54PUcewvhDstCLjOuLTQw3anKimjkCR3sDGC
e8irCcwg3dVO4vJYj3jTx+ecusAlE6dabirKr1hIf6oyvWO76aBb7JDku7uLskU78F22ZZwWNmOR
kVTnFfZdLn0wCQxCYK6DsnAg51XsKznni3Anx21Yw8ZSd8uATQ7bUECkHEmUSO5eEZznqzj2OTPJ
u6CFnfMxYgOr808OdS03GAAH1VzBC5RBkKxu65uZgrmTKmt8VsSSO+rukmE+H3kKnJ+s4Sc9/Q4X
WJbwgLoxrKPmnCGRZ1OFqGb2Sf8OGeK9BnR/Am5w1gqCQDj2+66u6+4Is2qQkIHLtkE3ooc4m/Si
LZ17U5Q8kx0TOOyRw7mYeOoRQ2sufR4x2EKKpjq41H1ebit/ut+HNeOeQ1fxYDa9Lr13bT9IVfE8
R2ERyQ6Sn2Pc+D6yC+XjRYz6EjtG6p60tHU2VxTsMO2CiHlsubgMi/pgdVgHg/0q2eE+rH3FNn0a
338Wljfz/UIiWTPNJrWoskoB2DkEl9wICkGsyj0vAvluT8TzYYXdEY5KJnnu72+g0nUegZfauxPA
SMWyFGg1WYw/JXoSDy2TEAuiXjyzmiH637CfHICycTX3VU39NqHbnNb20OChFsLU9jdNzyxV1Dab
ENFZFPunJX/LKbFrqgRLmIAwIUr3uIwTHQXFyKqWcbUPG5xObleg1ZiMyekRCtQmyN2pNfthreea
L4Knda/OsB+VrFDu+3sAS7+a/WlK7PVvKSPGIfqhNc8Dld3hVWFbPyR7yGSnIR51JFaZ8vocP5UQ
M+Bu1iJJSaKJq1M7kRdrJ6FUAy38C2yFjfHO9cRiooUPc9xD8pMLIg8LGvYbWhWFu3+/4B22mo6k
q0qm2fFpUz9+xc2hWCf6OzM2W7qzEHmSBTlG6KEGEv9vlJ4PbiJrnqJNLhEcBqCSb+FblYW16b40
IrCtCzERL6iEB/c+PpGI4xCZ1Syb9PQWiWsh6cjP/4Sf096+zrQrf5zE6owFJcFvK0Ppbtktp+nR
vm08o+F9njWUtrpbkec+c2nRLiiMGHl9Ot8+yQy/Tssze4I52wpkwn8m9H30XYjbUXb51ikpFXaF
UWpFs7JACWcYGV9yrgSD6GQlg1GL10shLhDUFPahTZLo1BNJhHQpj7q7Iia6FgGSXLn+XRRtaRaa
tQ/moqmnULtMacUZEbt28/70Jzt9TKQUBRHShdzzXiRxho0go3YP3+EgOhT/+JNXNoLZ+4kNau2O
DEt8nSaad2nqmpv6w9aJRpHxxinVN97JaXFMiAs8NEBPeKfxd4HeU9QAnUCsUipel1PiHPIB7e8u
12TJv3Ey8yJpp2tTuqSq7gKy6rYJYB+DrQWjzT3vSYQZxpJoHUB1m5WCculFomyYVL4c1u15mlUI
VVqqGn1q/kHCDvToFuJzRNdovpdfFd6UDtMfuHkwb951kZm2LJtpuOU/NfbnbCn7IWa4shZDWy4O
J/sMqM1dg+iDIFyUVns14Gn7L9t+I4qCiKab8c5XoB36r/9ZQvnDeToDUGuMmU5LMyup7uXCaHPU
U7Wsu3s2QOFNlzHIFm9L0EjKof3ZkXgWPDNtkJRi/1lACVC5G+0p+I/Tdxap5CNxwuziJbn6iQJn
J+itwy1BCMQnsPL9cn3PD/x0IGc7PnjvImggyfw0KIKbT98lG23En0s/OBc1oP1QRGMTBJ5+Wkep
+EhoCI2WU5EfylJDMFyUchsntYByMmyIpsQ/x1PMlGHA6sx6elVUPA7W3N6sROLSv6zblMA/YZig
p45Kag5uX9W5kJeqHVTX6JbBiXQ/VGx0t/N03MAPqQHVGlje70jKBVhg1rJz6kYQoSVKIT6bjS4X
dikTAoSV1grXCNK01FOlvzErZhjZunq9ZUBpxIM86r8wD5ZvszVSEDIjWtDM88uuIlv9ZyeDGUXp
AklKGHcHGMTvgMzI69Khrisw/MJf4Al7KOGZpvI6e501OAvCvPrPcTog3EYpNvrDgtG9Mx+KhRhx
wHiYvqmc3hg2Pc+8q3qucIrJsa9x7kgUncu5qHOc+2j8JVlB1YUtn44bpfCbWHAnTk10dCAjZ5GI
igECzP5c9qFpH0oFdBUaUNvCa3YSPQ+C6f+njC75iaWlIJH+weBsXYVyfuc18slzM7xUm12TxxGO
5R4+45SVhnx6MWgKJwFfY3WRn+TZnByr0UzJ/GLr3WqElhdkg7dziEgxyYrJR/13PRRsjx5IdYFp
1JVQqGNOKYMXZ+rRAG7zT3Nj0sox6CDM6/e9mm5woZMXgvQW2yFOG3MMg3aXTe5Ep4X4vPaFIpm7
chKkR3oLOA7N/RSBiX8rC5ZnSR+/gYRLZBOQqxS5jKSGkP0kfZOVmWB/la72YABnf99UkexxHwGF
KvglWEhptPpHJNN+BqSDuVfCRvJLU9JveIHDake5PhvhNVHOhQ1osgEZXztFXAjvKEsBNrwNMSwZ
b/g1GqETRo3KJsADCZW2PTdtEBdPm9gVR8q4Jo2zwgAhQGoi03BTkjQ0bIuG7zfgZLq2uYenUi86
KXI+EV9luchedgz5dczj8Gujm2yYkjFy5fIrhAav/sByfjVXvUeqAlJSBkN8ydUcbTuViFiPsyjm
maDBQcC0LxJSrUXT9gR9HoOFSbblHAVhiqP3wMwU9B58PXR9QMNJSETlNATmETQCi6YtMqfbnkju
N0eX7u5KOOdb0NNaNFUF5ZZCpHnC79sQu530FrlJg/joVCeRIE/97916Yy7EyzPGvLED6h6H/DRo
s+TKNLS/peKNknIgJ72s544DvG/Lub9wo+a1r1GRNDAXmzaem724LZmx246FTAMkzrLAawHIQKOf
jxReNRYgAa7HmtL9ALuhzhcIBPvmtz12lo8UW4wPyDNVZRTik0EcXlRhdwtFHWG+TXoqkqSY6iuk
Cp2+7mTNHKva3kilbYBG9D7S+fL1XwlYLxavhjRpwRdqxZYJBA4/NmV4aNneUQnTTxUcz89bg5TH
6jz74/x55K5vXvBu3EFYiuFz4JrVqxJJsuM14hmwxs2drM6vyKev/e1lDyU+Erw7EvlmAbzFLkAp
CSrqBHjvaBv/Qd/mwBi6zNiaO1n+5KE8BDZxh51Mn2Dk53B05NTrmotqR7nNf3bOIyNYcjuINeTm
B2KS85hlQc6q6Ithlmo7IjolcbVfCJfu3idIjJ9O6/A1sZ3+MxcN6Cy/bqKsgi4TbeBYvrybVyva
fVxiGgbTJgZ3L663+lznJFS2fDa5aT8pe2SlhGN8pj9whIx6z3t+tHfHyeQAfKgWDDFjJhwBeRi+
youvQbl7E6EArlDxvuqI/m+qRCDH6tF5yBBACyOhZpDFF5ziTHQftZq/P/RJKwzBk3H4II5eWtT2
qRJO2HYg03pJ62g5BkP0i4KFmBzYqranrNK11QHo3mYk64XUSKy99BMKxbVNBn6AVJ/rRZ4lrc29
H6W8HV5P171AgbHfe/DVDnIna1jVFg1qsGTRSk3CzZR3JjxzwvDqlkOsjFnruvvIzSF9Rt54u4Ik
MEk1oLO8eBcDKuPqgwgTDBCnAnrSHiJpnfqeyiqZyS0s2tWTr/W3ZEES4D6/ncL1xNOqrG55Dkdf
HsDu5Skj9qYuaGxrP3PuDYyt3qrju0TStUJTo26r46NU0et/Ijdd7cHQOetZ13dZc3Gb/IUh9aY8
AfG33VmVfPhYmF5gryKKPLmi1p9PSc9iWlqVPXAjaQCPNeIZAi40OjLztgLZQa1xbdn8YI5lew7y
Ti3nq/eCf8g5mNrQ+X7F5S7HOjqEuDoLVVoJYYdPrHaslD9mdnGlUv8qu9q9rrF/3USUZzbOywvx
cplox4iVa8ZVc5E9by26AYHwAOA8Yv+qGG1DJ1W8dzK18bB1cDPZE7MbewQw/sMf+QGzQML4EJaE
0tM+8Kl41mrWA/QBBK3b4psCQ+qS668zPsPu4HbnU6zOsb22Pv0jJnGoRb/+MUmkYktmuwtdFK1w
knozpK45CRMGHsHK/ilFZzT0KWzd0zABFGZBQk77JsQOjzg/1fzLSIkkkBklx7fmY2O1TgYvxwS2
AN6wSkUyG/pAcn5scK6p1/gvz1HsSkomSCQhuSKmQyaqRmrHEfiZwni/ayBSz0VaAd3KSdInhpaF
QLY5OG37OWpt91ALDD9cm16+xfODcY+o3W2p5A8v0CjSWBG8XVCpy4lpe32rSBf9ZtYcWKQoKv2s
ZGhs7CVS/EAFk3mqHqB7efcPymHEYAqHjxhFKgPdujbaTFoW8ILETJbJOqJ0Fx6C5XSeU/2MNr+n
Jn65u29WPxu358FjczmrkJZBl9RA80vH/ZWjqzf7cd/Cfj5lgP8XTOGC/RBVLsyR6vAAsLszj6M+
H8C9mK/7DONM/rUjBLeR4xoSyNA4i5YM4I3ThTwKNSrGNoq574QMZnJk8uNBrSRydZARmyTYURbk
PL2SYBoVS9A3oHmYXx8D0pAAwBeRAcvQc0aCU3VP0ZMk+gJkcMAa4gNZZ6EkaYZawt3KHdE+exAk
Rc2Shj5CncEmPJkBZ7Xinch0oeT38nOfarwUYq5vUbYSWztzHJ1AcwprdVhTS4kDnqexXFUzHwlH
mVSQSynmq1niq+cRkHv8PPYowWRBpNpDwae+zEDqJLfQy9MdZ9NXJhf/d/iytglWpfZT0Cv/Cfh5
UaZ7l5AjFhgqhbZdNGOOeHb4dkIIaTQaefIZORLqDtwBpycC6TBusoqD/0qosLh3aUXu8OYj/20l
FutfkzeEI5w1f7kjDc4b0dci4WVa7R4OnODuXV+eubSM1/Kt9ZXX9N+xO86Ai8KkTjCNa47QBEDx
0bdL/RzTYPqY0yPArHrRr4rN3gPs2HrGycIGkVzTGMt5QBoVP76T/dkiKYDZuLTdsTmHVFCaQ5C/
XCZ9s2+hLUt+UTmp8lKNgxYHvkeujDfLY7ojfGPHtZ5oDdFQ1nCjXF9OJNMFkoSqhRYPVZRqOITt
iKltr0Hw3VYtJl9mZBNZ6Rl8RdF3qBDTyRlJ5y76uOxpi1nDUvzDWl/rySytXcfr/LmqAuzEuhcC
mPKSIlIFM3tMrIpR7X471CP72bduRS+11wgk2I6AQMzl0f+T8Imo9BPa+7cORZVb0yw3FK6Rgd/9
zpcxq/MzWh8xXPmXVann05TpXKpntnfAJxq5ID5N9MzlXAmUbq4o+F1oqF34tOvV0A4ODfuKHxeQ
hXx3cpceXY2z39M5KPUPUdJ9bjWJ8pL335aUmOdoy2Hs8MKvX8rnTWFBFkp7usOrKOw1bo43+9Hm
v2i2GIrjp1HnDkqJ8BpnuiT/9Jx7d6CvKyb9DxLacRkfTDkDPFpgwYuN8rkfTzUSlyXJGiy4HmA0
2/hVr5RsAZSR5XFt2IkxAtYAUbnA75GojkY8kJ39IYf1KgocD0xid4PUXEYBo9aZD2gWFrVXYn7O
NWvdCloE5fbwlRXCGcwe0NvfqVBSlWXqs0roPcbq47sXDbdWId01r4D64Jsx31V/+X6/WozLVskQ
VI1t2tEH0DVG9cb58eGeBAdtB4b03HIJdZEHjap+CU02sSq9SyXO3anOrx0JAxNJS5+MejMKzbJe
ElJEf2tsja1GYHBmT0iSj2eIxQnoni702wxee66Bt36XAOf9VTg2zOPgF+WhHH/+iYmWyVf/avpV
tgvKdPBC83/hilfpzraO1AX2CRrfRQbIV7gfuiE8KqxA9StZE6g73W0+K6YJHN7cQ1Zli6UobxVm
Su7GGfMDhg7Q9Qtt/+WshRQpVul+Dk32qCRB8LlsVAw0M48L8q4Tkt8IENHiVvKOBextDOpBW4uv
BzMjqIEaS5uX7NK1EDXMz3kyRdaPCwNGSzAgUI8rL12ubQIEYTGRKMIdEONcTSYo+FpNcpaA76jD
XZTuqPXZeEb9j8OSrswQBMknP+Hu3veZorzgU7SszjFlmGogMEHt/9ybHYRB5tWcUZK5/G8/nIJe
RhslRMnU3EVPg76nhfX2oo0aa4CP4MuhfH8maWZ5FeVftlCA+U6NorAMKotA4dj2EDMT1lM1OvyA
zjVOOUvZjbLkc0ZR0bkv4pbtrbdE84KzbTZuyqTPxJxJTGT14IpFIE8et8JXnnsnXJpDaEYHMX+m
PZmpiUBJLb+XRMSo/8EqnQ+KLcx9l6mXRT5CO3KnzRJrBwsyFCGpilF7vEW1YFuj01AvjPaFtg+u
T+ih42QoIsQqtgw1AHWXtZSFsERIqIODt8NwZPQhjJecgF3L44pHAiPZgIxjZvBR06Chav5aWXdH
4ymoHikRCTJJUWIZjIHA4Fdu8ZGl3t3G9NS9zh9VpnYWqNT3tELoFdx7juHW4elvA4bLdCh46FCB
oh645ShQQwJv+K4bhYPg0y3L9UzGqzQhzOsArzhQqIX8DTlD5rxSMLxst5B/uYjfuU7MlBnwsMGU
msy77nNS4IwwfdU/ro55bnggKcJVPZXfqumW70nBRTcSsHK4a17vkQvQLO3WmUUnTtcfHNw+jm04
1aWIXOgLy6UbQeGAJFBs+5W+j9b5xk63i3EuEQAlupq6p8p6lPc1HAWjAlm4CMM94cHQUsKv2jKz
tnbQt7cSAxuHjVYfYx64R0j1Z8dm3RDYUu6zwz8YtnnxIty3/0zWVz4NIi0wJu3Idxwl9/pEKFmp
w/C6nAIt821F+nDc+7C8p+TW+bgvthEJ06p+NU4dq69ipas3BVwFo3Zs14F4OthVPK9qWDLD0rc0
7C7Bx2NmVDb9E4OM+f39gWEXU3mbN7+lQqY/V4ciaT11LsJewjR/g8X5flJBOCHGsAu6wqzip5bI
cD83HgwykMyAO+ykvUKyjX/AuQMMIIjgrwvVfz8GbJDizMgrX0JC1Nfb+lDK4mpxuf0xqpf3eS5G
gLCO9CbyhZedZSMSZo9UlZ+z38bQykE99HP77g+Babb0U1zKvg/kiWnnABpkiMQn+nY506xVThsh
K5l32ehJ7BNVjqChFKOx0vGQlrUrRPccHAo44grJylM9dRNx6+IyCqphUWKoxOuXLLJm88jO15yt
6yga8hqkBs7Ri3zY5hzetE8A7C7ie2bo+XWj2s9QuJmDHeqP9mFn/XKDx8Ce/qMK7/Buq8m19qgj
gxfoaWZXceMuBhtdU23Tym8U11ShxZLY1qXIWUDtlROTCW75H64gTXt5coLU6cNVjOHkOs7nf4A3
R+Aq00h/j6g2LTUbzNQzA4FOSz6agog07nD8U3I3Hyh0P1XfvVItsaWW6J7du1pICC2I9qdUuUgD
SHJRTw2Rbop0mPD8GVAJwXgNTpesPQHILVljyZMlaTxrON7HRxZumjiuovuRaiEVwaCcXJgH+DyG
/FU2r06T1tAkIdF9I0bZYxPZnPk5gR/sc91D9NQXTyZp9E6cc7ov6s9ehV8BxgYDgTChmkfwi+qT
mitchiImHCrXMWsSbt5t6P7z2orH9qFyrgkeI8iIJKLvBjxqqpobZihHTUFseYWU0pAO0cEULPY1
hdDRUbw2wzYCtE1BlSgJ0C2xR/5kZ7rYWwA0br9z37R1dZKwNl2zCpWEWMZaPZpT01adsJ5wDW5Z
Gt+P1Nhpqp1r9SAN5S81wtpAaoKeyIF6NGNRU+pZzOtmUlF/LCEClfQuAzUyXFfQ8Y6igMuv8pkn
kGbvjCIlwFDF3G+gKs1l2Qsvml/WQnaOXnnVSDTA0lQFbcjxU0IrQalCCKfZ7IwwySD34Ff+6ZP6
S6VmKrJ0VhrmBJGdK48OD/ok/k/YK+c2n+UCTa+InKNUFg7BMNY1u9ZMpCVrrAbUHMcJLlG2aE+o
Ne+0RSsZSYwbMEIM2dXpg8SZ6MHEQGnI7olwnL+JqfewWqbr8tAIe9IY7L4DxYW9Ue4z9YzezjDG
DKcJT0H7MTrVIdS3s++4tEhe5N0+R+uJtmLIuEFBdPg9BUzol7zlqD7YDuS5QZrpZABG6y0U5er0
3iWHP5TL4gi2fJZzkIR+QWv0awulhOpdyF9JqsYC8RpypuU4poDllezMvMC5p500WW24wBEH1rom
TfYD069DkgXNtupVV+4mNFRn1hMyreRTiLd8qdso2ubFlOXVu5ZbBjzFnvF6MGxUpN0tJNaNESln
aUhXxJmUV8lt2+GN7BusJ+RtEZHE1/YuGaGSW8C5rhaQqaYHKWBHY9pI3FoQFQGdzS8GsvKLtwC1
DhWGTShfLSrUTTIZrdfMjGeLMw/FFIFHNGHdk6xqy7Xak0taYmTAOUOwq56TRqRFY7W+r914iime
gFZmv3Medb+mF6KCFi4/yGkDjAe+rthENjFHIp4PT4Gd6MkPLvpvsOy4EKQIrws13KwSBuuc0h9Z
1bSl7/+oFKScRaRVeGVVnyCQvXjQnbfR6DLmQtjL++LF5FDwYvXY9ViqcBeosEI7BWJHI6Bz2YxV
AJ55YCGazI75jq3OCmmMwdXtCFqfAkAOTr6As6PBnfD+yYXBbjtt7Tg54SGd3MRtXVqWdEpSar1Q
VXpmvdqPRXnGZ1TBPjuKX6+UgpkrzqSScqA2CpSC4qgXCFhVOKahUd8xONH4xUPYBnuatCmBdWhb
ZRASwkfdSIuXqLgt0knRZMHczxDa2JDhpZb/Mfsfeo+1TINenIMwYjHGy8sU2FbcE6hFQ+2AgjDq
vassdMv/QTQRQzDayXIRhkUr5Pq49gWq4f8BAlrnUK5sf7baugY4Q+zdGGJbBYp+hgN8xUwvQCnp
r1c3n5tOC8WYT/kK+l3poOmfiaOInQK4RGZk6TPOirL6cq4E/8I4C0w6NhsrDCaov4ybU0ULbLew
XhuvaysnwL+98lotN71yPSrLkfulZkIg1AdoxGpiTAAuCxeDq/LYVLHjDpVgJYc9rEFwrmYA6wiC
GoVxdVg31YNCId+Z1E43YHl6jWUFuPnkxluxwtdX/xPGssodCzlnnUL72hPQO7JjQ8VqEcs2kkrl
wJ5HQh3zvuiZl2pKQPgIVR1ycPAct/gyvIovD5TwCw50wOl3YI1uyjFgM26x1hhOpJwmcm56CfWf
DiZlmdzpsslOMRranJ1UOnewL0ZhKRBUGbqRVPfDzXax0T+jjtnjEz5s1osZeCeD2VWTc5aM1OGN
nmd1JSJUVqIdlaIw5BvAha6FRc7EUKFWmeY4KmGTHHH8YvNBmXXNRWgXhsKwU85zr3/221aXAWZu
WGuimJfYWicORu6vOner1bn56Cr2oKkJXgwlJonM3mNvOINZvVohMP/VcX5ryCsc+aDQ49RutyS3
doMeDhCqaAqZhrS+2WvbdxYI1K+yYzLa5vPJ+Ugzv54SQTYZlUCHl+5awsWMQjvUjvL+4WPUNgJY
Eb3opK4iqLAbwVDI+IQ/qAumF9ZT+IAfg9xNfgm+mIevieczi1enwsKJNWa80crAQDxtr6hfHyZu
Z1h4Q9xL4fPmfQ2x8Oe9OKid1nCoBzZLbfs6YtzH8jpwOhrNQcWzZC4rLm/PmtpQ44QdPJFAftGt
umOWDeR1lvNWgYSOOMEaqC0Ah2nktIvKc4+0tS9RDx3RpxzP+ZdxXjHUUnLBZ53Ly6Q4k75L0Rha
lytkkQJbW02IygS5QARD0ycctnM9Ejw7bjyAXwvTxAhecrqnbh3wD/fON/rVA2o5VODrzEa+NWG3
X1ZcK8AzeDhtLpciQ4LRXqu2plJf0Px7OnLtZ2fj8l4v7lPabW3zwXW+pw1VOZ2mIcyh5STVyres
HF/b/Di6Xzu0CcDkhU1KNYYpg8Ss/Su20lmlWeXIeR+JVhcENQYPY1Eeo4072/68oQ3PB+OOPQQn
gWNlS04NccSdU99oos6ZLMe0DN9oz5VAC4V04j90FASmPKXpaYFSuIBiZSGIH99tWQcKzGhiRoot
TCWCwFMKwk9h+or6dwfFcqviE6oV3rW86ZWmHnovmkdlLBw01RnMU1zkkmVgXo9T/IuaWfcHaCYv
UAAHqodngMM6iOivS1Mm1u5KQcDIKvJEPtCA/CE/Hpqs2lvEH8OiKdExE+s7VlI/1LN9iUyN5x+v
mrUCRXb2t5IanY0+cDk8hf3b+po/Pk+LNhdwIWxTYYnlnGVxTFRbTHAEwW8FcqtuoU092v9IAyTg
xxK4EdP2wmbI2K+wXGtlW660H9YHexjbcNYIl/yrbKNJAnOkX4JItmbqsUvgQMRH+z7YKVExvm/4
gkHfqX9WxhYx+7rRdJYsEzuuUlRxffzQA0kNcUcFCFulJoV9BNCfyd5mkQ2hoBUXm9SyZUZM2VUL
tYbZKYowjcoQQ9abJ8GbKo5PN6CDtLVjh/lx0Mo74S9err1m3BWNOwfMrahn5j2Ivza0dcROn74o
XAyz34o+B+PC/mwXbaG8u6nQGUPuAruFXLsKPmlnFnoFEy53JVPe6gUFLgJzymUsmKbN/hOP9CDW
zENMwiPvzEOqEjlYqITsmE4eRoO+Pri2pTvg7GGMkBJtSJ7lP1jiD2Vo1X/jWa+0SuohEGs7Bpky
AFpZDuQ8aJfZDp8xVt3A30+4ZRAcDtUa3gxtL5aJ43O95mGphr6s7h11FKz29wV9cUmtvDG1Zr+y
+IOnTAPZ/Rm3NcNlKB/cOOtCeMxihRCqwDfVsDf2G0aYfLcqSdkZBE3bTpPkEnU0UgKckvKxXXvn
1WDaw+a/l6JhGoxA10GplbwZtvp7aKO7OJwSoZZwv8NP9FnLnaefrx4G/zEaE/tTD/3rzAeoEBBN
UV0us/hHFgLwd+0q8alzcVaqyEm8IxwNeesZFJEr40HJUJb53EqecwPBXl/aJrNmNMaU+8/7dXOH
pphMnLRipXWKufmgtVjL/YKGF8AEWW76HXkg9rWYd7JXJKGmxWpHHykyNkg9VVyQBXT23734vrxC
ce+yBLYdjrlQpj/KVpJD8r2gbIABwCyX2K8Sg4KEsq4hM5CCoWDUzK/OCJPajs1oOL4/wHAgLRIs
pfFolcrB710bFiaevSKTQLuB5hkmSA/8LgEbkCOuTPUB+aQjpk6F4z8xSXkePejxSYpcatk7bAza
4a6ut/wrTMvya+vFzOxfBltjC1foqVHlMKoOl+xPD575Irnrzdt92TFxEMihzJKeQRV1ac/jjy/n
ruDkYi8DdnzQM+/8VWmFdURIxOlZqNfPvBPF/XhRMBf99D5VrO8mHuk4tHKi+Q2l6dkDCBuN1Rl9
OGdqnPvh2QOGQtPq3oVdLiLh3hX0SW93ClpTeH4u3a4C51LPMH77PCP6ioeVlEveJHoNJF+ls94K
JHFUTQaH5fv16lhJt0QQwgGo4hjvb4Wp3lHAem1TmM9XSjBu01ygA590DgFalNxZufW5Z4HflkAM
dOs3ZNHMdZDynZSG9xCmfoP5+kYxxaFINqZ3bYA2EivHw4E0boRJiUAyKOBRglGH3KAr0h93mynM
Dz7DN1pr7R5D6RV6OxONxxlAaUw+4mJaOs+9378xvkbihfd7l6rw5dQt+quaS/dmKm3evoIfkgw6
RFhq5rxxvSGEnTfR+GA1BnH0SbkZo7/1hg24lxU3X0NhNeCv/E/CJYjmu2kTFZXzCGpr2OIZeVK3
Uip3ZVY5Vr1B+OF4JW1k3LLg1VIogWZ+JMSbxfOUcJicdIT+p/4kp9QXkB9xeHx20HK/HvWUJx1F
6teU2H/9zW5YEqeoyIYOkGYIQ+4eukueWrGGP4FKiUIHSQX0qeZs9+4OgzgjmTErBahTw6Vlb3u3
AhK1XTfhpvfGeFF4BPjz6Lvbs4riyHjb2H+SedMydKZDYOv/W7Z4gbnKPNwuGgVy5qfucPbuTJgO
wrl5UAWTT2+NdWSN+mAjZUwBz62U97gi/rQzijh7YwYmaFPqilrOjCcfdZDpZPNh4JX9FiCvu6z3
3VE9l74LHsgtjwYT5GGYFAWlEZT6/vA4CaLSOxS4HAMkM4cdFeWfOjFiZdr0ZfLFqr0DGz4h+S2o
hHq7gTSuGRnr23CYLYJ0ek35Ks/MuHt61wcNRxPJ5OAFG94iNnjSG/DLHbe9csp0YFD2X964pGER
jVXB3fRjzp7eem8DCFiHKv3QjiDXLXJJ4X0xLfCqchgTKfSev3aFOjMbMjNhfr0x2z1EC5s/FrwK
X+Aziupn4f0rq4HvWT3PcsuPFka5+W7f+3o9zJMibvLasNi0Mq2qCGC3JUE828zUJbr69eKzpx4J
eWpqaPs+pdhUd9hTjPE5GK2oKUzhclTA7nKaIF36HSBcRhc6M0xlL4i0yWU+4yYOFGwru3cAUojN
QFnMIgN+KxzLIv1HEoWYrgZGMScCKlbBiM9LRq+ewWq0kKO9v68F9tp+E93Fwp1yRABrNwHJOdlh
2K45qD7vPonNW3AyLr4XyxCsmtV0SNByDzulzUNFoqHttcDZqNXxwIp+oHbDctIwFfj51YZypyZB
3zpxS3q444A4zchjJl7gwhM14rexdGDeqP/Bbtsr/IxV/iy/SPN/BIIAMrCfY7C7NfDsSkAi7Cjz
w7DGndBgs6k7BH7PUUEbrShkHEHbl1qpuVJdp7dQ3j/wPrAXRPMLc9mCurc2KGLDO+zpYm3iBB36
BQdpFgUoVvl2PJatvid7fY996dw48dh8bxpEDFMKAgIuizAI3YEhg8siYhnOCsPD6Gas24US10U2
4muuEJBxS2xoYsxbdHpSK/SwbisS/BNwNm0+H48MnAwZTH5gdVrd8Zu0/voi5pe1DMAmD3evTny8
bFasoV6HalD67LTzN7qGMG51j6++NsfqbVs8NIlIiYXozlRame3fpXScPnHcMBk3uOlnhzgRIwQ3
7QRHBIDl81miv07kYwySp7C0FbzAsnKl5xIoM4qE+G6FG6IX2RK6XVUeCI2mZ9SgJj5IIFuLuOS8
27jQdlJVHVloLBiIEuv7GTjyvanrJyKwR4UoS30gBL9fPfbf/TEgbypL9lnVE2RInhbYsJnVavVb
FHGoxi9N1dMcdgClfWOa2yPjn3y5XrNxkQ7H/Dx/cobVRN+3LShtDS/Anq4N4sDJC7D8KeaBabcd
6SHBlSe5ApkXdq6V6Iw3/GUt/oJ1XTy8Mu7JlyJ+VFeQoHObxGqXirYvWQD9k1YL3xU9KiPNkk2J
QKKOdcVImM+qfv/qKnoZamkdtaKSNlwhhHV+8Su/3r08+wgjrc3Mxrhiml02tTO2QKSMimgTSrNa
KSggQcEwg+U3LOoKJyO+UUpJRD6CBiFFk2jVbi7rRw+1Kxc84o0u6KjPaPfMPEZB8u/lo1n3nCGn
Q8JAxdRB8zVPuTAjdpA+xZd0IEk9SBpZNUuchWSxvSvrJmFny17F435dxoNFZ8MDg22l+TU4evp2
pK46Voae7IMcB9/oMAWBgOEaw+7WaqDa7iVNmFAHUKPJ7SWPURqqZ7AsspkN3j0IPQ5TNu38Sf2A
cOicUO/tlSPyaaWLq0IJmSX1WLglKGEPZtBGt5x7UXtqrUOlx9esYuHYZwmsZCvAm3+5LuF5mXms
jD0bwlc0WFtIdksk+dCbHFHTpnnUFPCtZK86rVprELeAppCx1ZnBMTIojtEiaO555XcPnvpUAZSO
tesQztafndxmKAZ7RXTKM1Py5hIs2XvTr9e9htlFgT3HbfQ1FqHDAMeSqXpt0/aO0BVH/70y3mXt
mRmhnNR/Q9MNdaO80hHP0+iWBpEockwdAso+bn4hgNtsn2Wn3qjGKaOWL8FVgt/ep2uQBrefLyV6
qSfT50ngSA4/bNue0tzrSd3SiEE18GQ1DpYdXxULqf2tRaZGUJyH+KYQ8j5yrJP4ze8Jx8xpP8g+
BBEy1zdYaJci+nPaHuRHIAj8vmddVb4vVDPDYUPh7huHf8QSDUOrGJhU9SLpzXV2sE+ZkakowwiI
5tkCYBsqR5qrtvexhVUc/fu6U95VylGgLCHgzjEP5TVeOxxa/Wo7M2MKBaHzpR2Q4E8Asm3lrhNq
+UyAMrTW7oH94VF7ZSNDckpO47mFYVSdX0dxKqJAaVZxc1ObmlqbtiqzdOFFxa34cYF7IF0hPXBb
JBpaISm5AsQWanFq194O1YITMM/HekFY4JewbnvOE96l0QgFQzrolp5dGNV5Y9Hjategu4n+8Q0g
g6xeJf8av54vEYTwR4vC1Vdoh6r+jtTud6yP+1+jVweQ/fux1AULtr5xzSkD4znJdnfCd9IUjnoG
oZKLpRZSSQGIMgY9vFkDcK+LbCcPphRcbIKcbfd+omXQgwyYB30TfyPwCbX21+winotRywE/G1Go
Zs2ouItwAx1jB9uWRkfcvhSttSCzUwspHIMDg8v/4dQ/6d9n/0nSo0TljryD7FYmXxWBjcMDC104
wdtBd7YAhwsuqNKwcRygFEVk1n08Dl2Y7Vz/tstz8p9cxp8XtaKiKTiBroIEfuW7jg3/J23Vy4ON
XA+JafBMx/TvdlTSLIZNCagIfvBHRXoUQtDrPk2e/fkrhQLGCZ/Utg9zhgQnPQMRxn96ZAu7dAKn
sfk4drIsevziN/g+IPMQycPPIVnXrrf4m0ZK84NGrwJhUtQX90sC4+vaJ4ryuPHybTsZyk4w3Ais
yecxKGcITbn5su1f8atuT8SJ2TP+sUEa3xCWk1dNWRKAnYM8G1rFccYy1pRP5tKOxPsJTgLf3TmO
lrBp4fSzG7uwvLS6PBYz2SmXT7I/tX4HFbYC0H9g4kMcndecwNti4inWTdsPyfvlOdkHRO6+VDAH
9Qpf85yq9uXU83oIpzmkiBEShFbsytPmZoIFGBQxCH1A2lTX1EfY0+dKHQhvK5XYc5CXoxhaZRwT
kBJtvhKBDHfigF2cZ+RXK9Zrkvy3X9gMK+JqTk0a8VN4SCbuSxfWypCrSrMChB/JRAUsh2pJIaVD
aKKhiJO2gHZh9iEo62qtYqSpSlwa59ZxzUSfyY63EkBR2muSwd6VnSXFvyzhy8LDGvgCVjDCT+79
CXQcAgZqEX6eR3ov8GrBM+Td1BdTrZ+z8V+ARI0PQHW0FLy1xGkB3LI+oqc0urNlAca67XjO+4Cl
27nrYNyZkSa5xvCRe3FKIXA8XsmhAbTNO+7ofgcCdPyrr9hzTpMHpO1tfRi9VOQVaNnW3rOe35A0
hNL0w34SpsBfRk+cm2uDC2XHX69dGR14Lh8w5gdgfL2uRjRDStx84xtzUqDDgs42kLGxPY0QebZ+
oYA9SB+FH5y1lCdup4+Xp0Uck/oINnl6FGBFnueGv8EukOvVek33zOWQuXM77x6GURvBIcjGaEej
3dwqfdXywO4k9NT6XRZl4dsF+WroGgR4SWgl502C+Eejwq31r30nQ3JFDjAgZ9CIFmes430lDLfG
dNtcIB2K/RF3leMMlHbgTD9QJVRizspSpC5A+9nPW1nD1vvRSWOh/iytMBO4KGL6rwiTtxgqg/Nm
v/CiGN90XGLoHs/w2NLm3qY/DClM1IjAx/3/53LLahnUBmjIb04yJ6L5FU21Y5w8CUmDkCHoZyjg
SOlDBo8Ogruseyc6dPDcswKhfpFZuCCcWis0UNpUE/LnTM0xeADPo/xPocADSBz8RGbFOu7U1YkZ
4mwsDb+src7bQc0NJmw1CVMeq3ytM2cY7Ns1UJZSQagUHi1VdVN/qjbRdejCFYdiD1CHbItsJ4Se
l8AkP3KtIVdfshPMl+xJT6m5K3R83FgixsUmcUe4VAqAoZ94dP+NILJ6gwKVPJHJrJXR1KoRlKRL
LE9nE8VM9mgpPp6xvm7Zkomxm1GK7m4UAt4Dur8jGvLFBoJk5Su8UPdJFVKAzrhm9NOvl8IcEXhz
mZ25uZjMM45hhhC8jsum3O9ePO9a4Y0kxf3VNimXgrtuPXapk3DKgXg18a8jBdIit2xYfoFyjwME
01vuTK9aWUVHzcEK2sRn+x9DXW3fy4vfjzvZr4fdnz8ducvynu0Sqxh9M66/iUh9/0+cEzsTsVr0
wkWLYIxrU7nAwz6MSqlqSZQkrWrNHQIXxQ16vWecMqYBl5UWKIWSycCS3mRNekLHRuyrTjOPKEMr
KS5U5BQ6hKZTXHJm306RpA3uSr41xKrwLBgjp4VRA4kPCEpiWb1g9wW92bdIZshNbnCerta9udFW
FI5b2i62Qylk2stNoodJeMwIGuREVqyIQSbD+uZFzX/zehQZ+ssXCZN4b+jiAcUGf2ufNfDbZI8Z
52iVWTjH+15BBu2WNhO/I3jFbXOSQQJ1yBz0/e09raemswKY9zMXh38/tf7ki8v843BgBCSUuU+3
Z13vGF+04tJ6K6slUYGjpA5jCqLIQhHRKKqvh6OKQzz6H0xdxxPiEG6AU2h5ZTEU+1Sl6cF5EnAD
h+TSDomQi6/DLyqKDEHgZrbOmbFjD/mo1LKoMMXquxUGLtVu8bfOmRUQIvA2I60ozoRZMo51Fy+9
WillfZFSPj4BKWj5QJjjsqzwGPbbyf/VE4ONBsQZkhdqd6br+uxffs71W8LTbTAfgJV00I+P5aK1
xdjWTnf/i+QipRs6pf41ztqwEV75PfSFHGBWQFwABwuYnQ9PopmxQWbZoJ/GrNhFbTfZ7M5va9qy
fws0yFeYMhzjIG/BgFSQVV4zeFHxt1bK01DW4gsRGDoepii/MS0q6DqvOrSZqSoE/6wDKHLvCKXW
b3wCEGLtvCIlg8LfspDDBjzxsxTsGyu15hkYCVu0BD9fUEWs8xXz2+ErP5mOFv43hqaWBOA50v1J
4IZNlcMlBzEsIDFKDiddLwhNz46vBVoroo15v03ENm0HKpcA0eKuHLlxwIxjy2IvPVWWbpsjGu/B
UFn6sYBMLjiHzUExXV9rh+4hy1LlGuBSOZsOP1r2RYfFhy7FzEY/WpBK7+JvkehJdYXm15AMdB3/
Uax3xEjfjjLjYOdAgfBNjLQjCXyOJ+kt/R6LJRNdSflRiR3e/UM3NBdA1UIoi+CEQIvB6EiIHyhS
BHgYQjNeWO18tPDErH+QGnWyLNLC/dSaxlSADly7NJCEIcKhxfZL2DQ3LMLeXyUzS9JlRo45/4uI
j3pHWdDM6SY6VmBiuVui+OrJP9NcWhfYfqeoeYBAA058naObOwuRqbd8BMvfu4cr7L9rZ+kLP2Ha
lP9emcQLAKTDflrL4UcAUm5axVmvIcC3jo2BtYSqpntyazzvpTD9XI683QBDQK4zZV+TLY6VKmru
0trrysJCWBjiQKV0YtieUugqxjg48bXS8RJgYBQfYPQ2XcAQFKn5JdCJ//EY7DTqoeIaKc9JTlDt
OR1QWtQisH7qyfJY1xHnMXpnoKh48yzi2zQQSqEJXHsDf8QxzPT3Ut+rPKtBHSIhE7/E9yembmVK
UQzsDGYgGBSI+OTJ08pJ7ETipBuPSKL8MgEOPVqCWOecZoo96tVCOU4G2v52Kzr+Xyt3/PrazLU7
ICzDpFSuEBoGF3sd3XrhSYU0HyKn9B9f7yzRAR5m3jyLSUrI/4uKy6bodMNY+CvTk1yL6x9n+rEw
Y/Dga5ruqi5t1MLhKJ4qDPTTkIevzpuLPFDZRRIwd9xvNF4FB/gDdlK3qug1kpMoS3yq5QU1RbCS
AFpiRae9w3yKeFqCH7YQC3fcncqCB/4TOEz+1tcRHeIEhd2cr9D5coBLG/IKfpIN/jLzPHzssQU/
MEqW/MCngP14L8NTNv05QbB6j9Ot468ZSRjoeaK212xVdk/oHQHRrJydDlLCx1FY9qEbyKXlcicw
cYerRACurc9k5CavEZAlLap9s/L/gfpbB6g7zYh3w3tdqXnGAcS7BaJXrPksNmsnFeUPLMAmMjTf
C10BU8FXMS1PM/yz8yxJTnHQRi9Iws0kKHp51lmUfhkybV8FehcCxZnVyFt8UIHbVwIFS/gmBcw7
48VR20/n5jxQVO111WWHoH9yN14WzAA0QNTCezUjephl+ChtnRjuLCj8scz05CVdg8WVKa08k7hv
YngPkbUx5T68uPlrwWPwhpcnvQYc12Rm06jQLgqFyn3ahmJvYjFvfRZEUSWo31MOj/7w26bjhMkV
guEh61vack4vBtKquO5VXX2KP3/pJx+T4YZB3++1SZ6sseXkPwSb+Ij8JA4BKHplkixCBihfTAe6
Q7LUVtsjdWIgkgeBTTQ3tNHscbORxph3lEo2JgkKjL0RtqSVjfES1hIoMfeY3A0213DwSVSLO59M
qUieViKirPQzRJtrbQwi7vdKJL5sp7m9FBLuIs2XFwmHk1/6PM8+C16oakGU2Iy7LOubiLTWD0KU
tbX3/n4CpUh8XmzFRYimm8TjDktwmBYNC28/Zijakit7ayhTVvo30MF4o8lyhnGH7GU+Y3dGE8Fx
Xm31LRb9d5WSVQbHLzBemXNUX5qKMOqa16Dm+w8tVL//VwLtAgl3ZfYvNrytrVcG+L9pPmmTD9I4
bfTemf0dRFjCC03ENHk3Cu1ns7OWCs1HB5VNPOWINHcENtAk3zrncFPCKIm9rQiHPa+NYtIKNnPu
0xN8Sh/5stbAGYQTLkZ7g/ke+POkniTzHClSgwNFpg+J49cLfLa9+AZ3lmN0in80jFcaXP12F7ls
+wi/IOaIvniBtVkj75Aik9cO/mBJG5TPWKFJoLas6BBMpum1sVRzp35wqLXplWo1qpkcsjSnxsEv
ywOhW2XFSHjWH5sJBguCZpEliyyGRzXH0tmW/uV+3voOiE5S4S351JtAmc843WW+rPSjWmTUzTB3
c84pGu40H/xHaKUwR665lujlrazBD/OOZ//+oe4X8a4LMhmKURTydsk04KzZZ33g2zGD1kRP5YrR
ws3fwoB+uksJzUUxNsXxXxu3lsIFvjjdRhLMgrjCyL7WaqVPrw+R5N2QUjRPdNPgcx9rWhuVdlLT
0sxuL8VySHZNK9hLGlnG92f9qMu+cEvOFunGj0E2Jpzd/c2PRIjRh3YDM/TGz99x8HfU+325dPxZ
Ir9YNOnf1cgjMgOFGd6Lc6cpmYyN3HLGkwlN6VSxg7hAdxvYcgTR7a2w65C1V/ryo6rNb8VAK3bN
rovX6pBPs3d4+u5kwMlz7t+1nvQQg99hAaPs92lQwR0Erb9O5B6HgYdXxZmxxL8Oe69Xk18hcWEn
4N7Vxh33/l8wUvnEZhNXgOCoPCoQyFpkHzE3s29F87Fab76MdK/b0buUa/p0WEL14oxAUPsTTTDx
Zd36XR7zY/oaXgGWqrvHGsj02PpW8s/v62z3d4nXyHVu9ijjfvbfcFc2KL6edZsGkGZ6JmaAYOBC
hhLL0d9OjCzfhdcSVD7G0Y1p+sAg5AyutvS9gHtJtvqLXNj3W5859GEanV8YveeFbj9edC72slJV
giLESHhH2kh1MZvug7cWTg86V4zwOJeG0m/Lb+6bV7e+54jCYpuAkms8jeCtN5Eq4zLZbiAXQ/yu
Xrb4lraPwociTQZAV904/41VsdAgGDLOIbzRPbMKvBaNVoKRK8U0CLYGABgp3cpoWwZ+6zopp3f8
pp54rwttSJXfjIFt0V6qGYcQBuXvdhEfxZFqlevUgII/t+reaho/CzbdST0aC8PbFDmb2DdLrK5S
TMHFaIqpGkVPOM7OqMEzqD7yuKj2xYMeBCJWmCg2eOEZ5Har63cOKha8z4R3qCCjs6nCU6VdfUAt
kHNP0XjgPdRqyspOgwV6aBBVxgT83Qws5c/Xrzdy5X9LM8JRrQogMF8B0z0icDkrL53hKUha+xpP
ZOOyjSXmKvOcK8JljLghlk79zomNOOZm7hGJuEHTBTXJnaDeHzGzwTqhXUxmuzScOxX0QwIk/2lZ
pUM1YYe/3JWl6OM9HEf3zcV260WUjit6EHw4NO0d7MpQWbOGp+6doxGb2isPRV7P7/cOoramWA7E
BoRUyQqVeoiJpAHQoF7v243wiRxSF1fUcBisd1M3HGdUIASAjpccRXoBeL3Ym5K7vVIeuY9cDNfN
Xp6/HPekX9c5owNnpO0Eep7AarM36W7CNisA36fdh/DlibcSCqm3NMp9QLfUP0tNwLG0LThYA0JH
5WNgPmJbU+xCVV5p/ExnNejX/EnQIBqt34hHFXgfIOCCZ4VfrpKXtNYthMsulrWYiesYq7W82Uvg
dYJpiNYit6HN6j23DNh6KQF0AsUBp1F/3wDhCRk8OXVlx0hoVf2sTp5Ga1i5O1X1e3rU2jyqqtNQ
zBEul5KmhZZf8TJg7c+cJi7oe+lx9IceTXwKcczkfwnjQ+AwfZHHEcOSRGQmL/10UARMPO/hJq6t
3xx4pq9zEQ+Nk83ukW7+Tod1wRh2kP1OrM+Wknxzaegq4nxwiM7BPJysUnGmdN29sT4DX8nUjjY6
icdlHkApzqGUfrOxAEbgFj7I/POncciArRJTj/jtDmf33VkoOd1U+pOBO73IBtCaDsSTskFIbAy8
EtUyPP2UL5CiTMTESvffUsXga18oBI8/3gs8FiQYKPBnVPO+GCOR+prCV0kDt3mTTcMsn3UEMY9z
J7GP9VZPY+UDCXqnUYvUnqLufLvyYvMasuUvq08X6A5ra/cqJCPEjiccHW/hdCqsj5UnEki83jIQ
UpLazcCcP1Q6L6Rycr+M3YHxjKj2np58kpZE1QC7h07D3Z8RI7crKVHWj85uDGU1hf1MfNpqxoRY
fvLJi13MiJjsCOcKYVE+aZOQ690kaH7iPRjQZXBFv3f33zKwKThcn3ZOhlRXBcgpahZSeGQMIfx7
defxDYG5eZYtKvFXLswWvByI0Xw34QZoJ9/FVhn9hlmwVulNcRjHltCQkttrcbEmrrPI7QRloCqc
rqtr3dFgjX8XL5zuDni6xyWxMJOiC+z4RzWzeTePNKkvwbt60xCzSY3vflQWU6MCPLZOcgc0O3L2
/52mtb3rgJPPC7mwQL4ItGNsIVVaUU6/zF84hC0cYCajJo8TnOt6BNtKYHRMGf96eFrC8Dq8sKWe
cC35J1P95Uw1dccW7BLivfNEGfCG/4DX/DdHic1RdjdQrR8vkC42t+idzs/D2Dv5GhTXUjyamUuY
nAmcSn3ogZSAWJSDy6bl5Q/9Es9uRJvdbWK4prN/TFUNEVhfgn7kzpR3d2UqhK3O01Wk3/6hdGbr
/2K2ysMjl6rbaMFtdJM/zUDNiHoFWYvtD8PFX9oshmWar2+axSI5bcacNqGCsA7Uk1bmUwLwfZLD
1FALkzon8qE/n65c0JxkJFaghz1rc5BwWIj4FMKXpG83cBgdxFmVDATXSlGSYD+kk5kSJJkc1CNK
0BLGN8izr/fUYcmruQPA23qN03af2CXY4j0gdaV23nUIKGIdq2qOA1ubEhKqD/AeRrjZ9nf23rEE
/+u0UEUMVLMIA9G9n9fdG+NnBKo2cFEkH8wflig4I3KpKFRBlHGeXVCxYwd6UQQE1q08f89ObaS3
KAyOkvfDykl6bdnl0NAEZADfirlaE1SxfBViG39bYhZXI8UXBH4NS1kXNJR1Xxd56eiJ5oZrI4Q0
DjaNgzs8v8x7EkEn2qS0pEkF+O1RHnoFlLfAwS9U/cFt4cpy+WylTWhzKzrF0nsxuvY/1K77JNXR
ZBstccoQyTo8uux/SyYRZ9pQQxniOCW2/ISF1NsOqBo5lmtkdZkTOQ4WZQkDV/6ZHTCn+HQLs/MG
KZQ51B0Xot/dVsXu2DZSWxA3si6qU0A/SU6wRVydMNA/EE9Gnn13xt+vRrLB6uBCgfQ8Aduq3hL3
pYx7OEipyvGUoeLpCn3vBHQB8cIAttaKXKdocVrvH1UWb2ppBid0Mtddj9zdFf2fRB/n61E8VUnD
mHOrv0vxIlXBztfr1jUpiIiAoKgJrHd2VyB9Y9KBGCMWGgQgOKhvTUXu9TB8svdL4gOmkrTHiBcv
bj6AjAhnWbV/wUIg8N6ghOUTCZXmO3vjURVZ7zj8KBrL7DGkpjWOMrTnKMm4Z+QV+eTW/PK46IhV
UoSVnevihZx9J1Lvr51eUzslh9o9s6cnzYqAdsZr7fgoK4tG2vPFyRY8vFoXyNEgzBiAmmD5VNUw
GKFbyaaZSKF4PDMDz4yPnKpyOT/rVELrRaObeFdZbrhADFw6VzRgniHxKvAGNfhxQiwU07zgNn+F
5VwWiARQv0k9DazDhvbTj5ZepUa7TayXUwpJckZuTg5M0pq5b5vzReaccStcGKxZ8AZnlMlWmvm0
lW39rJ2GVeR1EnSWOJj6JG0hl54rlVdP6pTUxMvwdyE4QQhgBXb0tvtbNCYKxOFMQ6o87scj5KQA
tIliUon6yVI2X9GsPSa5+D6bburgd/wBSKCgHEO0TVQ6KPZc0CMgPrQzk8MqQyd9I3G4WroNXBze
+9zWgrgR4uqz/J9VXx/GDRGDrH3VmQBSPcPYYrP3H2tV314iwf7Bz2D7BIATm4XTmMDomWJWfKJV
NTs5bGOE9tojHl++iJS0giMRkrPGOLVCqC/JzTG7WY4ZT2r8B/fsxbBSOQtRyip58DBBJVgGdZPI
7C6YZTTaYPc/sS2PI089fxSboc2WxK7Zu9bLV6yN9GoCy7kBwI9yhOfH6AK8LE0R5GZ4+5iGuFEg
XafFIysCccqmzfk4uPsNtjn97U9G9lmWPgxvAj+YOrU02wcHpmEruwYItsYmc7Ra91Mj7l1nXymD
WZuF2QkjECuJq701T80VRXN+oNAqDSbHqCI5q9kBfm5hoKzKelKK4ZSSuSSwlIsc+06SWB9EC2YN
idGHQX/OYC4wy20j+GA5oeeCtpN6DUUXtPup2Uug9SjH0VjjvHM/RwKFlcFkfZxW5ySiioRS5KVe
kHvNTr+jcpUcavyNzNEOBSz0G+0kYLAcOqYcaq0DWj9SiPktnFqHrg0FNy8C8VAjfAttsy4mqrLC
bqIcg+lmJiv2fvtXwJG8OuhywqfedR0tqm8Ap/GInU1uTZcXr+cysQ8c7s1TfSukvkh9b8Sdcl6r
wanj+Kh6nqF/sIdI2m0SZRqT5/B6phurCh25dy1dpLRfR9Pupz0sksq7QWTUFiUKLe8U4RE7RNNH
D4MwByes4HRTygGEwqk3G+NBoxEXD4zibj0oc1d4/WrjGG+rQ9cgDNhRtQy0M+qjYVoal/ez6MFE
uvHrRi7HNefneLNYXug9ZVBrAXYo5gs5+O/OUGUEsFabg8gBMHCaeJ+Ld4yFfpcWscle4cVoNBTh
lhwjtDnGANRJw20VF4AECXLEaCKqOAMDAYaVm6Q4aX6IG5X7Y4lr2QNf9Z+AdQeeaebkpq8ibUpe
BhqF3SKhO0XtAxCf0VMScOKlHci1p8tcVqT5yEJG1spUcB8QKcJ5MB8Fp+GArEwI0TdEBxX1uXVI
tv/M7OtwuWntsCRh2r5bXNgrAnF5a77ri2H2VDgf1hCvQiGYDgFmxyaTJDvTqG48VQyK/VDIK+sx
281VoTFa3LbV+4DDoPWc3mjwe88zWhsr7UWVx86dnUk7QtqYr+t194LrzvBgc6/oZeUTOeZNfAoq
qbbIoDFqAAwdi0tkHVVQ8JoZ3xnJr7D49P+gHnsW7BkMmCm+xSHWqexAX6SNazJwqsdFHbDqSbdo
20JrWwpv0yWp+Hliby21J6wqdyfwGSnt7mRifPyxmaHYTTE+n7PhXGkVWyTwYsTMbX5iuQkuAnRZ
HKTz/R8CP3ZrC+h69o6FFHulOcH5jBxtPqkmPCvgqdq6iRhStqDAtWHkytJ4YR5jBhnnk3mQ0Zpw
l3RTWcQ4iFv8YuRBKTGyT4U/WDX6mq8nkoTXY7mIAAA92ygzb3Il9GPPyQgEgIUeCT6BIN217xso
gWdZfoZk3crm1jHmETzy4nJUfhjsemKD/2wjZADTRdxtiZ/SyllScdQSPy1ts7wzhcvJNbQzunlL
k/Befny9BbrMRsFuxxFO30P/g5CzarjhjM6BThjV8f1Bt/c8D1Pm9rWwlTTrEUx9eYsQYRFV1SNS
nDMBl+3mKHTr+d4nKiwaTAtp6cXJaNovXFRmBo+Kun1rfK3Yjcqd04UJET/qq8nOwL1CL+IT/p4i
wUegXO9C9qGn0yYa91sQH8XanPFHnD7VTQzdG8WgJztsAA9R2p+EmtQ0y6hL25SgwVXcU2gi/Oeq
sLS7ipcmom77xzLZZ5OWoQ6dllp0KrWjUEtApoZm2/Td+hCZp2cKYD5P5Hk/OxXEPTceNUb35WM3
M0ZG/WdZ/nHnT4evyewEie0/96uxA/YsOu/uwVlhP8nXPnBgGL6/glf9OxfSVLxeSdhBPRWsxxpz
uK5nE1H3mCePX858HjNkYCVJpCn17IngugarUKSjj1GUHw7ZMsHO3QWppw81m9D9M3HZoi2zHPH9
p9gYOiQt0YEgO4UrNTTGMG5R8Ym+t800fH7kCopgmHEZ9nxAqikUuMnXUQemjXWMdeV37Zqd1WcL
0uyYjHxTEKidPWFxX6EG0qv8vjZtkdLOE6tpaFnE+IQE6tDC27G2agnxI4Rjz9Gp5wx5cp9Ptudu
xwqy4Zp2M9H18WP47h8GvMHMCNWE4v+vWpdTV+5IvdMSMObYBwklbniKMIO4Mu3TlC2QJG18gjBi
K8r7MpGh7f4ZdecQHO4ulgDeyUuSL6vHuOHFpO6EbXZdWLSZX5FZvpDBkWcsfmO1bZWlsJSl9Q9x
6r1res4/Vp+Fu3QWYM6On8lkDUGajksWMdWHPxkch51S9u1Mn+id2aRyAuo4ayRZwe2OOI1ATUkK
Jto2a7j2VIZNDWWFfl3ZL1uvnseHsMahHSZ7cGzai66HcO9zoPLynd9H4BLxiXfHqvIgVvtxICBD
2R9dyqZ3rhCJLuNyHh45tFtrH5Jf9zRth+81CRS0xzynxYZMTcInZ5eC41Uy8fGAQVen7r0oq+Xg
nesYSd7INyLyGBuK69OMO0DweoJw6KT8+jZF3DvPap986ZGjbyJu998NZKbWOaRrfKMEHOfR286u
8CSIx+mkD+w1i/kKKrBZcISfrmQFX90keYPpOKpB5g07x5bwx/qT3lexFM9uPCnNH3RtrHIu81gR
V2ohFNVMVqP5sn0DjjCCVUP0falmILNG6rEgD6Kj7olpmMjMaLIQQOR4XCREVAiaUSmHCxv2YoHa
4RCeoLeEoO/Vl0GDS4N7CbYEPBkFrWSwQlu4ru+SzxqW2eBpXwqkT1V2d6N6Ej7U1gxb/VNoF5jC
4hpddP5Oz4Vx9ygNUL7t+885WNb6RpubkMR62M8kUJiYQMEBJTM/fSqoJu3qGyp380EC0A1ObQ4P
Gn2/wXwVZJfHRAc0906tHFwuu9sIvkVFGAefkebukZLHFKqyYHJma6oTin02LKLCfHA1R3AxyxHT
qb6huvXB1KeLW4d+FVEmEOeGdAJVr6t+kw93miW4eCZhVxrT6rEQLRHVY5OPI5aSLPPGFsl4pwFf
LCAHGnhebleMY7cvFPIMMuyVRmX9qKY924HEsB6b4pywMWRJ/A62z0vWet/0jvJFEnP+JtQtr6UR
08BbNg2UWw47u/gJ/Eho2QaYgjPekF79H9x1To4rZmsqwn5bNUS3wcTOqgqx9msVK+GO3jUGF7ZZ
UiQG2GK0LWFFZu7ph0j/TwxKxWp4i0jEtfA3/JgGdTVrw4tWpX24O6l/UilPrKTq1IuVdtPSJtwJ
EiT5pXBlJ5yhV5N8cTQlR8YzSY96qa0cuzTlvmmPGln9JpdCjIGnt2asJWAbNXTA9yqNElk0vw4z
e9o7X9yDaRjAKa6WzHmL2HKF2l3q/sbaVxOPHI9o3gdU3187E2p9Isva/OGmCJMeq5AQ4T2sAG0b
IKfS0F4qOn7NQZ4QoesZ2ZTbc+cYO2C82hRyRvNlDLgD8dPWu872qZKH8+o4ygX1UHGbfAQBb1dx
049SvqI7equJFictmp7iPzqsnJ53aGOnwhgb9lnFU9vjU+DeVB1ug8tTkz4NALgEUVnKftT5fDXS
dt3xQhUHXLu6vh0uFePABCvZIM3rKxUEr4FqxVYyYl3avI6mir+8cfRp4lzjy8ic1V9A+q3bFoVr
DvwvwUs8WGlADsY4wSsJLxslQ+ySSYCffHs8+TPNrjW9gv1DsxuS3EGOxxhMGFy9WlcrNeaIwY7W
WzYbMKK41bbvJicIElQV6apHAtSu7yIxwKY3XH6u7pIc5JU2AJwuvnkmTq9X/2/OpkkfILQcCpXF
+V1inU7z3scqM3uwk092K8QPk6WCYbYsBgVh4oTtMI6MRsYppKrNAZkRJGRSUpTM4aVZc7R0NIM8
ZnypmGjf6Sll4rsJDdWIppDFqhWolQs40CcMkOasRTmyZsxcF98/33XxbHXRqsP9CptHU2VkybjU
4NymHMXUZenVMxDgkkke9X0rOr6yJV9hw5hvwDOdmYXSHIJdsTJclFdmccmv0EqxwONoLqBMUwJC
d+ztLoOT4zoK+orwMWqV00BHBE20A3QbzS1sNhGb7CrtCc85/7/hvCXov0Wda/egm9fvVXX42yj8
kaC9nZdQeCovW8YO9CdCoBjg4vmo6SpQOd2yakd01TEGd/iEY8UsNdzyRfKdgpH43ZUH8OA3AkET
Uizw2jnu8wVqJ7t0FSp+9MpAaBdtQ8sjCXPIN5MQ+/HZh4o/AKvWBLDbEHK3m/zL07i/FQeY6/sX
7BOCHf2I5ICB6zge7vpF+mi+fRDUoe9xk46aTXR1f4yWTG7BdKyjiM7ykWQuL+IJSqdrqAaIhgpV
H76VBlMGG2gCka3/Ix+b9moq6o5xtOoVx7XmF9WrTuyExP6aZomHijqSXy5AyN77XqZqRofdJaAD
8CPYQjawlaxCYVa0tcSpUsj4DF4zdGl7US1vCq3GKI0OyrWbAuTdbqEOkiVPnAeTVhEksiw5Uzl1
3kp4vYdLflVdgL18l638M4gKadqWCOfkEtOcDiTl2+nwkmrS0uh5PIrKDrKH7LQogryz6scyIi1G
wIiVwDMcY0Xv/Y2X5no34DkonwHOl0O7A/q/cpGR0VhjbX0ASTY8tSSV1FH6ZGolB1yDWXSEcO7w
FKwlb1ta48xnhi5Tvkp3WaLGa09HMHq7ELXcuGibFnvMEeLR8AFSFBvROhk/GOfm28t9b7/Q9VHj
whMP6rr+I+1YhQyihgFgYgLPE01y10gxeDVuXir9k/wGdaCEuaSBPIo3PNQAanaHUv4odTqYApV8
zZPAquoA1kUFWalH33HvEXSoaD9xeERcnYS+a71Z5snhR0Xxkk9bKacQcN+iJjIGT7yO8QGC52R5
6PnQTZtxdVZs5pVbeuTcUwxVLlv3U3MM6HMDm+YfBjZ5jd8wTkw/gR16vKRPbrWRJuJBUzJe/pqq
f0UkHMmsFYYr3Zavr0ZOnRjLVmAhGTqgcry5Rhl7opglp3j5bIRXUdbM7nScwistsSdOrhMcu7oN
QEBqtm5dneLMMyJBCwdRbu5FBE4bE8LkDSj1Nvl/cnk6Gz4OZZSEMjcUoJkq7m+8cKzavnGE9fXu
/IDyaAqEqIn5PhQNk/AsYUniAZJqcxGhDNhFleCSMpH3sGdGNpxrlOqj8lVX7O0AiZRxOR0pYYFa
DgJT/QcH4uBDfqOhOQ8Tgh+yr/A8YC4ZfygfLWoJ7K5JopnpCA+hTdmUJQ1vEiGadfgtcAiyLejF
ytult0kUi67QKLHglXAQJ+CBBnZ4jbUBYUSfN5hIIC5ZsV9gzrsrtIlVnZPWa2RgmUtPHbz1m0Mt
PxRPImP1LnyTBaY16CFvyQkHHpfkD6coN/qWnKAw/H4WefZwnhkeNpqLNL7CdY7Oy5Y2bvep3JWP
7nebpQ3PgF+2uC2qV6skFV8Ro/FjDfscvGAUqUrcN8Y7vapmgbYgHArGp7eAbg9zhQHrjJdOn7dG
RV9P7stcfPcrDrUQgGpQ/lbgFFX92klV0zaepXHQ9tQNmDPPqZUPsMp/ji5/m42N2Urp5F3IcDj3
asKSH1Fq0NDWKqpwS/IXkCsLaWCOWWDQr5W6lyWFxH/hLTrhRqMNrmg3HRoYo2gS95NPiGcDPmM/
VrSHwF/7ouGul1XYRPf16/ynnOJwBgkwDecHR2UoARzuIUxWj+AJ5cZ9GPoiuKKVmcKQ9+Two0tx
LFkxZzbVyL8jkyY9nEkO3etzZC/GuUxLzg3sfF8cM5FsE7L72QrbzqHeOHiuH4O80Dj2s4fX3Wjx
0TTtO7mP/Ptnml56llRjdLUnkV9ZyJGdDks5IpJ+JrGX8Cf9I/elEcCWfrN/bl9GgzkaV8jtRzX9
QKzgowHLUPUx6QsdSZv2gxSIqBGQRKQ0y3LJTZBpeoJvDkaAfep6N8wVb5eSjpTisYFtTPZR2ybB
kdWm0jaa1VMsSiky1tpuLUvKhylG3lAmXDKY5eSFCVmjUZLwTIQhmmkCd33WW3HxZsb+Sk4ejW2M
bS0UUmug1kncNj88+KChAJuM4FtLFHki2otL36+thUBNUCxJMx4I6kwnbn/uD0G0sF6Om/NEj7EW
7iuK+d7Ja2nFRN1btX3Z5OgzP20coTB1PfcVYT2TUGjknkFMbsKGPad9+O9iCaho4o8EG5P/jssq
GhJDXQ/a+q/vMN3r+8/80keszZSgXmyyz3PrEyJcmPnE+3j5cnRE224lMkBMXcxDtL6DKqlupOD0
rEjQNNZ67e7hCvXVUrU3nUNycRkL1KSLhIoPCtcRJcGzsd84YIPYh3gFyQeCcdu4HBk525Y2vVlL
PLEwuMaAcFqFiweDayF1Owi6LnKxNcF9W7tMTGUUa+wzphNlaHAi9P20VFC+j6GI6oRV6S8p+uAK
gpZ5+XtQSh2NuzNJ8sR/5U7u7E/R8VMRC4mCGpWYle3XY2qWFYfx2tezqTKoP+0UlW6p2T9K//zw
YOf602IrI0d4zvig1+0EmHt10jx2WR7znTy+Uhfoo/aX74uh6WhRBD6kdCw7jVzd0xtmaTAQG/2t
cHiklFHXh2XcXlPdpdr96PXOPObhYWI/nfOgEpuOGaVay9zrjBWsVOqu8VDiByMZuKuYtWsw35xp
1ORJ861e+Jy2H5AMFHkB8xMFch/KOFEKrs9HDaGjsqotL3scVKg3PChyW89ZKEWjW0J5GsNh0Lt6
xzLw0XjJ0SV5Ott4deXfM9j7rs/wGqftoweciu7JCb1AHFPsOZgskkhXfbAPgrsZML9UgzIlcO7W
i4FdJ5a7TwwzS+xFzrDKMhdvPvUugNks21PYw46ZWPo60W59il7KIimlPugu/MUb4oU3kFJQeCLa
0B6BmGyk8ifO6hMttRKYxwGlDARroys+wcOVG4FRvN/7mEq6BKzZG40tgl1sAhcPqvhl5MBH6y6P
1tiaiedb80Xe7q3cnzOrKw0NYGs3/YVwPhpVzzjOEt+nbjVdU7xIuNnoqinojke2BWyaprnUoQ9c
LTWq9SPnS4A3Kj7uJvMBXCQQXtWAHFa69UIlLwMxiS8py0YTJOoCi/ex33q7ae7WL9hytI28QzBi
RIAbTgFiTWlAgxh6HAYlwwjTexwXlmtw4SygUdCy4A/ZQM2a6CYV9hh9lVlSziVnpYdiVxSGh5cp
wOwyMbYxkGwR9O3AEIuQ7d2DXPvhlmj3hbz72ZjFfLBlSBp5oeKBXvnuIyR3bvy909ajze+yereh
dpXfrykGEJOg641X5D1+n8057m2Mj3cIOc740wKOP6WOo6Q4zWe4wqC8L/Zn8KCD5aORHrxzulcD
eFjeWTke2/Av02DIpYtRCqWVx/NQLa3xBsSjFiu4UHf56AAr2q5pITfc9l8Nf74hl26/7O2x9ca+
HUIZWGOH5toezyztZa9Ve9dySnrkxT6sDTWZYpaTeBekL3lhnTSf9n/aWyJYMtMH5q5IYfjkfy21
EXgRjqb4YOKLvEpMm03MNb2gwSl+pC3IX5BO/e/BIzrkKxEADz6vg2IffAuZP/opKw1eQWCLb8FH
oORFAqXTJ4wAwIANHua87HEfYhYA1EoDqjlewERXgEAL4ExfQ1JlXW3lEJwCjgR+fWLGa/y1EHma
3aQrdM9EoMFl8vgfrL4826BYMWieW1RAxTAkgqRYiNrVBqEPV+b9ma4+0Snc2P7hRcVozInZuX84
6TOrzab/PurjF96RqBJ10yv18Fhu9M45Ynem49yc+0yvk1vjHLH2+tJXO6LlPDNIBV5I8DNtzHs5
FttZd6GrwqgOExSWJOLoq+Z0DjdajCBYEAhUiqm4NWttFXuQgsoYXr5uS0eX4teUkzAqe2EmJKnA
sLuPwLZ5B6+vnV0+UD7c2sqiNNZNeq5TaQpktS8wwqwWkPdQLMmpvmzNOfh7KUY/CUg0skMdpzhd
PjeI7oqA1XymkOiHn6L4fBib8Hh0vhAnLFWHPCsHaNozTqMy4zwQUxjHZpwlT+13ni+ZFbBLVXwZ
5Bg/a9OT9tKC0l6izWt4PmaE+MiaAfYG22PBsd4lPA+j0Fxg97fSM6a7go6TWUFrc6OftWSWvCxc
tg+XgIlxcdil8hbf+3Rpdn+ZZT/CZI+lK57LC+ppuqSms8jluMDWtoc3fr3F8VPaIwXk04GmqzrN
Qvyh37Z9ccxLTgNzSsbGd0wnbgqgUADNg/YQPXw8UqNC22ESBApEuAsQIAgnnNzUw+CUTdHYKiJI
hhM9RjMXXcVDfGSzk7WqnQcMF3J3+2JwJTFcngXioNjIH5pGr/NGp9sBfVaoNH4SyFlNnPPOPRV6
o3134DemO3YVbNMdAdq+pWzyHOCfhM6sGe69+t/3kAWdWiS9XvicL/UQK0F9Uk0+vUWCWKqRRuAm
SVu/S2/UDVK5wE2337Stzg9aGfPteEoxi5ikQ6LNV4tdjtRmoKckH8tKNLrLm2ha+9sLiRMcgqSD
GKN/7XRuXbrwsVcpeS7/alzwRdrf7uF1OZFxqzJaBdF9zK7aAFkQPFiNaE2aW2I4P+7k2Fl1dQt7
pKVdDohqFOvnWn7zFNgS2jl2bbQ10hlO6rXPOl4bdOsQ7CQ9Hy0TE/bSK5DFbbNEWX+1at4Ko3dY
NunCtErul6nqUdTPU07KUg25l0rPNSNOwzgg4rtd0P3MSrB45D2ccHx/zhrEkdpbHUiYuZmSpQDJ
Dweg6iH2wrYVoolgh20Rmua3wT8kmmK/1RDzB7IvRiFT9QgiSoSWCDm6CcF5J3LxKkzX2B1Ph7ul
r+/ZBlTre3jfF3sRS08/JhPOHkFMq/CeGUaAbeeZQ1JvgIPun8O5NPP3O0kar44mfyAuOZBNFvMX
/350dt9w2BC32AJim1ZUM+bN0TPC+dxARG6S59i+UV9p/bUzS9CRxyqj3J3t+khRfLV87cwcJzom
nwQNhJflaDTlDImUlnkHBKATHuZbcE+VXO1LuEIRu9syB+TvqHia6Ezb6jFh24oZhbyuGqQk07YI
Z9MLxvENq056PNcvTaT+yrq0oL1G7LOe7BuZmHYxrSp02EYKG9iiYmF+HdFVIxEWkRnofjUzVwY9
C/Y9IZ5Gij7Fl2iEodVsZNz2DGAxc9JPCI23L0VlHWxf2S8yrnzv/71/ZT1gp3PRaP5/AlDc/T8+
G/jZcVorxkyZCV95UbmXAhaDq8cnoTLP4aspHQewJHFt9IDJGECObxnm66s73ctuAhk6L49zXe3p
HflhvSnIS1OUtaX174wGt0nlmfXL9zc1WJ2k2xcP16X7zG2OrxJxIFwZRF22T/Qfp7fy8eLCRReL
Pf5jVALjX9XzMGayuANjXgJPIMTS18Aihp8WYC/8lsap2poO9HzzllJTf5TkmQ3r+ttdRnRfBXze
N7k6q5btmyKSZ/niV5Ly+ETUXLnjmDabYWj3dMR5Xah/31uPfIQ4h0W4vz/12i/jayHPdCdnwXPB
0kizUC+885p/OtH01/MF6PAZO5syRVJH5jCNNYPxIGv7e0hS5bWvTOAVP+mEcxqih0PlOTZ6NJ61
c1LXDtwV27s4sTeNS7UfACJOt+DpZH65IWausIA43VJKtHeiA2OYseqwENdHRtT+MBU4n+/FPXcB
6kv/Tfh8z7ljCK2rraQp7YbIh34NhJDZyN1cnpPEjQdaINHnlsPpMjeqzz0fc/M8f+BLFkroApWh
CpJK5UJsIza6NeZtaOHkzgciIgE3aDShWrfNwH+TxqguMDTlCa8Vb4Kf475MS9xMyjnPGbTslEcW
hLsmx1lWOW2tIhPCw2fvNpXFAPc+aRohk4LkR5mT9GkLz4mq8IjwctHSV1Cv+HcLgD/Z2i+f/MxQ
I656O4SdWdrrN2tn0F3XIwUYPYE87DTZKFXeVnDFMoSLU3S8ZtaCZuaDllISgTL0mqpcGJwdo9qN
eH+9ONZ3LenR8VXoDWE1svFvsoAmsLpqURoqqzakaAFwiJsFt+EF3IbsigJyM1qVLltjrXmONrVF
ncXo49s5ZxYjaTHeOztqkxPBEzPXMf8vGsIGC10qgYOxVSZXN2/ttV3vdTkxTEG8dbVRT5NkXFNG
m+BUyzLT0GyTElTszkCnBqx2aQv8xD8KJ47GLfN+ZoPTXxtZgQMaFwsHgeRXDxUbUmABF+jbpQY9
F0jmAlgieg6caqVWQeJB6XQlEo3iGtjaC3hgkcCt+W7Qp1gwpxO/Tgz5xEpuLtygoEKh7x8Kjsz7
m3fprqpblnT2t4NRmctoG4EW9skzsFlrq4TKGZUmvLzzFNkUh9Gst7H3vdup4HKy5okQJk75XcdR
g3eMEa3ge/nDLWsNFzS3WcRRQGBBLjk0V0WoywE7s3o0T2xDG09W+SCzfMihDMgz2zHfR+0+nr8S
bfFkLCWMksaMdtRApfd7/76BVKnhl9qrzS2kK0x0X3n6umdo+azaSpfThmU+lDI97sKzoVx6eFSC
YyWLNKwOa0DayO+cYO0h/SLpwuRGqLlnB9GMOc7vT8Ox4ZZj8VTnSL5n1OhEjuQPQw+mCT+MkUF0
hsP2BWbef0Evtd6xJ6J4FzIO5bHRFd0dO4aP/AjNfrg2lGWpCjIwhjvv+TVzY0pEMDDtMd6MNqdv
9gxq0CFd03NQVjR5cIKr6Vo1PxGgkVEtqLh2NgXTS7SSP811eySBGobhjsaQyKeoSdcmgMQaGYAz
NGOqufkbRhi4MoJVTFoLssAIAIi7qWOcOp5Y+a68zxiRjoB1SJSXZDttNQoK8LHdAzr2ee0/KA7X
Jleaas+vBhCKSTxf/8cuJsYCwtkAQ6IlGhkHEEGqMrICAAh5IePJflF0mZZIHsUVZcIG1+bx/0c9
4yLyRBIAIqiaV0Y8pw0iTwSNOsNS2aA6Yjyjr9NNPzW58zuhqMT41MVop8oiyK2xiAVHteHbYFWM
cRb3mnFNlOkMG72a9S8MwAp6pZaLt1K7vA7gva3jARn2Qp++G+H+jEutoo6fPSGgFUzpm5acp/wT
C8OY8Xg4RPPZEV5NNCEWrTimotFKrvDwasVFLsXSUa3SUzFTj1Q0enLb2pE/zFbPRpYLvR5oU446
fS/s2T2fu6Enhk288KEQYQa0oBhaEctLliTSIWgvhQqFEjwlQpKgGijGWM3cpYkCoKg5qGLy+TIi
cOVZ2x7MYWaw2QuBG97BFW+oXAke8YVtm8OgnXTalMqw7hPGm+8HfUH5sGFwETVwAnF6r6d0TBX5
B2231UUC9x1veyZuxw3FJV0ss5txloXw5v5ElhoP7dhaJCMOWwFczsww1tuvfl3rQ5R1vmtHqzoT
aWlK2ZWc/bVjNg7F6rkpcs++k0mEVCUU9qwTUG4NuSHqqAdluG9s3kG+XiKDHU5Yy2i7N4ikDc4j
Rzg6j51ZuWXxaTO5nr8Uc3EvI0niSbsJdbvRVLao2hExNgwGmruhWCk31cG44560BKydFsLL5dcq
LSIbar1zNGrTX58UF3r9dxc2r8J1UOXB1xYr50Ow4yYwSn68F4sZL8lBgYLOPVQqamU67xrnvjN4
ZGcVUVWMa1id901a8oSZUW2ZZAE01hzD4qSQauDlbEs2/2EIii9R1y3kaZZ92fx9OJuVhF+QgFJ7
zkmN9oQ0k+9ygDJg3o/hWJYjZtg4Kw85WnbLs4Uj5hA920MGxq4w79RNtoO2AHgThrFhg8DfVSKf
0KACyXOOqoKbTpZPHNOak9DbElpXW9qc1abhIk6NKdwZy65Y1cAU57ECh6/P5QVYUWgX5EHoNOdi
7V1z8GXHiLD9GolNgW788igIgHA9HW6u1FxX4nMg2l7dAKZsBvjFN/b5MDXp6tZP5rF00OiB+syq
P4CAUiW1ucbbUN8V5Wye4IbghV1syDCp1xJT+wSKcA7x5BWBe74MbtVONNyz6ieFB4A7ih6C4Zf+
sGQrc+MtovST0ir66/9bzBtmCFgT7kPyzt0n3xBnMnTfa1gfpoNpSLXsFUbDeAvJI0PWtp1kcXr7
RoaHGLzaXVYwi+MOBIgm5wBWPALFB5vBtB1bmDGIGmHFcgENg88VajyR80baJPHCHFhNsOu/XVeg
+x2Tr4AtQiVp/VkUuGZsyA+DgkVwW+9eDOaOC5mFxxjMaBmgIJOCKXOM+JeWV4kFuiZtfsYAi2hU
ohFiJNNf8IbKI3jv+0KC1BoL1i1/7CLi5PQNlOGVqAQaYuIGnKP39CTFe3VHrxRKR7H9Jiz2Ote/
FMWpiK2urd1sgceaD0ZWt06qBBUq7bD2IuqpoGMWFWyz5JeRlN3YUhwXWkcibYUIXOq+0TlRiI80
c+ep8gcrddnlinyCSKhcRVZnKQlrsTF4+7VghbIVJPtJJFhfnZbD4Gdx/8tgmlfo7W30rvMzIlDd
HCIXTtAiK00Qug8Ftoh3C1Trvpk8YG0fm0N7fVBkQIKtJTJ3xHeuzLaLyioIdSp0aHdqJ4xjOOk5
1D4Wix/24feGWkbfmBVqeR2klKT5O5a7vIf9Hix4+KB64jqm9rib5A01dvCFEIm8kjSHifAlbAxE
YRjvrqHtviYjJwVXjLPoTZb2XCGnan8M0eAeu2zC2EHV1WMK2rk7khN8GxwNIU3xWGNn+f2XBRns
vbids0pes8J30/hKvpradrX+xXQnNcfHiZeYIU69/J6WuUCUkVAKBocYyTzEUlaxXYC1REdImeQ4
CrRU5HRMlLPWJX68RUkVzDo7gkU22SU941J0MyGdlB53964/j40hcQWtx6c35JWjSr9z031ykCEQ
Rdi5Aqoneu7Ro2ClrfPv/Ax/Ca7HpIg7OyHh8Pk4X5YwRTEE1eksUzmPiPF9w/2u8GCGKQj8ZtsG
qYCjkgBA2tm0Ak6Z4waHrnKrt0eFt0e6ugFV9zpLzghln4/EO+s+cYdeGA1cVAxJ0Wq7k7mvbJ+u
HRSS7cDXshDDDFBcL5dN5TEQrX2msw+AyXPI6F13uKTy4R6f1K7FMFmR9xrUukZFX3QpGThoO/Bj
BqJ9fSGrnL5oqhgPoBLd670jnrZ/+whE8IwdOT3Q9L4DI1Z7Uam2+HrD1mEWWrkfKucP53L4RTzO
JsEOw8eomANymvKPXRLJ7GpjFGHrGJmJrShkgKBHQndT3xd5VaDgbqqVSpsFm1W7wMv1lyc+eong
2/StZjCGzKGXyrfcqsobGG2fwP5Go5LzA0HOsN53bxMOsdXydtEpMYY+SRPSJya12IlppcJNFCq0
K9FzHmJLMLK1zeTVAcZFqBZ696x+ZMaoJrlD2R9Mil42qFYggxZV0rjwJRVlv1ZRBvpUOYoTU6bw
3nCgpLTIEs7bbxfvw0oNc29dHPCWzCib/o3v+0f4QA9OF3gNsmQxBZZ7oKD4lpf69+EJRhZZyzRX
ndkTAWC2BZdtpsAaeRED8BSrw+H1q+WoGO6S5LT+A/OZKXSzbZiogArEAl/8c2ivNhHDchhI4Dey
WEADwXlkvmfISXv050CQgx5dS8HyBRoEmESjPcth1lTvXT5nEs7tsXoAvSr2PYXNzYpNeq61vs8w
7UZTmlkVYewVPUDYKIsE+jfV9yDEj7qGG+fkX4v0dR/T1syeRSporGYNBOTiT65h0m6FtDi4aUTr
Sd5+kn8gRiZHrsUE0Qf5kI+OYSrlzBgyMcij5uLo5JIIBAmnbjONWs+xZ1gcT0kUa/e43eEaDA/L
bEPvVOKcp9pDytsoOTrBewsidsL5VSBwj271R4P8b6ms4QygllmeU5eT+YcuLk9PbAlarciTbKhm
VGtp8wrfTt0QUbYKM5wjCrVXOddnXZ75lGOuCsTADCAhinrerDgm1f7TZrWTYkV/X/VFUsAEKIHw
Gtk0FUfrD8UUie8ZmK8oxjdaktw8kocogP/VUFnKWg5KKVtIhnflqx77U39w0F5MgFP7hPBZIQMs
hUhajfM6yT4KPzc3CxfilY5hVhLZY08nTFW6Rj+kHfLeRsNDtBlFd2wXNHqnQsAhICHIhjGehbC/
hc/A3bk8FrRW6me0hSKx7FP91Ayx8LqV5XLUbMQOCkMQ1iWBVwy3DkrFbt/GjOyPnjgciDBLvoZS
fvPn82xXYN5W5jFTJy9xt62C8Au6pUmYSnFbetEEx0vLCPYecven4akXr589I8yz+CBDH/IhrdEf
j3ggbx+9OSCvq9m+cv0Uc0OvFcQDtrLSpCk6i/h3I4yJjfMGwyW+cpTaISiZkJcebhjJuqnxpcJN
PQaRqi/+xhP8lNj/RRCVrzV4MKM5VakCOnM0IblDU7mZ+onbJVg7kIeYVm3OLeCO8IhBYM0/CSw4
NzSS2sacSWBgX+A1k0aR/PLDmS/t5lu40FFOoE+nKtPziybwakpOkWUBfwb3hG/rE37etoRGGaE0
dN+R5AtQMwDYt7NJlzt5hsDkkYSQ2vxdDzyNuJ30A7zxqM4XKOJHRWdY4nsYcAwiZvmnwkKhHEq7
ppIv4pYaDM9XBHkaj+GO9JPCpw9s4HHKR2IaVuI+TGxSTflFLvcJuY2b5A6nvj3khWzmOMruZwcZ
nvqE+C/PV5D2H8qnuhTULjMiPu4W4i7KCLu46b5HYwzrrX4APMf4MxvGqhLzy3QTtN8Rwlv17y33
x7BTtNbHAUgu6cDKG9iE5peHi3uYBJ2eCrtfx2+9U/X/OpbTGFkFdM9AV4kaXDbKEVUB9XSzp8VZ
GNsSnVqqiDOwCSkPj76hY9v3yjtpGqIRYP03r01X+tfnMFeix1TOyNMt7DMY1JuPFBA30qWTq8E7
mibqOaNR6A4pOV9lrscpULslhf4qIN+4Uw22lwAmwregI/MiLcgBrMWIkmiLvQZ8TQMiC6RTfmTD
OrSYlzAyA07gfLshimfjAjsCrjr23INtGtY8ievRelTCmRao1N3VXaAPoz6NyzZVSqpzrpt2c7W8
/7dncDlc26wE2Ggifyb0FnbYO0VeScO3eDv/OqG7NBaxeyBk835XZy0LLD+ePpbyIpYvOL+cz65/
IX4UvTc1/p40W8bZ7uWct9pgYvzWzTpnDg0M3OAP4O+zmrg5hEhrRVCswkisvlpHM1WLZtadRHqC
4GBPN6QAfqYyurnJiznqrk3olS/bnUsT4haDnV+gptedw6Uw+Oj3xwNduHXmoje77QzjlZY21ETf
QLDLJyx5F3tcvytMseoxQSgINinZQbAU6sOe/NXajGxDq0agB/QkUbiq+7DsP4QXw2O6m86RIKzt
4OiJRdCzqsL99nWpZzp3HrGM6BqTCjQG83cRl+UpdI9CqjLJOfFyiG/xlCp+OEFMXaVHHAZ7hGur
5bEHu2a95EckXsGj+mGhEhg0TvEbKIx2/c4TE3H03vb2EHb+nEvqQawcSG1KtUx4ZeDUcKTI28S4
8hLUlJ7eFw1OLz4T7LV5osdy6Pj+UyYJ+X2XEMjsCdBF3xqe30nM2TopkM2TvdIfk39lQFjPYcfP
JKM1UudCI6tWQW8Ppx5wHRP2TkdyCKc7zsBewMp3GxeJLEkQoC/AQe/2bZCYBsA7oCOwnNlmnjo2
e7Bohv658zqqrwXoaLanbkkc+fn5bBvQ6wP06wshjSUYHSmNIc0F/oxH186cTIjy5OPNve3MxaLm
AYFni7lfgOl0tV/TEr2PPSL9FHp73+4DZYiyBpOGfoh63Lv+rBpXQICvc9ZHvACdvRUmItIL/lq+
QzzjyaYvT28RWNS1mTOrQ6mqjDEmqNq50mdvN+Ny6LpScX/IQ4DjKH0VTHUh8Ek6Z8VOiKZkA9Rk
eBTRrQMvUiNSRcwcqKHfFZLWUBkJi/6gNIO9JhpMEZaZUUXzoFetcgviuiwUmESFdG+Yi4dLvTOI
j10YqCogzkCZEVrkbKlbQGZ+vAW0OIifMXRlgACBAYkCe+MKi4wAzC5UTYalm71JMRDMUrMG2tTD
/YvpH/IrtMBO5lSCsdudbq7fuF9dBUOA2b1hc+4bPJD8p5lMxRCXRGOSmKYbaowCTJtBzgXZhZHy
Ke/7frMfzE4YvXmKeOFf1Ksw+thISvI54O+/IyoGs5BSYLuLCSQkn2ocCP1rYpawG5AD00SUTbnH
mFMMILgXqzu2UKlTHSwN0B0M9gDi9FMApguUrHTlvnZN+Pl2rUiRHR86MCLJjNuFhPsyy7Bo2p47
diM1ZNjh0nlVEXG+/tH3acqa14Vmg1Rmxe3FWTpyvRn9akUt1QSfiVR7muLoXoL7Nr9rNtc3T8gZ
UFiZ9GizdV2QX/OYop/wKqzpSzQgK7glWGZpEiKh0TE7R9aFzef0+LQZP736BSM1BYwnazfjfTF6
BY80qjcsboMDtcfuInBQEr4Qj0mfpd2yEuW99DQkqZBkPku6D58JEfvVTQfL6MrfBI1IoKbSteMK
jX3H+o8ayGl05r2SRc9tpZGkc8awFuEea1UN0Esc5zDkSrMdBsWmhQ14LE6hzP4WHP9rXaWHwK1d
1v81ttHmjix3caFBUElWElGwyOCAYws+B2tMqgdsK/Ib5/7O6p+0uoZQWKk3T0L/Jb/WEHBMox8o
9u+awTRRrQwsbA8q/ENBDCCqnD2xBflmNMZrak+spwKQl6UALe7zmhhcyheNhHlZtTDW/ACfxSpz
RwAXQDqOS/xlDDfnk+FYPGOEPjSeT6UCfkz8rQC+0gm1tphta1D/czijVHPv3/+JOfFoKOhVNTCp
QU0kPQnrFVxnm+4vbgXEy+9FU7Xxf1Uo8sV0zcG2/gtR3RTB1qtPk0sUPMddm1vaeOoPX9bIJoGf
y5DWEgDVrV+uC+jW5anL+bm93IEyBiMU/nr6mAtmnyt6nobgoIFuflTkxG8kCFypQjUBWMsxeh1K
mgxxdS9dulmloZhjEtELIjA4WZtk94JzVxGKIPCSiLEdUqjdnqG61kkXYECTY54kYF3UnygBslzl
bZB54L+/N+UGY5M7xq5hqPJ61asyXeDdZarZabwHVoLuL+qReuJS0NDihBw++3POh90EvN8+HSIa
OxeZ2exN7ptJ0QpEn5LA24iRwAuqWbqv1aBZ/Zr3PKVtfrcvB+6g518eMToi9NoSh4Qn0horGNjf
55orHiT/j691UJkOgUDKFcPvz35shOLbsi1GTGNHbE2MBnKn+elt51+lSbTEgoQz2Jk7bOB/90Zw
Gv6U/7qbZ/NK3B2n6UJFvjAcjlCpoWkw6VXN4c1JYkiqNUPi2QaMnLNLO0q0gHo3rY2hXQZCNA8j
5CZPSmAWCLVbV4n2t/2r2/9CBeoOR/gfNRUnL1DrLzYgMIvl7lPAa/IYhssO+JeU4e0wVpkbPXnX
K3M57aTMj93ypKcvgktFpnjwY9B0QgN26gLWG+7UBJ278Gwa6rM6Od33XSeYxPRxs+kP8ZUXxOQ7
WzTArPBuVQqt39nVboO+NA/TBuIp1Z1AaCkJl+fuJw1+jdy9VZSXIa75uuqPmXB1jEz2WzQd35MS
wOK52/TAsjdlwfShtdKkT3AQwAOGiYGOc89l3YEJwlPV6O+NaOlMYvIjDtjHizg3YgL2M1aMhpN8
CR4ONsSxp97f5x+7IkeCl32b7egmN3VzXbn3blkKLELCX2O4vOYeT+ZzsLLwHdYskwjztlgQURsw
Edgap8yFiK5KjaMx/4t5Ry4aPrsQavKZM2gSURpd4jDdoj80rBLJ9bpu91Kbuaj5EjRRQgAet3eI
KWdm/Ezf87PLYe+4BMxCxqRQyXSq7kFTDT+HuDTo8UmakFaWPpsQm0rDzzODygHbviAvzDV7m6xv
dJIFZtf0iCrMOAJAKt2yZOmojNneqM9Cdarto5dRxO1RSwo6CF/zY+Vjgl79xxj45DxmnWNQOHmz
XGIcjIeGP4kPKFHEa4Xht888xfjLfIthLUmqXgnbOwlr3JLLVGzXAThwMNXpE9MBFnte3B1lTjGQ
bcokaUZiEAO4iC8wMuMA+nOoGqxzmaZEB/T3kqp7y+YtJdYJgYxkXHF42uVti5n6MIu5YDmu0t77
TrygbVm/Hkvq6eThairDNU1WuzZ5Nms6yP/IKwjde+pqYtCkvmJj2WO74mfGahmOFIPwIAMqfkz2
edL9VbLNqhhEqifkLdE19h0DES5mJ7gy2ukvDE22s106IX9a25rN+Ux54nrPWxa4nEcJyOgRwIkq
7ei2c/Tg1OpOYBLTjrbGf/Z+wPQUtr0t5YiGk3XwWRaJ5psV6jXiaROZ3lWcdxUTz2hkH753GFqK
HkP4D8qJu5v1jhyTD3CudhUXnWjuwPCpc4QNWuE2NeJpAs8ZXmm0/+UmBzV8lxWB5EFTxLbN9mIf
MXM29lFf8oy8QRCVOWClxpxR/CVv6wzv8FecxSgFGg6589r8TNIOZYJe+vSKBvbOv76xJlXOrrsm
Tulu/90FTd8woFYc9kTvt/izdGe7JZcvo//8JLCwjrZbVWWNkjUjFUy8kZIVHtd3Xcy+fzGxiA41
s0rFFhz8Ve8SyKVsXkyjTf1hI6zqQ+dZnBiKuowoIzI4v6iumVtA63UTI5DYekuiK2VV8IozyNAt
nambfJ8m4yivwv48+JWPOEcfWd9cca6/iUaDtKxgsKYaxUQDHU2jPuHh0EFt7H2yy9uAwiVDs5fk
PXhMBauCfSo9v4ha9aPVsvzmQM+RaxVZlrknBkVeOhZkFV901smZn5HU69UB+xA6AtbX39mTI10V
o5Ldnmthtbo/Ga78FyFjWvng/6okWYVqYpzGxleOHptbceyY9mtgF9Xo9sm0h7o8Sfns2kf/Adzy
jxBlDVFBP8k+WpX5fPLYkXyj1Xbwrfevd4kKgIXKmFMt+OMMSSAFo1d7bQDZdEkR7EqHupeFSFvu
NUliX9HEFnl5BhO+vKzH4CQEzGNxoFYh/oCrP3zzUxESKE0zdciAxvHfF8JwQKBHWXT8imrmxvXa
SXMKfD7cABrlqPH4uYSyunSH6Kig4nmeskwozExNvbRXRMTdgzE/RiIawcHyUctV5uqF1N4QHmNF
vmyBvCHNdybJzYcA7kxuYUtaxocNLCSCvRjUBJtz0XZoJolYNbtF5OQRJmb0w0m590NzlrKj5A+K
G4SsY4KvUem/w7XF7c2hK+neH2536z5DYLLQRTarVNYsqY6l72CwsXZUV3dDYHExHQ/yY3QDLg6/
7D5+AExLgt+Ysuf92WVnCke585GkzeZjxksiPYF93LXRGts0tRDHn437Bpi9FL3bZdPAoPMExz6w
9pMF+n5AGLo7ttHYC0apdhu6ukNgzZiANyd+HC5McHGSV+OVQBsQByNlSqkrh0jBNgD2XM0ocZas
8FfpHM7xIw2XlWtBLXMHyCcAQlr3fNqaIPgoZP1eWT2O6sEqaKtB4RVQm3Can+Amy3G3OkxqpCSB
fC0uptA8GQca0a6yyq3ww1JIlY3bvFQ3B2b3fp9ZXtgRMmXEyOd7aM9vNRBqBCCWdL4ofmVqZM30
j0xKZ+93g5ixomeOy57lwWcfTcmhuW+sy07wOAKQ4fzWawMWrCeDGKXR2meHllHO+t33x/+0t1Ms
t6jxtBOD+FnK+9i9cQMWXcQn5itJ74GfIZK/2kwjper4twqkeZ076+hwBfVZX+2RUe2GSN4jMXvO
G7wztmkSs6ec2M4tT6HJ2cx0nZElndqTVq393rtYcoaj29qyT47oCJlcVCIXNE0t4ZJS61mmdHOO
l6ecRWYuWcNNht3bIvQKWs1ltn+sbdWstZPy0nQDb/sMSyBQbMDk86ts6vGHNe69ewC/HQdVo1Ob
iBiBeNSIr+mEQ/k8dGDJo6rz0Q++RrIXXc/uUXdu5yKNLWeUJ3/KYeKVuXL39M+qSoym5upUnvs3
GPN/urADCHkUiIYdB2OKKs4czOuVD9h96H7YOTieNoRRSGoQyXiXZs8IMoFhUJRBBbmpMmE0bR2J
QRSTEZ/GdgImgrHQYifHnCU95uQoNyCYg3W0cBoyd1OSJt3/0Jc6NPE0wrgSqijYDaYjDeFbCOiN
zerB0DSxttEqO9AmN+yzbgapSOFJ3x1I8vBmaBVF5ymTkPLUNlPlG67Bi9S9THl7SinQuuxypEI0
IFbWCAsSQR3xaPhM5NAUOtyAn2VdcP72l/qFS/+RhUqLtHzjZKaLxlQJGKeqtuYSFU6ILIWRlHcl
cY/48oQyA2ERkxZYT0OS+bS9+hSRsQK1P981wf8hRjqHSad0Dz0VwippgI3aNOa/EpdeEMVdPPgl
lO5jufV2fBOj2p2tFHdFUzDom97rP/f1S2Umyze+nMPt10h5nMbqMVFbXuZHJ8NmsnNep1FWB6VX
3TbRM61NKQXFmuBDemIpPolZFMM9uxleowFzeUt75fLhCYaF2Gcbo9nlJsTmM7Zte69ahfQzWb6A
52LxnLGwtxORj/ljChToDdNlRvI2J+eu8OtKf7f9m3AMLe0vnGOrckJ5JLv7Gm3cbniRW38LFqFB
WofB4fxXVZVsLNmjyG50kWQpvcfsUSlcRTjXIAhu8bQSIAgab44Onil7YjKL/cq0UbAA3ED2va6A
I0Y9QOWsArdvpRKthekc1XK66yjSEWfKOdMmvYvVAVxD9AV2xED+W37c4NNm6vVB47lybdW68W52
hx52FjF6HvgnNmpNb/WtzECH+ITevkf/KUYxu1ci/Ee5lfc7nyRcp7JTjWMltehJL9toJ9FlTiKg
SPWHz0w8a+wWsIUqyCl8JDowu50GjmIGlOrlcDioCgFRplC1EzHZPUEySTZsWY9pjJH4pnIbJJqm
qce/sOgHnjMCOft5cdRe3hw9WMitO02CQdUcApAV9P6OzbXoKaGwY31ujnieSq7oddnRQcH87nTR
/EZuUUznDmZ1Kdn5RF5xthQHYO2uAErQYNm90vMgumMZh6G47wgNH6zOyhlOvZNrUg+7gQMZ7OPd
V9EeVeWwycuJ0JgBE3zTMCcuw7uh/aQ1C5ALpIIEq11olkCctzTSKsOJLn4GLc6XR/a7f2ufOP0h
gFHkqlK3DNCMuT3b54ewTYAv95D5+EfpIhEhe/ug/VrWDGFodHXDivzDTFosghoSfohEOTSx6Ygk
rPHThOq9JB6fhz8gHcghVLv8ObFf+dWOoGbheiuDBVJKuk4JPi18J6fDQkf2ASslmSmPS88Ibus3
0uhF0vIE0WUeZbzCM+FyL9co5bWZyfrCqTkeDxrv5spCFDJYqY+DOU4YX7HW+6PKlrpRBBgFU4P0
qVlZDXGgJclXi+BsqXAr+GhZ/K/Tj15noLqisq2Hz0gyOstxoAsZlb6fRWzOjtudlnrZLkVZ7dvM
mUCKz7lcGDC/qqgKuUKhtyYqhFV157sZWrdGvZjABIAiVa1E837EZepOrZas2wdGSv8HUm+l0dKN
WkcQoOqNteQmZiMvfY8iIOHgGcuTcxhILGwwgANA9bgqNDTTjMLmRXltmEjjINKt5E+aQFoUjze5
qc0exQtZCS7kkhmVLI2e9pQwtIa8gDthtjxf/ADy589S2F0bFNXKrWO8H6A58XAGwxf9vurnLDcM
xPN+4DCxKUJocoYptZmuPJWPbBk49D+658QTH7IyrIBgEiLLyRCnYiEsnwrislm4Q/sg9T+CD/gA
QHgxWBqey9smCeEVBzBmla3RQm36m1PMWUYP/oW+cWXdu93vNd61Twygk2v2MdVhVkb1dTiFDNuL
0qPwoP9HuuNvxMC/6ey2a2YcXscRQn7UBMJEiSJ0kNEql1jbQmEQ72c+S9ChvX+e77L3RotYIrvm
Ao9mU9eZ1j9bXo4jBAh+8ZGCaVsuv+M9WxvLxjWzh0s5DVI4nCBsGq6NhakOQuGq0QMOwMgLyAVp
49OGPT+YyIqrHr1vk2vTN8C4ieYD0VJRMjetqJN27/blm1sIJEcRnMQQeYRr70OHWS+J/4QSWH7r
bfBzIkIpdWQ5WXV/1NYb6qiooiEQQzK4DrUb5V0yS8vX7O1uJC/QbvLg7DJkWGv+ao+6rZibdgH4
3B1oFHWybOmoMtIFD48GeYH7ecxWCb6O10T1vsSeHtcGDWf+Rz9pRbBQqnhlpv+MUavcOOK+iNaT
pDDCzth5f7dIrH1XmS0iZLFAwlHTcPxxA04jVoy9Zk5JVRi2UTWKb8JMtBr2aK/EbH0kedVPgq4O
v0WYGqYZD+X7hOrgiIMasZgDRbUn3gFxcNVmSkF2+hxNck2kwPVZRWtifD7hGzZALmJY2aZb5sht
nASu75YSwcggHLW44yE1G6iBD6EXq/DXAbC+DzdLaOfVRBhpfn38oEmtdyuhzpyW2myPmKrz/o7l
jMbwBvrzAi2dmj9DQ/nUUy7A3P/9lArPy00hkOA1oRvAFhPxSW3v92mLytfs52mBQXB9aj+eeN0d
FSPZJlRqJfTfmhGGcRCBGb0oYtaAjDj35FJScejhlAkXfe9RK8msCYBt8xdGile1iBpxGOxXZdft
9Liz2kpravD8Z8+CV5NjXABR9hVs+e9saA8Hn0Ra68XNCTYXyTB97d7i1nPGI4nESI+5UklPur2Q
IgTEnKoAboC4IbZofmsQ5lA2WXQlBcmlf8KoUobS8FurwfJJCTJOjejHt3ofuIs7QWGDT8tREwuO
M5iiIOggECYMlofe6XCskrbMIBWlV/meEahvShG86VaIxD1kW5B6VM6I6CRTrkTaDwr989/E6g4X
TTFzcGs/Uw5h4HQONVSYdp8MQwHjp9+b+9nAnkgGCGAc9ZuxvP45fE6PVhfUfB17SCrJ10Z3uBSu
oOuMMoTsBFpuGiPMK1hv6lIK24NMVJFa0ojkrc2VcuU72q3SYLiQvDOktenRaKaTH7mQnZDB5BQG
NURqsIeBmY5NqU96Zns9MjDxDGmmRo0qq6olVOHZmEzJQd/3eWicX2ElUIR9xDuqx26likn1AHhy
11hhOk6t0yedmIJK+J6+yEOy7tgJLVxZXK4CHcgaD+a5EWMe2B0jhwcMm/eLDazDyZY8SFBRBlJZ
1DVdh0ccBWuTo7g3tzub+MMMBeuZPBUAjF1PxA+mwHYCiKKH6iQH7TEFtjNiaYCn5PfEpIk02MFf
y79buiW7uNnP/3r7YooPd0xZUhehJ+EwPAb0HFIuIUiXMjFJYvQh5z3QlsXHIBDnyPvykhhT2H9b
nDfpCFPVVwZoNj0c+N6WdFIhk6hs4n76cO+8AFf1lzf+BeWt3+7RNhLIFns8r5nKnc6FwaJy0L0r
wFHEOKW9sC1Cn9ZzympESAV2r/bjnDWdhAPWFJRDFAyZEYJqWw2WIozGOrxBa4pBPU+2A2fQ83/8
eCyzw/BjXB26RAn3j9hByLSQuWNRSkRbnmyuENFCKoEQWenPYWORusCHBV8ZNfDRX09umlXEZvkt
vOSwNeead7eOuU/ZvGULqplH1Sn4LGKG7GUQWXt+8IchgDdTpbYixPVhOMr7TvmkprNGGxIp2yRA
icrC75Uf3pNC9ikhNpy8S2UbtA99XqDePIlHN4vPxP6cbSORaQS1awWNn4AX3+6si8RnliIiuyIQ
8oIlMBXqCJ57xEAGBltp6VnAz5OuXIXbc2BafFkGIkYUdr8XR00pYw+NlCnsjFYmRaFLJuTdlznp
mMY2yV4ObMvNrWggKBQpr9jpC+MSH3l8xfua6TrbRdyAyfjAQLREPQsp8qCeR/eXP9bJatqE/hDX
IjJAbJeJ9/PPXJvGKZC0KNXDgr7ZNRHcOhVaKEFZ9tEmRc9uFh3Kvey7eQyvK875fmEHA8gQCsE2
ZjTqJLa2fD1qaOs2Sqs8MLQmpHXF5ARQVfrl2I+VKT1FZO6PIXEzuHvdnhJPYQUK/7wl8irDpt7N
wibE71qs1b5hCvP2x8AKUfLyvokL5VUt2Wchgn7j75DfOS/owCo4xWDvoOZt7UGRR2pjaDpU06q0
R2+N58fBMOW7BAhAMxB+b4vVHuyNSD30y7Ku0Wtgj93t+JMCosq0WrKjlJZq6OaRqVC1doHNtHkI
WT58aFHr8GjCN1O8eMaYdyIpggohD4GuZwqndOF3Tmx/xQoQqmsleNmN4kMyQ5iwZvFa4Ib87l3z
vOEbfD16Y99UQj5xkgb+yqbx6auEzTrklCmKC7DwTdpsmPLXT+Yp7iAQw0pZsEV1sUMCtQDMJkGo
XXeYbsj7H/wNmPgEn82uD1JW+YtDty1M2AYRWA486v8VoW1wajlfLrghBlswzmMEToMLJRuzd46d
GvGCScLAHgbgIXiGjReTrZxmflbDUEts2vCsi9YB+6WimsCSTFCLMpVlnNF0I57vyl0seEZ0Dm2d
TRJ5YgrEX9atTgXSr9jATy/mnmGq6hrSkDKnYhcAh1wnGP1nsecp/+PHrkZpdTcAy8jUzRaB6Qsb
1kN94eh79SK0zQiGdWTfQd34TuINhkRUwnmK6hbqVazXVlPQ3Cksc/uWFU+0ZdvwtzOM6gLqGpqP
gpb80FHIzSTR5moIp3Rpv5lbFuZQteIUFc49mDA3BaRXitsdf0ZNnm4WWdaeEtzCfo22dFpNaxjz
VxHhbb6rRTLCuxqcYc8gXXloOv770Nv8azDGy5hj0wiilcI9dBlM+oNxuW5l9gYhXJCm8xzSr+PL
NjJpuONoPBTD/E539s4pkAHHMGSB/Jtg+0VhR8F/bqTyNwCjiQGbvZqwT5iP3PfLn40bYuerSxz6
bqZRTO9snnxCqoBAmN2jYXDdL60qgqQmHE1QsvHJj4dpyFLn6AbDQ7ZSyg8lL5Sh6a6t1hG/s/TR
hSQ/S095flJysKmnN7w1k+ZyqVr8ZBltOEPoye7izgmu3ETjdyKFjYs8T4D6w5aYEGq9QwHh+PFC
HysyTayz95cAdu4fzqSWbZGjZmdMr30bKnuvCiYMkPh4Z4zIqzgX3pDaE2r1XZ6fo4MQorCQFkOU
z6cfR27jmhvWUo4Q9mwty0GS8a4qlNFEfKI0cUhMslO1sW3wAlKCol0xPgcmtxTpauq8CZlJAERG
tG89vxPLton4kKeI+we7zx2Hu6DtdXYs1u5Em2JHpuTlLs94JS38HvVZaIJCbUCRhTctUrZuqsR7
B7EyjCfVLbpTZUO4n/NzeMMkM/9nXhWl4Z/XOTLpG6En9HXr6GuBBJE/FNTFPCva2nkhokGwyrPL
BkWbqauY2wrCj27h++vDtcceLKI7NprOjeP+ndywOkP3e4ULpnQrW0v5BJcZ/ftwaRnDtvQpPWJ+
geMOpUEwN3LyPjoc7yhaj81Es06EgvCOWVJMlVJOJhADSyDlgohUgfYfwBw3fgvlfxPO9HmMn3gm
c41BkUDuH0pmFTdo7k2QzxV0oKdo08+1rzDvyR2n7C1Q+ZLkPNMIzl/O91vG+KCjr4XSaZscPIRx
mvcxpQus1UVR5RuY33cwNyrgtYlXgON1Tl4RHADm+jtwYdeO7U604kPVBmqzpuG5USCsctFNBv2M
lNDEZmj6FF+MZPDFBXk1+E//whmW6NtOcnDkf1vUMR00Q3O0i1bOk4LouqqfdQLuC5HA/BjBE9+2
csWZlwVLfgpRktd4rFrC+ZqK63hyt32d4qdT95YwQm0l3ZYXbykhVIOiQlL7qzMmbgmVT+QRGMHA
+Tj1dnIPIsmyxYvlbMRTS+Gc5UZFu3wvIljOdFaSXHXVfFpBXkGlHC2uhSDOVMx3Ep+YCs9cv8ho
OScx8XkiFDEu+cxGFKIbixmad1eqzLdOeywnD30jJ72Grtd9Z4Wjg5aznGhlaaNlbI229UgLTw8x
/XYM+cBPPng83Cim6gji9Bg39ZHmh1xalT8yfAj2pbGyaanmG9zeQikkjGMQ4OC1k8NHkKQLLDBx
e1rMDP8MK9Qx+yG7tvNKuBryjZ5hwxyDZNOWm65568pQCeVNHaPQRCIUC+xJfntM9vsHxaFdF5WJ
Z7xKdRi1gM9Lz734P4+Qdbn2AMcg1kxDkxD5TKcMbwFyluxn+kJgsQX9mWOIKiEHphacpNIBPwUS
Zm017Xl+/C5Zeb07H2uzi/bMj3oThP/4+BDf60gg4vmick59+EP4um+dRI5n6c6ZcZEfq2KxVmkS
A5Zu4wFeTNNOV5odFYGFklMzuA0g5WYpeWYUp+dvUHHOtV6S8ANkEWQKypkejcavzgZ2k+nMFNBP
y0z6G/mIBfrK3b+2qPXQS2nADZX1vWi7CD9n7Yjk8DREg4WldkXJQmMHfZ8ziwgExLwzKSL+VUjS
sGaN7sRxYFbuYmbWkU4m6/lkueBP3IY0XZ1OBVJv1blPmMmJUNbCfIkEYv0mA3k2y+xLga/7monr
Ds7RD6J1ixfkqPGotbwg+tw2w5nllQ/GqkxcROVS7e0m4ezsvbuyUYs3acknuc7qhtbAOhRZysKo
Qqq4SX/VJc27rxHcnkgmNwPhLU3EknykxeBaURMfpvHbg0g/SbzoMvJx+7Yo4h+K9nWlzkeG/AIv
wDbSyKtwgJf9WngXwYFfybLMIWwsFrEaG8uOLE1xQYAj+juz7tCLnRHhmax/XCHVR7ev1vg92z9f
bMmUURDxn4emN/jYSGPra2W/eyes6+NTqSD3cXwHuUcQpOO5LeqzLoyq4I1EtQPf9q5nRIk+Qyo3
lFk25kYh1WdzHLICUcB2RK9Zn0g/b0+KbbVx48mfMPuMCawnPjMHc8UWh2C/aZdCiaSuxQTBuQPQ
zf6hWJDxiFxlpd3NW11T2NfMEX2mNOTCdk4VXDv3HxdPK6Wvlsa1gyQZSpmXIyQWUpNfi+6XBAsp
V212kpXNKseLxwQWABSCgcpVowrqqb5k7sYI6OtUwvJrQdF/7ZDfsbx2C7Qo77yMk80Np1LO5j5f
7yq8JuQzqysnOzSSuc/9ET/EsyhNPN5us2TCnbAr85/NBqOW3z6CKD6j4ApfZ/cFHVyFaJykIgnh
Wi9gH136T22B9+ina+GEtfrywF6SMXR7c6VszpV8ALRLQBVMKWpSkK/7mKh3ndGqYZ0NxcsZpQop
TcmxEAOB4sGS3fnDBN9uoePShRhfOndd246jtUc0mKXvGwkkXq0LjWW/IZH3z12TkjbNKAL+Dl0h
FDQsu0DPTieBjlh+eZw61fwBMD9G27jD649y4PDEKL9j1Og18uUFt/EU1d1FgtylsZreGbRRA3yp
qwWq2DRquU5dE9v+tJCvpw48d7gtTnWJx+yw/i0Gje36KP8lItMcaEMpCugvL/roBp+m+dDpnWv7
WGJ4Gv5pxUcRLo5NrP6Il9OYl8P/XS0VAryLNNE/6lsJTFs6VHiYGd2uB5eKyjITkSmA3R2jyN9t
5oeef64tfP8mkmwSmVOC8gFUkd3T4CSudyeUbmeFBbjndx7UEp3fokS4puA7w1BDbp4+PaCO5UE4
3XfmAut+24/zDutgsU1mik/W18oOTUMrM+tupt84V9m9tLUBg3rgW9KY843NXalvATy30iqPL6to
GX0iIvUhhFquihMGGRLXDhwhH7ZGA7a+Qo9v0ew3DydybmqXB3rNF6ozXujw/9pNBs95c5NQes1c
GAQ8LNBNAXKdBaX9Bywo6PYWZScdwQPl8TvuJDDGJLTSKgfrBFsLkCIlgpxNGwkuw9Oc8Mf8my5m
wZQFnVJmvoA/69d0UuVj7FSyP3L8ebm7L8NtcUTjowC55bvaqJxnBKQ08bfSmutTyOh6viiajtrD
v75C2GH+RLjwL4sx1RexI8OUMgXkBLN4beYstaMCbMvumxCn7HFCy5LaoXQdWwLgbSd3H676KThT
TgI8YE1SMmr8/H+w9CMD93EICa/q/w32meqc2gYfVwNXM6y2FTWBuhDliEWd+j5PrimNvKOVNIjz
0cyJUFS1ZDjlBqjYm8zAL4QDOblIWO1m6ktlr0Z//TWVxDhLXB5T4Owa3lfvemcvkSHiYkRrz7N7
2T7LAf/gW2Ss6OLSX6Ur6BPSKWqRYgagY3dubi8+TnadTGsLwyCSvUyzirl/Hf1zRYZtEJglf45W
5q1IzAiJUJ+mN1oW+rh1uPlnGhExOV+6VGN6+vC0tIuXX9qA/2mAtHzEZtnqsMto/a+5F1Y2vpsb
IlSq0HcjQBhTSEphhIVsE42hc8IOUsDnakGRKByesAOFndWzGqr2w4Sb52QG7xktcjopzi8tBJnP
OMxAQ9ZIdZ9p5as+e9NYRsA9Zinr0sqJQiqIdrM1jq5PBOlihN3EPlmnqtx/4/vOCW3olTCTQ0H1
nTRpS0buFE9XIZOeQG783iQAk5rJhxs5IbHRgQgUpkFCTgUTLW9iQpVNBezXBM34erctJa9bh2Xc
jsBPI32BlS+xVycphSSR6te/yEceuj4VUo+ddbDcHva61knahd20rkNGND5J9XPfGUbYos2OFHHe
AX52x/Is1j0oeweLAvW/5rtIa0yf9l0IHbvtXj8w3xoeZJFJaqxMGQgOM/ECijS7fbZOJpKQ8j4j
fhoOqsDWy83cdRryItcdMhbnZpBvv/L1Rlm2gT1a/+VmnTWoz8E3YIASyb2Ed8dhjW3RLzwkNAZJ
YCMCh50Z8Qx/cdeIeAPeI/ZjAZ5TK/qLskvoqjbUGMrc2duT9hcYR6UnjJ+dnQ4BzXupTV3ky1V2
YguMJSd9wGhEu4U0QdbXjjQeOmr2U7cbt+29aS047zhyOZb00f9nwZn/yU7Vq8epWwIcTSx5/bwa
9tFWlrNZaXEWjDwIhdaa+V1xXtAfkKbFzX7Sfb9mHMrZMy5qocHGUqgtmxTwNz0dXGJqHI2rEnU6
hkzcaIuFTE2J1m9zotadGdI2PsOh6WIbaEp+yvwz7v7mvsPsyoAsh3aDURn9IRLUZqYTnmyJdKrJ
wK7x/TFBUfKg3CEE6gE7T5D/3L0Ass2FA37/7wNmR4wKWeLOoRcZN5fpGA++Tj2te+zJdnYm9Bjw
Lo7wO9vszGnCq3FekJF5BsZzaEm7p+hEavYKtMSMoY9oqsHBE8d8pvPrsPfLjl/6LUuluFYsdbSs
DQ9WzqqcH9h6NyG1lU3gurqzPgI56z6g+rMQL+DBJfvJFMDcd3teOjQGYVKBdYirlS1ekNqt44Ca
+G6zl9q6cBe2CgZs1mjHfomCfu9Fw1zMUIOgry9OUr2/pnZBLp3KippB6zIFFSlrDIgBPrc/lVHI
ASwtHfnGrsmLiisP5DGAmFqpcwqhjHwsAjeiVj8q5xhwHV2tbpo7d9Z9Wh9xAQxXU1LOguRmmlSD
4xEsK37wMvlNKi9a0nUEWNMfCo6F3h7SUVTYasiu6QCnU1qYgPgvOEaWcefX/sJqjKBUHjF9BGtV
KhFBH+/Zsq+clm3j2W7rg0kRNlnCzbpnwu/OWwhHKGmRQ0qI0A3KtIt4Kj11sY3j9t8u+nYddxW7
NY51cE0pQmqGxDvOvLyxP6lU5cMZPrL+UhJ7Y/jffhDzHIosMTgTOggL8DC8zPjexg3CVX264Npq
xehVThq7ItC+hJmh2m9oBDwtZsDEMfKghcDSCtQrum/uJc22+3TVl7VvZUlwKE0KL0F8+jVjS3Df
AKEprZBUGCGir4sNlZaQFEwZ3uF/egaRCOJO3fuG6izYQwNNRn5Do0Mj7oyRPU7sgYzYf+o9TcEi
B3AgNnJepajPXcvBCf6SvqBDtR9MXBP4gkgLBEtuyd3crva0fJJYteTC8+j1b1dC8xju/uAzxGoj
O8tETU4IVHT6WKlA8qmWVC/9DMObiQpbqf1awYKmL2WyljqdZ8VOYd7Luzs+HjQ3fSncDFEB/ar9
R1jT0MYrlMpt0f3CgJxxsBpKhnY3S8sAWD3n5XIApb4IzqmuraTOO+KXw5QnCop3vjLC181vs72A
1Dtg2N/Dn5CkWH5bvwS2vHjzU9CQ79nePC0G8M87SYwo2cToiP6GalBnmOECqZY56Wyvg3uPuCZx
PguwLmSHpkRBxT4jNwcHNkHFRAdUsUjtZqk5FntcOa6belNeuLZ1enWEYk1Q6I9zWpK+Tfh4XkD9
ztKoNOt6fsNS0Qu2JE+nsf3hgoIItCcH8Qw5X4AIf8dp2SpOQU782BxF0JCqQGiSJv60ryHh2QVJ
bxMkk18Oomel/F5mBBuqiM+T/iFDBt0bXZtwidBhy7cwDw6e99H0MbJZEYO0ijUZJrxtHMgN8pHp
cc70gp9LI9Q5g744/yq1CF6lLrw5VppxNE5pwb6A8u5IAXtdD9AEFz6vIstbG6b3sAIi8YKu5iaW
ATPaYpvBeBQdi+yqzK7qsCIdt7vnmk8JSy9b6FsNBTrqnW8JWs9jiunv6vls0YLuH/AKHfFBPDms
sezDmYs+q2PD4eQpHFm6yVsay6Lk12MHFMoKXaGVXfSR4qiLLBkegncby4ccV7Vh+GMvl30I0K7H
ZvWjCQC+CygeHovgQtqOMBsPTXCD4vddY/4HhsAAEjD2Xq+8IE4F7Mnuc3jROv4ng0CtRegZrern
S7fXsRweiOT+kNgcuG0bPxciOxRB+2yqElDONDY9JIjf+y2ZzEImKDXsfnSHukKZfMwL6ksPt5ks
Iwg/XQDQBvSNdcg9WLBXFsBHL0xs+xTtE5Cr2leBcmcbMMQIeeIoo54CKuoY/JFOpfodbVySCZFj
/mHGF/XKXxn3e2zIzrkqZ7xm59+cLxA8Czxv4QZDozq1nKvsqUH3H3CKKrwZzKKaowEQE/iILwrx
cLewkVaEAooxhtaACMzUVnTiHL471CjYppSwy3ImJDiuOw4ZNWDbKSn8NBVy+U3HwiUz6fJD0Ooo
2eTn/t94+XGyLKb76syeMpw/LxUwioLxBfi/InpFXdnWZN42m72LLElEe3vzSm/lbv4UNoZyUBKD
2ANjnJwpqQFs/cgVHfK4vy48TGQIcCXAhjVY6qgmHJXEKysXOP5Rd0TZVG/lDlNmLa5Yjyx58vdB
VRq/zbTbYHb1CsNNdlCRgtbL+NfBFTosXIeMlW13FSgIHr7dPaECIQn73s6GJACW4fIzoMPPpuGd
k5TdN0O3cPa0iLl0pQhLcSjlOISz+dV9XOEWZUFd1YLc1FLOIVavOaIJcDgU10Omec/rNEd1djwu
UqATQGMD2dqZx1vpzwWMO0KJPhyglYsBGdheSu6w/TifDZdooIf8S1j5V/V0Y6KrnwhLDY4rWjca
HjHQIQ4+9MkS+uUXquvhvN/Y/hTYhEK2pxfz6EqI7VO+PYiY0ftH2/882PtgRqdLqfPbD9TmcC1D
QTizFPIspbs3+NbIrbpbw98xxtJslwAT9r6TWzMjzoJNV7WH4c1J7XEdMs46ikI6W8cUchTR9bKy
X4T8c4n2aEqkPCUvA3KrYmkaepTE329kSyQndXy6EniOXLH+2Q1QsK+bAkmUAU2e21koXkBIy7+Q
rLx6gd1Wj0c3bjWZz9meE5YsqMoF0BQjPBgWww6+/Prayz1hdHxq8130qBSpszKsSpNehDZHkesi
gqbzAb9XLvKrP531diDX9VP8vZ9qio+GsWgHtzbbwoXXNm4sRvxysqJrEu/PALGHbQbN53lqhLzw
1TMpILIfGhgDbYUPlmLQlhvrXIssJJDRurVRtjiwi+K1Ba7GJM1uWH/wLzZeSgrRMygYstfHAvF/
oD2aBMYi00zKEeLhgr510DXbAa4Yk+Xve96goj1KG/n9Y+1kwXW4hGckkfDfMQt9A2NZ06Xmuebc
yKFl81vCz+Gfo9YvrjIYhLJJ8tlnCxtgaEl6zDAxWguUKSTCwTVL6w0n5EIgCewVEXg7OxUTZ+ai
D80sL+60XR0c+EFPkfRTeXilbwnFQTlD7mR+VJDE75ZnFsZOTx4GVKaMYFmjbt8QYioNPLQhoDaA
jbF7pM/lK734SO0Hbpf/kD5hyUjaQIOcBL+gmp+Q1BpbsZCA1yvchm9V66uqXZEl4vCXL0faACz8
YzIXNuMqJslsiIhOLYhpRcklu7j4zKPA3EB9Eh2urTlcF9l8XiKKeHqVDNsfXQlUSMIO0TqDBHxK
B2Kh0lkSlshVewfslEJoQfGVe+q5GfsboFC29QA0r0T4hvTAG3doHRniz8kSkSofvwOdaFyWV/0c
tHZ2HbgpeBx9B+NVrbkaLxrWy0k7asjiG7eewylLpru2h6Qg8fk8jqdM4ZPCuSTDKV4L+aPqR9CR
ZKUm+a04c0xZxVom+VdHx2muQrmyUAeyIAJGViZCaLOG8d6xJGmO8+2s1S+KpAq4dI7Qh5lEeDmi
sRLn3RTGhSPrVFVX23RxPXaPVWfld+kB4ujAwj6sTfbrmZ+hPadBWLpBYWJ3MPbjATdUEZS7afac
EnMcSqq5gfvxCxpRq+FomzgMT7m8oPj3FQU/zbQBJdN7GQX3o4zlaGk34R1FJNtNRG5eni2p9J57
bvcTjFc0EYz5miXsJykZkWmLh2VuCkaVX86vBFCGlD1RAFNQuBtefl+0nt7IMvTrVrURDq2Ly13J
U6xs6ZTfOjDg0ZJz6YGsKTiN1rd8lEBkX3qzsY2JZuA1goo5ClUZBw7x+Y0XnHJorxoEzUsRSvS8
aD5txUGOJI1OjPu/Hj2b+DSUeen3LP1LNOepSm4TRyGY/FHMpQ2y6GSDqSKD/rjOYiYIbNn4IbW7
GDVn19hdd+RIZkL6An4M1s/em14ao68YkBFEkjALTyR3yz/Bzfshxr01MROAbUoo2EQ5B2MrsSrU
PM6E6jSn62cNvDaBGZ3Kw13PDbLfjPBvJDV8JCbSmNJ7fJgdqXyHFnRTLbEJlr3kKTU8BX+F6wmr
/x4rf3wrztGbwmXTsgcyu/b7JslTNYTnZb1DCK90+Qga9mBa9yKEnLlxVyTkqW8hnGJFl46tr0Po
xe4/fZotfLi2wWWn01Xp36i9rxsm27wzf09h6YqW5+gf7R8RXlWUF1HyjIdEYGh30pAQvsUjOxIM
ytv59eqkRg8KO6dL5dCCg+mEOMdilzQVEoJ/1WWOSW3TNH157MtqrC2Q6y1Rgzs665oSnerx9FF5
k68HOEpjOrZp273tPkN6VW0TpVkuIYgWKv7lf7a7grTdweepoe6C9hvd3XOk6QAwXxw5uR1z8SV+
t+u7oaLh5tuDtcrDawIdy4H7uHHRAJF9Oft0NMdsMm8sfzf+D3ipdAnc/pQ/sto+VSnSdVY2pBIi
pbBh6mboPfY4lHV57ZS9Gu5uWToz3WUEiJfs7iYfgg42hxVj7EZpsDEi5+bQch44zwXZABunkYbK
hAJyyyVStgMPZbaFL/lMcvZrKB7xaOnd8DWqvt3Rplms7bS5obWHhB+l+7+zt5VRUnJNflOTEMPO
qCdEECyWH53SYpbrfcjOomrl+tthhbCKYYydo0OUV4tKSTPxCtqww17lmif+mc3yAux0FrqFTMdJ
WeOCu5l/Gw9eFRoc11bl8LQXs8ZfrCx1bP3ZyjNrkP4y/7hPcbcZl4oGF1s81FUbwFrvhWVGXjrS
h5ELLmVtpBjt88na/9r+/2Z8xG8nwHNaNkTxyMHxZ9l5wk5TbXe8EUUfvgD/4kpA24V6HnY5KRkA
E+T2/0mocq4jrtLnFj/NHewHItshSDKfa1AUGPGF8En8DOVn76YOvM4V+W1ajRrVSVdJVkwcksW8
jOTyaP26J1v70rcLqGI9EzGTn9npthFWBfcweajkj6wrg52CfqtbIR/bq8mRDhR5rnx8tbYAunqe
/Og9VU2o3Oc4V0HzpehGXH3iziiQ6JA+ru0gGM73v4/9Qig8Ji8z+1n9f7p005CVfPqoMVhrUPPA
rE1okzpRoB0Z1x+u3ygyDIxWeoWqev5ZwXiSUVGtjRwSL1/13zCFkxQNK6HJ0Fjtk8lFi2H4BlSU
B5nLa2HD4RO4FVevkp+bJZjKQdmZb8K0aqvta5IsyQjJStYBir2TcHeVtoMmI1W0bXZbEZziiHqO
Du/1+/HkkCzrmLsCXePfKMgQNLjOrTjejvd/KL7MK7dhTFgwn5CdG5ncqslhbQWbm0IqO8JCS+NT
ZyfKbVqp0fDrVLeo9AZb3tx15vtGHnWDX8ooNkRUXW122HFrQ/S/0nlLAMkdK/qzvisVFmG4fiFO
Ma/2NJT0+TGGNCzkNfhs7JlisrM5Dp2hYKWHhDI6Tgi2cOeyJxBLKGVj8jKcaQpOyKr5Zn4qpymT
6Y7NL+1lv5XrqRUOC2QCMhB+UHGiCE0kXX7vh5rlwzEHRv337SRBhlOK4sMdnsH85x7XaGWTVGc9
PELi5Eg3VOsILBIwUFvGxZtdHEJtSba7rH+skMWiPDAdaSNcSdmRHM9fj3ht9azlt9DowgOtLZrH
JcnIzt9i1olU/XP06DZLVYzIRBb8RfMvWF4BIdmzzcsGn0+vx6f/vbGHbmCn6zt2HwsjUe0d+4+S
oH6pBRcRU3ICyUqABQGJFAUb7ol3+Fyz+3xvkdKHsjylqpYsH33l5DOXcUxCCrvOU8zJ4QBTdf/s
oDFXUgmhqv8UfzGUCJFoPgBwRLALcFbteSgTJuacPOf9t3ckGgWK3aFEdMar2ciHxHdhxH+QFqTV
8SYy9Jk5mLSKyiRKOml2SmzwFqrIGrZcShdAXhkixzHGRX3ikzzvgNBvJUCZjgfEFXii8IFgIZQu
Hr7gpKxm9LD+1XV9Lo+uDsLg1KPZZqSCqfD45TAgjyKi3tRhuE9fkC11yvUNnL1b51cTQA0YDOra
x0OIw8TFQs7bvKeKSFUjpZUQhIJKT6MgMa/e+UqDhYzvG3SlYOOSxTLRPUXJSeXJydLsawOuZV6z
99JPabEa7st92Hl+R2nJJOsNjTcuZ/7CXjR9LB6Dnu4ZypVMpnnhWX7JBN0due7wT+mdmg1JXw0B
JS0qox0CeFFBS4K4fQtqPu3qXruIPfj8yYyZdiIZrnFLMY4cyT5MW+4pvQgP2knMRBVcmeBqkMtO
ZEQB0CERHXctoiL97d6qEM7djm4MfE1BaCWlDgj/L6454sflLVg4YzSo+r/eQOHaP1z8tZdU5nqu
83dHNfRJParXMQzncHMkn3TQ6RVPnDzQxN9YwllY9tQdaJpPkjAhPfc/i7gfORarO4zdMjklo7Iq
XAvWdulNcgW3wzheDVbfPIKBWjh8KQjsegEqnnoaoXTNtqnRXLY26Cwni4Nh4DzuKjfGJtUnoBIc
pYoAnTyWG7rfnAhPt0shTOkoBArv504nbuB2Rmry5qIKFdKtr1nGXHZ68+uo21FOeCoBFb0Tkyp9
nPNHhlMP2PYmbwC6QkzqeHjmPKHCHjcLRHO0OBAlEhyn/ycxe4FYbLgmzjzte3EAZjVICMVA+wWO
Xcj3eaAcfcsY4WJn97Gst/4Gx9eaZGbKk1H8KdP4nuOzmDqAi10se7K/0Rgnc4ClJsbfJoJDwTde
oXRO0lFLEvNdDXaKieZ+u5OshxOw2a9UEONIH81Z1QHx+6dthRs4Op5iKjn6IknWoNXHBHINaF4e
9ZwtVbgzwIa0OXLMzAKf5FLV2ZDnuWu7LLSdg8DX6I/KyVsTwWRRkOS+QChMIwdNA1AwgwPPecB9
HClgYoOzrVYR/VbC8bZGXeAXy83DsjXlcNnWp4P+ZxrNI0G7u1hwlCoq+Rx6ufgQN5QLMsMVHTit
mi78rGezCA2lMhwqzPLsgqy+3j2Sx8vfJAcmpL68wnKDlW/ZCMwtNAzQtwG3rgU7dlrA+vqR8L3u
HrLdPigdmxP1oyznBhmWENCO6QK1/rKPUV/I4ibagedMR+xwhBv3Ys1FYir0DroLJcKrysRZLTAj
Y77CznZcMXcE/mPMVTiTBU+dYdSo5or9uZqvCIw9ylMtUzO3PRp9T+NeNACJ0wIZBZg6Kn5apSUt
LfqgW1ExsH8raS2jv1i2j2icvg9UIdEtgxvZj4fQYW/l3OXm1W3WQXH+7UMeFY6YN7/yk0VH25Vg
Nei+tzkfHIgVCleFpjK7xXfTmdK5laPTn0uxe5/h4VIEmDYiHcNPXpqSkPaIgogSxbPzKyY5YZjC
bNdCa2XbJy6so6qc9gPfHkHIWWZ01lwPeC8sSV8o29dg4yPZ2M7Ww96uPP2AA7o/gtyLkBUrG4ql
wEILhvTds5MTp2YDAa5AI100fv5S8can63zW7x7xHJr1CjipYRhYaX17KH5yqthip40mfydDS/xZ
zk6e0bqLzaY8OPAxPgkIimQwKbooRL5JDZriEOz5w17CVBYsPizm4HKumKObLfx/LJghQlOok6kg
3BF3K2FhP3Atf8emKPA8ottr/ixjqhuH3sKpCaNKqbbQw8UnhPrmhsovx9hot7L+jYXJyDmUQawd
hB/MEuD0yPFy4BlawM2AdGquKxdU9q52BPOWnjF5cTiYWZpmqgs2pB/pN4MIkTM6iOcO1m5rJepU
uDkZ4zkQ7hK/OqDdfm6dzIBiqzi+h4sWsFvsrylAkB9adDitXDdHhfeWfi6N9kpW5WyVN7QpWfJk
8axE/EwjXIATlE7pgqncp9z6clXC32FrllU8kM9Is37eZyRdmtZjdsZXt1h0o4Jnlk+mXjn5l8kf
PIvj3PO8TfI1PO89WbhjfnAWwFojrmtR1Z6tYHAAhoiyRzsse0wiBO9tZPhn9Q/A8RVJNXk7MiGP
HHtLCmKiQJC1HEnATsD/54I3JLBfe2pxfMieMP6EWU5d0adMhE+qBE5yAHuvvboMW8HZkwDR6/Qw
FPe9+JAk9uKR4reeFlgo92/V4P0gAV/kxjUR+uoDwwtJC69ylS8Ya4V7iyKmjYJNPxTXU4wJOGhg
aoSxCIaOHThaIX+PoedAee9mi7UFas0zy16RAmkvGzT4NUOBYJnt1AlXqDzwaBczfLt8gS6L1nH+
O1W0k+GGRkWB7aQFy190Na8GWi3ZcJFFRgme0QMhaxdI12+nsjbztTbJDb/4M/jEPNEkvLQ6Nn04
vfKXzEb3BF85MvzET+ElCzQpcBLhKQUZutcq7IvBNOAuXTYpyYI3ypIxbWX46V/b+TopOvd+aAND
IcZCnDF/TFG53b2By2nU29CHodYD6w1lVnpx69l8MUK0zwQyiZLyx8sDMOREbgDJqKBUaHUrDiJ6
kn2JJQT/rwoSWU6wI/OeRrfePp7gi69z8aEEexWLPNqySZLQGRTh+XR8eHhTCXwCFOIyHHPyg/Se
NlMpRZTQgVfHKe0K8+WXuqMMgLJmLs5rlKtU7ZQu8QqSs4J2W+EqFfWKrObG+8uuTlH38vFmtUo1
oCzWj6r8r7ZlvQN8Q+V9z+zAAWjdSBPolXKdRFiIDp/X3BhkOh3v2X39NsrCnqDuS4V/fahtCxGG
Qm2exAGVZzLaIRCtV94bA5MUSQYMuh61DCl1WPa3H+1NLGhy2AcGOPStPhCQ9xAh+wYAPf9OZofk
AG18R3y+A7TTAParqU15URo2lGZ9eezyPv4XFymFBUwjDWP+F1dqyiYj8/G1xOd/Cvz/saeWkelO
aYezgD3pmNVDTqxuGKuWs4GsRHg90DfZRrT6QYC3j9X6Rm0Yiim+5zjIu8p3iDdUldLCoBYjdzh1
O8YoHcV6E/6odYdkgK8Ni5yXU1Dt0uZ8T9GG3pgaLTzDjdbhUGxXFyADtNDRe3OCUXK7jCZZjrZ6
uij+ORi3kcwrHd0UN67kKAHYtTA13hbOb7c7SESSFZhqjr+tHHXJrm7C/e1GLa+tWGT7cxaAmmIF
ru8DYjv1hnMdPwdvAiTfUrFUlSOUA1HVH8YGbi7BAA91hv3IiodbiJLOL8QrNXspAQ+WBwAcTqdD
BHHDd0haRVa6/i/kUzUjRWFOTbYc6b7H+JY623VnWwrN5lMNcLtusZFpqzJj+sYmHKfHySTkW2Nv
rg4a9HuuIZHTWCe7GL51mYgMYjD+IDQREh6xdbqvhG4Es9931164FhKh9IEQzjLQYWW+xS//VHPy
J9/HwnT2LuGJY1a1sF+XWKeOQ4tK+rZSCvg4IS7DlhOJPVEwfDo9V8LsKq77wQjV4V8fgj6J5gKx
z8eTvQg8+2O11duLMt3s+WwwnWkVhsHfoeqMztvIMuIIbpgcfAdJpsbFB9YrhA6RQZHgW7Br+K2Y
hhcl+cjjPdrr7xxyZDhQfnpWGpuiSuPsnXY7CAEUVWobsunaP5rrGXX9gbv0pGirAgo12XO8E/Bm
uMO5MLwkIrffevp/ov68ZqjJgw9aXJ5V/+3w9mPcmrPYRu8HoKlLQKfXd8mYKQyd0AON3kYmnVMh
yDZQ8ujS0kb3mijlCz4NazyFbycT179zjaIL4YJbqE1nEPfbY1muQ5KNhAbpstpAy4WfdVcz26Vv
wO9UR6opZZzcKvA9WVJ4Gd5OUiStV1GiiUi6IilYgucMZyAQkAuviqcniQ2BACF4H/XojHfrkBdt
N01xaOW8sEGwm/6NjYVy1PgG3Oyuqvy+a6BnCtUoKiVG+Cdj9/sKS5SCT8gwZk/ZqoZYkn0gbsaO
fitC0aIUmOP3sONvQC1wwbrfacrND2cuodAh4IDyfxmXrpAnq8fFsP/bQ+O7KkMuk+E5Xpnp5I7B
kiOTg5uXJko83eJhOCkOkdtb/aKCDqBvuFopXj5pJJCVOxPHuC7J8JpAU8008pe/i6f+/o9Wq6KX
G3sy797aA/M71sveIKE0kH1BlB2b+magwcx1z+HaePnismn8uUOHCrF6MSBU3rAeLgEOKqeuY5nD
NSw+XGH7fLwmaeOsxQ/xV3Yrmm7tRvUz/yUVayQZGbHbo+A+mCWRm67qXzb4HuySW8bAvKo7DI2w
J60xG4w6zhvevA1BMMDjRxuvDtkURGDOU4dZkPr1IVpXWEmczwpWDhQhUg/zs4heiC95BDykPqn6
ICeYuDiOOqQi1IF88JI8aW0M8llDVKcnFr+Jt0mW7hsqDPUzrwzjfEnZ6iNpHkfacSFuGl5/Q8RI
5FTWkaCJ2yj681jAjnEjl5YfeLOUF61mU5wV9XVCsKfgSslNhUKFwtIQfATZV5mvh04wttvS12uk
obu+W+/cLFebeRfIzdW+wf1lEp4cLd7+5qLBsbYTWeUEpQK9VYJ7EWAagN88DWK2JCfmWI+n06Ic
b5+aHrHvgEVMw5yhXGaoYL5i9cWUIPcVP6IOG6Gm7Fc+7hM7wT3gq4SaxBwonql7DIO+gG5o/oKo
ndSp/mdEpx85tFONXxNUBvGdtTuIlYce3nlnYsubYRmr1xZY7ez8aE0dZCROZ4MPMSaAeKjYu2pv
TQ024YMKx8CFfz6KGk71XvydwcQItd2aTlIi0hnF0J93U+4znJ0C+V6FKfamrc4AiI2IHlvxiWS6
JVtoisY9nBiF6kS6s6mr1QgzRluMDW43otwknIruTI/wXXZmLTgfltybK8yQpt7Y+FkJHwPZWpLK
bAql6aZMujr0xxavZxo2UgCH4G1MbMOVDYYnqs5IdX/B177X0U5OolJIY9/ZkEuGzc34YtQdMHPt
5eqhvGnCnWVLziWLvGTJ+Qg8QI2vs69jOs7MxR4Igjrm32gZ2xB4iYmyEvUMMzK0ypaZG8xBz0l/
LMzsuu6Naq9syZ2Q6JMPSZA/+hpm4MrDJLWYL8n3D6UMroGCGBx81oq3BYJewqnX1wGSVKEFq/6i
2Vh+5LCdpwgfgwgfFf8/e4RXhL8tRZKw6DQKLDXTMxzlH/QjmUb+kWUDInLVZeUCPlro8EGQPOf/
dlQPMZYE9CGiQlh9mSRvGg0BSpa+/jUqTilGRKs5KDN9eyfBGYOvnC0Yl1zFYmJb7tQaSIxLOkFu
RDuM66eNlSV3PlfcX/0F0CHpR0JKBXp1FCrYRrdLXt+HdhP433T4ukLxuDMcStHAnQD8Uc2SNBcg
nMnw4d65DMd1KXUsuIttIj18vSW3XopOMfsbo42QyJwIUL28qcqrMsGOP5VJnyFVVYzM7jSWH2J7
kjRWljkgz/7hZZU0sgC4Nk/+AnfHa9QF/424QVbr2sMTlRKfnZuVzeHIgDDTeGfFU5OkfOVvN499
D/TgBF52CUAqbz8V6099u6d2LMWAKfI+wDKFjctUeoMekdJTNfdCv3CFkWZT/U4ZefM6dFy54QZR
AOoEoz1/0CVfECQIqxxl3uSbjGqzbS5gN4AQMvcVe9e3zZqPpU3tN8yW7Dc81BVxIW/f6nWrCxwj
vqNS3TDCREif/bGcyB6/ffP2C5C3wswuRY1XO/ehrkynhPEPyKhTwuiEDSOC3siJBrxfR0wnpaBJ
71g5yCkx1PJkZd+cK/J1LUhO1A2fZR+WEnE9qNVtiCFnyMAKoKqcqE6D2x/5xc46nZdOC+atVAqp
2rQUCIYHiV+SYxd0RKNGqL+m5dH4h8L8vxw3TPW2wyhpy1WCQuccg3pbJxCfpEgVf9NjGOnnd05T
9OcqKwWuq+0MPLhvAFgrF47v7B33spczyM64uIdGrXnC6PSrjBUj/brfwn1binxGa8vvoAvLPx1f
INZkChHgSdB8BcxMV9mv2cubz07cQ2qEwYoM0tbM3HsH1+I+p8bMsja1JscAMOlZulPK4ZZkANPL
N6d+Tk49ZzT6/B+kNwsSQ1NUw7kF7o6vsmajl8Vsnmu9zxUTLi+MHJgjoyS75bZvUN1PPzWtLN8r
F6ZX7FWsSkdQjkFMqtCyqiMl9uALT8Xgnog3X8zzgk45e/K/nZYl5lOJ6NQId771UF2gIWJMBuwF
hC+79NlCwfSfYVpMoxdIQTQMl1vndIUpkhhZUqkybLGon/dIlLfCdSCQFbd7J2Fl1w/4o/nomRcS
5fZNGHD5QrpXAH7JjIaDsrvwvz+nYE12iLdQsrYzBKkWgDMGWsRBx6QC1UthjNlmk8YXvQvK4YDr
TxKH59s6DObwE+UdfL8OoZYJf1OQRGoMGzoilS9DAIRwRQNRsJbxH7ogQYczz0ri8q6zE27yop/3
hSdTB16mLCXg7xiZsaS1bfQhxAmruA2mCrHX1xKqxkiifkuLxzzUx27M/P2J9bn+BgsULpklg/iP
4tv44lWo5ddxfDh7m12X9XeR8ShPVGNIoYfhw2FN3G4UDihEAheNFX+tw8uMimda5ogUd/aborCm
KXfE5sTomaBCbrh15KlOJWN69bp/zMD/NnJNrSs3jn64QR1rnuxS+KSW8O45YUNRN17RjG2EQL4e
YUxVXZZJoipj4IPy5shKFdgRYtSCjStUP/30AtJMAfft6rgsIisQZ4jbRgX2y9kV0OP2y5E0m355
NKeYGfnpU7BNfDBupj1tZxrv6hnU6wwokhotxPR/AYFQ/wsXaW2n8e4Ro7SwMwOdeS2ZtiTRuRlA
558nHDoWG0KAyOHkjGC/cS8AY0OyuHCpcxEA5SKT+kOFPDXTMCHDq84iD73i0M3KUMm8en0ZdCA4
XWdu16n88IFjRHKUVuX+Ki+3IZ6OxgkYVNZ1SMDCv2bN9XWqLNzuHQY0A6PJ6GAheqTlulDlX7e1
OB4JO2hD4u43gciooFsPkGpPFRszPride7Opye3cP9sY4uHW4AISwpJY4TcT2TXnQ0wYz4px8hxL
Q3+k55cbAbI/Ym6K2iXU+Mm9Z7sf0WzMbnWVWumVoeToPkEEKFBT7kDFEU08eH46NORy1dOTb40D
pL3lImUkDLmSkmKt+d2nf/ZCoTZeBHwhaDWMBV6RM9IITUVpBzEBWLJLqO0LlKA9U3voIZe2DBYV
zrIUcel61wiFMBiJvz0m2UQmQf7Cfo3vDZjzTQo6tu/xNZt0BT3hju7JhhyCpJ8NazPrJAvi+/wS
L1NMOixD5Oe8aX5xqXTB6+FVOLq0BOJfuOc2+e6B8h4oUNfc/tEFTfQExCIBWSRsyapcLZrhmoum
1bABikeC+sDrsPQQUngzO16grv2MAha3JksO42l7DCh5moP4D4Rqj54lKz6+cTtttR5O5gQlwC8n
hMJDKLMxAGPJYTrVS9QPmqWqwyE4Up3FYPQWJOtOYpSs46a0TesGZQaSgVJP0I1VDeO5GRCUz5WD
qDDgAkJdxHH9lEC59FVGZ3gamZLOaG6pGcJkdWIpFCTjf8qnZNzzF037MuEVqWY8ME8u1woWybip
vmnojcMeu8Jm8VxlgeidQ0IYSMUba2uw08F9mH/RyUhiOGjRe8vFGjAsU97n/ltQuSqqMkHjc6W2
tcxehXbFK+iO34vyVKacf3dqJIC8Fnq9qqooPMPzqFdbUYQceX3JZ2GFO5lskgaIoEZf68mH8iNQ
LPC9s+LfrPJH0dCgk2K3u/H4QOWugbXr0mPvOc2SVijFeMir42nWbMwUHxlgUeMNS/nwPjP9BXO0
LVoM6K8cNFV4YuvoZxBbURYRZ0xWGX4I8NgaPakjlv1ymnOylbmAKX57lgqtir1PqfB8qc5fkkzR
CrHD5FkfJWqB2LUOLc4uGxl10bvQVchgMNyuA/MTjcmo+iXC9KqrfrIl1Cx0Lknjl/5Row0/WUQ6
JEzEebdbnvPUalGrQ7QsVGbViu7UEw0s/m9LDtloc/lPkGKDHv7PRVJrkCmxzLcoqXCk3gNdFi7c
AWRFJIN2z1fzGWcQHcploJmtzOFevoSbhPpdB+cjdiwXXHUVzlMKzJMyIl3goAyyNegsZW/AMgCx
ZYJqJBA0VqppBKVMGzJ++lcEVK73q5k56rQdtP69P92e4HKXkF7BZZmoejhy/F5dS0/JA+oQpJa4
5eI+RpU2PRwKs78X/HLyrYOXdlxEn3jN0LrJuF/tOeYmPHeei65xYLIViKxyJutEUwreyl6/p6vj
pyk6xuHaaqL0Nm2tmkpm2jA8jcjnoOGIxi0gRtvYUdwKWitAoLi9+PcwWJLwxSGUrzamS9FTIFrJ
9jSMNBgg2t9jeFwNzgGnkdyTACuRhujK0V/f4s2ft//QOewDGOwfL2SzBSzf5Jyh3N7JFIwamgAG
Un7RyOXAiRlmvonEfv6Q3abuwMX9Sz0KunADJxNc1qnhTxwpSG85CoLz8K2pPJvI4D4nfHlvCBPT
7jV7BgFBPVjmEiFZVQkPs8D57Inn+aWf7w3Bgq3ZwKefIlasgjqJvnDUje17v6zERf330NB+kH66
xtQHPUTEtUKsy2N8KCC0AE/0OHarB4dzkr/dQANk8zP4bQ4ND4niS2J0g9fYkqfsvZxH9sCHPNc8
Zp7Mtfv1KBf/mkXaOa6nGb46yMI+PjiwoWvRlXmvioojzz+wxTLIdI9tj7V/XF4NeBfomRajHxOz
QPKcMoMRfQPsdibnBwahjjD03Qa7AgPm4C21TEOjw53gbYNSk6Pk+ONTjfUGgmC5v/d4OPi+u1G6
fsw4rsimiTXBHEpjYHWOG5sHDIo+Z7uxDtO20TNbsVU1coqSUy4HXahYc8vxfaHaa90g92mZEaFV
QmZqdie29JxNrGcuwGrukMwvNFhIkirwD/oovg8XxDeyGcGA0o8ba8qf5J/LuojQL5CxGIbF/tzK
PQDDKwDDBfpiXngDn/ySyyqUto2xJnuycJCqt6m6dwTyjIil+dy8QcQoaN2LXdFlwkv0qWf495ur
iAGZ0/HMfVwjbev91R8KhG6S7Ke7UnOpWommxKGT2OmXIkxKqqd8SY4ICXS/e0JK54MV1IIyRyJ6
zg0o4i+AKFew2iR2mpnmUuqrSl247UUrsXrbNdI9cch+MbRNMoFqYE3/aOXBQTMQMbIhQZ41beBQ
r44IYsNjAsTkF8ZGh2huc5EaAebzYYAL1WvVlW6awcG0JUDuHVZwdfFl2Tt2T0phxW1S56/18BNc
GPP8Tnc2hW5Q3qc1a9DvNs36+LGKiREU2Ma0OfV6MO/iDgaouive5sGQQqYX7HPBui6uvKuvir5u
65wkasqPPj6XAxcz3Ex3ZgzTCEAs7Vbeze2/otLuUMB72tGBJhvtS0ULbnGU1eidEvS0RCOBqv6I
NMTqXVNVYrTdE5F66aWJ87wFUDj07UjINJ2kwln1CQi4EF6nOImO7omIq40JNwdBE0xuag2Vz3zR
GEukGVzZ9LLre85BVNE2FHqbsn8kS16DdUsTczLfl2WpisS9VzooNGQBOdtsFtKScs9OJJVA2Np7
n/gUqWFTv22zKmlby7fI/Y2qxLI+FpJAoiANZfKwVR9hLmmIZnzYRu3lzSVwq/kCe8R1c0sffkg8
sbgZhZaB0j6IIpBp5F3vjJAS7W/BOw46eAqQIE7EPdCZWaHsmnuSfPSWwVcg97oPFlscsr1mSMML
u6op0gXZjMNCaromPwcblx6WiXAbS5+AW/mpJpz8eyJm9espJ1jjebywSefQbj2QKolzQGWC6DxY
Yr1KZVTMSt/Vu/KR9k3OZcfPsLw9Gk8vV14qUzE+26erMZD6FkhMDMpXPDhd4mortc8OI+0ozGV3
HtWywSEwZ/T9wiARKKmTUB3q5xItspRpc2THqAWAs8o+oetXIDyaYCIcpZcbEsIoJ5r5zijyFIpd
mDVeeDTCYc0rxfT3EVuiHWCHDC/iTKe9s1Lsie2MdvX4JA8BmEPdqrJhxjsdWIf43a65YJpV+D71
LmyGhqjp/8WXEqOUfbIqF6+MtCpO2zwTbNnKENVSz0mHgOkpLwk0hJ24FZ/7haSjY3uWxm9JKpo+
6e0GZ4s/xaluXcxV7PBswspl1xrCdbSP/h2Ejhpf0284Yi7ROzw91LE18mTekrtsrgIcOSCg3N+G
CmVmcZ2MXrxEGuc+vwtC3YcHopRUIq28gw4J9OLM/yqHQLKM8j8YQD/aW9sDcjY5I09hoCgVlhWE
R94BOP0gD2y/mxYNx9bUp9h9ZAa7p9YLJQmDdPuZKB8JGFvtqoRBnlkxdK+NyXouaVQ6BS3UZIdA
vyrl3H2lQc3mrhynX0UDbInWeBl15WtvD9llpbOH04vAjU2Y3A0R5PNBz0i+ee012363TGLDYa+z
h/YpLOgyL9ynhyH9j920ntzzISCwdei8kmfjEInInWaKPR560zecB75rRbJO1pk/SZoCJfpDmGr8
MJ9X72WGLIBa5NRdp3U92fi+pGhLMIigb9MDtKQMtFG5D3sStt3ndZ4UwHpKFIFEAPxcGiMmN9qE
HcFUGGBqZXLuBfMlBLU0ry4wkaliVhzfrT8mOkZOifiB/P6Mek5uY+CO3u4jNpmg7gZHSEoSFd3o
cZTeGFjSKc9OwiaUdSIc02EsSExzsOtWGCl6hRhYzxu6yAqZNIhApdZh4V2VKODysW2o+Yv5PxH8
irenk8IkoTDg8KDocUS7UH3Y69bDiffhVEzTPDc1ErcsbQLBZv3kLN/06v6OWF7RftZ8kioKmqed
IjvFnQXNGOoHAIA7YXarsrY5e9BvlXvMCB/tco1fjJ2s8mCpiicQcDHA0FeHLe2riK28Ww7r2M38
I2J9gZ/yLEZY63XX2CGP9/z8dKz2aAcZJSs5+CanfnJE1QkvY8Jg6kQeg7bZIrU26Jn33bi5f510
yV1tNo62wV6P38BQF4oTEIs7FPr/Eb0u8KACgTmQIKzLGuj2O13/MUCg3FODoQUOldS1yCieixbv
fhxi/zKWz5vbsVIuruTo/HjdA9rKtKWwDAMJqEXMezgJ458DxWMvaeeqLTdih5F9ss9LPuKaIXxn
tsGf4gB6RrwUCAJhEmd+gMcL9I3TDuvBEfNrJ3AQfJUp0FLj81h6vas6c5qUW7mLhseC2d3PX1fG
5SWnH1qJkNfbHgcKklj/9xpiTgoQ5FmACqd0aTs81U/wHIRCIoZU8dCjX+8QrgzVeUPSQkBMtgqu
ge5WifC08NuxpOsQcfEphGOcgtS9tW6JdKz3jUNgt9sPzrURdIma5KWQ6nZbFQBsi60/Lr0ziVBN
GyP5l2aGQAWc0wIGslRgoCAmbz/tZC+RnALOJuw2P3/uQ3e8UAL+rnhDsJrubjbUlVIzdyrdhX4r
ZQFohfP/0MrNTHBNA68OWriuYiLG2HHSl+a3Ke3o3ZpyNVVrQ1Cm1Oz/EpncXbNuSdlzxEi4FX2D
94SLBAJTb9KPlli5kDmYw27Ox8Q4NqCvGVQ3T/tvosgBa6xWLaNYLfLUtRiOcVRTyJAzGB0ZxjpH
KzCo8+YcyxJg/9aCI9vYOVZ+m076vtq/dVL4sZkK3HMYK5nd9pxgdZMIL7j6saQu6g1YduVYhrFV
iS9FASJt9cUgEJIhQzFfHzTbiK34ZIT2JsdA+W/ZWOmp6jAB6eqd3OQG93TRZEjxPEEw+oemgKEL
Q+5qhvmh6+md3IzG+PimUlN0YtGfQy37DNdiXCIDzwmWgE1btqnD+rKvGgUhJsgULjMkc1r1JfuK
/Xiy+7KIjl1v3pqLLSn0VrbDZvQy1f/DP3OtVRMGKOWlyCuP9vaqn8DvQ7beQygEL7dg/vHP8eXN
7hXy9+R0Eh5FrSEST3ZfixCQOxuGuw3Md6+ARlYQ0ma268tUK/qGQAdWpjpFgJNLueUHpcXm9mPI
xEeshcVwWF6amVlaTPD2+2Efb5V/mVT5lZODoDUKGZZG5vHT+BGkv7zmmHMmjgpmszIsXENBTKLr
IcbujeNZfDoxHXpNXmRX5su1ISYeYq5sIqnGMn4HrTZozhne9A1pCUJkt/yb78nBltg4zeao5+TE
DxalyKzUBuBLvT3nSVAcO1j8lIJQW8jYY6V/5n+/VBDn7paceBaDCFqWEMJOwwLQbVqWzMWZPNpg
1PZNCMGpkJhVRNukcBBv9Ftk/Exab3nfl3UUdOQKcHn501ZiSQVNiof8aCzG/ieozmPCXY/ohbbF
SKYlE4UYr/73U3g3W8dRbeGag6R/Bo/2Zo13crJQG5tLDQ7N55EWC7r3dj4tNzMHQ321NZ84BaOL
InZ34aGkQcyG4mobaJXZhz5tMa7cdekaZ8n9OvLx06IWvLyuKX3ZANJ/Znh4QIk7eCsKGX02WBTo
GOZ1hzddw6pU/sVwzIrvc4clIgxZInnivqMw8r/q7lDlXisR1vzQr5QSpjsAApFG7qNhAIFRZOc0
UPdYleWsUrF51WhMQLOq+DJQAzT/r6sqJke1CYHQ/zHz/aH/ztbJCRMTPtBjXvYoiu5lwE1sNreB
woLTQ0OC9nm1YsCwdNwpb+2oB7MNIzRfNsJFNSHhx+LHwdcwZsmk/6SkZUqAzau/wK6W2Pr2UaI8
5iy9RJIL35g18roo45vJFHoUZ2H/mNHYteRHdINwCDPCLxyKf/DDDDM8GVW5dmk0tnIaflWQO6JU
HeUDaOGS7GQpkL7ocX54s6y83tiMV+SWpdf8Pt5LGLV4Z4OMRzKzNZn0jlyCYMzJLfqrgRhQQO6L
6MVVJUmow1HB5A64YsIL74mYzHYYMz9CxGbbOY+X7W5T+AB4tDyCPPrL5frvV8gz8jF5QnqjfIgN
GEN6tzlm7cX0NFJZWCiOtIl6toTMvOgAuaJnZuqefcyazQuvdvbc7N8uoRRBJAKwSwyBaILnMR1s
kOBnCK/pi5ukcsmMYAUMTEDZZFCf2lqRajcnWNpyqHFJDEl3FFWxrliZYtCH71uh2rZizcHCFm37
+4TZ8iH7TlKth0KMY1db8iLwv3A862q0+k1j25No0Zsn6Kae/HsNpR39LVd5XGg0J+7OWokjUJ3r
/g1I2ZlTIxztn3KInknnBFVaVgiBEjRBL5MeFxtaXwPbKCfuv7doYwx9tQ1mMKL9kQiVNh3fAkwD
E2M7vkTOs7IW0klR6m5d13LsFtjWYqATMXOB8rZxB+ghE9yEzoZXOpVBKiznK29I/tgZ116E2AjS
ApeuRbUcA3q0R3zcKmnAJBEGDD9IxWBBBfqB6g/QtfgigJ4or2D6Yt6EbSa8FRSX+gGxhC4rvTr4
A5GGaNHhd4MTICkds8yhh+LUGrP0Z0KxOSBTANPqI/HtBDHzBuXkHKo4k17GhwJdkEMEHHkh1RAr
JXlJSZ+Uns8eMW8mHDyrkef0t/abeAUbevsBYJRaJPfdtdBD+DY59nA9wLJsVkr5F550RFsH27/N
HscPeNHyl9yB4BpYhcydRyf5GNc/SAE3mbHg8cUk52O9G9itzNw9TPku4IFMO8MYM08R25cAj6mp
xqpXN+AohaNlDEQuG0GvRiP/JqAWQv7ms+RSg49XuUDCOuBT05z980/pzdowDv+TrEPtJaYhoqYa
s2so2lvkVycNuo9VNk7EXzvroNVsEdZTupV8IPV5ERSYONZHj5PNRk45A93JFlnqq0F975OY+Ixi
WFOD7FdTlLrcVD8tqL5mt9zQawhL+AEKdgoH5M0Zovzc1CAWP7sCbeWDWDoRIYTaPDr3YqjS+qVq
y5z3MR22LyCETYKbdVEVRZ2qmVZ+prmNpTjbHJhatz5/e6omBLUtT+OZq+xf+3rUHtrNDqdZpBbR
RuLDAPP3NR0Z5vuLF0es1crFXrNDVbn3XNgY/LzRczn+MeXVzeuaKM6ZJUyRe9z8CA9XWFMsdplA
OLhM34ChvxY6teHtc/BO4I85VxkqplP81gG3tPnt7MO32zFjFhA/CAZS41JvE+7AzRDGdBRahm9R
/FCGYGeQmfga5ErgLOFopN8d6YyowwP65eFSPywr2N4+Rd8+uPvDPX+ERu4ZKixFBAKuULljQHTF
0yXjYpZ5LlO5e0WD252kbd9dbD1p21l04IDKPz63NpCrbPHx+Jy53/T+G/EBqQh4aaCsFu+heptc
DOHEUk/ePcAUQxfkDEOeEvYrThYxOl2ITQf5riFA5gwqZT8wBZMxo/fa4TmeH7V4CSYl5NSu40ll
kaIQilGqySL5fOc6y2G/n/YhzAmi84tpV1EhidhQtIhpTmAUeqMA7JLIs0lbIeKiIN3VndgHEIMC
jL+3cG9QYIxOelW+9Y33+PwH4MNopEXFInEjZIXlu2rsOz5uqQ3mVL3GX9fUi9DJnWKFr9OcrOsv
PkCg2Ma/iLKXmexrmXSiRVrd4sNy1+2oYAVgCHdUgEpZa39Tb2tnWh7hytDxpcIhXgjcn0AOhUt8
7GHzL8pXdmmMyv7HYcIwMkuHuDzUnu2DpEMvW6fcPVKprBT7FaERuTOLhj4W4YEX3RB0hqCc2zw8
rtUP+TbMZH0K/hyhOUnkQDGPYTgHI9YLZlVexUCeUp/dT+syTjlL+Ktx87/ygsODRZCfUhgQ8npe
vCMo9oiozOQWuuhKhggvy7F2JYo/K/qAV0rgivepmiyOtp2UoZJ1o0Cp97ssh87FQ4wP3A133XNj
t/9KDq31jCO3k+HijegtlEMBCkz4vZQcrJp/PmD19B5EAduuyjiPLiPe4nngkLn5D0S+3llgDMlP
BDRQMempOOU5ZlTa1Ln43aI5m+GEgGkaWUTJpt7XyA6evudvblBTaodgCLs2RAhZfI6tkLJPPQ+H
/O9meWVmSQlErhc/syVcNap66r4G4MICer18NXcsogvNB3ifi6cAYCvPywvAFck8URbGKAJ2SYoD
vJycRtKkacJxqClbdkX6cn4o7CuXuICeyhnssLEOW1xv2qrqwRQaQBAFFXdXdQYSKz0I5jkYB7M2
Z7AFDiya59UsXzIMnYfTQrYHwXjOXg5JlUVNGzi+2S7ZOkcuo3Uio6bIOFjoxJ5Gs/YNhO+YfFj2
8yAbPBhFruVxDtNI/zJwxzb8H0I/Ctfjt8YWSnv4udb5KF7HCO61OdNX7dwZxM15IfXpSI+qrwcC
30I7C8Gos9OW/gnY/WZRBZE0sZqAmn/nsLU/rMyUkFP9Bj9VummD4vTmE+q5Rzts/I6fF+5AxOjc
0AqYXWeTzXgfKoSE4WM8PPpLmI9uUdCgLja0PBF7nkSQFBJaKaHk//qtTNa9n5XpgW00yRCTvCYW
JTV74TKoJPhMCxn3ixBU4OlgPEoJXVEWEI0ihrpPQCYbeOR09K0BD9N8q/8wOahndp+Fx+zLI7Ds
YuDNffcVeoz0Fa7U80w2xmN9zcv+OS7nroPp1IPdI+R1v/QD9Q9BtpJW9PCKVKaVfWG5VyXyGs2u
O1rmfC3Cn+iE8q8GDhJOkyl6w+zt151aIPYIIOCzbnzN+J5ZQtJFpNxk6QIzCICNvvF6psDiVdZI
cr08u2xNax5Qa6eF2Dkp21wZ/KF1ehsbMSICbYD1EW0nD5os/xLm1ZtBQwsS8ut3RIYo6Su2mQV6
SU7V7Udbq6pwonWFDqJ3wcCyW0t8LXGnZGxv8UeU6wuvCYXL6sVUdIAEWcrVMjkzr+n5V76f6M39
8moWNZV58ixr+syIj0Wcr68Crb4Tp4tQ+GDCV0MkZa+sIqGSFlLXYX1haOvyYpzZV70C18EXYsc6
k+cOZOcqsZYzGwOLWA+7ZTEYk4IhBnBdpFRSEWYU8oauRXVisfAUpzG1IHE+nyK+hJlKtAxlQYsG
fmVlkegOFX+U7D+rWP5np0z7nA0Q1UCt6aj+NyDBcbeV5daGe/d7kbrO+pKJfOPQ7Jj2BB7DArTY
6SRJbv52GRHkMJw52eRsYtUQgvnSGZtTUgmcs6SsSiaTwY3McuVos8+1UQSI/XJbyvamYK/JqX2+
8QUI7PBMAAn4AHvetF9Tv586vlJBJbysjvYdbHX1z/02M4qOv62X/R0HmR7G6a9eCLrjZ+o8bRmq
IF17/v2IR7yo0yum/87ECydrBmJsNG7cvqeGKT3o/nyACrFm83Mw/8ea3rJnh5TOCWFHUaliftWa
3P6zxUfOPL6scMyKlq1KMI4dP317qXTIml5U6uKRjIUjSZt68WmpsrgLjrkWOP9Jzb/QD5b832ex
HrTlznct+vczUzdiZhm+6CSWl5/k2wTwZ1T6nVi+KNQhdx5iHG8ansh5y+zmNoJoSLSb/A3oh1X8
qoLs8qpmMVZ0rXLB5bZYabIDkn+sLVlDGT4gx6MQOQjcF+ofGH1C3ejXqMoEFkVYqs0uRQ/u+gAn
dmDq2MJLMWgXArWtvptMBKQH4RCNU9fRR50+yWEyc1ctfpAp13ATnZq9t7cFCR+lypioU/1Avwjs
unP5ihuo29i8Xf9uiO+c/YSiloN0v26RZck+Q+yPj63ZbAX82tKXC4xPJQhxMymcABQqGYXGH00j
+ZjW8mkW6u/yOkW2D4fOrOjZrmFMSXV07TbJtgV6cRz4i6rEe0J+mdT2AZFiVuXep/B3+pSJK6Oo
5WNn56Wb/FcUIa8J5qj8BblkSiwX0jUhBLAPvOZoVlAlubqGiWsoFPFeWy5dRmQ+N0XNswmuuklU
bURagjK1sLOmGKF/ACLJjHzXBQCNvZGhHXD+eZ2gbGAzY9AhyVqo3Xpnd+OvPJjyhKW5XGQgrjJ8
htt/d05hjcOykm1JFccJNCguWUTNtPvgSlcJYDy4B43nUWbGYG1pmxnbJd1ixuoLE5saNJZhHPmB
32XLvU5V3KqLKS7fTiFvzvUdhVwu74hqh4+s57Bqkf5xboAEqnLYFZ1MxIrGsiO71KtoNBrPiSkO
UXv8xkHE+ZnHSRce+XAkm+lWso3FeRSFAgYzhYFn0yZ3sSULIcnc68RiVkRVGUMjNMCS6MrDdKJk
kChf6HtK7zfNdR38D7e44mmm1IRjwSK86UjsXvps6+0tY2ANPZan2iivnn3TiNbQCYTbMmpBpToB
jndCK5em3TxBorpiu3uLHfWuG5F8kvsnuLoFvxSUiTncBq+k1D6RiWSRHW7iniGxFlsLeff7PSs+
l6Zgoc+EMdyrM05BfFESmiGThKiCsIPDFgRox4YKge2+lzpFMefwglcRkCx6xvemAEv3HT5mtEkj
fcno1CNO/1betyBE73ykccn94gcMbb/WKdVJXTILKOotZcvFW83oVvLl4nfg1M0BecbR5S51G0dV
DVL3W7npuPxt7sPIxCvU9+cSi/LfAJo0lX5w28I0I6XksAAff2sJILWs+dR93QiCmVgzu6JUwm1F
KQNF3zfsjD/zTo0JnlMC4G96/7rtlCS9Bq9vTvyYUfz3ZJRxDUyGo2R0+Nt7I5R2Kcu5BLhiJv0W
E++qjSlnqJzykDau6VjUAjrF9/njvSJO6Qi0VKtuvgejj9L7g/tYpV8sYONTjeA78weiWIXB7AJn
SRIg7084CwOpu/yzY/CZr2UUm80uPHjINnK2nkH+RbPipfn77Q6bkABAT2Dv6sC4y8TBTERUibxw
Ox/KBsJsRD+ZFmhZh5y+wBvZcMXQXqfFGdvdmw8B9MRwXUpkWT5g7xR+I3ERsBwHp7qnGHqQjS+a
FVXElP5V+luMH94KmSnLzfH7lGvUGaEhtzRmJfxEUvxbPRgcqYBfnu/VOu1lFKzMb/wRZ3QAA63h
BiJr4WzzIoJ3DS5lqVagYSFPHI6DYG5i0BccbSTdqKLHvogK9f30VCZYJO1Vzywo45isuK1KJqPa
gdC+eWqCAvotzzB3HhaXu5m13pVriBXdpD2xSH5tcq5xeeiNy/Fulp3O3gEn5xxIOimMaUZnc1EA
f/Oad+Tdl2CYf0NxKCz6ebT9G5U3TV0lTfdDPoVHViwyK68RaO3bGS/oiHUo0IVt9uXUbelaMGDO
cqI5TNKeGzQoCPXTGO9fBW/LyGIpaMNrWmnvU0/NgsQPeC+YhuuWT74sPvQ4JedpBBHPYgBYFpV0
KMnSzWHHnHqBWAbjDtuayZGOtpinOp5iPl7nTLHGhEjMC5qoipC4c/RSQdPq4DJTSjFvQFDGRJy6
LiV5LoWgXcfUit9K002ggMwY8/k+ToJJpRKmckmHytIsjFQwwwciaDtZwlokvDbpg3aFM+4mgRj7
I9OXKqqaaULAKvF4bLebuqNqt9myx7dhBZzOQj2kG7Ws3WM1DVWYCYy8iB/QBKS0n30tbxcw9jst
ThTq3us73bojMMxd4yHzyEMq5qsDznjAqLH5bGuf9FbibIjMHTRw/lHmvKc5M2bcl6BwSrX4uw9V
pDXfMV7otIdbxHo3MQys3/J0V1ZZxED0JFeoZl8TxKgBG84b1FjUzfNJl5y0xEZALZwDCUfDACpY
3D5oC5gNBF1AImWi/+Ve21GzoEJPAmYBxJS9wsaQkZWbA8zERUOMD8+sChTZ4A1BhLkNoom5+UmI
zVuknP4of0ekzlhtjrUvAWSpELKhFaXpvTjXJBOc0hYbGfDAVC1604fuh0xFOfpCas7GBp+EU/y6
PPjecTD6UlZxyNbshkkCAimJgSLF0foSklEfEjc/Gse4I2dTzZsj7+X0qPORjbnpMSAPuWDh6i22
a6kUwj/q8LHk5Tkv6HlgHhMC/k5neFB6kq0pWSvkIaCpYfPSTdQEMNmparYDmCsgSyPkU/0jcs+b
/Tgal7Y80CvLiWyJ6qdXzx7UfY8IwQO3QPykS1cgwUq1S0Jb49ZIGKQJ5SS9Vo8ArOklRRqlC+HW
7AC7t10vYEGfaK/ZX70aSAH1Gv9bBPLhqFtwLjsgwf4TFFPGzhbk7SBIyHceh0DUZTKmB+wUXWvk
3TR1pgl9D+XiHeAdAEqZL6FCcMJobnGzNL/R7k5vyWlS7HV+4jJhkhlwqLYXRrUhOAeT1I96TFQC
lYbAAv5JoHEb66HJlKcxWWdTKYH4OKXrPI8VbWWHlVOOY83/scdVKCwBxRXIf+d6vR8VmDakiD1T
1EX+Xlli+0I5ebcf1aZtmC5sQALlCjtqYLPW7oXTd5s8gtcRLkICk/d8JGX5UJqv4VawlA/Kidcl
bcVc844qiBXNOuLycx+bxmV8ykUwtkRcXYygheRsSv5XZMVWEVlx6dyTS5Kav36KdaQ66wNhuyQK
GAhXVf88qEBZAx8ngV2Y9DyN8kk04X1SdfDVlLOh0GVcJzDMNOfTpIg9VcIuKOvSQCFuuZiFNh8m
S/i9xPz966fupgOrk2WK8aXSqtkVOiT+sapJ2rnnhYXYXppZeMSl8U9cnbaGkv79tW/PshwVDbtH
ZFg4r7lA5t47rZ7rxm4M9uTDZ6RlDswXakLKa1CBvi7YoasNbudyPJSUh5Y60zJv1zYOYt55ixx/
7foUGD8cErAisGpk0E46bPhkQ0WJLO+pCw8ExLg+V0MCE9/vy4or+Dck91KYh2mWHtSNU00aTfKl
xeZFpdYTt7ocRnNRRRAQXJekbJUEIfyiJFfxv5x+8wGgfgIP8sQRQ/0ujEdShRXohVTIgrMvX+L+
SzLF3g+60rq5gJeQkc5gWNjaY6vipBy6soJ7Hwd3JLMFFR1ar+fR5ced3v8ytp6bYM+BTNqenFmC
LJuYjUY+0AgGQ0h8loLOg8Q13nzQSeR8hviEpNdA62J89Fm2dNzNhw9kN1iAo4Ffcag0C8kcxi04
8e9ErYnGojVT6IRuFdwKPaqIWB1GqjDD3qLkJFk7EMQhDSiWn5zCCPu4+AENK2YwAtSNeEyAL8qY
RwfCFhOYg03gg4FRatOPLjDlh+W04PpO29kTnwaumQ+E/men7g3QLLtHcVPs9BLXXPeFA87dLBPr
N0Psl4xPL+R9nWEpHr+xMjmFbtpRk75+giFfINzOXKoyvLPYlNV1EdBL9R1rL7L1b3H6Ssc+8qtp
kyQzWw6LOvO7hrm/sE1JjjDBfR+Jw5yZt8k9AtAp4jROFLdHIS+876HGW8rGF0ICf8su2c6q7pm8
zcKbNL1nQF8Jo/4gRTaAsNm1KHssliNYkyk0C0fBwmauir9Rdl0n5Sdqll1Ey52PEAFy0nuQw8o1
VF/SpvTFsbvxO5NOt2QYd0mEubETrFVrfDLjQed61xeAO8c/wtNS5qc1IC04tie7Niw6gnDYK2bX
wpMwhLNfsD5I0GhUwKKKmPEsNCPDWSqGtXZIjZgm1nzR4jP9BsQFj/zrqfTXKTf2DRmEYYllURao
PTtQxMvuLerketcYCz0R+CQFcAjZo2O8eIkDlz3JxlVE6XhXKDRC9UyWcFQp8XU59NECXvQfJPgq
QLcyD7mgaoc2C0eY0MSAGCevdIiAVs3QGRIQss2GsSSydwwtpdXneRmQWj73gVTgUsurdfNvVmK9
pm0U1QNdY5tvEL/HZtNrCzJnXjVk2YVH3DONpDYRZ6PF9G1MQ8WvbQba39C+1thBNWQ2C4LKdIjG
21hcU6DE5PmAGDJXoy6e26p+Rz5yqSB8kqmEz8WKb9KRNrElvkcq6n3j7uR32Wr6ow/5w6yfZKCd
9SKbT1caK2UfPm92y/qwnTKJ8+FKvVZas9JqXKI0A/D01jWBsDiTcPKwi+AguTEL797nWkjYzLUC
26brCIaCUcjsjjr3AEf+J2UxYezwZCMzo+sY7+cxRexbATwd5YBYrYMlnt5bm2IUg8DR6z4roe0q
H6pF8k2/xsVBu48gdAI/pdtJV4evxR4VZ1tEpyJWT033SkNrok0WKti4OugebOBhcGvUpfnkZRGQ
n5zDMUZ1p78/ncHojb5NYEwfGRSGQZaQj5aA+OKLn9p8aVrScZwEQWs9kgApqUQdz+14ykoXwoYi
f6NX8tya1+CGFcxHRyJFCLTO9qTcEkmwsL1pevg7qjHweiYiBMTLfewO+z+kLMVDjLiOuP5h9gBy
pBVxtebavARID4sGmFAFOWneOkQiBk9yZixsai6o84x5YqsmnP8JEKx71Si8+EfzunZQX5tMwVC8
GLAoqoFGbKV3SruPs6gQM+hFeGFJX4EboNwPD5dndpx41P4njNouAmHiO0aB9w9u7wogrH1zf9eo
v04RgV5uoOYhbU31dvs+bICKVbeygUhu46BQyiPd0SDD7rDukoXPu8Ai0veNwlowTXjgY1ogkpTW
JxYylblgqP8s4/fWEmkLrKqdywC1Y7j5mazBwLyQTZBeBHRev5aF73eZB8d1YE4QWag8MfJVWWfQ
u8Zef1Y51L4S8vzuOaOvD1lPOtq7s4N/cdCw/PuNXTcUn1CUBdkOf2bT7DstZ2qf2JxEPU4kA+ig
aCgXqchzNel0OSLFyNNa5A3o+/Qh4gd3rjq5JDHvgjwM3n5wTjIy3/WtfraYn3W+3RjPFlBFnsS7
5j4UijS3cvA4EmXj+jflsN+S5c0d4c57xTQBGAxieDTirqeXRGQCLQYUPI+NVEIDKOFSIH9M4ZL2
mjnTVg3X5ZgJpHzv6a9e8LSNL1pwX2SHK2NFC/Wn4TtfONvyFgzwik9t3w20hzDsZaDzRtO/zIic
HF6pnSLoJXP4OTkTAPPkdE4CNaxqUnmXKUJXNE5tczi8DC06S10+YN61Ab2Q0Nfc4V5jwE9wNQy7
I8H9Pry/dGTTR7bi8gFem1O+WPmezffKDFliDTGufd9i97liJ2GjmQ2qfLR3b/Z0LgQCzraw9Ck0
wXu5iG/aVg2Igqai6ziDD/ciZpEUmpW3jA58d1qbGqaisbxbZoPJiYCwHBf4+Mv8gOpJd+cKScg8
fkQliqCyMjRky0dG2xT9gBMyhwqSnwF7E/nsNH14rGxqJC0VVcBytPkxYLkX5AB8eq2hNmMqWrP5
xEfGD7/gfUPy5R1iwD2nYo4//MKZYEhoIhKAhKZt0/XuNKqlKbobbCbs5nacYXzvRoyGDtS6UHMv
/iBbP9AvlxMKY98g/LuT765nJg7YT/f6vSRNXrxq1J3tbhpx2rmdGwVyaRZ6CinYhs63z3ejmRet
MDINYUCkt9oIeMoMzPgwNebMnSsc+lBCM84MzzJSgr7iPD4Q7Kur+9M6vp7w0c8E1j8ahsGZIc/0
NnKuoLAlyEj+cy8icpB3PFFoP5ZuafahkEF8zlYLIShQ76hfmr4EtEHZU2J9VPAz7RxlP2YEh29Y
uLyXVTZF3rfJkfECo1ykreWvVZMHjGlj6N11l6R/oPrgCjm7zm3fXQLoItN/VkxzW4kYSt9IFkNc
kA+6BUwv3rAKUDkl9lviKgCdTrcYzLzWvhPlzPeqKuT/S6DdAPK2a4QnjjH2NhZh7zTYfkRw/NZi
GwjaSIv3JdHlrymslzkW+3kxFX0ZCNIdaokgLVPVuw/W1Ciefu7RpDFznD8J3Cuh5/89UDSk7LCm
NUF9XOJijk3GpE0GHU3kANRvE9ysSrlsXd7RJdys6n5FyZTMU2G1iX1S9NZbcJVZ9DtXu0SPyzTi
wlOKB27nAl3a78YGSuSzRAbz7v0R9GDhX6celiWrX7n+U+281AAm4RMyZxcBzXE74qZ7a4CVUcLb
g5p2Y8uzYY6EIZH+c2Grl7zU3YQloi9uZg2bQz9QgR4Q3WKrgxrorovF4WMi6pt3WGv/wn0nfsIq
ks8v+5JCv3tKmCDdW1Ns16xcBY6J5k/dWtqY2B4hJT4ZBJIvOargTHaSo3FtiWCBkNQji6dfHeN1
osGoGbl4DgNLp+M52mOXcmft4Mld5JoiaCEtw39cAUe0dqgTgQ5+qrX5pBA/JRh7W4m7hxzjmb3/
SQPXwmArI29ZbVVURixrL/ORFc7y0iEMer86BHtJJnrwIsHyOEKYe7wkhxmyTC3dTAWOjkJNpFoh
kWDwZVuqh5dWbwJlc/y3myl8cymxHQadWRmrctGuFf/sk6w+D/vKMoUVd0o/Ze0g+11umuD/SInK
pGwnjSSbT7azzNuYrkYwKMzSfjyD5soBGMFBu+XHi29OKx8cgdx9IKrid8nLL08keU9qnTcSoRX3
uld726qj53+3U+T0YdG4tbXizXtf/kyqPyI5VGrLhpxBOBIZV8XudHWaoLc/T9mAAvtxj0oHEpqD
JRNkDKflOKNcfjdKJWweJ0j/iEV8f954NxbKmD4t80AnWQfln8wvA1u0iUmfBAGUF4QtR4Hr0END
cv5km5UQnsRRxEbzIc+XQBpvoRg+9389eLu6pIN/9NaqVy0f4d9MK/UIbVyMvBnT2k6qqZ7gRbkK
r5zyWUiQ8Yunxem786x1AD5nX6zUBEs3CLrD6egy+BLrqQLOp+RXF9DPRQRwbO8OKwOljQ7o7IkP
hSglZJrgbzQd0cxBHVMQo210Ne5vUyQNROFQjCf7igshW9OWjfgtBTrFc4i2+q9jaLGNYb6YNgsd
BIf9167jBGsxE09Dvnq7CxJQoFSK9iX73PjS0vdALLFN9FjqktDC6eWG6Y69S5MHbxP7vF1A5gq2
VZuxItym3bnOi7pow3wNPf43QszvmCqOPeSBJr4wgrCI7V+2PDImWdxBfiOo6s0NYFuancuzxzrM
f4B0XI9bR1rc5O2uthzOI+NjcvEnZPIngIGpQtzx51e9fJs8+t6v1+O4Hmnz/2/QKt3ni55sff7G
NRNIROZgrQZg1VYdiDbOxAmkIWE3Cf0h8RY+IsR4DrElfEFv2UjplYTt/71BwcLTfjd7039SlQza
n4QNeZz3R7pMt3icOYBpczXUw8H5hqdQddigudS9gXtTBsJYgWFUfQ67enAYLQYd3rEC5lcV7TDl
MBkI0y7zqpLoKhEChPFR8S5hxRwBnGst9aI+E1zKnu0tiZMPnoNu0isHiuFnlZUzcvowgu0eeLhN
ikHDbrRR0J0TU7egovZLqUZpOaL8xDYTZfpLKJhBRykQOqVdqe2JlugK54+gjGw1QhUgy9LtB+ou
s3R0R8spV5OiQ7FOsuxg+HBHigAb2AeTE/Yv5XbZ21EnUlegm8JJEQEWgbuVSUUwAkIr3hmplDLI
/gf71vwFDSezXtChMQy6nVWEfP9QUIYUW00H53K7vIxhiGP6tmBopZShwnsozRG7crlD6eCCWdrc
eZQEy3jiUAOQcQ2EHUeIuZrER4la2T2wJaUjO4TfrXhvMfrwxtgqUShqPhOwcqw9NKKhiDBT+Lyd
YZcYFmFJmLPOXcIO92ZXr1FuWFyyEpkMYVL6d5PrjbaI/VewQDnSdXeeqnmtkwGEcVAZc2KGDPbd
ASTcurNV5ax7OlC8o6V7lI6Q/gLoigaI9/DH/sqdzT2vLScesnoEq5kgNUsnzWDmN1R/LI5ZQSAn
ps1SlAkT3l+sfe7mYN5jpRcsAMJ14ditXMUfxX8YT+jU43KWJsjs5jp2GvU0RbII8YKpYqyJ3o0B
IqPLtiAKsdWcbHdIHSFd6AcryCdRng+PJdschQtZYqEzSpCsX+SAKvgRMpCj3mQeHBQ6XGc0JzTV
TKRTw195ZFPoi99LvET7ZjktelP9DkjGf81qXJfAy2+/+hGYmMcRPA888OZen+nuBQkKZIIX3G0u
sULMV1hpfD1iqfQIpz+HUlVIYcFl79Lx8ssh3SK1C8en8V/VhcrynsjzODrQ7EwmmCjlFB6Jknhs
iXyb1i9J6QR2peYGdKE/QPlC/UgDnpdDYTWTcVboU4L4LSZmpZM5dU6T2XKPA+emgZHDOhBPz5Oi
AyY6JInL1s2+63HGADXaVEiQBBvdkCIgwADuueBqHgDGUOx7W3qbcOxYfQmuFPr57xLeT7eJYDF1
W54YmnehohDSzV4P9lyLi06EjGPoG2XYd4hyFXLpGaKW2z1WVErX8/kg49FMehyRMrajJXXfUGgk
oUj4WLu6S/CGbdZLsi9nG0dXzopBLekM9VsKemvD0u+Tp8SBMu5BHoto77MDzDIhAz7jDwRheOZq
/zBb31tm0tLrtXKojlRBlIJ6lZBMAHVQ8F7mVGk4fwm23PUu39PECH1gnhVe3VUgQm2cm64bulM8
i+nscc7GTkoQwfya1cfsdG1Xe5Tx1in7lH/880QUHjjOaLXz8KNR9Zj8ITDh4ZHDgDP89IsYLtJx
50Z3XZU0vbDMAuKDn6fZb+icsJ4MGGfqleJN/j4ayLF4ATLfiufb2bfwdB+cw/178CaIdHkDybF6
5f317DjbdszYHaoZ//Ek6t0f4MDFmt27RaBT7SvHqPh1aGaX9Z3EKhZ1iLUMy901UDscKXguxDns
7EFIhJqFCRCdlUd7WzIh9yaOYqWtEEe1NJQo7L6j1qxQ0UFDI6YXrON+b16Axur5Imf4PRJsRBoj
0V9km7o8X6Cp44bHPMvEtLq4YnqE56B39UCO8LvN4adV7QmKggDUHvHVAyJb+siB/mYoVkai+Qa8
fmNg0gwUlSX5n/x1ONyFPMZQQquccRKOq9ZxkW60J5CjnaoSj81UehHGF134kNjOImoWfbZsPT64
KoSPshPfy/2oH8XhMCHxLT4PZfSBRrtzTrrsJKE8WCDySTxn3KS/0agoLzgI4b2IjFZ+y3iIQCAH
IAmpXgrmqpc3i860btKj108iEEnUsGWwI6uCDxv0ngW6yv2lwTPrIzi11lEiWavwflxiXW1er+9g
lxKAyw65ptIhpylIBfsAI4rAbSTRq5ycMcqMdNIbjpz4vB9yHQUBmsSUtycA/0PTkNtE8TJuz9Zt
h5QAGticOZBGDVW5+Bqz8nIl7RCJiP1hpW45brvmWesd8p627h1noykTJndvat+Likv4ZmjSxct1
asHkPrNiA2MyTHw7y9ujXBJBo9U6lR9gHKZrOlk9BP05TnbhppSbncy+8jNC3xaqctAu+zitsEOK
NVdHXqsQuBeK4OacaYxPvANvk15XYCDgCTrnm1lZMduHGGxdnTMgkEWjLZsd7RutjlRAEMxcGPYa
tlVy7mQmyZx4QOy801RBFCqDoitgPmuBKH8SC/uIZzDIwOfNrofWG39hmxPDQJnlS/YYOA+cXjFy
0wiR7Izb1X+veY+OpQSHANCOyVzvmN4UzRlknau0A3WhHMCzxNQ8OG2jilQl5kpI/CdIvF0je/rp
WGInQbriEqKHDO1cS2AKR1pi/KWsQ05Z5PPsT20KX9kaMWQRCIq1KQdO0vSVCGingG1qzi6pBs/p
DzKLnx5MRJSrf03RWvNFQ1kGHLZj+rElolHe/z73SYOtdc5fLScnJTN7vtwEAL9wYIFqviVxGN7/
UbkG90yKiBnwzTUg4ysHkj1+QIUdjjgleG43C3FCAfXETCH5dVvakNcoP3UfeVIUvkB3soL9/qGZ
zAjig/U5Obt0/S7SKj2WFZ/1pA4mlFq4IHGinWqZcgfQ3a3DDdQ8sbOAykaj11c5kvNL4iXCwmqs
nGYCr4vMBNDcFuImqFvuiNzNSqJdxQaytJmdESpWbwrI3+qX55YMDrnjyAhQKWDIfa5yA7a5Wbyb
llO98UKHm2F9wZjk2O2h674FzFwbxKpZeX0VaniuRBJkTiVcPwyBXYwtINouzaEPqNqrBureVcic
HW3DyRpCcYrAhiS3D8h0RzW6cubGbH3WSDuuwtN+U6Zl6fP4+7ao1I7YmPJ4Vx/+uuAktj9oJj8f
lAWqdkgqo5psRgyo8817SRKoHVInIU/ZBMlbpmHhPdNQYbeHdCPjEgNINgi0LyZt03s+xcsblHwF
IXCLlRznsZEFm7o7U4maG7Ekh47NxXWKPpKoGqTgu0zbysTefE8DtMta2kef9UNek92lGWkfbouZ
vjlAvZicYCySIJq6jOO/fYNycM5fStE6BiUdNhrOS2NYT/EcdL+Fy8LWDKFp5RDYnwSE7Bc2gxTL
y/geTKvNY5xihiVsF9sJ+/yv3GdyT21Nxwp+vPgzEWpjAi3V1gQgnJkGnrwc0yztt1PgNW9pWuvh
pFLpkBpxnTlnWn8/dYN7mXRDoHMJ2yNwPIdmkG09orXMMKbasWHkeE1BbXKo8HfbAlaCR+s9e7iV
PMOiB38ejNi+/lJKIvR3PAJdOt32iFMbrEal3wA2ZNwR6Wh/qky/a5aby1TrXM6PfXlcImAacONa
86fCeVwF1N2a00zpwjxFQ8WvymUL6XQSfNWC4HPu2+jL1G/u3/1jdkXxtp17GoBFgU3qhiJhcJbZ
PMSBR+YSmyB97t1AxX2dumTNSU3nA64Fyj/LTt/eS8VjjUjtQc5CHKWHfFs+aGZBN+XJ9IWQjOIV
vl1JTk2++MPslgFetzc1Rgm9y1nvpjklQRbGkZIUo3aZv26hFVwg4wzdz8YdZ2X7vYozhrgegusJ
mMAuTZeRmTUEQCqb/iyMx2/8olt55NgXEF2MYo3mFQM8oaJqQRLKTXi9GB8YTPywEJkSJNrnbyRh
VZWQL4tFIO4vUTzR5bV5c3k8Vph/Mzyr1ye3tm6G6Q9Eg3/1H8ZSZGV1YTMm4oIImZMw9YWD8Bmg
t1IdTnOrV6kdxVJwUMWYLaBziUnsp+6hHBknVDDDCxeJwnWgNT4h4b8VUKGBYs9n0ffiVNwxN1XQ
wOcX2gwXA/wIM78qRLHw6cda0153t64WzH878or8LFXnJC5yFIatB06I6QF4k758YCkqdHSZyKm9
9OZ8Sxr3E/MAtyxE8WyPm96MajpU9Ca8qgHY3OCaw54/7997v9UcLyUm3sqztvPmcbvXK9KFJw/G
1wlpP1SXD672xeFl2kOcxZaSCk25Gr6HxiLFFXSv/hoNKaMKyz1QOZSyWbRYCsmnTwZG0az9afTZ
0jO/4I3uRi75xAvZes0PelkkyX+3dwnYZ/DqHpDuoFCFK38r9Y2YwYC7E6c614uORlf+NUVvvVTH
/4wKjLqhus51B0patvRYQsbt91bhhVn50rPxfKDBoCM+rEn9WyUSikTEhLyP1P2PzdgFTNY31QZs
o9+4VhnaF6Fz55Kz2tvLyjCE2TFuWhiZoDDRjX1LXwr0z/YaC/LanmRBUm0RPJq97VKaG2QNtmeH
b1YzcsEpd1Gfot0biX+tBsPnASknDpbtzH6Jx7Js6LZkjxeW2GeaX8wHxLsYgyt34mAPAZB3jN+Y
7fx0zW1cwXcTeeK4d77obT5z2eTahQppV5p7uSkLhh5/ThbVkELqdonKDpDH5BSaeZEgPa7jCrgF
JHn9AZuSXNqK+AFu2ryTcLznD3a3I4WxdPkN8gagMd7LfFE5AUj9ZNLvN0ZQuKOyesTIIGzRahCx
TnstCy1WVp3/o+oRcirSYI5PJU+0ut0Zz9NB2X1tBWUpecRoUW2YxTV+aHszfr8zhyj51YqZaixb
vnZhOIlLqOIZ7p1TYu5eew5LZv3N5bliBrkxsBGM3uim0yWjT8OnFOfkOxmLXRu1y6XPStfyAqdE
z0swJgGua9osdMA9mcNOZqIcRj1s7n5tT+E81vmGxPoJm1/PkgUCE1e/dLsIWkESrl2ddqlOR+5r
eEWi6Z91ut5W98WrG6DhxV/Od+50FXt5Wn565AK5VKtVIbUrMHggYew1TEzm5jm9hZ9JTo7JueG5
mOp++ByLo9PD32pneTeaHn8KEZueSl8LTnvfp7ngI/jD5K5IB0VPyP0p+XYFmFtpKZmolh+NXbxp
3LdIbRKH9Z2Ck9JIbxePt0boA0Rg/olFaTN96ZGoOIm4sXJq4PcIbdyhqmquLDrqap5fJiWZZXfw
68v9BzmOYTapyr7SPbE0YhBTJJtMj0tnrfn98TjgWYOYqGqS3Uk7W0fAbyIWcdLBNAC6ghkjOB5c
qW8n9ctg5wjdVy5RYmyk0IUET40zrjyRUYe1eS3FvSXOetFg0lp63BCStsVdpNQlNwsZA47ibCJ4
sJSzgzvdw3pTjGrZiMwrV+zTtFi3Ue8A8CbfYGNcIA1731dBLUXcITLsWj71qWT2SMiS1CZmNwOk
P619z85O2EAcdwJZZYH9uKIlLTQPfxCl37HTHn5rbaWYydjXOpnTyEX6jg9MXvRLY0m2BtTr8Z3h
Uet0ueroCTG+rhssS2Wz+wsbeNPX66vZF5ehXPBdTAJnH3lRIQ6yp/G+f6fMem4g8DpXVlolc1nj
d9OCEDQzpNibAOQFlYhd89j3wJplLwWkh5G2eGNTHjmedLk2SfbE3PN930tWWOjwRkDpHk1lubVc
nF+2Gx+PIK/S1tIRyfO0GRiY3Oek8Edoc313XslNXyMbxe9I9bJCU/WZJaajLlkQ1TQFLGB023Rp
mExnYY8Cpd41Whk1tH4/NSP+Ud5iebyYSFOmcf21nSCiZ+D7iYfHmN0tm7MVikKrK5twS0BvLzIe
bjaiL6RnBhfSpaUjzXQlInXlHpE8p0gRDHdwCAYDWn94qF0stzlnNLX01M7vJM57Ksj2jlypE08C
ctGWx41qJZuQ+ehg4lLLEqrJjXGYHtA460FqN8TJh9m/K4uzD392h5Z8uhmm8Ica+UtUIvMfuHSB
hT1eBrZ9WbGXJHu2FDGkZ53zP6oAgjlGLM2U/IYvNZ0NmW7VtDhQhilt872qmvK0y4W7k4r1Xdrj
z6iXQppmMPoAfGSnVPLpfo6/QBTEBCu43hTXPwzObgTDWVeufO36NXRL2EzETOoly0FamasAvi4z
zjVn7VZv5LW6WCwyFLFeAhMZCxWauCabRGd2HMJTGNjKRGUeJA5XguvbZz4AAuZkDBdb4CKkCPEs
VKf2lG4CaLqd05HznFt2YSsQmS0O9Pi4nPCeMPx+Cde5JWwCSCDX3VdF1UDGtlRWFgFKQhvBWArM
xhdV6st4HcDmohs3QdJPM6PDcYJuEXHqXMOStZh+sC2JI+c2/afIMA5CANgCLe8xMrMezgDh9JRY
kJGuTY/s/ElTI7IFFbIfP9Q3jG4qtKOAJlSDKaqPCt53ZLYhQy6el80ul+lnyJDLlo6nSCvRI2Jt
NQ7Lak/NEwICFwyFk+TEaYIPndy++bRoOuR+b0+gNsO8JymQ2833Ivrq2SMVQLWsJ9B8IcbtnbME
JdRAxEJeBpLFPMOgieDIzbTDXPQsC8KZAvPATlSzZ2EzGHnl8wzOHH/arda/fQa/oY9xilLPKCn7
NU9V5JmuyodL0STp58L401FVy2UFiSEwbr5HMx6Ca8QlX7KK0j0E1c1UMaryG6fMPBbCqoTbLSkA
Mp4VvvhaFOJ11HqzoUUsCbifTkT4qO19f75JrYY4XxSzwoYlckWUzRiAocbKW9kF2wGONHVpVkU5
ZiXObHQOYyypU+2pXSRpLqSy9OWM/tY2JjIqGOEU3ffE8zDxM0X2sjsn+ni0krhBgB9KPNoDTlR1
WBWPcTi3psExgIkycN0Kn6EZRDtMn2r1NqH7LgRiyyAkai7SwiCXXJS6exZc3aU7WzKDZc4tPt2+
Zui76pizAoZ6xNP9mLrae/27wrBjrwKbdahi4i3gPWSd1C/LZchjb7swC/9GpbIcrN7O6YABTHR1
GJzhZyBLGRmMDGpCR22I0PCjBZpMzBM9Jr0yYDoCVfujU3kplaMgwutYAj76TTCXjXnSzdSn0sZ0
1rgKjAHDNhqk4/6xChXPFpT9jdql8VFrHyGQSk5znH34mLhATEq3qGPMCHGo1lM1sAR7ujZmxNsZ
Bza1Q5pJtI/oPYanJHkNnMNy2uDnq/IDfWDF/U7Hm5kykDD1iHRP2jCvqfa9ww1/zKfr7vypNB25
Pjeh5EC6wQewSeQTA6Woqo2nMXTQX7l3JFtoCUUkhYpaTB3ceoMN+rQcgWeUWNm5RBIoXqUqt3ax
e7xzNDA/PvXE/49J22UKNB2BiW1eFOMVwi7ALCMUxLbmXYhlZif5JDczg4LvDiWI+MjWCjyIDOFO
V0788HNTPKFfDtEu/eP6vEs67ILgXBZCI+1rdK2vxwTpNVE5/INpQ5X9wmrIk9NDkk7B0Cn66V/n
Bt/kd4K2P+RqBgR7dKskdVnBLeL8+l6Y6+5NvBi1IFCNjg1GE7jXbR9vVYymY2BMTmlYKXR3/r9M
QlNZXTbc7YXhW/XyKKSD8BCxOvJITNxwzAa3ZCdD+agnayzNZZrcua249smijoRs3YMT8QqZld3N
Cz32b0nwhlpVK+QVnaoIaOD4XZyuiNjPYDwxkXAQzczPrHWxJvdS0Wii7OZ+T3KS3jkTDRegy0NI
y26XQbVY+bW7HHOaEgZtHFpIWVjbTdJmZ5JPK6UvL03Ml0BMnpPMinzj/FFmh5tLycY8Tp4zLM4R
vEHIVEefuMO+mE2OGchYDwz8+UY0OAZCpvsiJubGD0dgShw1SjKN+G8s08uHpngyLSIaJexR4qKe
wDWAUxO1FM5DjzPCl6EIKK+YljSym5f1odOeuYPeGetf6bvZhcWX5yqjiv0jSP5xhbr3pC7x5Itu
qgTnjXQ+ueASvCskCDbFuZHJ6U6zL/RYry2ZCBk6TyhhjlzHojSo8bgoUO1aJNZ1dmaWDYzphHXI
BhPqrwkvD4A2c6REo6zIlQ3eDAAjPh0X1z/ilobLpHTkIsum7FOppWf0m9XyZ49ejwgsRryxr9QD
h48A+f8ZMGTzFcAwnsiEaNdgkZcjRIBcRK5Z/tqBFchLl74sdxIzuie3BscDX4fiVuhMji+BY2du
t5XBKvLrU3gIrMeXjL5R4JnvSsfBn4FXYSfQpYsOyu+HT5NFsImaVXw37Vb/1T/ANoE+sbGlSrb3
VucNuJnuHwDoyfNALinL3lFptH+s2n4bl3o6gLybSnMq9XX+SXwLou4YwQeqC0GwbRPDxBigTxqG
fwcSnjgOB7fChZBYExpEzYcKoWNRwbLFGAELmQO/OR3gVWZvKIBL0PKCp1ug8OwiXDMKUoHf7TPM
pKrsxei81sC0ImIyMmIfaJJHHxqEsEZcMcyRodgxbNyhr5YaXvZLcHgAoZu4cN56daflstsHNXoh
p75llvXPC4PSAocJoaoFNbiVgQtC6xsUvzFrOFvIm/MQLwZIDaG6hkg/mvSNw9Nem5bkzUZq7cD4
eD84k9uj1yZWL61LiE8H5fEMyg3I0HqwxPqreWukFAfHffp20+XqhUjP1+FVk1wcasqyQtXPsLf5
amPu7g4dCVG4Q9RthLt1fQDvwCDT1yZs0XCwp1oIm78mxsLCdnjyh3E6J9oydvlegtk0GvQwrpuP
0IKRrIG4Nz3Z28fVEyg5uSResfjQEYJ8swPORwJ5UI+NQbjPBQzXYNIuSPPlwJD7HTEsz3ahBl6F
Ppx5CLY8PX6fPw7oxItyN5mft7t/c+lOn7lGcOOf0G93JJSBqMrsUKWbqhR3jHQBhowWSRY/sI8N
gr3Ra6ZwIY6LH3oCO5/HHOJzILqQSUVDpdPpUQn2yL6bBtAOgqDt8oPmUueac60INYLG29K0UdRj
Jvo55HXWWqb34JaZ9tDPHmMGDpfsuLV8oUGKrq5SLUMhznnuz/hyep2m65No7LRA/WG/SXTJl/DS
yR+51ZUzIDdhIxrSDOBgHO74H2rdB13HSGXkMGHxKobORMH/0Ze82rd+zjQ1iabCgxrZDSG42ieG
O7PdVZht5UOa6rFFGSSngPndA9qOIT/DhJiMTjtHTBENye/RWeXNCUjkbSgO+RLyJMw+85xEqCuz
9bafg6Qnxt4RL38CbIT/bL1+YNB0iTgJLXhBwv78wvoIqPYc5x0K7WbzTGlQ+4S0YR1Lwyh86BP0
h1Un/wW/APGUJFXzck1fJ8Zn/bq2CMV4G/S3p+zkQMvFBUPVVBnJ0CdACNc/vDFuL1gNZEbUoU85
uqnYFNnUPa5UoC8pxKjZlNoL5Wo5bqrB1RNr2LJ6++XYjBqHBnmICXBApaVrrCeO2I0qVybONBFF
aTpw8+jIZ5uo4Fhk9e94LP4IH7h+Clj7FtUdp/jt/N/hmtVEsQ0RmtDbDJeHFXi/ksvkHUWkTi1e
39lS+3hJsX+fj9SWBZWfqXvbKFerE9QBp/sIDyW4gKoSKY9piedC81DseygprLsLh8qPnvE8IH3S
mKR2bUSsASsuL3f0P85/4nDcYnExO9Vj7RoTGXoXQhisL7MqVlp9yJ7nvAxt7ljsbVK/zUy/H9ai
XSzUdJ+zvmqg7KSmrzr2yERnRr0HoYuWgJwPFg8GjYZJaOgsO+Q99vgU/sDq9PIFO8IYvpu56P/R
sb1UkQkaPwKdAK1lZ0XGa/uYYobIkLvqbD1T5JLv8mvg7ErhRooC49Oze2oeGuoX2/vyMzywxDku
NOLcuHS+f+tQTvMmZxF1h4lxjhXJ7PvTSQz0jLdc7+h6+LRIobuKDH3F4vqczXbAyevVxHTC/+TK
yK4EwK5zN1cqyaULYGrdY8hIETEX1uFUF/TDLrahSg/2KZOsnBj/7zTzC0+aUhJOYZX2NnfCgOHx
rASC+GeozRxiROVex0RntCbrU/lX9tAtgHcYgK7r5o5/wFXq6uvV+Vb+hPAdVnT+0vlHbjDmZyGg
7k14BD5Zcrchom8ELbkcpqKeFMZPBWetVU0Aj7B0wcsxK5VOf4KP7f1IpagJu+SjoPBNn+xjOozI
f70S9Ldaqy+mXqVcZ+qHN8ZnUwNR1EWyTszhn2R1SYwzOyfceAlsH6RT9tJnhN2bEYrH9uqEmk+2
KXZsx96qk0ZqsIVCdj4APigAncPKDQJoNrBiE0nsFTlzaZgAlK9lCm6ZZ73e9BmdcR7i12K5WloG
SS/cyioUQ9OEL02XGRco3DF9F8zdONPi8mlX8xPmBqlZIuaa/dPbVd0kt9M7uZ2LVMhVQvw2Lt7M
YbcxvfH1OJyr90yO3inVNKVbFuXNpn7CdmZ/MG/7u7CuS6syQP+kXhes7d8E5AHBaeq1kmTtE4S1
s7EJpchQhlQJNPqmqFuz1HifEW1e+RiLKs5zdJSkyGeZgDex/BBNrRk73VhcCWcU8SjnySEeHuPR
inkh3RejetZMFTDnfJQRyJZR/e/hpat/Tu1aWsDkOtbsnsYcGv+t+k+mpFleWE45Vy+D8iuBJI8P
aClkm2JlEbj0t9OBv0cpdtd8TunQgvzPaaXjXJ6mbMOiN6sVZaXY7BRli06xKqpyHPxt6V8xUcRh
e1Z4GfAKwYePA7ePL/lMXG/s7oSU3Cj7xPnnp0SfvrPgeDjL2Lh7dH4RtOuwAFFDEmt6cSdRn8NI
KUlYiZ+5V54XExuZ2Aj6ZIXdAJdvkyzHie8aZut4zGSYxvCzg9zHuv7v1tJ62//eytSS+v/74EQp
hBXdiqLaT11Ue+gwR2RN4NOvWpqTSuPRH36a6BdKSBHo8weJwm9GjAKlyFnz/wC/xXYrSkIQfJsS
3zyY6iei8Twja4E1aaxXVx3is7k13JV2/MNyLcw9wm3xTlJKPgH9Of9LVniI6YLtyHoQu+RyECVL
5dLkvTtuwJJiK9WjIlMCh1Kr5YYdxTSpDYPL+rbEJwIHFsM/57Oa+SkXpIXoG9aMNuhkCzIwZ4az
onskvnmT4VUaHTFVE8Jbvj1yCFG3eGKmscLXedaNMdSIoPTW8lfQ96PuUiMFb2gRtv0NJBFbS8eT
JXlNwo/4VMCDCQASoR0erDZEyQkfp+J1sNK/PFXYni1MRpWX17KSd0zLp/5owqjq4jlg/W1CQAQR
tpAnC0DU/h81yGIPhrPul7Tt0gUwdgx58LXu5yEJ9xCjacg0gCDoBOkZyf3FqsJRPbKR+fiNdNRG
RdztQj0TtwGyLPk53KaA6G2EEy87pKMGSB31Phn2vFgq6QvgnxASiSIJTtE/7xAcgSmRZhKEeqp3
/c4Y/z+RgNuIZUg/KhVmGn9hbf732QifgHbq1xnpVf7SNY8HnSkcdS8Mi7hxuad+jCHMnWpdV02G
qH4m7AGIEls42Oo2vILP0OF53vAeR464Xpk8/1UKlfY8O3J8nM0w4c/sEG1LDhtsa41pXxdoYe6h
RneQ/e5MAmKCQqPtDjGeXu+Yz35zaBGugwiG04dgSoNIBR/ebxZN2eP7S6yAFqZTkV7tKe0+iJa2
wFlqBVxWEAq3xK7y5IFm/0usEFrEVwfYBjT2pR6Bhx5g1F8vMRSVRf7IorbpCJvmVu/V9weqN4kB
KcCHCB/7nDt3tI59dxpRzVC1tafKLHcR+3hOictrEHmfifLdJUoHLuDODdR+3ElDuD/AxsClqAuZ
1yX2963OyBfz+Y4Vp2EOxBOn4CO9Ziai224O7Pdpcthanauau5PvFxhUJEbRB6eUdjNryYdjCmrw
pKxpOpnNcbwuus0njkhTBZcOkeE5ROcMzxSRLfS1sPhA/aph4jF9QuiYFrWKJh7XdngvEm62oA/A
Xrsz4ukinnq34naS0G16kJ6kWe2xM3ZZG19BOoQ0hUr9TMzQJ1JZeg9HCNRpxW8SBt47/5ReJnrK
M1BNND0GNW2KbERaNjlOabwF6tOO2UC9w3uL5jCjcu6V3Z2dj/sWJvQaJLr9UWMCQhQd+PKyTxhQ
HzcQXaBz037Qh/5aOpZ+aFB+lntB2+i5RDoEJmzNT82sAVPFSha/nO3hkFJYMaeYI0IpTS4uee74
7g0jRTVMZWZ0uWB7YynzkYyjtH32xsxcBTEgM8YYZR13B1DGhtGX/aZ/X1SNqTs8ZP/uQqpi7BuK
Fdl0rhMaOh6M6vk8GXmGSUnq5lWZDg/HVKhQVlpcsrRYq3Sm+H3v4q4jUvxhfXVAjs8m3chE/IkY
SUWnCFfKs/hDSoFrv+DVgtzY84WWp4z1Ae4NuaN8TxAhUPYsPj20vMAy8WPLQByMaPigE0wuY3Sq
ZA7B+fghyCav90N5Wm4jqyUr7tBJi/w768yGzBJco8ofZ80MccGD+rKdpl7rNZ7tRc2DENcgpVTy
fCzv7qBz/sWakxQ8BrBVLF4s+5xkBPBj3BSUss68MXUfmZQF+HJ4Ox2hI8byXs6O4sFL3a+iItwb
ECGY5uzr/sQmE0/QS8QP3WFKd+oc78q6y+Fnmpd4ZzrxhBwhuRZ9DIU4e3cCTPER78UZ+YCHNIYk
6225R4ozaCzcHgZA96IxkN/HUVyH6V02SHlCcuMx+EU885QIbBlaoXNCAaOW7gvHTFmP415GTOiY
cbDpjcHWxvedO9SATURYAoznUwv18hDoXAvSKTQUEppnK697/D2ipoJKBayiybKbM++bVIrxHImu
RnebYOxjf/DcgJ47DFCCYt80oU3MVmf5QqOfMB3KYC3kQ4FSxbYw59RLY38R9Fo66SPd6vhGp1F3
K+1Cnk0bux7kMl6sWrhZOe/MuhEh6AqmYvbh6qNJlouCdDiA1wtRgEC3L9GTcKCBDEan8GHljM1K
AvYECgvyfUq3bZiwqerfwKk5UMaLTYdj7vzhuO5P5iJH25yg2PcI6WHMf1hzVmQSDSOU0aWCyjn9
kBUWyqOK8pbjeYxfWqZJpAudagcg9BAU0RAL+kTII3zRU94HQAQWu5UoZ6Wx97n9YG7RTVgwyq3+
oU7UQH/xth4TiwLF/MIMN7i/dDlBv8Am7Iyy1onzFVauiU4FH8roYH8CCTxWBiZ0auLhhCcyNjpi
1cl1Xf6QnmuB2i4jQQDCKhhHbGX2Ict7gEftb9g7UZv55XjCoAKnaW/6KX0BpA+5OzoqvTv8uEx2
fPMerR42a0tOU1xw4aZVhFNe0ACi/5TrUrruWhy0gFEtEwBVndHPTch6SlnqYwRHgSTc2pW0jJKy
2QKjNlEEQnExwXwE0unvpKr543YAcilCb0ZKAw+RLgWzaEeItM/zdjQqFkG21+BLVYGKhVqk/1dV
xyP7MeFbmmcfkmLZR6fG72izfUz4o2DKHwJ/F6aUAhJYC4ENIhRhSmSmV+Xo2q+nu0r3Bp3p4NS5
Epka+muWQagIa99vFjbMQpmRseKcvSq5aX2CPUe9/LiWB3txb5f0urW4+M2rl+cHow9NYwPaqMNu
pfHIYufL3RjZNRXB0nfithXFdoF8fPU5BBHqhjqMWBP4WMh1gCBw4DPkpA03DTFAJ/+95W1GKrTk
MmfpgjksWBEBoHmkN49jeX2tn6fgpZWyxdShXz4QNfxa1187qedGbKFobUTLobT5MAbC05Bk1lOi
M2mDX+rmpiGAchZXJT7/CKzTAI4MeQwtD+VQNZKhBjOaf7HcW1gYaQlmFbbRjjw8FCk9/vQ7yXUN
n8WER7nHiQME4LvTwgJA9o0R0aSE4e59DkyyZ6n2Kmxr1NeOe0UjoRhLeOD5ZJyoKGYmTPbIGfhh
t7FcR0AtTiYcEKQeietXMYUl9Fbvof9A/Rzdj52M0r88Lt56WblbfP9czDzI9727ZMPWMNoYTNkH
sJLwHn5Nc6+2S8gUZH7tT/O0flEmgzAx+AZooRiTTUDrOef8g+mtlYMB2r+ociTIpqqK+F/2VHGM
23lUWX4OYl3VZqtgpWC1QPnCLkNDYNQceiF/CpIu+Pup+er0KP2iG7uWiPqPVA6lmd+HnTBSd99k
VwrQJ7ryG0yfpe7uaHPnWlek9PWl+RmEpBH3Mdvwjm7K/N9cfNq8ijF6D0q5ayMgtYAF2vCgmZJ+
EbhSgnGm4ZLdPPZqwYlYL5C2El1wdkbf2N23PKK2n2ahqjt+/BfkyuBBnbFtBdKJKzvy9PDJ8Vpd
pUaJh2ZiVTPykvaQuJHUTXEyuvWeQ5lMViuTwOMaaNKAGmRGiE6Kc5yTnZoV1WdD4tx1vzoupWo8
Dj6BuKLYFHdMfyHMd2zoT8MduTE6R+l7QQ9CthaJakWSrLwiGCvfNOeB2nIwEoMXE1cUHpg+QKBT
XGjRshX8RxI7QrTGNzlVfrBhvoQbgTmN88CP/G5OSXlxxCKAoTqfRfu277bJX5hVf5YbVLwQxJPM
xdCXcZLw5BbA4obFJRW3QLXa/zihNiFnJDF2yPDhL9S5vSTAaXex3a4LmJv0rywkWpJC8PPhQyVL
oux2V8DSM3L2b2Y2DieGKIK+MQIZm7VsTFh1y09BywA1lptbOnc5RL7wB0RzmE6m3z2s1O1ZtDP7
pCgEG1VPrLyVtwq52W38PIu7ai7tUvtQdcTjUWDDW2g9PY3A4pwURZrLgaq2VNs7bIbPxizxfnqY
Ms97YSSHAtzpKnh+u9QbOAqCliDngS75UhM2vPLSKuI2iIzdvHpKv2rrK6z0lVGnpSYyfBaqqsNv
E4Dkgu/ITZp+RMyRfqBR5OT3PI8/ZKowaygCFtJtfxon01mtzVvv849iP7iGb9/3tsrjnxPnTR1u
NGwToUohcQY9dI5mKDQsPMC5jf4agH4RhNJdUieBp8PsebQwVwmJbdZJWElbQ9eOOBBjX6CDSKhp
EmqNTjs4cnqh9z7rCPvtMblvSk7TaUdFjMst2MAOFviO09fRIfkJjUyLIfKPzrrMWR0WAUzrjds2
VXTbfdD5kGvAgcADpd1W2R0J0XnQXGzs1Vvmy6zKMdr18YG62E5hUS7Pbs+JwBmB8nbkNomjScqS
Esbc2pnT1umYbq+UOx3TWVHqt3UomaQQHmeJzLtIFeNUIZuOBnPvVymI6zrjfwvmeeEfCT6GugAZ
DI3qXIRchXmlYkGapANHwOuQj9e97VutsIJN3aN2gGRlwih/J9K+qsu6ueVYTPwvcZ/X75XLMnuW
osttHF4wQ/YUpsuQ4Zt2A0RIZY+3F6j7Km+uzmlY6dV81RYVn8LfjcaLg5dLN7NGTc8cKuizj5xG
cUIMM/cJA8aBIieDOPVhie8OOW+LD23wIfknYKAX86j5rE1os5NvaBdGud1Iq7yTuBo5ymV6zTuH
ul67Vtr4YycLdMIxoE42RozdKEPWXZOsgp95nxexgDrRJmrnLW8NLCECmxKp/VvWBf1mQWrc8X3N
B7wPSIK8O0SepBak2EyiQwq+fbPncXdd3YF45MNpr9d+2FE44XFZRL2vY+hDh4KPQf0XKT1Rmwgd
vSRqMfsTGjrMJnKtXTvKs26xLPKjpMb7Z39RGG1NdskPMSzC9Szk+Onn56r6PpqcDGIAYCj1weCb
Nn5mXg25gkW8LW8VKu3wEC9CyEUTmNd9pFBxn4v43FierB+XO715z7PcMJKoRCIbmJd4Hf6wBRr/
CcnBJ6wzN9IDanv9DHo4xJCLrOsuFktB6KuqD3Q2bnj//BbsPQzYormZ461N8jDmFTRi0w+ZaDCV
ZpL3f9qiJ9PNvhH37EyirASgCwJmFjdLnkDebb5JZDLTXT9Y6z7icFxXBhoe7+g/V8O3PuJNL8Tl
D8nDWOzfXiBH12hSqKA5hVDPSQ5Apv1iciNMiytoXlj4krqd6EgCNAxYna0/G75vR/HtmJttZ99u
/p2qYL1bLPnXLjoFghW3/0wbJ2VoPyf3ytMduJBddIME0qX6giw6bOzPbVff7QFyvFOCnpqOvJJz
E78S4wODugZ0u2V/ZKe1LFoLmdetzBC8tAbZJvbxWRswy/Kux05SMpiTLIUnWRlzhpQhqdp4KdhL
HjL81epY7P9T0dLS0MhQRCLD91Nbbvn0IbS5dqDux4obITqqzer+qjyLTlX3e+kfIjU3Fcczc3Ff
O+lU2yI0tsWP1X1z+yBtAXpBIEjv9FriqjK+9anrXiA1pK5JP/aTvNgRJm9/a9NE+gNZFr7f7bG4
i32G4H371nCx3maBSmELy1qQnK3mWX/s69jx9QT9c85AoGhrMtrVr/k14F5kRTHO0YEZICVkNpAS
US8uLkN0/dnuncOdkrkAKBR8Id4bVgz7fjLdMMxFSb/NYka4f1si50dw+UOwe6Ts7ojmFn3HSJyE
hjpcZjBcxnkuvVVgmCdphU9AqBJVgQ5OEbflfTVVeyI0w1V+/a+olXfHnNB0tLoqGcOyQ1qCNfdv
l7R2OYh7irVsEl77x+Q1ykFS7CLCHmt3UOurBq3XBYOaTIKrgoEWdFaSIUrLmzGzwpQsDIH81WNH
Tm9PWZuFtBWLYdj3R6VspGyvHse1wMDVrJS5sKzP7BhqysIeFfOJU7q184IO639y8a9RGLlXXuHW
vAcPd6Fesm9WdlcZtZe/X8sgcLbrmV+iewIMow0HqIVZwqeJ0rmxwh+ng+Erm0yWxdV6dekY/F3O
9RdXrAJAw3+fRhQ2fwTYKzZrlIdF47XI04Unvw8AP7HzFVhMvoi+Y8OOTpteB2R3PT9yYD0OGund
qI1bldl90dNPVgku9Pev4Fbq2hir57XJu3GM2AjFKe7s4z1c8GlS8/nJ1V6In3VDJQaR4J4unloE
ACIcrQNzxEPi9qeMjU31RRRKbfpZx2+4HXQW474TMl07RMs/LdvioPX6QOjpoNrRRlqkA2JitQrp
0BTAgNFOEWmReVhZlFjLodmsNzlvJAhV3LApxbOD+ChjiHGF+5SnkVG5BeEI+cOqdhcC2KXCCCNN
BcWqZEUndnrxj17nDjnEZLnrxpo+JV79BnC1DvF+Bx3RyQcSJluhtt+Ln1f6aUEjp1+5w2D+ZK9q
rP0sACoehXGwfcpm6gIVJ7LoECm1XTM9u3UA/HxeKoL3/Mtu01rIS4I0XVWwQhWI0dP9vLI04uFP
i2wzbCpBJqGVZ1br9QUKOWCE5qdI9A8wub2Y1cycxdL/nefhe/Eh4yEkeQ33bgo4FiOrlzuRT24q
hflV9ihyT8sy6mF53ks1VG6lhpE9Pmt3iObJdN77GUD5ALJ34WygQ9A3bwy8AWdDJt1Jk9dtsbZS
XA4R5eO0+puPgNfQ5SLIq8r+sWNMHgkdJ84wucyqYOJKkrf2b8tE3pSla2JrzqZSLZdDwmvIV1lB
tsQI4AAsWcQgaeVg85Y1tkK4GtKmWSTnpPnd/rvOi9dPO5HYi3rivXYVDTzrfYe3GltjStkwDJgN
pHOiMKh89W3klpHcxx8Cot4mlVHSarPO50uDrcUikCmmnqOmYdUdTEZThheQQY8yg9gHSago2MXi
TOsreFDeZ8THvnY9xGLerE6P3X2rI0g4jY/DVlZIeT0oZLFF800+9N5BTWCaISYl2EtTi9p31UbX
q93oGUJ7D+BLgR9E5iqW2lPuY2aKDQ+sG+oTD9bbP2GDDcDqOU6o07O+k4gPB8SoH/4dSSqGoDvU
UvlcuqbkMITU2TXbIWPz6f/lKFmPGjAjIfABFBlaJtjpRlFtSHiDcrieIuY1mjdlXKTydH38h7ok
ojGgJJeAaSHVQ3cE12qe10NPgQ02NvH+HR/4e9p79Cxzen4NktyvNNaptXFFcWdcjNk/I8c02S6n
Dg8HZS8duI4BgY9ixTcI6EW7WDjDW1YLEFw4FrqYSzjdc0FjE5yF4BZcqPyi2Yj6s2rfMEfaypLU
wikf64CO20KF2ywvvNhKEqjt9zSlAJSsKztOrqAamfwAEy3QwBK4RQRh1V2pIX9LFb4JDkIb2OvW
YyTu3Kl84PxPOhBr2AixD9yOIYDR4Gb8V5lducSeGYDJroRQwbSaYD60lFVnGgH+SbufiTFOBKEy
3rW6oPTp21/vYl2tDps/r6z2lmYEqgAtPGyDrJ9nR0gnhmMOBln1gKi9fbjsV8dlyT+1gnP8waB2
1lAzsYWkFQDZYwoCcMTxeRF8o9ZFP0tixTHFTcEWmPCkZx/MpjNAy87VcuJ28eKEQMz/eLtOGjZ8
KfCGHtasC+eGQVTjk1eztP4K5aRO0xiMHVvLrctBu2ptIWax/k4WISZnR5+Ak8yhrPgTYNtZBy6p
chQd5uXmD480CIs1co0zrIwMJuoj/RjXbAXwv6IG7Loo7+OzrnM3b1QgZmoFXQ6GVor4jvViHX5k
TMYdqHx5ReMyr8syxi9Pr0C1gL5knhPYl0eWTOtxduVHzyj6tkfnEAy+iGtdXfn0D1bJzx2lop4t
MfKDUKnvIcWqYq+ZKsAEp1uBWnB8dkwxgPzQthdvFtSwZ7bZorrj6w+TyKotxN/IxRk90DWFk6G5
Z0it1kPyrQsAnJ1D+pyYq2IOqv4ejFlmiKZ5aUe7apYmLebbdLqsDalbkGOUaNe4ALAPL9/uVo2h
lbuYqa4rfbtvoP2prvo36s/Vfxf/F45N10uimhQ047hTfUapvmHeN59Mhl59UUDyVFZmH8AZ/gxm
XyiNG/ix4BGAXZaRiysFvZOmNvFaGBGw2ufO/7lsamPwDMae1+dbq/dPqjXn9ddNXwLpHhrXiUSx
olPgz2hNRVbbRDhE7QITAnooT4U1SkPurxKVsPywO/Xyl5jJ0cxN8YDslEs8Qp4mhRsIPVgVIyfh
RPxki+lL8OdKLlAvnK5UgJIMyaVePrKWqOiKO1d+ZcHQ2fE4Apauh+p6c8GCF6xat/ZNVhGmps5j
jCW2Jakw3PxbNpmfTBB7dZN0pNM0XUKx8nj59SDwXBL2xSIDc0UuZsdnijEBH59v+ab/ACJezyka
9xo5dYn0RtL1m3kacHSQny8PegtTpcYne7FIeAaWVhkp3CJ9D6c3yknyYG0NQCgUpMOtWuDaNRck
etVFbSc9yjUZ1EYUevekmvHL1oAq373WF9nQlSDwPt3e7aUvIBYP4u9Lg7lmcO7EtOKmlUJrmrUH
rmxRHls5dzxX07YZQQDHIIIYgtYY9xuKSlCdLIp0hQ2AgOhEvUvJXB878KK0Xqbw/fwFNXsynjEQ
nQQyGDSNZbiMrzg6JwqL6wVN5byjRvBNwLC/sIWDTKjYtnuwt+8cMU+DMOh7tYORMVQz/V5A5Mz4
n99FaPHiTDjTtVqmEn/bQoffSPEYO9zwqKGmumj8ojJZpVQsDJ2heNiMgRHE/zAjV12/vuA+JOJV
qPK2wfezzbhwHGY24LODFMcNxAvYKpL6SMSGmQJ27VyIMNCQcXgCM+LneZ62VRYN4P27Sa2IxZDp
0JB1vgVEf6DZd7+p2ZnL7l0z9W3fJsVuTdUyMr9vA0KOSYTGD8jd0mtoC9qzDsq9rXxQdoqD2Oms
BLMouwIXMwNgJsvtChavxVBBceezKs7KP6qoHfqb+M+IRJxzMS2TUuGDXakXCmnfp6S8sLHlqfa0
ilKFg2H9pI+DXYRzC+q+FSpY3UBuvP0Q0i8LVP3x2Y39ZbPI1P0N/kUOoKob5DilWsxSMVAVQoXX
kooyL5iPlcjG9Jq3y4ceFqqwQpCviipBZ2O8jEsNjekx+HHdSwXK8VddsEPOtn6tQDPEopNadxiO
c6Qr7PG51bfCsZId4H/k9HNDifgtf+8mv5QHOl2/r0AyeR9ilMyKZNx32YkqO95ooqIVQuDGsDh2
9D04GdjiHy9Gx0E3L5//a2zvlOdLzYbJCFETvB3DfNK+37pwmGbX+FSHyRlXx7zDNSllza0UCge8
hZOcaovaeuAMxnO7PM/ZioLBK0bIZDK3YSiPEmYU5ic+/BZ2BvVzB4Obx0I8ZGbe7RlE9jzAf5iV
En7/dEsXyMFF5+XSt/OOMdcBu6OZD8E9G+cu9tEaV2XAR+cEr6/UVb+reoYKcCdh06j7xHXsRINz
lJtslhxEYgVwmFFYwrb8Ma8C+23DIP8LiLd5JlO5C2lQquDT32JLyoLFDI46DsMxs/O3U9oJF+M3
r6K4SfU5R1WKbGwiE9SCkuo3wrIZGhVcA/TAb4uw9PWo3kxKiy9rO4k1CgeypHewATORulFnGnIf
BZKGQyGDgXO8TepcOD9m1d9GbHot6lsTkh7giWBu3fJN9sZzahUD4Bwjp5XksBBPedMOiTteRRSe
LN4s5KGU7gcav/xYeWT68wBE3azP0oI+BBLwLJcU04/PgOgSISWqzcbb80LP/VOvqJcVj+rxoEHs
jt7n1xa6lYQFSgRM7Svb1/hQsKIRY1eZgsDpUrUS6bJJBYnDU+7FnUg2/fbQi6YzPIWIerwboXCW
gwMtnKJjzS07w7WDmcdzidp/JqGuG+xnSC/MqNr8cIeYWAMiIA640a05pV60FZE30gcYkgj0/2EO
ewTCQBiKCpK9RKVWyLyN39qIKftMp2uaFoE8oy+2iE7WxNkyYlvAr4CGz5IE/yuEtKRqXvTkWDG5
ui54D9u1CDZZ3PAlESurCjvkc1xGxDQvzUX/OYpaYqqGug4w1NA9XyGiGQ/Npmd5fICRmS74pHQe
ruq1E3jFkEAwSB9HkXyJvWOqhl06OSOe5sThdBKS0/iNeXlO1h/8BDG2+CaHhH7sEiPPXARp1DHB
3A4Z0knN/pu/GqXSXfiQ6SPaQfsyjzqLeLygdUoHBMtcNMJDg5nEbhSWWz4D/0vdvzCOPulea5Rl
ScMV6dyUOyI+xmlWIIPPC7lFrMMuCPqJWepdSxraR+qDWGVMUyrpEX+LT6Z6i8wt2SBQ5KZEex5Z
AWATP5PAR87ESZOLY082eH07tjLAf0pd8KvVvoA9hRQgukmpQmfKAVKZ2vSu/nJWnGbQIUSaVOIM
SeSqBx2H38N7jaJaph/CBDB6eUzMSITtWSK0jlKvBsADaAYfjGJHszTnHavONE+j19D2npkNzn48
qJVhgVxTwK8Jj74DFI4HWOB5SF4JnEklA9KDov9qSl4nr29f9WmNbG7AR7MQvdcuBu9PLc3yhPul
48zro/RTKlkYjinORQgpTwp/LoJpVusMucJ0Yb+3+dPPWl7hcbdOhmd31un9qc43FjTkRZ4qAKEB
gPSHGJ/IukfwOgYfp0WKDtlR28BNkIo1US4+jFX7wmkPQVxkf6Z6XTQjjdBws7RM5IZDPWYaXXuZ
3sFqUougM72FnVBKa7JvVqlYJk0KsB6mSL/OLixH/pCruEXEKB4kmbBcUWNlmjSXT8SSuima/GyQ
jSOvowjKSTNj8Mdz5iwcBc+uXofBywAGbyxKjkR8152EBzSEy8iu3/iM7MUOwve4S+g9NacC9j55
ZIDygpzB231nme3Fn/vXZlZeAY9hK8PUY6syk4bc2oMteugw6t0hmXCb0M235Ifnxl0aBsGmr1iR
o027zrESQW4c8fIE4FHFiQcbIgaxC492zuILxdPLPjSlk937jDWdaUjlyPbXeqBGsYLXDuHG0SMm
pPi318wDqW+CXUpOdYoK9gSifZwSnx9ZqW+9L6a7Q38vA0pNiYGhoFpCFpNPN66kIpkHXJqCRv5O
0Xpk+mzk6j3MdEzQsdA41UrWJ6qMGkfJUvgnHvjsQZ8wtVnX9PwYiSWmNJWLKpHdWn9upkx/0IQr
ynIpHGYvuN5t3+ozIRH+O325tssRxGSTlOaQTmk39YGmqkqGFoUdN23zNV+wJoRRHbRvpIYcZPt6
SrgxOrOe7nLfDnN8+peHv0FWuvpFI7o0Qh5D14ZsXQbX4a9X9OX/heBIOhSzp30j00jlX9ukhIyl
274l8UVAM03kQREJU9/amfZEhor8kGJmuPpoIZTujKXl/SSNMx9QTft3DJE9OkeC0o8ZzCtpUt+n
J3BGNEAX7jI8vtvwAzlzuuSSRL2sBTIPNpi3L6RtSn+NUZnyiH4X8VGK8vpMBKq0Cb8waKBwYHTz
GRSSnWw3mL4kq/g8FwSEk7zR1zXKXX3CpkmDLNvzL23xn5Z5SoWrToI/BaQTD0U1FbngUOGL4BCn
8n7SY1v/nsMrUuG9erSTkJBCXGEBQC4a3rN3dko7i1U48Ci9IwrUPKzS0bQTyvJzkFBsuoszqBGU
q4VZ/LJKGnCYmRwh82mcwenN2XQn04nt1uwIC0dNpNvioxvogkQamMZ4hqQkC/wTV2aiQq+oQ1Zf
wz51qsU+WLZgE5MU4n/q5osnOA/8OQerNjbW7PguEOUBntFiH9HYoTjpf6952405W1j0DNGt3B47
hnVw11S85MKvovWmcoI85R1a2BTH15IPUTAqBwudthxcbVmV2uSCy63x1goIZgiH48o3KxUHCdOW
FoThzp0I1EEBxrrGYhD1SkX5DhzRsboGQPDjXdrMGTJIa7zfmanTLMiogYoFgZChk/+gP0IFyyH3
58CoKNMVarb77g4xxU2ElcPCpGfKEmM3eu3xQe8/tZFEZ2VMnwmc7hoL9V1PjqUeskVa3LorM+RI
FM1R9Rm3GFDUGVMyka1rDwd8q+oLyKI25ni+cC2yUs5Wai/xMpwW/zl75uSsSJFrxjdRvkzh9WWf
jkHjW/JevgxY4GeyCRIMdoJbcvazujjM+2PimGyaz3PiVNOr0e2MarSQEUd8+eFMDwZBSf1gRT52
nNviAoifMbub2KTOwcyUSGvhJRVadix/g94ZzRc2TWzPUcM9X95YJxYb4huADkvo3c9BI6q1Y7NI
7KAQnue6111enBseLmMbWMt1QnbNvlnpAJFw0M2cEW6d1bzaVIqAssSBmueGbaDk4sOL1rXEENRp
Hyd9hGm+CL/Feiw4zs3PWeWfV65q/9Qv8doslcuCIfb9OsawlB0tjfH16vNxQ+HLoyOP/0x9SsgE
utUj6WS4IQ9+d9K2+ffBTDF9PKKUxR3Kz4l+EB6Ra07OHXRrr43AILp9/PBlxKmycwCMFRnl0m7Y
tauLmgvdL522YZtEvjOrCffsKt6twlNUMhUsC7M3uvkmkc2xy6Ht2JGa4JpXWGOi0fo0TOOpXdfe
XCI5n1O7KQslU75mZUY5AH8TyqAp29C2DM3nKRInSHtBRipxZDV3clkR8irlWvBN5AqeYDMFj3f9
4CLjArwn8bVD77skmUX9yxd1kYB2Y8cyOuGtDr/KQ7gm7PpkEX2b05box+fuaMT0aQcrF4SuTXf/
A6SqniF2PziflrrQ6a5F2ihMgGjpAOkg37O0Oa59mM8rYFwop12WRUbPnJvWEcKSojCemfranAfD
Oepy3CghZKjTprGbnk4kqEq7pVZGy6IY9MRvjOGJVJk3jDTCX88of/9TcNYf3MBPhikKNAikNyKe
KSenvnV0ZOMq1vnRS9RQ1Lo8qJBtUC/ivC74V7PONGPEReQslJko1urp3bPnU/nyw4JVUvMBSxjm
2S5/ysY0BMN0UEVSQqIGSJjsaZJ0/B4xPHh75MxI2wzzYoXkDGNBLVYWmp83hCuE9ZHQZiqMAyQl
mUlGHuJk6uWY98JWiFEh5qfGf/xOoirDFNTJQTrGll5B8Wf4ofn7/2ulYMVPEv+4ZNUA6zAAh6gt
+2E/eoRp6MzJBA1lYkxa77SU9eWhpY2rie3Yi7vGixMrO9DbPBydeaV1SkiWgNdLi0N2KJNeBmmC
wv/O167VX8HLqLG+k6TmrfTze089BzPQzvMe4RuUNjHrVCcolXJrVgVvv826d2TgDoXAFQYyY7tB
Xv4JRErJjt0FvdyLQu/b8CPYT9zey4pJo7TXA+SFeI9hqh6U3+S3+hCHXuXkZJLBmONzwEVBiV/c
quqLOFzPqivGr5yZ7U8zu6C9uHOvyTyBQ82lktmmeYf901sq0BdcCrgCaLbZVuWNZDfit6Slmd+V
F6fzS2iWULgIMd7NfeYGABxPY1L0LZw1ncflQ2+eDbkleLpq/bbVuhX66cswqGOqDtvmBftVgp+Q
71jE22ETdNzfzeOh9CdOm74eCVAvxJKHdjyrcWl9BDW/6dmuuxNabNI7oPfz70rTNuVTWHSL0qI4
HMgh08JilX6ub7nFHGruDsEduclYIRPoOpxDCgP35UpIgAHOvVHAcw7isMzhJh/YEw7PZNANx2DC
KPfpWXVZt77ma9DV++kMIJI+s6VByQewnZuZ2oXyt7lUWTkkdnw41xjTW810WNMBlvhBsFKT4hPK
4e/a4zYAy2FgQx5mypG5pTQT3qMHPSAkXFmuL7t3HwRsn/dxejzGUVQmzdwpnlidFYO0RHoGPgAx
fr/mJdnSZwZQu1p49deae1G/89gT5D2s6J6V9PMl856fkA/YwdxkdtVa3RsA7t87Hsour9Prq1zY
R5fPk9ZmgqhOALBoU0ge8dc32fpYpbWyl/d1zo00bSq3S/9yhPgHK/NknzbrhZLk8JKGy8jIAzAL
K+QCa5s4g7PE/K7rN5pn3bBQGKwmqPeLOCbTxlky6BP3orZjPfsTF80Wp785IHOQM1qzTRkldy98
EMqn9tICOPNV3kw1WHUzbFXtkpHrNC9V8HBGDV8BcdyV5XWJClXw3ousJM9KwRbNu9GmjmLBYFiG
JAckV7FKzDSm5nwRF/PsSa4wDH3c8iwCSITKZqKLEg9zU7m9ulyqCnp75NSTXwzHq0J375ZzrY5U
de+hiqQ5YLqLgCvbs0OpAodFTJUqz0S4czS9ovvWbby/nO6r1TEpM9WlvHr6uvQn67KsdDCMzDt3
qykkT6jNEVOkuWzzJTJFZTw8KmPqFq6/1VlQeYDySVxgB12vF+Tklgp2FXm9/K0XkY1+qldzmFWy
nw3gfsIa70nBkaHUWZNVgyDvQcuqWQWCAExyGUkjKPb3Q07IizMo+DjF5a/ex2N1s1TzPbJzj/KN
FznfZCDQ5WOvcD+pWfdhtZW4yZzFNH19vanTg9Np0ZAkKmMaUg3ScBW1nnRxKQ45fE81+xwn+YhZ
JibPyKJ1B25v+2gPcsJ8/gM/nqa9lhDVE0YtvkDIrLiBhp5WIsEG7bAh4O/Xxy3tYabeEvh+8g72
U2GFUV7lBnM5Y4mqSorXB6p9GSCb0cTFgkWO+y0y1XYXiTmJI/c0UXpRJ0v8o/PfTSkLkqEGV1cG
kzp17CCNcBOmmFTtyfy4S712B4M9Vlad9Y5zp7Oy11NgC5W1ug1Hea9lirDfb9KGYrH+u3ZBnyRh
8BJj2Di/vUGKKauoiAGbDCea6RR42UGCYqvGG4sAx+/PSWecPEjwM62biaKDkmc9AhzaqgEjxXxN
jAOU5CuDUYTtnrv3ftYmhi6PDL1nPtxHmbQ0z1mRJGa5I2IgzEEd/SjY7g4OoDYAABXiqduqimjb
fKbRkXb9Q42oRXyvzYRHVuGF4dQf0DAISNr+UQgYlak4Hm5ApT/pzxBptAsSva1/OKpSvxs7P5du
x6oiz5v/8jHExMNJmEAzBK4ps6dZuRrHcteWYL+l9JQfgKNXujh6zu68jLgYmuxhfQ/YlHvZqwxR
YVzAjh3iTTzP44h4b8Avc+cSQD++48bBkf6iva5zMaFbubK3lOSGIZ934g5AFslAEd4exCyYSeju
WSe/81skef4r+lSUgYD5hVBSJma7pqHPgkw98HeLY3GyiF2Xrz0Ku2wTdqtzYfqGznVWv78x/evj
D5j1JhkM0V43EwaYhe/2l/qTZlsjU8BYUKM4g2uv2JczPiBxKrjTZkds4Js3aAufKUFg7KLa0BfC
MAJHDK4Ns2SYl9omSimxIJSPtvd3j719GW63CtASzoTFqD6rY0BWLV9zqFDLpTeWifj3yqO/Gja9
fBkdf3WBrJEnxRR87DMe9IuODf2IPk3+nUFr8WloEn0jUYHN7QBVvAdrJqwS868pHm0gI+iY23/L
/1bdaxvX4buASD0lrJNVV2W7XgH3oa6TC/1G88JVPfHd0tv6mIfIdYrLvezojwGh+9hQz4jlAF/8
YlM25yA7wkD+LVUgSH11wQPxjiro2RJR7dfw7UsHbCZTdSJgsU4tPQCMsX1dTLEzVUgiQZgBKHaF
uDIqNzwLsPu8bkXLtJwCmrw0ZzcQSkEAIjSdHesWEFscKBCelcimV6LfsGT6PpOZMlXEQUQbk/Di
NhXxb8ieZdb9SdbDdYjtwc+35g1rRvvtVTq/cJDv0rddkIWvLkseRolv9TWeFFTDn6bz6g4pvFr1
ZfGDPCpbzbyWVJ8FANQA2R+2YCQOcSdO3wU6JQ88cAo1jhVz52RkAbNdk2Rf/4La0Onq9EDbLQbN
Xs212YdVxOf4zJIXnkAcyv1DhusHD7sbDJKMmkaMacpcanGxqvD0Eg/UZGY7N/RdM5CqETQFK0e7
FHZS08EnTqMJkQ6JA2QsI6bC6H/45ORsJblnX+gSU/I9GHE9ApqV0EXJRrtihBu+Ontdpnc7dEzC
/wC+rxb/3EOD/kkaIo4p9KKd+aYamKVjEt6/t9CmmQPfVZTNI+Pptw9iqrwq2EWa3ihQ5q4rLWlm
A/BeOChCssVr1N88S3C7p+p+FtbNFwSdQUM+trAqKVrpsJYUPfvfgitfpkW2SV6hl/IA4FAfHO0z
dNn4UN8JkkUiEaiJC1rHo9aIvCGf4FTQwSAVY593v5tGHhDMzlPfllNpeYBK9GFjephOhh5oEfIC
KyHVUNSDQfguX0SW53gruJTasKKq2qNDFawcWkByiXbibjjWXu6Jt+1iTs8JQvnaseQ6I2v6hZ2V
1yW7dOv+Gemt6qMea9qtef6mcxweDJs6I2CuzeasYg9SNXEHlVLk4S277kcZ3Shdm1Nj/PIdS1Vz
yKfaCzUdIsACnV3MLjHQxB2FouX0Z8MLs75wXDkpO+7hvisUE6VR7sbDvC6i1vSOaEI4VVOHV0Zk
5vhkDjAIV93phIJbI5fPUNI5dXuOz0ZMZ7RujQy9fT/3CMM/dwK+t58ntywXRIr/wGhAWldlBRz2
WgO/reqT1XJjaHVihBoIvGP4SXAm/njYU7ylrP1nZfVy8hALG++ChVagyVagL6UXIRk0oTh1n2Ja
hyf6mA0RcGzHC+3ovmMyfX0zpjnO3p5zflPBqI13fQeupop/0K+M9QPfm+KftFteVHKpmXJp2T76
I4hhU32NN7gE1I1GxkrAh5nQN0embc0jmqBFAF+cE4IeYqNIom8P1nQqVoVaLQyMrm70gD/migTr
ust+rwBOCPu1Lv7NPLaVN1misCI2JrwZy8+Z4RQpSOd4RG74WBuDMRI48fFkjS0586RRN+V8DJpG
uSvC2al8TAaC4JDpEofNlX2hu/IWntc/KGRHEuRViAbZRw9fR0U0Vt/8Dl3024VjnGtx73gsEHmP
7Lbcy6zrD9gIlD4u6HxyRaD8h1rpUo/x/aj19r8AmvqfyG0qprPogT6cD7usR6/gqQkGBjnaJsAj
0q/0DHN0FgUEbHJn/Iu/lQwZPqDFbfVbgxylMy62Q1odZAxW60K4xOYRvupJPtwSTkBVwJJMfR7D
LpsJzLQ0s9+7JS9lm4uIoTq71J1DI65wm7Z387fj1Z1rSdXcIuc9Oybw0QyAnjVFbBCIFfYg6TK1
DSdapWIUa8emlg9GAEUCpxhsi0Jojp1XqZE59beJoZ+qOV/Q8Hn8HbUa2nWWPshNEBx7OfwRGUkR
XxeLMgphOKafPJiy/UXYoobTKKuH4MKeolJLFqHGCy9E0DTNBDzV54fusHFTulav7L7vKlaSPl81
Lr/cylWgFOF6zSRLDyQo4BSjx6VZZVAj/ZGByZctavny469hGIG1nWsErFhO/Dt6d8dX3ByaV4Bv
gszAuaAjFwXryUzZ8O+5lkFzQTDWtfAXLMvPa78aNhN3YWewu2JUXqND/jnulM/5CqnrtXNXAJXi
jzEsy/4HAiGTcf7wxFW3s+tTpls1u/txkA9d+9mJ1lb3SWIzba1W2i7d/TMPsW+sJ0jXp1WuWKNm
II8eJaCnE8qgQdHI0sDTLp2Trdl+LDkCI4ezvrtLPnP0YOlb7ZSH8+BiFkxfjZCiyKYp22vQ+kG5
cLIuzP1iyEMY7CDtl4/JpYqagmrMLPrkR2zweXT2w7ig81EsN7o/0uDgsCD9un0fVREIjcMnrt9c
/L0SwB3cXLnQnSEqNIAnWa/nrTPw1WuUkjU54Ez/F/X910AKyivFwiWErurtqVWwElcSu/rdsS66
2zJlFWTpg1bLAleOelbHl9aAjFU6Wlj4kKJ66AZZGYHAwklj/w7R7OaCJ0GnsjiZxFEteDJiDIw1
wa/2xuElgcAOq08NpRgZj4b0YHXqpMInsS95Usu8ZbFAF5tk55hfCHjHknDnh7azgIcG5JfKsszP
5qdECtYpuPMsswtVoFESFksaSMXqD+qbXBiHxooNi8sB3P4M9xeQTKmyADRc6oine1Cf81crhoG6
U+zXNyK4Dl6NM9ha7annvdrUb07S5AWz4Ekah2qo2uXIQhq5/saIetEyov96+F+jTlt09nEcAyIz
ybQY/bO5kva8nW1b0kMic6/AW9waBrzWR1npF5BNJ9IzjXoVLlRRGtueksAJ+ViiUG3pgryPf3Uk
xTuLkoCYGeeXqO8z/SgjwDE/KPlsZrQAySB/Bqhz5tNqdWPkhGId7CewNQv0LxeeBafmIThuPHgd
wSBCaqeC4KMX5jBY2c8ACbgSOYKRMz6vbEPrfhXmqQR+LNojmRW1UyskvnvU3ErTnl+PcxiYJ/Fj
GlhiVKu8x9vAQO1nQW1e4NMFBP3vaPkM2qpR3ONynSOwzTkMAlZpVS4yZuf5h/TTTCRs1hTx0DfS
wtVt2vXjKYmoCe4GcYy81345xCFal1kND2IsXjuhxLKJPy018QIQKe316PpmHz+YuhlDxfIhyzHQ
IHJO6+gE7Qm+Ynvwrovj+JeIK/iE2P15+UkOofWIcdY2VvbHHqO8LRjRtxt8en2Z9/bojWVe+CRk
Vpws+KBVlvngEwa8j0PoH/8m+n06Phwgy4+Ts/vhsE7Z03TdOQH0BagY76nHxtD2rqZzI3EVwi/1
6lmZ204uNo7F8VwtKzv+wvHwjMTwaLu2PFVqox7ir9gSbqwM93irfK1OdqkC7w2/AxQxUHnEHl+4
rW1K8ro4lAKXWOmzboTPcsVz1IqDDJh6kyf8MF+PxF73z5Gve3Mb9OQiZF3sNeCav2b5Ig3PKvQa
+XLbfofa/9ahTSMBCiZBVT2nCf130VahJp4CY8k7m9i0ClBHiAZoFZOeFo/PGcuvRlUaGzuFdhlp
zhCdLmXFPE4e8oTQT5DpyXO4iLVwttsDO3wUs4kNYU42EuzJd7BlbdfUCfdw7JUoGs+g+PGgIA0V
G83bsR/saFLgNj8QCds3URybkImVemqMe3E1cLkfLg9fYZzPQNFWkO6i7oCXFgFkqXtZcJQ29s/g
5TWTqtkIg7+OHZyJgWEg65E5kUP9CzA1nlzpserOTIKqeTepDHcdY7xN0usIo1GoXXGzYs8hRDM+
uY6BF61F52LKmYxnKEwrLtOG+tJ8unlPN/KUv9Rm6gQcvDGR2j0DKM8GwksVSH0zF94WJb4MKMVL
J3DeM0ZkH+m1rZzTk6Yi0YBo0XGrL2qUMQ0Px0vzouOcpjxHKpbe5HpdBg6FHDaNz4JCyNxKdnbq
lGzRhMZBFWWL1K/daQg4VFg6mTly4+Hpgiv1QVUAiCLomKwsW4Nx3TvS26+bAK72AGHfhsAnhM1N
1k2A7MXiF8oLIPxSAbGOazCJ+RXQFOBd8L2tzdMcwDusQagfbovpqbtDQFLM1JmefzRN6hV48CYN
SPtywWy/C3ZN8HbIPxgJzXaODWreHSmA9aqRLMlZkNi/6LPOvgqllpFElEiHl17QO65lNTNG5Sqn
mxiADj4n/X0MyPmiuLXLtEA/db4qKvNrvFrM62QSpTfylf8U11GOMtYKFusTZzjFAO78qXL0IBnE
Lm43Wf6aJTLwmHlvmo10RTcSnJ//Jpt+TgjzXLRmogEuJSItZ00lZ4GPHSLMhBL5LIffxX0Afp2q
Pq8ZMu0d8PlxmzeVw86l18QVgi1Q8NhQLogD6SrBgNi2mTnvcDwstI1ak3L3rxabRep/0xA5aNFe
Pc2oMdzwThwQdqndM/ncHxbjh0Mz8U6wya4Qlv5Od4UZhrL20C9c6CjBZZ3kS01ctlFCJ+lTFvz4
Srgy2jwlzXuwK827AKbClAH1xPr4a+9N8a3BRDyXu/CnXhic2bnJejM+Rn10g7/qRVGLwy4HTSKa
47k6BPkKpM5PkgpgAZ0tLCfWUvX6WX8GrU/koLmzZWMn4IgMIB/mtZgmzuPsvLbOZvVRaLiE9rUd
9+4+HhXnjyT6jFL4kRLS4GfIqA21croGAaeVWdkFWhW3eNIyPdkDyha+oRuIG9yGAA8ifzyWyu8G
ON8ZypWumt/sK9D53c80CHd50q4zTzPnIV8bvVrLuF8lKhsafQ/W6ih9OkK4i4oiE8d8dniMSb6o
lEa+WKUZpP5qIHceina8103M+M2/bPZ3PPqgdF2T7ueh/N7JVSMVRXBebGJaq71bDtr/36m8J27o
bWbnHBHPb6j3ihXBmTIp0qNjg3YveFPITtjDx2rQyUUgvU+BlD1DJWV/OvHl20gNQqYunEMtXjvH
Ftuq+vtlO7ybvWnNfS0RMGxNmVTfRPKkxD+muQFU1VTIIvMV4Fr1JOprxR2Rob+zb5/znTaCchSR
NG+hvwMkoFR+ocCRGWy+TLO96Ak4WidW5UoWv6hpsl3n6cWfXtYxi04BvjEqxQNR4/GraIgSDLkQ
qzLmS17Q+Z9aa25IjhWAjHW9i3zT7Nj2135r2n4doIDUOG74Y5O37cEPJk3wyVoaengiLX0X6KzO
t7E+GMEDl2hhLZXSjgH9zrX4DtrsFoMXz9/oc5RXJ7gSjz7gyADNvqgNHB9n6q50+fwEWirKHL07
GSfJwsaiAGu3AmGJo5jDeWiunPZTkpj7bcVPeOxlbv0/vfGkMjlXiTVcHPlvAv9vqKnbK0kaQol7
l+spiT/4oAVQnzBBYDfnZa1vsVFxwScnWcqWuIxn+NZPBdvZ4/pKKsMeU4A9vOZI0nixolzwxEzk
8KK1zHo7XX0z/iriYtv060JQxNpQki2s8X4RMbHMZg3Skgmd9F5UMcuRkAxQLzzh/YeNH+EGp03K
SJc1WMfGCra6G7U9fnQ6BOkBWXT5IcxZbFpolZMBgh8rA7PArZHCGIMC5OnNqx3mnNQBZfvJrHiZ
KBhxhlJ/pBnyBk34rhPFNFoljYRuL3jfOmL0K1bxKxPTRnb1Y8Z+upw9ZQqj5E3mxJSGAUO12qqn
MPE0Mb7V0LJFHVAMf6eYyYhktFkLmIIDyeZyKtym6fQipMeZJXflRmR4SjjYQ4eMDTl3VPjDaVJU
CLPJPfxc44K3RKkfKRVxuY04lEn2z39wo/R8oyM3OhMF47ZTi/kcLS1iIzrCA5dQllQV/tA0SGZt
43E7iNymLGxWA/J2jwLiCjowp5SmZNmpGP1lNQEmCGaSIl+S/gq0c7TNyFZfOcMSw+WWkidp6ZxA
i1vvtxisiwou4Eb0td7A5w/qSrpAtOKqPFcYL54w/+ZSa4/aTyIzoxzo7fRlTojcb8umQtEBxvwP
d+ey0zei+JTrg0HcDzkN4EkSTm7m9myeq6zuGEwlyxJ0dLD/f+zSj6ORPCehitZl882tvbqcwGl0
fHKhSFFfSBWOAGUTLUIe5W44Ceojhtoz4dGPhf4/VWV9jy8euhGzMtIWrwyUwAiyrhQHFNQFpiKd
OBbisUnw4XGU9/fURyXpw8x+Olehkq0lukym63ciJDrZRqdltLTei9vXGIqYAGVhziGjvLB9SOPa
d+llNZGUNxgYr0UbTlJgocKwSLtzqsQuaIzkR4+89VlmsFwu0wRjNqrrm+11+SYgYNzF16cHv6el
dbaZGkENNbCgUdwvi8Q8wsLN1tsKBmWUE3x7bCufnRho9XNN4XisbD8yop5pH/0N8clyYJiFhOyH
Fg850LB3cG+D80+IMnD5FkV1PQBIWH+KOttJCWXvyo03WrJLfLiCjcyPzquukFb+bhtTpHQbpcHb
fDK3EMRO6AXOLta08gpDtMrov3oEgGmJLxijAt/fQTg0Tip5A09WvQ0KQcqB0SYtuVA0pn6c8Nyf
Ad+ajTwW5LfysevI9jebp86qZc18nh5svCx//zJyEB+ZuO+4ilvyjkDFT2VtwjzU5guUvQIcpkF4
IkXcD3MuvgRMQzMcFtPgXnjlkh46L0xv1pcE7iHqK8Ul8pfBVCIxCSv1Uzvp1TWBPW20OX/00lMW
DtnOT/1InE+1lqjpxGlO6ML1GjpyVpVaY1z/+nnZdrZk6KqEkn9OcBbYnfpnfTriTN0SXBvFFOY3
fPnfiTVXiltuqkvyBFHRFcIlSGwe+T6ULzPuhjY39hZ88NPS2qfNeqyt65D9CHzduRkGEFxhiN7n
XTfzSKyVUHIFFuvZWwIN7NvD92F3QzkDR30N4BY9wLx/unhD5OxCoTb/tPSbW1S+Sy+coDNE7K/w
G84KMOameukilplx3Z+NSXrmVMpWjFl6X3ttXCAzlMwrQrfs3X2FZLrX7A5Aa9aiwsbMlOzyWSzZ
NvkezOkjuAcAQZ3N5Hw7F0rX36kOQt7iElJHeeQKAjcIFv8T2KPFzTZVeytQAW2LbcQulHGjvjs7
ntGYDp3+820RsMg/JWhclpqJjeY/Sx8yXqDzubFtLL7l/qs8K7AenNBCeVQQ/xc/7wPJTMcBYTDD
rjCg+jR+SUDULtX0HgQRAhKJYEi263L5cmJkMP4jX98g6HIGm0AhvzInxMpxBYLjdcEMp6B5a0iO
23tYrmnZjWv56OMJX76s9G/KtnyWphwzifjG01Uw/74UajboiUNKFOcmL/tb3L61r8Gwx/QSmGQa
j+WGPe47O9g/VL3GYLgcvGSgM3THPmlxCF1KGZkXO27YVnmUpHBCDAOZxxo1+mJ/WD3AR6+j9BoX
6oYnqNX1pPnWqLiQtutsR5AugS2fbwDJ3TD5T9KhXXFz0HDNYdGsTOSPnpcjxljD1av5aZLs8lYT
UWSGjYeAt3O5B0fSY52b4PI3Y702BEixTigTJgvAGYfBcsAg5GAoUTwE8VEBpX2X7qxfJlwF7SJB
yOsW4ShnoKvYT2HXmqcf2LFBcKetLwphZF8Q5wjsSy6A/EluDSHpNAQDgBPyfRNLznU4r2Pyx5PI
K1+nJG1sPzVipy7zn/S22/nBJLAGIDw1gTs84FbCRwsPKPSdzf1NIJDRsBMyjAqqbWbb6OSUo6S8
eL6/OmVafw31ncYmImp12a6be/CUkSoulHF8SZRxXE1uqEoZE5RY7M/xwCaM/CC+5OG+nUoyFW2m
+aDt27ZgiXjwnizHu6AkQ7YDlgvUGdDCrdzmCcU9gKBHqggGPbjlg6RWKp7uqRQ101un9yxLUOeG
FzAUjhT4kezco2ZBqH/6TDi6FDrDYt+OJ+jcP2tiSyhwE0snwJ6Nfp+PlKfvL2WUdf6GOl1N8iJW
P6hnHTY/u3JwOGKcI8TJkddNhH9dENtYsgofuFkUiracmbLiTBVoJp28l1X4PGeWcbvD+IKXE4Nn
UBnHsyrE+aQal4Vzp0OK8XUnTPc7VNsu0JPt9fPaTCtThpwcvx01tNK4y8c3/92NlrWEp6HFlxqX
FGohazB68QkKfsRH2NfKNexZkRDVjmosp3mbY4l/mIta39lR/2xKUpNow4WARPREWCl6A6t2miKU
Q6/h2N0rrhYZIeilBhQS//GoCtxDrJM2AjCdtnvut6riHKViU/kzIaWMAbZm9rSRgtbl13fkYbuR
1P28tM7J9XNsY8TAPeL9DccQ6pkIwg0WyKXD2satiVmWuudfqsDoSMXT6GFOqhsKmDAjOGqEuNSe
99ICF4aa0JhZxLxF6O5h6UW9wGxtVRXY3HOD675i/4fnRjHAOXkbS2lUkDFcyS5yptigRLRSltxm
1PoEgjcRFLm+XTHRqjp2MbgIWD+r/AxJ1MSQ38RyDgWrNrazUSCvOCo6HckkAyRtGle0rECCEINx
QULALSK8HaYIocELok6oDmKRRT8NlIsc4tYPaF3hYBloK1f2RbqJCxkFzwwhJG+aDr2Fl5Sm2eTx
/fgr1cquiVan2Q99jA0IZRhvmjO57Wnx/F1CBJ2nkxkiz/cuLGxyEzIx9wgLdjkeGEX/0aRdBhEb
GJwr/zfNY/2PEe2CuX7ERMoLEpNsF5t0a3tSfHBH2JFNZGt96EexhjqYlGbvff2aSnpdPCwoM5n7
ENS4Z8q7CepkBtxb8jVv7jcK8qxg5glVIf24ERVeTyTecXwsxv5B5EllPzNDH1NjkaB6HeP217ko
jIM0lCVd7poMS19/l1a0On2aoCnTmZVBfpiK5TsYCL5oKXKxCrwU9J1sYpjxuTE5p5jA4ZCkBMj8
XGPSbVuXWhNTlda/YwlVVeO3l5KLfXnVCBlKRHdeLRrSSd4eZ8K92sGR37iPQol9h41nzskt0Oq9
L6yuVjB1QDpMFRcxlXw6UAPWEizOP3iF7200pE62E0wIH/dj/GWqnPniw1APiDwYPaN0OcrkxAUv
mExXVNrTkajKI9PGJDJbVnxI9/bdSTSvGJnXDP8jKR9uKP8rsLE659lcZJxlG1CshYMwPr04/NIB
GyxR9jn9AfY1dyLNXRssUNG/CkW+VxIGDVSPLbIC541qAcGEjOn90ND4FyfiNuamMnyOHkTYTWK6
tUSOAGLxLIFHQbDozOqLQr71Szqans5uIAsLkinll0COcHgNLNCtCEXcGtQxYPHqqBGtZO5WQyIs
AtpJZIt3GrrP7yUhvDpUiNHqwVP4xfQ6by/Fl0tnXYPh9+n2Wq6lLcaGxy98TsdxzWIRiZqIGvML
gjFMCKxuENIoiUDEVJZ9a/BSSRmQ7WxZ3IDZtWrmP0yxardH9wf+ZlmKBdBS2YOcaQ9YlLfhwPcl
LmCxQXaoFf6nZPyrrWbxIpY+D70ErTMsz91yq/FCSuZBPDJ+zE5I2xcf+u+C9ABU7rm0MzJp4aBw
bbPkP49/p0WzvS+v83IQygYOf7xXEL+2WLlvpYMGG01y+DlZvHsuwTIjjsMNXxBsHOWh7uFDFzhD
lbfQsz3+AiTeUCpsP8EQ1z/6PSl0xNhxjNfFJtRQCTsZMakTlgI0g31epSUM4xPkh0Zmmmtgc+nm
9ZzztYQF/i/ckKync7QiAeD1HArobqYKCQcejidkmTuRl4te3aJrxaUp8I9/0eKzcWOZPbRDmLdk
De979YikqkkaDrElgU463djyeHo+D9kY4X771FGvgvMJqbavOWmwLa/eucE21EV2JujPe2N8GKeM
BpWGkt+WmVwBHG+PFJqXLGPtsRRJjXkmuk6qS8sNuzBbOLTtF9jINLYi2FtvIvlMw8tG82yDUMuZ
w63lzUxVub1h8PMA1XNFeS0UvOggJPZEMJsptsdVYjNpGQi41Ms7QtfTgWITKpgQvx1GB+zVrIRn
XA/RFgW0zNFVDS/QWrGWpaofThDdvsV1yQeMSkZY+CoqavmDcRBVyfxUrD9PUtaAFkey2KZIICi7
VfD7rxQ0+/2MT7zjUMaQNpYwN5QkyrAYU15wvKLHFmTXc6ADZ/8d5Zy5QAbQWMEAjrybGZb+tBvk
+xIxoYoXK2yITop90fX9awdg2Q61vIvr9+b/BoH/zi3BVacecyDyCZzTezFWCozXSSQz5VpBIAIY
G/BF2ke3lq5ZVuP1r/qEzhnZOauQwsqx1s217logQR9sCK0nmEKLnpjSdsY56JZPkkbxRj3ox5OO
e41E0Y+rdEQOC2E5Mv+RCfJTv8ci9dK/JD3MxNqF58qOok5dhdF2TK6CMyGnvMio5VNFuResjDzO
oVyF842EAOLl3RoHlEHXNqhh4hCU0AH5hA0rcDt4Lu0v4Y9WQAErfl0QJB5Bp1C8JPadF0VXJ2oO
bDMULai1fGZBWktVxgHlTgsmNDv71ijRAgkutfMjWT0j16Wp5um4mVioq1eCE0LnT7u+5Olgd5hF
we35Au9yoka6R4is5ZiqW3XFcywQTLGvJOCczyNKbpdi5bRIAYalZpY1P7NHCOOOeF6LJXtRAzyW
zFe2AXxHAuDqC8dA18I7rWEEg1kUxZc32Kuwh3/0+wxTlHh7g0O4yi2WmdJed8zkU8hwkNUjsgCf
kRbaNj7/7ioD06e0d4h+YMThuzYbH1yXoD8gKKlt27v1tM/BsDTZaGJhvpoY1eIcNLqa2PS/WpXF
or7B5h9doyd4StlASG0eO821BfPnGm1dQSauB8wGBx5HZVbPyBdOdFDm76psi2Ej25JE1PuZLxGI
th+jNN/SVj3eIFxv1PX6i6Y5I5FBiK0zg84uV+5xcc5Hs2ZhK3qET/hEMtDui8C2RGGqOSqL+QZu
JgXZaI2VH6vY/E/VMKhTNcyYrfV/pj9BJQpv68MPkOVMiDVm1cBPusMHQmT27/PBMVzU4fWJux35
AC7ELLuLghxLd2dGkOeiJU7GOccKo8um8itrIzxuPCM522okHqrGdSGarKwpftXTksY/ZBMo3tum
rb4LpTaW5G+DxjhdRzbKe5qnoeO2nZzl+3xJs/fltkshOaDHtso5OB3r2E4EvaQ5Bb1c+bqwAQdP
ueWUjS3rteQ8U+tCxw2i37eYE5R5bl7TamBNXDyKfyBNDjfaZiB4gtVk+bkTeiE9bCl8qdVXPYiH
0pgZHzss0AETWpHnZEbVAFI7DQJLgB3MKOYJa3+uwVrlWVxzxVr3KydMNyCafqHHasOfG+db8rl3
aeiR7nkxzp4OfuUBD2Eq0y5isMkwxXWOi5PB5x8hzNhEkaZcInpTV2t76dX4dI3MP18DRQaxl7v3
Sk+2nYQ7A+BGdxdArRXbxIEcoE1cvwF7o9misJ9W2UP70Rt3z1/dlNKkmfOWKf/G5eGPugD33k5m
tYs2jRxNv/AT2IozMw/0uPGdNuN0tYbKy1ATKtGRC7LVz1rElDqTYKCp1SPSg/nsC5wz12UwvoNt
yynEjl7Q7R74ZQc0A1wm09PZpOXNgAQHNgEkZ7mllPl0sdtHnizQKh/Ng8KztiPOuvRAOfgxfrQh
db8bzmoDRjHRqPyYbIsHBYlp+MrtYZ/DLIcHms64yD0qSIEsPXn6jUoFUaH6bLo3fid1oKA4eNNS
5CBOpixrNXIYeIAUJ0tUODdNqrNvGA1Wbwq0duK6PIz0T3YOeHLPPaG8pvTKdEoCkBD6Bz1QBkk2
D1THnZU4NZbSMPZIcawZ39V6wXlcJ33bGy5uvUxXTakwQj5GveNO1DrErC2riIiGDJUoG+NlDKOT
MEeENWoO9nG+ass22RvQsg56pK6tqx58KDVZYOpucrWEsXsMAu/jJM3FPogGQhFLe9HpxImmGu+/
hqHS+xIwWoN8L9tQD90B8qovLOAGgGreiQD2OrUbKILJGaxQudbiwL1P36r9szvJn7ijVPGkb2oD
DeNYeVdVvHACBWEbzTIW0/aiFxN1CG+u2Z8Vd2uFkn/MHNVa7T7Lmj83jx/GA2Lgtc8eR9wvMfiW
Daqd4NePC9gG50/pK8/1oi2pSN9rd3rshyB8alQ8sL/US4YOmtweJBg5+4tIovy/Rafw/njOXZ5s
2te2EM40OkGxWBC7fBjXl2XO34dafhUspBgx1DocU5W7ydL8AgTdzoDd+47M5y9yUtvJAxYYOCYK
EqCJWLS9YMXCiagMhJMFQgPc01bIb62YNlDP7XlNOQ0P2z1dtYWFsar7c0fybtbxsmmibpAg2Wri
cbOMJorhuCudmj3SQZs5N5eJUDvTPoXgHQpECJPUaFRjIcqMViV/su7bGK5MjQe7cVcPSg7aDToD
6EEDbwjU5iKaZlW9hJj3Fdsej6oMrRAl5BSoIIakOhJG8KNvYiax3QoF7LPcQIUjb9I3Y7YoH3P8
WlOmHZwVJTuDaR9NNboFbR0LeppSFwYq2AeAKtogt2mitwXOjtY2+fzO8pRumvGC7KcTV2vMcX9s
peOYK/JLc3KGbyJKbEnNiZdCcqRGt3KxgQTLdDmivfkK8RSvV5nDsBZuaLFfmQSjKaOn9iXf7O/y
zzfkQNrYeI0k1H6HJ7EJq1PQKiIY24nzimdvG8clZD9/BcPB527JDiFs92QaCxUxNcd7BRbXDdBn
h577slt1cDMCLOQ8BBhoMqx+IvndLwHjFT0UzaXm6zYnga346EaXhwfDAoo3gSHpjEIWSYmbu8nv
izG9m8n3t2lW8Hc7VpIonnL5SSperFkGs90jPldHR5DpyjmlXgQMbMVPjHohx60TGCuvoobWlwEV
l1aos3WrJy6dIuYcdWwXOMLs2GUxQnAZCHNIS6pKGguk+jbprD01B+STaKtAczbBiDwJgYljc8IN
p0JYGk+EE3qmNX9tFteFEBRdvLUH1YV+JFDo7eew74sqngx0KClPx5PA5DUp+pOD3GL8nCvVL3jt
SPPqHFe4Thihh0slhRdOLo5M+5hIR0M74X7gsjv86hH7mOpL6ErLDnMKyC8d4JhXGGJkQWeuLgJf
RqeiSGgKj34ts3LA1BJ4+40xBnWLq7apqwGTS3ITip7CVTlNzoPMhfxafkIlE/qjsMaUE7wqV7YN
f7RhVogD3/+feu1PhlcCbMIcMee9sdkBz09x1EPS121K45agWO6nJkcFVBjJHLzcEEg0uefDgZBa
nO3fuI+/QWzoyxVaum64JFvcrnLXcdtCYrAdbimIBRdSI8KHAiKb0j9UnVoe7xxJ8Pmr/S1w6nQI
zlKta8gSmsdCalLjEE9QY2DPAoPWoczfSXKDwVQxts30wAI3qjz66oMfTgwj83jR4M9jRrbWqd7D
jzP0/bxuup8QLsI+LS02pg6IJ/2PsMIZyMD0BjeAabZiO0iOI9O5kFiMIAGRTmhK1dsupnyVr1nH
M7QMRRAQNOKvHQYMa2/wm2ABw+5QdnMOTEgMbIoL3gQAt1P4nAqCfpM9befH8b5aA20h982mqTcN
8ujG98w9u3DAYy6Jcj4+j1MeZgDKK+vGTcY6npHbXswEmSif1rdMTJ8ETluypTTo08FORWLCw6+S
saycYHW4SP3nuV79ZTkkJaCXpPt3NbrER2Wld73ZEB+oRTjqlP4KbzP268vQUtRG3IEM2P1EwQ2a
NvtyhnziKbCEYXb0HG1gBZOkHEL4zVlRSZ81tWSTvC6lTLrzHciUaniDDqDHyEwap1/ZfdopDCLF
9wB4jGBeh6uqiDqfj0R1BL9UeLGymJN9Qvhxm3azV3DLyAffEcXEiJRA9FZN2ulJK6EjReDunGO/
l1n9tuW/+pOldqQ9q1dxRvWtHTBJVZ1IKiHdconKgm/50Y2+L5ETnh1yDc1es9qT2VRbFN+suqxt
Fog+qr9rTxLWnWi0zxSlayLxP+h0SdesA2TtHPsBMNjBXrqM+/sp5CnFqj6JR24mXAtHrkyYhaCJ
jAp+braPzPxcAGanYxzor+R0QKPgpY352bXD3KnTrYcon+APffjdvmfX2fu2knWgQPCTt06jsd0v
KkNcl8Tmk0Q4Y0LcfFnh0IeppHdpxsei0gJg7tmH4mIjtTzUUIzikTUrP6uCUohXFbRX6lD5SXoN
nNRohIU0rQ4xuxeJLcaSDnV7U7o0piKTjtMf1neiucwrspI0QcRHrXcA4aHPmDdpcF//CPKjyMnd
hX2dQ4lt+E2r0d/sGH+eV7QqCPYjvU/EgWBPLfEe1MWU64CUJLjApOsx/lRFOSSQRWyrQFB6vgPx
TWETsbWA4lHoUhIsoVmWNMWbcnLGN724JV0D6ZU6OlIrIrWy9zlphAeThpxWOMiZTvPcyH3RhjcX
iBpu9sTPZtSbHPamUQSf308PBvpiPBFUtxdSwNIaktnULtxc9/jGe/V2I5co4PuJAfCiLzPRqs7x
Q0XQqKtw4BEKVO9tRem5CnklzlQYEh/ZmWxm8KHqVOBH0kdCV3DRxUdyNLqImg2fdJ/Nyll8DzbQ
DxIpADldMnzqqLjFSfyFAfkZa2YoQ3G+tYnBOClOG98OwOE0FhKuBl+lg5cAHL94USg3WYPNzu+G
s2rM4saVQ7XzKe1Ej+eOjjvN0IEc2C8Qkk1jtTPgl4QTmtu+1OssOJP1Ya2n0B3XFu/O3+YMR4QU
rtGx9xJWzSKGwsTI0Gb7I0MenCK/KU2jV+ChG+GsL5QzJt8mGOU8FcvZHgqunpVMrPNrWBvFlPRq
0AtP0NwH/8me8JhAPa/4SrBaYiBHoMFo5l7fzATABJ2rJrXaro0GZXFkdJGZAGR5IEwkQFNHmxLk
0Nh6Sn3C1g0xNm6aXDH5U3jEKyLk3QdC12CqVY41NJue9cXs5N4nRr+xsZcf3PqGTGj4B7M4Ybx8
CFKNT+LwRUxZrnVLF7co+GLoiO8Ck8IJEt2LvvqCraNfXIB6pkn02a/R77N8OrngaYbHBepNNLyO
u+SnvNUfzattstR2pv5jdDFtq5H1JXKH6a9O89fIDNCvlW1MuJ2It+I7MD4UpHpFtZAOWgQlDjff
7Wt372wAIPbpmqAjRD5aAmqnPNs9SjF+26gDtbHvOAjyZPQkFyO4PEVRbsWt+xmlt1g4agiwc1C8
1HEbdmJ3VIFCxeKWKTO0ONylzmO/TPrAwrf5dzYvnUq2HJQhFqDd54LUotfVPrGHRmqXBib5JWVQ
3hMGcYFmd1QuIDFInhqFxJv2bByv5W5gE0Dx6VJXvAuqwT5auJ76o6w0h/uaBuSyvslDm1+VjtwV
5u4dTY7mqA34Qi8XW4dENawSRycOPMruaw/EyFbgAhriuGnMKOe3SLp4nN5HXv/4zWt8Zo6W5Jui
ZyE+k1+RzVbELvrAR3xJ8820XFzojlgUR3wTA1JtNQyJ76PyFieaIYPojZwrULhFh5cpQOXStTrK
qQ0zFz28GhLLTw1DfJyN42LK+ME9CzkNtCcokut+ukeGYnBrHcC2wYHnZcHrY/Lg32WCv/FBZZYV
VNOwBPzMezoKjE0/hsRp5LEZlAOkEhtA2V4LaApKVZnpFpwjm9kD0M+Rvdvr3ruU8kOopgpKnYqJ
FTPJyEqlP9K/JbG1RL/+MIm8Wohx9/hRjYBDfez5gl3U7E14lj6OivoSyqR/ofHTv44fYtt0CSao
Sl57ydJ5t+b9ftUpQKF03C1S2C/y2uddB0bhAHjMfOSozKlMJ9p6I/VmIWUE3I+ESr3zpk+C9H3T
IxPwFIRhj0TnKnyprqv+pOiCya/jIoZJnpYpKcHMsxlLi7qFNFLaPAMM42fgS5z1KNxYBhyVlvZu
KpbpqYFg7S1SnBgq1VshcEn9C/MNPfRXHfTsEqnhIdwrvlIvZ8p0J8N/kb2/V86sA37ktLsCweH6
wu9ZmrFRX/zGh7Mt4sFr0ye1EyR2o+f5deqCKViFLYjef3fQ2t40ywEFR1xxjMMIoZkqzdd1+S47
PbfgkyU6NmczJCIGMafPj6HA5SvLOrLn7gPC4zuXRuerEfX/mTT2mu1uDsVVdvxO5TvC5gcMvias
eM93uscBkkH17i0WLoJLKkFL79NMGFZ2r0DO2n5BpdO8jnADlMV/CRuhWQi0snssk7ZWpeUySsdb
7Zvrpn+ZzFQIu0OXU3Er9QJKvywFYrVE9ddEzCXWsuJOJSYM5GLMkej4x6UXHLp+f2veduFTChw1
BjGeOk+avroUvN91svV9l9Gj6yGIoSV1Mi+VwDDbwAz2fsG3frsxKyQ2h66GvOMQCWBbvUddUHN0
SkS97byqvrMVyosTfBcV7ppCqLXjd98+18r4nhfN7Gssq8Hq2Ft0sIcrQeslVcLMmelGZQuWoXwX
HbMTLby4q1CCrMi4KM3Wl7TlJToUQUz+/XZgblGw/bFBkS7bZw49JTegjam+nyZuS8WYyH3QPxWs
rMMQwg90fjTHQ6cEevHMc9rM7ZtzyRdKhq+k45XmidWNZfzxJ5jJphSNoycc1YJLwzTVQ/CdtP2K
lvDpgf6cwFmnwqVqSTTE+93UtGKy9kxMM0vsATMFYaKf9a4/I6ghN0jWK/blAn0L166xgfj89YfD
HsSDXGTcjb7OADOekEbuiSlYOGff/dnIkOxb3XhBUXwHp/Q62uGEwXzLnU65cNe0DHP4UaVSJ3W8
1GNZHtuU/XnHRwVk/RQhnITXDTbnR9DaFnAYR1NzaE7vUIZeus3GipRZxbTDQjdtdjPBBna1PplW
CN/y9o9B3aCKtzmNZACnfJOsHRv1QvZ5GiN3gn0pd6O/gJUPsX2tpL/ZM1tYUpaORTdEpNfMVZ2n
h1rG4yqRXDjzo5ur4VAfdojpiqwQ+3MFqcWlqONf+chOhw4XQ44hz1HF9Zc3fUFAZCZ/3zQ6py6E
Ydh7h+y1op7srNbdYWCJgyZj8Trq/zIp5F1PBblaLeM+eE2uhqEqiNb1HUKlAD1sbAK1VxXlrKEz
8vbuLPCJKMZaJxaKiqdSl8W139m3fuKvHJl0YHI88axnj4SXjMyMPRiawmRRDwOXFQ7XCx9JP+o6
wyEpRDI2CoQrd91VmqfhtKtVgSCnODM23MfbdTjgQ1yk1J9L9PQplHwDIwXueATgkehF7I7WlAmK
6lMdA6tLwVAnIjWO+xmmVtLsGn3kN84eBxUW9uBUBI5vFX1oDmz9d60nNNtp7r0wNAgeEqGPU6t5
pWFpep1OXaDZgQ61yZaTWTOY3TSlbvlYeGfRhfTc2H4Fgfi6mUDU7sPf9QbaO2e1eyZQY640rWx3
w7A3K77p9sIGNSzPjD3S5EXlokxlHvMVqX2TEmlc4RTfISBXXGHCURQfHGskc7GOLE+o5cCONe3E
XpChrGqxJdVdcWnJ/IoC9n0yTVNXFTiE6VUNjeLCgc1KiKkA12SUYhJ7IjeT2uvTqBFn/iIY8j35
R/TNLZQq3OmiNCe4kP+SzpUChZ7ZhFkKoFeVzPbpYtHZgGbOHkAfV2AZvxFdnfm+TeHuE7tqS2Xg
bcNOI1JSCB9tRAjUGhF9NjkZYcgnHZmzyNVYr7Ltl/yAl7VT7TcIB1Px2vyfBnf49bJjBgbCvTOl
PoLPrDKQbGbXpNevaunnnsTZ+hWsQrbVh68E4X3qnMtZBWczpCLWLNrXu1NaxVnanE2fBMYX3xhD
q4re5fIvpmcKDn4BJOTAfGOnq8OG+zAK1Joj4g4+78cH13O90wOQDGvVff4lKUSDfccnUOeoy4Qr
OQ/yWsmEz+mnHlcQxfwiTS36587KdsHjWdSIIuOXvIsUSt8psBf/Le7w9CWjjXImLvi5bgv16sK0
k6ioDKFKu8vuvbMU3T1S+AlcY/FKVlgr74/tOLsAH8kGGdxRGeLjCz0/Lg75DkSo6A2rItHVTXJk
8gy0t1pQ93Bs6xw7Axq3oxfng+6oc0O4fQ6U66FLu7yDwHei1mD8V2dUyxAqdxwaGf+1769YAG6H
fBUWaY+rfm5P4PlBQCgCvfM2s921Nab2cq22QzQDYYNJif/YwBMqqc6aTRXLU1xDi9Y9Gx++K8ap
jEEUL51rqBN32KrJnEQxUIf/+7LfUC/BL9qBNCBXkGL+JbZZAyme4pS8ebm4EXBv8QDj75nlHZlt
uhzIKUK7++0Zdfwtow29kjcIk8DPM1VoDv5SPV/xF/mSswbLl0PhRmloI29u9mmhVfC1DGP+XjKQ
I9sJWaewcjx4xofoXIS5td3beYaMosPkeduBN8YdsjwPADj1OPyq6JOFYrlbyI9qAMjzAb728HAp
09R7pmQUAmThhKkxasdU76V8caAzLCTz/5Op4yY/+gF+csuGuDlSy43IwJT9i0s9Ae+DT1j7NWeA
/dWB5WTdLjcP/kWwCJjmBTZ7G+IeMFWBueeXx1g4IP3YAhNypIQuGHnG5r43lZtobNvIUk8P6qhN
Mv8NEkEK/GgCqwQjvG1iPnTL8WO9NwD+yUfXVaIEWAs0nchX3xujX9GyuxnYQbYYT522P5zXOKjY
mq8R8yqslL9hGg0K/6DUEObFHFnfo/AHqYgRTl6pnmtuz2QLsEmdqM3YeTpcVwYcno62dl1XOPBO
uxEEoQiDClWV7QYL0FLL++x9niSZ4lddnpQHgf7nH3ifHSK8WPKMchu5M6X+EcA/NI/TEokPyNAz
rzI/DPHYH/D6dEzKpZPFjERVAVD+KV69u0Y6YMyOos2X3x6Ct/8areqZGbr8NB3yohdhAp9539Al
jBEPY8a9K6GE4dDGFowGW8GwC810hfHLtU1/kX8+zcD557wRKitAdVr1vTsRQqsuz7Wi+NmejYZf
IBPegBnVCxRIVBhLPkN09Fy+dQJZpxOpOuYEvzqUWY94cU6mOXKxm4wAuED4TaJw8TyhP25qrtii
WK/8z0B3I8wPtcQxvFX5eqUATF8/j3O6qhzHALpNr57LP16v4e0OMaeGdtvKh+8Ngd37R3CM9X+l
wxnu7bz5M7JvrK0Dz8BDi+Tsx36Th7DqsIqoxJ+gNWy6bRgGl/Mi2FUaQblAMgSfyqheAXxEreqk
UpWU6UcdsG+Rjz1w2gHF2K80+YROezvIOn6XUg/pc+oqXxHFv+c7UxUmYvfrxHuO0tplfxcfNQ5a
Trbz5+Mb4HshVWZeo+7huTqqM1Wg5myxtPS2xA9HQhj8vBU/v/f52OA/HzPyyDyVv10C9JfiUTru
g2m+UFHg/VFlj/muTP41OeZwy89LBo0mI+YXs3OmUcl+u/u7RNNRyBBe8/j5C0yyK83CZKrfhXQb
wSO+MO23em44K111idWzgGBbFiev7GQyEGRhq0kpJw264Vdc/DvNLG9IG4oEDXJPPekPTGmrUb3q
x8Pp0pe8d3QwAqj8csq5RQYs6o+n+N/Gy75ztdU0MFRMtiB6ybMnHP+hC0zD7RFhkoOPWcv9uNk1
6p55EQWrWB/itzH4HsdfzPbh1reqkoCMpOjl2fP4Kh/uNLCTE+572xLLpwq6Di4/fs31dj57ovDK
P1y68zekUQIVyKXZTKEhXJW0boa3iVrZSVFJrDzCY4maaQLtDhg+HPR16WPRSWkAM6VFAMWorpD8
KHlzuKUFoCe1FFvN01f3wEzlvjOz56XxnqFQ71XwuMTrZ0OBVji9RjT3qN/CXd7GZYgmsOj9QIBI
YuJezVwHlArCmNabl7dOSCWV4P0LQMXwjwt6YG0HKA2bHMMWFKFkAKAIadicyWgIXJPmkq/mA141
PwxUy9KKbPIs0MRziOjn+Ms+PCjhcCfts/nX6okrAC1ztelxEHMu2NSB3mJHmOX3DxABxwhumvjo
nV5h4gXv2r2Ts0bsfJto8fnWS0owGwITsrlM0S1SnFbvWVNtvtTv0vqcs+aJzUNZszzJbbhe03kH
UJojmTBjraLYoJVdwTXWvRc3gVqU96vYuCI3Zo+g9x+6VOqj0bMxIveG/BtM6IHvEMkKGv1ymViR
NH0qgqNsroFytEievQu9UZfSzW4FS3UDQrHVtGGuBGVuLEXB7BMeVtpa3mS7OoNO0aV3tLhUJiU4
F/3jfsUUDh6SwZTIJvXF5MWm8rNPz89sT6cwAawLIF4deMx7sZmM4IwbJrL/g7pQGRXx/uH7Hg8e
4MjNricWjbbsr7zUeIold7aJ2Ef5tDuLAp8FToFuD20am7gLH/db0vbbw6yHdEUebwCY8r2VJbhb
l4fhcaftMuhjDZ7XYssgds0+RZV1zOC/oOxUP8lpc3g91ei9GLWhJNSw7knq9+mjvJxyfRNSX7j0
+cfHZaeb0iYZcBqBHxqnZH/ajfCftGezyhmmOPI+A9o3D6ZcMimsCYhLeVjNor73T0i/FZnaPh9d
R5iIxZAk14iYG8L5CbMjlSeCTgba9E8Iw74Zu1jmryvaA1gsKUWJPmtwy8DwwwfdbNn9gbvVqLsW
TbcHSym2830txNYpcyxaEK87kQlCmJlzrTwkB4Z/FNuuVrKONzRmqybr+UDjllAD+diaFeIgazDk
AgSXpCUiQwHyqc6nuTPeLUXqwy1Dw6Fdd2l1O6Rkf3EUKb0x706Nkp6LZ3mLt+fDlIYzfCDxfCpm
R7l85o/kJGvvFolihgwgl2s5O89MtFBPB47EWtmOVzJ+NV+RQL7vsqzUHyJ5X71s/mZHhrcaGGyT
VUK7bSzUWGDnhXpjUODU/L6WXRx45ayJS8Lq0QQ6VcqUneP1GfzVJg9SpGK4X+K3PtUR6Y8xKvHh
cqilLI5z6BopqOsY9uygYFsvp+YChg8mEJWc/uNGMX4zQFNNNEEQjDrnesv+Q9sjS0fSs5OW9ncd
Zukf57J/rHCP/QEVge40swYhmC/eGB2+rFgxAZWk/EA9HPLnDzXfpQF6Cl38Px6bpd5g5VLt9fVq
0eWlPaSEpESGj+2z5J2Rf0uv9prIgjxXzhhak3aCe2z+HOIr1bhnla/cchm4Y84rBzVd9NUcjnZX
D6c7TAbTzDxucTAbXt539zFkxn6Za+ozAkX3RlOBzAZoQV0dMWrv3N9Fd3uY/y0p3LhzyZxBbohy
3bE03yt9wzhPy13yk4ekC0Ev2ZTbv7v7w9ppgEnf7Uft7Sma6aH0fXMp6yYFq85N2WDMJgDxGa1q
gJz8tey5r1LPjFNE6rhn0PpJWzGDJev/LPgZyHlpnhb1N+zcn8cVkWDXdebKC4XwIZLNW2xiKn4R
nehIbXDfcYhDm05SaY3a+aqxd0vZ5HYTW9J6X583dN67Q9xiB1z9sd3w24BgvbM8rnVWflx0Cu5S
KcbVx+JRgrv3RdVz1QnelCHWyHvmy5kjWe+cobjl74CcYKI/LwQZ+CYsfhb8ONnqc1jNLxGeLX+S
x8hbOcBPfWjN/b/eZDMCup1gk+vxNQ7pr8Xl3rTw1Mz3pSK3fvBhwXJ/LKa4q1uXtttvUxBSwJJR
1rkgxBSdPNt66mTTd2glznUaO/fFYO1MB7DkUApkxbymDFnm6t9F1cd7YP82u5x2zMfpGqrq67nC
uwnuRu1URj3sGU+acmflpxps/xISa2ybkaeBTjJy2CMry+SWujVoyjm4BZ6CcsPeRLIYpwoeARJO
Hk53o/DXkEEyiR3uQIQQ96zjaZzUZDZdmz4U7LNfWj/BTY9tLihc1lpVAMeDS+xewQDyhXP+pxBU
Rr0Wofzf09fZDSWQK55Q72Xwwg3IVBCUyPK9qexvgoQ8dAN5zCFAhu9m98rRjNWQSmS2wT4rVU6B
Uv52rtabNhTk3K7oPW7I3KBjFUlcj6sx2y03nDW4CCei1pPJYald/QJdugv0G0rbHAug2V9fWQV0
vxlI7WhAFCLESchSIcNk+sDHiQeK5j5jApZT10SzAF2B0+bsGAWYaaaxDfhvzXSoB+M5t6IGbYaG
9zqoJSKkfVNxveK80xXxGMJbCpv0DdAv+869XlURrUpbyd73JWelRngwEdB5p7mJclYp4G+ZadIR
uL6vlbc/J8HW3LsdqVtSdBlUDRcI1beQLYmB+o5waLHxfII+CXeycazaDhezNFYSyJ28xq1GluEA
BaJj0tJA0Py9MCGx8iLRjGNm+Ms9DMWHBwZUl3xyCPc6OZm/bjvsmT49rG0YLTulMM7IaMYUy/i3
aQYE/MVIZddeRhdK6emKxMQgrQxWP6XXRetVx50ONb30LWlclF7oomXNBJd/dDKxJwGZYmVxTGYc
3rpZK6qgYb8Z+AGgUPy4EuTgHnxHQCVzZ0gbd05yd9mb1a1/t6XU3sbUXwG4Pcs+JrC6dR/iZ0B3
jKaM28jL7EwaEmsN6i9zVshrVXyIZ7lkh2UUuj5NzevKu6f9/OyPHmKkHWiPW2dhTtPM95MnWc3P
WS5DZioK/SkkSkPoqOtPNQLD9zVExdXO4aLvsHu78lGUIibe0YUNQEhTibFabEujFjF7v2yhzroS
pRbizfMwKJ8myFqJdC96Iaiw+Rd1gNbvIu6N5EwNrjuHSsBrzrOyfV77bYV5g/2fmTtCS7PpZvcM
FAf++AcW5YcneNdnUOjkfgOZU7Mf0IfupL9r7TsZsnQPJIvpGX6jt6o4xhZ4LMFinl39nuVrHdC7
kF655LMle8ySDCgTqF3pLZJ5g3lLJpjZIuA247ftuaFHN9JgAt4GGdLzVzKIhWnQ6uyHOevhmEYQ
DhBaegkrvd/GruYUpet7c2j3uOvkWs0reNjAYDMfDZZQZFGqzsjf7X8jUoqYGSO2zwngiFcXrM0j
OJ4eedncP2qVRKt9qV0sXsrr+rO3esKBQUgZNbNZCah7xEojZJq/JW5GgLxd/5gMpWSesOT+rLII
8/ujSNenxVdbv7C98hj1EOr/+jppQvvqPjZD8wSC5Z7/rTDZOu6lBpdHw4xVwltEYSBigoWdslMh
AgQoyIzYjaHUSJBtfWY22VoS2MdBnsW3xjngTNF9UAzaiHzJtYaROgjGt22XWBMj1QejCZc6vfTa
PHfsH8bHD+WksncLjNl8ZidyGjcNuuGDNPa+RRnKRzM/4JXF7SMHf0ryRh/pNNz+LODrGJk+QwEa
gdIb4t0Y3oc9gsu9ETJdVy0TOsIwbQ80OyRn6Yxm1rQPmwWm01hgzOrQ+1o9PbEwZQakyIzBm+PT
I9E3qwrhYBRnkVzz0VOkbra3ot69G/KA+Q378NO7OLwfxnQY9HGdXJurn5Tk737qn2aYDlGSxCrm
ulX2DqSRR0eUNYBYiLvQDqdd4Qt4mOCpg8GQ19COtG3HQtvWyYPQwXCidMxXxGT3SauMFRpOxhsV
gD0fWJzvJZtYkEVi2Sd5S+jOnrZHOiX7PlGf0bn6KwD7BKz8d54RLStGjccnDdM9dmbPyC/0SLlN
SJqtCTr9z55yH2ZftvoJRH/fTMp799ChU4aHlt81C5YeFATNnBQ0Ktcs6QI9T91L9376ooeQlVd8
Zz0fPcj1g/AucU7fOC6MfqJ09wbS1JyZaNH2PaXK6pL9CFcrTw9u3vh4pGo+Uk1+BFA6Wg/o/K8Z
KGA5YGtsd1O7I4irB14Gjnk531DP6BGdzIliLxJER7adlYcLQA1zYvAvujOWwWywN/mNaH1eGka1
ze+2Pk3O2hfwKgi4RhBBg48B54E5gSaL/4o75GmdsPxsRKBm/xg4FROdbh3jbW12VusjGZfMohXq
Lw9CAgSVKt5lE+jkgWtvyeU7oDskh5QfRfWuppdy9zHPiYgM5wV87RCaHMfZg+DRgSw/X51dEvJb
WU9hTO8hHuKyxl9bqQ9KiHDO/JC2J3joz6MdWPmd5Wz4eZxSjTIYKDpF8aDH7077kJH2MPygKLiG
0b8zyrIG/+61bgZZZlVx0JCG+qDjrpqrKr9K8riyYCycWuQ74RoomX0/oQZJ/3S7P6MoCNLV3k4M
8fgUJmBs5GKRY5vNsYTo529xu0zAQucFpeMoBXl0cNsUYu3e6MVkLz9EjD80RQhaXL73l13pX65S
jyQryMVUMxAaXmCQ/gRZLwLLSK77dxosvwJOjxiYhSUaPjc/1YRkwAHIYW/gW5SUygEPgClE9hOn
so5O/ly/JyzZFFLwx6MbNqkRjbTZq8F1cdj2DlEVdZdKelFBzkKa7Nu1DMkkCgXl7j2xGJltjb9+
c1JtjGJHZ/AknLu19ANqjwl3rtfa+CzLtq8mGN+e6wO9uFDpXJ0sEZxDQB/rlQxMSKK/zLvKVc7N
vcCVatgfX8UT+WNl6IPXgyiRQHbfuveMY1+JEqWvth5D/B5DnaZYNg9ccOGTDL0ac4YphpVnl+6/
sO2x0+nY78vk35VgBJnOmt8t27Bys2LJdM4Ycd0MgdKI4FbBMC8xmgiJ2HMHsztsBwyg55LoJqrw
TTVX8ULYacz4IOY9+nE5Lm36YjOei1iioff4Z0GxvIuYmXfS4E//B2cP9VtaBvhKx5yub4wq+9Nw
t98Xei2CszHRHEP8Fp4kHwizX9Tk/GldFK2WEQaEx1gRQexa25Kk0UygK/cqhz0uqq5FxwFZiTde
p3G5oOEOIfCidd+z4R0XSsukbQEeFlGBPX3vn9ZG8Ok97ZPlvarmDv1fg8eNQnzybD2y1wMJOw8n
tFmdGyaAM0OIMtyGDJkt5fy4wm5PPexNglKFK+l22QjV4vh6LgGZbRlIVtraKTyViCx7QvnLhZFA
DsU6olBdVj59nnkdRHR/wSSNO5ChihqOLKcDyywBIWeOuewfrPdNhqkYCoEpKd6YoypNYvob9Rk6
vVQhIa55L6FomJkug+Wti7wzzyJfHH4RZt7tzjZAOFAdx3ZT+WhT9niJ26omeP2BoY9MhGunI7XF
3ubX1SwyZxzMmghpOvxEAG+OBad7vO/Xwz+L7dFUUX0GDG78PkwZhRSftav71q2Pg+Zc+7d/r8Da
sznYLXslJ5YW1jXXyz5cDwmIu8u7TiFFNTxoroRBOf7AvObiuCFFmfugJn3GUMIylecZGNOZUtOC
S8150ZuMAah0+DK1PLbk1kS8308pNz0iIBeTml7CFV0Vj15eZnXDXrMQjXe+V3lPt7mPvWDhPx7t
GsMneIsM/jaqG3RHMGPdi7XlIZyQsilSu8qQiYvOz+sWRJCmU65QZ22Z/PiOVX8QMTWRyAhcnNK2
rJYxW6HO23Ngl20aOyx+VHLRsxFEdhPMyGMwu47FMJ8ANZ6Ugi6COQ3rDJYm7caIDX0LGpdII3xO
HJXNTGxxdkDBTdbaFe1/jhMowkszwJRyJz7qsKFHL+pcybDff5M0PsK++p6VvpiTwrFWzZ+W3v32
xog2WApGiaHK0hsZiPb7pBsOT4dWV/Shy23nNPtBC5rfNZ1G4x2okViow8CYHbYW38CC974G+Hl+
Vle4cqwddMTqjUfqWEydyNVPrulEk7IK39/SFHeL3WTHL9k85iv981SFwF2LbR/gm3EyI8avIiAp
h74al+wqCjrSKg02+W4xQf5mepVuFNrRzJbAsLJANYczygieyxIZclIS0E5bv6D0hsLKOffBGb6G
hRngk8mbMFWmrx+O1EQU9kxybOgSKrkXaJB5csELc8H79bMA9A6M3flPnbkX1TFfWu5LgmZsDAHn
XSMhRqSSMEi5tWNWFZhM/pjfiRPUwiDF0K5vyRkr6ly60fZPjB+jCxRWH9ksfxqlb7RPQ7Lg8SvF
7nLtCagJbapaC9XLkoJkOkEpL1mVs2DYkUXArcV2Z7DZyp8qQRoHscBNSNLkN7gpiWxrn+IN21+x
FkRw/e4jCKTqdnqfMA0ooiBfxaxQEwT+LDQN+d0NNka8rGcRpjRAV5E37Q3HsYCMuKmDqrS9DPc8
XokkxR6tQZTRbbxOf+3YgNz7Y9uaSBW//T74INTcZGuq8QffHp2BCFOAkI3JqyxLuwKvqNEt1j+h
MQz9eP/W5d2kvxTVRmW1kkGbQPr8lU5oze3C7CzLcMzCYUvRLg6xhaXm0VXWJLLSPtyRHbcTUM8I
hnrH2RqnNCgjKROrF8k7xZiNb2InUQE8q9ZvJIFM+7EEFVCgAn9tjPlkJ02f37OOFO4FwSadFiBa
WPfDTjUkyXcPh/zO40r4fj7igiG1Pk6YNeucRnUzxWKCMk6jkj+6apo8k1YOTa5vv+iDicfH+VI4
OrvuHckxe63C/d4qVm7UW7Xw5BkYQCPzgzOhmy6UT2JSkqbcYqtRMomVw0eA6EZ5qBK1CojPRlym
geMdqTR1NyVetOszFD1Ln1Oqv7XgNIqKGt56//t5wlGzQh7CWaWP6gd7SCu7gnrQj2fAjHzMr96y
ZRYsQ9/YdlCJNjyTlkJKekbsVVQQeGrLgLhypq/JmVTbVKptKNfXk93JG08KTMCNd+t9hkNnqPUp
lllBa1utK7Fd/d/p9hEZ8pKsrNn/BhdSKXZRey7ngnM4Sr5IuqjpImFyX7jVLjPBBe06AH7cCuPb
8Ro2Q9/AEzjU7kMlBGK5IyYPfDSd7ev/7l7bmkTWx2DRh0pzO8zZOTHomcoyMSReIDw+MVWsql2c
W3zqJ2MCyV092jxKunpB5VVaReW+ogzlB4/yyFULQTSLwNsLCWI9NsBhNsmxiMjqmsTNDMfptwy7
vOxdayyJbR6tlhn3mCtyE4aG0WRdVUM2EgERPYu0c/8dGiAGo+8rOa6xjBqaPMkaTbF8Lrl96BUN
9U2/0p3oOjlKr/NrQnKmMxY1fu2mm/6CiPn8JqLWzf07r4FD8kHuA7WhRhwsqUCVBzS2MASpBe+3
iL7kpptFM7kMaTgeBYmcgn+DyPTfhgKYaG/d3Xz/UOPrAZRXV2nwxKRVXfaeiGcbZxAQCbKj1bMs
OW1KBfrJJXhn7VeejLkwxJS8EeG+n8PpNadgNLx9R90PXSYkN0y89VF5TETWFCLnP4dJMwbCZZri
Rp/Lt/HlSssxcsDPdNuX5JpTtgmxkRXcGr+LptSiWdkJ1dBMf9+VLc4IA9KwJtyRZAvj2KgsSwQb
JtzMrgNafewk/eoDVBOc8Icrpye80T9DUaAblG2gQely2wCSuQMwbzfde7zk0LLyuaK+Nvlqhoqh
M87RwB0t0mAzk0GFJPBjxAqH6Mrsekjdr04PUtOeT+PS4mMqF84QZBuvL5zTqDdMoTW8FtZ8EEoc
v9MTBlTSFSMvNaa/xR3843uKG18mQWqovFm92oJFDGXVC8ghrnAmHlWztk9cFNI1xQCzgUIvcpT3
oY8cXqT4bnbNRs7MbIyWlM/dzmVDL/GaAnQMA3XWoSiiZZ5urJoHy/zZbmqaIiFCc86pVz1PBkVD
eCmI0fnyIDGRdd9FGkYoNxS7VsvxfDFxi2C3/L1xXN3MC41brHAwXaZZ7LkG4bZY/Gt10AjPnXUj
OrZcSVsEhN8Le7T8BblV5Vtr0NG8hj8DKYa4iQqpj5JEKZeLfX615gsGs9Bu+ViOkZjif8xCQ1yl
HO76+MYjS2WMHBQ1jN1zfLJlmq2gE3lZnIFbSur7hYFdyT/pPK08LEjjI5LbEyp9UrvoteH9WySv
dMWQ3zXzhocIYLqVPwjAtartXJ7vKswS8DVvXs2aIrUads4KkYezzCgji3fmqqgygBGyt9WDlYqS
mLs5UJ3V27diEj2f8sUnw8AyYHVkOCtI1rInihsTbOq/8SyjVMHRhtr6tPHQhPVwIFsbrCVZrk5A
S4CM52/kMfy5kUNdUOXFYQZQfTOFXSzVKRSQ6M7gWLm1GNCB9e4Wmkf6ZSVqMBrh36RFYL5rntFo
eRDL+/OuxvJkjIXGkVuxUh4kjdIPr+I3OwFEhzRcqjMEXl4lViwzCsWXHL66om7zf0nN6eRgAILZ
61SvHwXQShiHFxletPT3Yv4aCOT5fT2eXiYvWRlW/V7ZdfKfKcfhxUtKKPKmY78NnzvvGJD4A9hh
xql5AG5ce4pxdgQe2vFh6m0tn1VT6OPfV7+pUpMR7OTJUWx4XQRZLfwp0mOfiB7op4z7R/naQ/lp
F/AWpwJ1wqCrW8nBi+94KpiUr1OTnIuhGDst2MpOfYVlfiYSuNH8smOWUn8Thj2/VPg+d2Fjm8fo
9GQsao8MtoigmJwE1ZCfG+56Yq/faFRFGT6YG603GrIiV8gQ0+k7BHEKXU3RvE+ViqLvSZ8wNisq
ho3a3Lf5ScuQRZyrW+Mir4JlsxtkL+ockPOADCW4A8jyXtZL6Z3sUQCk5kvAsjr67lDi9D0NZhlR
hmUQHyIfSxV7DX//2IgiiQSxd5RoH6nuUxutWhJ2EnkMGLZXy1fj9q0pJIzL3TMv8qxAwG3TJvC6
ae3+uu76Pg0WP0F9ywrM9UW2SXmWbTWUbV5arUgdq5SG7G7xoQ589XW5gNs4DFpfIzMG6eLwxKhT
1UdD84vqxIwiNgCdTdaiYPEMifnHbsPasuamPCQhVFOksyg39ePTn7NB13IFJ+lLwWekH2vdTaQ1
7awYrg8ZBpTj6HD/0GSvlGsrS5k+vzEv5/oGo9uHE7/FEaTNshbHByi3QZh5/OMTNyCmg2zbjMxh
Tca1PRDxgNZW/TpzagfAUztZpqoi+Ga4w5HLC6SztpFCuy0fyH3pRl6z1hZOYcS6P011jbdlrwnC
fM9/8UWd94FjS7XfxTNc6xbRXF6tvXrM/GOpA7tjxlYgfzXs2X/0SSj/uKTZpbvlvpRmyxHybs6y
tQvGxKPw4ZnLv+83zEexFcNqqnt9Q/YW85I/4WPoObAR5GhEMOJUB3pLQp8weiDLilNlOUckg+qy
ddeycWKlgGYLa5dyksMHQ7+gsVxH+siS//lwQpbvUboldx1eiq/N7mNQaxMP0gJhGC8s5lccxgLb
53zn+f2oNV3LouNVFAgMtS5v47mc5RVnajEs8WAKhAPf+PjrOEbuPcj47sReLabufQmMNx3s8e8v
nCVbHQZs6oVbdpGU+x/e90nsqcftgIIPji4v2nto2NogtQLbeDXutcvsx4Z6h4P54eHKLDnHi6xo
O54zlKvYiO8CXv4o5NjZrd8By873mp3YqnWTbkXLkk7LzC58NC4HTu0U4rXBgY44oCOzOEHeO7Nn
t4cl2SzdYqNzOV8xJVmP/M+GotOod0ssj7gf6LYyajzeTc0jhbr0x52Qn9jyd5mm91KjyR4Ed3TS
OouBsc94yP5xokOEYOkFP9wjpkRyA33maujiTUaISnxQLJoozUHcLoXHXUyEeq6L25/ETeW5CuZ6
aaru9nBgMOFPthPo0FxRGcgpvC9cHL0LjJrOiSBBILRwrjgA6c8ttstgQGBfMqckN5J55gI8D4rU
3xCgPvlIXonwC5V0WqzjYDBywUYmBnIARMXW6+gbE7Zm96s1YpmLvhiHFtDYT1gue6Z8P2sB2dIc
1t7cJz1rwinzcKgB1KYexs8eywut/Z+oCUXw7+7a4QLXoRECnv6PUYHhMn8Q2NXEvNDa3Fc8ewlz
AnApw623iL5vWAsnaPi4ZXDyLCA+sytVUg+3DI1ju0Nf7ZQcwrWyS6NrP9ZvUupWk9t7+WB2CZbQ
fXwmYE/N15GfZS7IOp993zXy7ngCLpbrGPATlx/S5lAleuuJgBt1Y2o41eInj6ccOheW+6vh+c/2
zW6GFIIsK0/ZHbcg2NkWcVhhdyvsWk2GwGVJ7CXzwFMPo29l7urvD9i+zszHyGlf6T9AlbKNyjdg
TQr0P6rGc6hMWOj3P8zrIKfQkDPO5ooe7W/TbFMwV+Mbgbu+qx2Rr3mvj9NCyDvrT2ZYZWM8p6fv
4HJE7hcmMheSojUHpur1r7+uzwJ11z/pupAodUKzGDKb2mkOObg/HNeTvPPxIInvdibZUPpBjhg2
XNAidOUc3WlswQ7g1eI35Xyxuba/kPVutS1wghgI1ObYT0P6jkXughvTKCpUSS05kQd71Zl0EtvX
089+uE8khegVFH8lueWgnMmEOU4V21ccVgqAHiPJMP4RD7kFgYEzC0nVtiJjcPp9O8JP919+hLkR
R1l03Y244akbsilj4pHzRISDvctSn4TuRjWbWWUjzycGDTvY1IvjxvEfWaoe5hD2mGjEQEPzsq2o
6bBc7OeT+FXM8n/y8JE/A+B7NdYPAcaeiwgv7LDTvMoPGAsj0Whg1C9f664z5Rq/pAALr/TOJkhn
50kA50ZZFAJYJj/lQKwXPcLiSkjwLrapXiiTdbAnpcO6uz+kfIqAdk7N8mmBRptN2tsqK0PCMu9l
EoUv/pAsrLcshaxvWscPnCtS0e2vp/SW+Zjmh5fm5FPEWdJbPRbpd1Qljh49VQ0Nq9VjDtdhuVch
dvfFLW76jFvV/JgtzwWZVxmFKjiFMZX2qUk2+eecwuZ2nA5IASdylS9VPbqKdK9X1Dd6N/F6GK3R
2t8FrHTe+amZr0G1LcOE3AsrGg0MH3eE6j571a8N/nDmBkeQNrgtLm2Clus0d/8T3wVYvCIoSaFU
rJJh4Sh/r6tSRiLhJpG223Q1b3nfpBtoEeA8JmL1HODzMZbuxIBXbzfulohG2c8ukLIR1ZdA6+IK
U/QHfZ9Smvv4rCJxSZBYC7w8FvLaWnHrkmevpcCzqtXA4E9pBnISQeZpkRhgw1sc3BaqNQ5dnWUX
aEHB90QDYA6Oau3iqpglqF8G0L/62ZyyhU90XzpVd2rrOMJy+4w1Cosya2axCBHjPsNxnakMK121
KP0XpmIJ0qZGFc+rMhjuFo4X/Nx8cwjAJiy7jWiK4vAKWahnOwo4h2xsBR4h7B618AZSZheuUQh2
PdO/EhXgZWLHUmZaZIfmMBl/pwyV7DVLXZiGgubbozIPHHOS8/Pnzsk7Y/fK4njrLjaxBnRWI7xX
NXbgUo3996Ne2eeP0qbt3PB0OXgr/A0MupUteL0VXAUrYqhB6fmVNzahLdJhlJEqGXDTvLUGtN9o
xpW7siH+kq+cRVZ4PULjkcEfzMln4jipxu87M4JRReowdvXmcKBjKekJ2ok4OIvpo4HFxz4ZxN4g
QR2GJboxgAL+bwVNUlf6G9F8CR/f0ZR0W/cT9Nijprl21TdveyN64clo1BbKBMcdAwrOP91Ga+X1
z0+FsNKkbNKXVShaopKmZEui+MK2b5Bw8r9+UAnL95U16ZPcl/krDMFWYeta5cy1VR/Yfp9XOmf9
dtnkW3jBkcT8Z1OFlG4jKUeY76XHRf727K18JHhKfhg9ybET3fPfP6p1Y6jwcr1hbFNP0h8R2R3/
bdgSVcR9Dmz39A9ErRF11LI54iKX2vBr5iOTm9YkUQOhj9sELrZSkuVLvocq1LLJ0dlV15trgZMD
hofpg5+f/4W9YKNJPCtR30EFZ712tzfob3vKVgE3SW9u9y7ZxJbRMog76ufnAmV8nPCGsIzmxFvp
jWrpJ+zvJLuw7Pw5dd+4rdQA2wHeVybSR+kxbtKtia/be+K4XmJsjGZ8pZnfTPgUuKRPsLZqsUUz
kfidBXxsSj06sM+6w7PYCOfa2Vw6FRND+ERuD3MShriV1AviEpf8H2hh6p7jvAmdxsg2KdPUiqHR
85aKLMOYXA3jRrNxFtG9BbAueZ1Mx4oHt0pEBY3ygro1i5In5cQtQPwRrnnrXLzT3WCk444XoLm1
TKxZSVKVX/u2wsY2EqAqtuVJ2OtvN5QOOpMyUC3HK9vyyE73SpD1q8PR87vfEA2atlk34h8TZRnA
nLW2JwUiIVQ7mITT+kqLwAf/mE8CM87+o37mumR0AtGCXdGqMkeS6DHGINNxAK7ip/+yLT1ptlQy
x+zJNVLCE7ZVoYAqit7YaFPDamxNnQFOSmqRbxgTlSYCZlZQ3uqUYOLakXG7O0q0WOpcvSKCdur8
Qr0/Com8F7cFy6pSwEfvDjHkIWjBb3eWMAWTqzXICLgccBz404B4KxNTrku6soF5cXSX/yy+E188
qSfPaLPIt53oslKNvAhg+ELlqCUE54lQgFJ6smh59aDV1H8JmMYm3pLspKodM74O8B8WSChqkatZ
xGObmKoK7B/A1IEKfmT9Z9iuCuLYKph50jBT78CFjAMMwa6A4Dj4ipjM3a+uUVUgRnyquuZWDCbu
bnULjz1hgnhnZFMCE6al13AjiGJyxSKeJPLbursy/YO7xFe1Vv714m4k9XBs7YZRv2cbTvmxzASj
VVSyjuQ6yZ2l2VmSNH/V4pBbP6inJHL/0rjrY+MZHzwKYZLmQ0GzXk9UAduR4UA9y2Rg09A7zcgl
2981SU/2Qmm1bUoDoy8MqLx0h/5wsW2IQqUNppPn2LztcLLRxWGJtUnv+gMjBHbBWrbY125otejb
Iml/EUcCpEw/WZT+myKOEZ5C4hn0rCKGhJKTVkcpxKXAFYTe/PQ8Rk568EDzv5bYbuxNOYmOd2y0
HpZe+Zx+hIslNcIq+clk+Rso3BO+KdZe9yQ7bBpVgOprhNVcOP3zrUkL2n1SdGOK+c355LQGX+yA
Bn80whePKzz5VL73BHYAFYdcSbTsaWVTGZ82X7KXeaWr8qG+eoWH8581plgTEnh35KUN0PiidRP2
CBoSyttEpPLVfpdlmaA/4FFKqj5Ap/kqjIHpvkj2wQmTHCGEQ50B8PGar+hrfq4e1F8H66izHI8G
tTt+eed4+nkP0+IuDyf0VI1QF+TBMcZWi64pSai30a+B8X26HwqoJ95Bs6+aixC2zmw8gqG0/WW3
w+ngqepNniEhJLxPAYzcu8CiNsrPccM9jHa35ATuGIwEoYjTsZFTLfdn1PKCaI3z9Dvz51rUnTCl
ftDZelo0powCvvZGmipDtpthdG42uW7tht40ayyL2M+jtmMpODY7vf6gLpfgmxPTWS0zTze4gXdV
AjrUv9aC8VMJpruKmHBJr5qUCoUzWpuPA9JbR2cjYvWbN2lmvgrvUPM2Tub+N9mEAW/XOSAm3rFq
AoRME+jRIuSnsrcqnkIgQ05hbtxC+GfexglqODVGLjpJ6Mt7C1L3g6J0e4K33Uaebn2YHJ6AhM4u
M2rAQBAFFuQdEXqnEst3oBV6E5HHmuMSvR2rGvojJFca7SmGG/o5xLnp9Fubcp2W5s3qNmmz3kIQ
B2eArjycKrs4t4VjcJPC0bkR9BZvisq3v/KlQ64qn/LVgG/vu6NDsA/UYHyXJmHCndhfXCdt+s8v
MGko9PW6PxU83B34G9gGS0Xz/3gGZnNNeUZlaOJDdVN2eNnNbJeX8lvEcv2Mhu19/7DkTeVc8FzJ
OnIIrWt7i291J5cu8WmQ8OUXUAvFti7fboYXXSNRG5c8UVxpz0fzgYWswk3b65r/fjgr8XzIzo6f
Ooz8JJurb1Eb3oxRihA1X1uCVDaxRS48IlbaOwSxOUEJsguE7X7AZuI0RldFxn7JbUjcATzT9a0Y
4bz61FezcX5HamNQV5oMWHsVqvJbO5Yga+A89E+6gCBRwkgEHhgh++jcIT49lrdWT9WQvnjzYQvq
h8Ov1vmZL3yaDWYNitDEqWQzpG/lNaD3oUCNr03wW+F2KBK0Dk/pJUqFglqZw2KEKm5cLfTrPXaE
MVQ2M8h9F/i7FBVEbpjU/NKeZYDBLy/76wXsvNS7AAgUnLt0DkBJ6AcdIqdSYlFbEvdvjiRrklFh
TgmepKCMobTcWjx63Lr3oZaBCvrVAHEU2r0wWX6tDVQ2X6TyzEc/bNuqRc6PLWYxkjUZDhnOq5vz
xVzRILdbuR42noQ0xPbGipFytJtZX0Lv7MS0ru4hxVJLeUYmaTdSc18tfJsqbSOd/bQlH3pAtf7+
Vqd3cLDNzYtmcFBnC+njWeojlIaTf3n9Nc5Hes3DVNSdTifqfofA0Crjm4xL3UVa6VtElrNLCSp1
Soh7/sUCw7YUcgogFMYyKpIv31IFfUvbcVcP9jxLjOk8iR2gt+cQe98yOncWrmsZ770/v1aIwFbw
4tQntQ8xK5PtPvQMSBKSmbNEzd5BGS81hjVcyeF+AfdL0XH+qbZNN4foE4G+79xpp3dTmu4cMXwN
FiMQxoQa3cflj0ls+gUO7gHoThsIrfG/NLVtwsvAGbIt4hWdKDpZQwdv6oaAg+gE9z5HS1g9Kkcd
+K2m5wW4bI5VjLuSLQED92OY8TV1rkx50QZOqGFd1XN48y28vvU7kjfuOh5xzLJUjlKFhmr2QyuF
9qIWef3IjhTm/OH28dtCOEURI2PYxWWl7R0y0RSs0RHPzP05IpTiq8tntY2foOx0ebGapKD7iMnY
o6bTEF1j3QsF5itMQEFY9vLELycou0Dcnwby9k4PwerH7HW0XAOR9NtTmI6JIuKrHarY6sLpQD6w
1rVbG0rYLsg9KNek5NuVry4p+fJeOq21UNNZFuTNSmw2+tsLiIT70V1X8nkjja6qlodwW7ufMqQe
CgnP0mMFzQBLIbVcHW5nNKaAZJd6FrW16O4I8lIiY294fQ/tMhOXqZtOw5rKxITXhGVvb8mVOPkP
K6h8HSOoB+1BnpMNU9XtxzK5Smp3DZ4NJD7wl7AEQEfhp/Jlh5+qZvrM3AcJLmJRTQQwT90fqsHh
W0KIyda0dO3/nUqGDtUQL6E4nGZ7Wu6mMRN0nVEHV9kzUKIm6295MojxHTZRecm+6Ud7Au+yOKOB
Y37ZoLaUCgmTcuMNBsnaEQSAQfTi2p/OuvwDq3MRRbhbTZSMHttH2RqCpGXjjgdtlQ8S/VVB78FD
VM3C60mSFlX9B+1D1AtArSYuW8L5/0CHIMA2TS5VXV9eO/9UFwXSqaUATm3H92eBogjNxDdHo2We
TwEXfOXhMwpib8w+lFdlkyOlfXcI4xjs0YWDmL4dFpOcFeFH8j1HVo2xIxiQHaOTAL+e/fhgoJYs
a1jgL+xOb7ubx0eV6npZY6wsKQ2kNzl5L3tBT/TiqYMF8m7iEZX8gLpCmn2u1BGYtNKw2xPeE2A2
3aaR4EMtVbEoGKJiYxM+LqbPF/a4JjazcjyMgHWieEMFz2hOHD34NGwSZiS3u5qq/O5Wg+jCcCuu
NZ7QbYdKSTsao/JiD+iUfTni5ZOX5hzX23nJbOGtocwoASuLslHIA1r4/LhO/jMtP8KX4UfqCnQH
gFTVciMJ4wHJ15GU0BSCupFsygbl1MMIvJhGvdaWo48ugD3nonpLTZZmRg1XfCGXtBYgwpV7B/yq
VCAAxbcL6rIZ2cnLq5VoMMlprUwLX+hNl0aKiqTg/6VPTNfyFSKn3dI6RIOWBwtXdSqifnChKR5o
EgQBxCaMgiKc+ZMTJ4Y8JjM7cfI7jZJkXucadMjSp4ArA8545yv+2J+yJZBAaMhWn184ML5seNcl
n7ooDjQ2cGR/Kif5azK7G5fdbuE7IoRyxLYXDePuQDggJowr+C2VR9s247z8fmPJz0fVVeHJ75sz
4vDoLvRoT8I4xRbMkgUJyRYR6I4V/QEckEMT/l0L5haK0wYpEAimiTOhR6x5ZRlguVKXgj/Bsnjy
pCD0dLekcIzUx3sHS+vRSABsen939UNw4oG0syoHNDPtH1m6fLHIbKulYK0LTK+mVnjuQV1EuTce
IZy0QOc9wgx5zQAq4uhfbnZKjyCVU+ir52IL5R5NeV8hPslHG9MCFCMUtPW+5i6rUpeUSURsblil
OMH8RTetIpPJnNNQXyyDNJhvCbhM/f6Ww0K++G600X4MAA+SNsk99OY3r7ZtazxKwBUgID618Sap
zuoF4QcAduAyqiVHaI8DgX6pETUEVZPeYopFiVBSClMK+kdxKEIsu6Wo4CQaqU/0kF4XnTa3E5WN
C2guLJqBZsm62OsBb8oEtaUrW1B9DDu9wCK1D9+zspV/iE4vfo0JcwN4qlU6jAmKKzq7yQ5I+8p+
4uEroTeWUUc9WPaHQD0MmSdQM9z2W80cwSIV2mExYs2rcLXpG9HPaQRimaX9EmjizGr4JwKiUSGp
i6TFzaZLZh0/OI43/XaI7Gd2LXCX6vegz8SsCiZOOJ8kILpExgTmAeaTtDcYf+m0V0YQfFZcb+a8
WMjzcDYdfcgukLTDkbs2TsCN7pZmy5SNPUDeOSJsS6VVl+NUVD1/C+3E+Xs/eDr/JheH6L9XH6tk
osV4e0KgeUN1LGXtfze385T3eqfukZvarg09xIlUSPOnSmcbZPsbpStaQzsjVyqGrh0yeKp/2FBj
OsDwVU9UZ0BM+H2XNyU3ejSy3rZ6cHeaxY/gbShYWWsDfsP0kGikVQdHcE2bP63FODnJsHAXYxMf
mFW7NVppoxNepWDYkz/wqUOy4OaDCFxrGWXZKy8ethCBT/gJCCoQEw+QV14MHvMhWBbD96OqBXw7
tK9MdRbvPBLXYjq1THYd1O4o8x9sF6up2yVLlLNFyPN+vPeYaXuCCZ8qwkZ7jn+WHx+Ja4Grw1xT
W9wmNf/POXLrkjqQRNWHuVf6VrCwQF5kTzw0W083E8XtdyTa2SjgQA5qwizxH7+NwnuSJkQXx/y1
8ISPfz+baPomvNJpPLIQ4paqisKcMUyDbOK7o8LX89i0yngKa/PUMYl+FtNRZ5lv9/OwqJRq/lKt
XBJ3dr1AH1TntFSImasXfC9FeukfVoVPk1ra4s7ikd3TP0jooxFg25wIDIrTjzwnqvoBZDhNO8L5
CpQF2+w+rcLquiiCH3fpJbJiXwVppX7PugtAc9nB8X5CriNUHeAgiE/98/csp46Bns0KU3OHfytI
lH6BPJUYztM0BrowKrcKX37knRD3h3Nf3vnNkouGqg3D6enFZDqTeqOaRUiX/IH4zwHmMEqCDPCE
DM+5C2oluGleYrJVCT+KnuURutxQ0sNq3K7kbi9TagWqUd9Y9FncMMQQzw3ioi7Lb3Nxy0NO4ToP
F5EmJfpjbKCawjVVvx7K0neja+Cx0w/+mUstr6+qjLAswgxoxLKyrEP86wj1GFGfdRY8st1AA6up
jHE4VlNW+J9VYEjAT08meBvTUQE+yitJ8kQwe4j0jvcl7H/viUUn2sbZmMHhXsf68EynAJMj69WH
8yfQCUaudO1aNRcUf8JBlb0nfl63Sc2IWM5V8pHe3H7qk5vYkk5BMt0FbLPapXLo4vVLpBdrsT59
d+HFKDIS4o5KYC3H8FHS4IwDJSxrH8KAU0kADgXQSawb/Ea2xeZo4YsGzeezk//NNz8ew/iRo9Cq
Nv5lJCC9qO/QWjNyhFiYoLZMQdH4ZwSQT7Vge/jjunEyZfJHjRcqxsW+IvGk+7vE/yGgZ1hOQzae
cuuoGDH849WSTARbf7bXNcv2TWfbXEVJ2bPnhRDUmkXqJa0Z4PYOOT6bVtXakmeFSF4/2iTWf1xZ
8+2ZwQaIiafy+DwyguVAlxA8KbzVr3TKRtuE6lSopR981RE/XTP1fy03xHEVqz0Cz8wqbluNxV5N
OQM8MKhXt6db3cLOR45rDebmkqfi+TwSu3/9L829Rk2qnnuru5BsBw5tZ1AsctXrZ2vtBORLwra/
dhx03eMFXm6yfK/Fo3T7BQ3afTa2lQBsFm5N9yvyAglG/fanr+ciFXfx9Yd1XEj/a2ahvTVESOpt
7HzxlEBdsBq961TKKHcVd40R031p330wwu7L/0Ohpv9aGE5n9jH/pvZRGqZDG8wh4Ae/1BqfkK1Y
WOXEcVsU3Wmecp3o7+K8ke9NuvJaws+97nf+UeOzrBiffS0AXiLNWhVpUQ9U2eR8UowMTHkQ5fH1
eJ0aTN1+wo9GiaEhQWrNvFY49QZoC61hWAYblVm9tXP1huia83yiQ4mnQGNTPL8s3MWV52GK1aoa
q7VYm7zwBCBJU1NBQj9KuBAhaie2XYE2luWUhmsKuqLNcbhM+zFcJOnaAeSRL0oLvfYzgHnKR4Xq
A9n105zhnLIi+LKBBmkXMEP77IaJnAyy4tTFYyNJIk3cF8b2eChgLZw/kVQId9bi4xchWe5DHth1
XCqrycD0q7mNXWlONQScwByVwhGfLuRJOmClyDmccf7YaHDOI9dE+hVb+hrrNpfd9EIL4x9b9GJ5
vL30bsZfiFhmdYZaPZcPoE+NoKMPPWl370qFDfKKtjRy+/9KRoQc/FCUsz2TSyw6l8i3VTqWXDvO
oJ7QZlsQVopgt+vCtYsvpwcOXglniD+wxUJ1SS7Tp+69sl4QHcTkIbcVOaWQ/6zTRvacY61eXRDi
wP3FUEcyqmqogBd7IdpIEso//Ej0RMZNkDWCfM78Q9lW6LoHbXRGW7v8XXBLg5dqN8frT6/qgBJJ
30gmO8Scp4Kk6q8F8ANs9K0kvRXcisj/Gs0PLWwd/LM1LoTn9BQ7+1yPcshoif32PJSsWS2o5JHg
F632SgPtVTMGuhMstQoaRa6Ni4QJVpyEXbwGxQubqqpITIdYIKy84O+dzdvTOxKnYkJkJN6zoMxA
Y62BqLwIjRD8/L2y+YbyWz/xKdviWh6OJVk92qqc/fBaGxTUmD9vNZkWrpT97lqbtbbYVZln/+0T
xl8xgwFDGzCwd1dnUeFkFXYHhts7bmyh/W4vW5hv5JxGSriABhoAsiZtdVRZB7Kz3Vdoctf58i2R
P27NKIIJVt8M692FakML7bXOl74ywO3JxKACnhfK8ehuVxI0pcKDdvELEaO75O1A6eCIiV+mmo6F
/0WrwI4DI/9PVMtEe0BabnMHhdCKwMVHcTvG4TKqeIlwT2lCOqoC2ynmY+UhpFu0mvX6vzySsFYL
klUl5Nab+WCOcH2m3iQ4oU5MBNXyd6NVQaMpbHyuuueodh+drJ/wmaqACrG6qR1yfkKHOKjREpWM
4jqS4YdsRSVJgkyXoFms6QEQQAaas3Yt0oSU2Iq8LV0sSuA4tUAX/IaRjp09/oT8ekDHE4pJur6D
GDXgj+IEjDwRivJaIqgJwD7++KA/ElJF8i/8PdRiNHLEreisU93hroCMd/l4fb1JAhXI1fC9JeKZ
yZX/PTcMZp6NEGevEwj3/MilUTOngTRA2VEPsAtAzhGtf9HevtHB17h7z31LjaPfdTCEUxi/TnfZ
AoKCJEGU2SFjZIoGAbXw9JjiRd43LhX402RnOTzSLF/7mlflReezFJLom/S2LGrSn5FYE6TXmrIv
Fh1/CyTuUnIjM09wTKO5cY71L33UbPRTjRCyRUcLC+GOHp/838Al/JQXhSmKiZvuVZHi4D941YML
fCl8CqisWjFRCaPHZcKpUIIxMOaM+B+WPISfERY964a7eBNeRdMzwcnTtT1+ka43IPAA2ag0akS/
js7VaqouAMhrPHbgjq47f9Ia/hx7PVHrkzy35pg8Roax8nov6qB8jhnA70OHZwmIS2YELWYXEvJO
GYbDDGdMqVEH658IYcl1watwT4oXUQ1QYo0Rhx3TO4kTKTNtH+/SP+OA1WOTYQjZyb2D+QCCKldD
e0DlqR2Xt9CeN+9ttcpE31oXLMtfk3ya5r43QUCQRVfP85Mv9Luxsk1K4zvnAnzt4uD+sVPAFYz1
5+6CmUfNolhTWPow4ReNuH1X/7eHR50229vWLnxz5Yi4kFVH3f6ajH5FAtTq74DJsX/p0lORKhRU
A41+DQ6PPU4KL5wIl+DR8wfgNV6yiQAj4vpeOW/H7AjuMZHOWS6tGi+BWaiH/9DpZju40frUF+Kp
OaPyaxOHYOhfVIREqIr8ndFRpRzUeuPV2HhwD2BndjDF2z2jJmnrD/oEwKXjtObp6i4M86NAM0eA
pZ0wXLtk7VOdajjhbarEIuSX6wYfExfej/9sNWLEVZC5MGVCjFPg5/+ONkL8FkF0oOq0UE/4iuub
oDr6uwQhRiELXNCYklNsC7o0UPFU53tX66y68l6Y1fHcPuc21h4eSMVFYIAErU3+G9Xm2u2hZKqv
mXswymvfnTtuI+hW0itmybLAp0Mebt0eXFkynIz257BlhKf+ipBRDqyobDN4a2fw/A7UNQtymhwh
1kjivWtRl+qOZTRzNJeUWFDU021C/j+IxOnxcXu7eQt2X/TtZNhbxIAtbrfzwaJtQZV3lLGaKX/i
gNyVljJHWR+33hJiZaWoWpnjbusOU0VbPJ/1gvoUTXb0YP1c/84ZNf7QEb4RHfyQLImgCOXkCRJc
/g0pO3Zti6qP+TRmuaDb/YoUPdLBR70cxX5jkqot6u/PWrwMvwk/kI1ElUUHODmVopqWXSglF/Hj
G6m/OYxQ7toPu5delXH1BADkG94EX2PkSV+t+GajxESJDNaB+ibTCQpe2OZqMJ8ZdaR0mFBxGOlE
z70K9WVOMRB+pZGGJwMZOZs8Ys+BkOs9Vltyi/X/tMdcNHgTPPCxFNxxOeiEqdDQcXAS6kN/OugV
IrMSMMRnlOxu8vfRzyWt5ylYQIRMWJmzcUXWiIxhqoOUFCucm5xgPl5VeQhz/06OkCQWR0TgqScc
dcgZVrw4UD6NudYFZwVzOvSbeE9+9jkkoOApDOvOoVMhNnc2JNG0E5HyAcIbQ9pL+t0BPO8QPIY9
4p7LdXzHCzhB094pOR7SjIAsvsOEFdwKp93rjP+fnjpLi2WO0A75+RZL45cpnXuZu6R/5m3BXsA0
a8i9GQv4uHJz7r7AOFYekPUzTA1vu7hevcocNsIp4cIF42t7gHMIKKCt18+ufZkLDvwAsf1P3Yne
K7RPBSeBSkcfLX460Z98A6/4rKcg2jAKqFEKhmkKK3Lfs4W94zpGxNv4bgCWEOqAp0v0di01ZKFc
AQxhnHQlhILQ4xliBusF+TNVsC9Bj5UMVpLRdyExItnC6EEJ/6Vmk43IeQHOPQedxwTzi89f/GoB
25tMD0C65l2C3EFW3t5eA9MJTp/tPTKNG6EXq3LTabD+r+3tosR32D6/vFqolWEVJRSteT6onx6r
LPrXncIi/YT0FkO90SdU/ct/UWgNmdzNfjwkbH2VAQDIQuSjWBdqQgHjhCMwJdcr71tXumuf7utg
a6Z4w5JS0sT2J5XEh6gWQ8Vc5eBsialDOVaZfcya7KIO2pkjVM0e10hNL+Z5mT+QPP5qeG886dd+
p3zcOcR8fggj72kklDvxmG/0SW3QHY0XgLE/3uZXYjVdtRvVRmnf+iRIVSA7nT+/PbsOGzZrsRrd
Fo3GD27g2T59TREtSZYEk20DDV7YixeIMxq/45vF5ESg6uHi7UdAM7I7YfG4T1Ogyg+RQ0PBG5L0
Rq4gq70xXclB3z8ZEAaO48WZQieXlw6ILQxW8kbAwczY3v9ioWR3ERKMA5q672EYcap9k4hFSgoG
2t39j+Kyi2Q+H4085xQTiPxQPkciyWdutRhNsowT3x5sk4v8++WfGsMRjfFfNE7Heq/3D2x8wyey
ViZfrCB6I7dBNGCWMr1Qv4KF0TK2MmqNFvFyLKbT7hM+gUhdHtsFpdhyn8L3WAh5YK2t1X3D0Ylp
RojFrB/9B0xF/QZiPa6M/ttx9wexWlJ1sQdO9XbgYKLesuKyeNnlZga77OwGL3b7QnhyrdU8XI2m
slbMLqRTpwv9g+492iWlTg1EPdNmuswe48T/bwKrlw6Bv/mn52v+71hmlpVyEeLdKJ+/kCoUSTR+
LdRnSKMX7QFrOdel5akUNtMP9skNKPxHAPrnml3ZgbZk8AoXs1seKNhCgqhsOjO1xtDEvn9cqrCf
BPN2+XaDjd4BuVFWfSvYSSt8Ft1EWNYWTem2ErsrvIayK/QgBAF/7u2+Bq8Zk3+m89M9WchPa2ps
5W26EGkYcfah8fv+Cu9V6/t/f7FuJ7gd++8ISlv0YI3FK1cqsOrJZd6GmB496LcdnC3P9VwecbXU
SHXNf14Gz+N/emJKP7aLDKA03rcOE+xXHFzJDnqyaxvE1ci7NJ81Yw2vpotUGsX9FCZNWw33EQkn
3VR63joWzzPdJD/277MszXEhT5WZZ5/frHjNCvXOi6BXdrTYMnIUALQCxH+WQkrfB9A5khZTiVbx
frTbT27mqIAzyzPRCt/19mZkDabdvf1YG1nebQNbvNETkXG50Lj/F8USVce1Fxgto8F2936T28TU
OLr/vmMllPGDeK6d9H3FBrNzSR8QxV4phjjKFLE4Ab9e9lpHeNofTjoUk/UZD2OmUpRIjR/Yebsz
RBVIWg+fYRQMBjpEvBSiAS5o+Z2/y7B5QCH/QP4BqG/5vAvtS557wHO9fRoF7l367uMH/zxNnUBx
2QcAQrggQETzQ2XDQP2k+N3Bi4FDklhq4hcKYJKyqWFPysPAJ+1F9pSlS0IZTjzu6NDFEMqle1/b
b5A/KtgAEC9+nznZHGAR9W6tUSUIILvhNDXNJijufg2oA+mAe+4moNs4soW4tCij2jj5mArVriLv
/cewETpbuzvOPNR227xltK2nNudMuWbh8xcgLIVBpnykugfH22ntxm3vzhzadmW9HR5JlRbWPN/k
6QuvjoKMhqnZx+Tu8SuF2lZwbxfeuvRsY4PbW/1Yc8mCmhxYMym1Drvq+huOqWzZioECrYCq6Qii
o/eKzVk7+uy1mwdDl0vFnnK2Bl+Ry0ymseTCaLNMQ0FV28p4biUQPYIGJwPGnf8EUYDMCc1xeyF+
//mfyaeVNx0DGj0PIEP0Fph/nWJY5VbDdKyZ9uQ9SzmK6yb1RoRTnMrKWlqI2x1WuMyu2AlrGs0d
MvDks8Vfa8/ueArB5LR0calVYM8jPVWq87kdF1gTod8VFg1maCFhh1DENfeHeyQdHwf34Eiyut+0
qkKIImXx9eu7ImlD8ksZ9Z63hjVjfdmzgUhqx1dTkk/750lgATNgw1MyEPbORESCl6mR4ACwY1XO
Oz5Ym7CYrdL5PnAc2f1+OU8LOuuxBh9O6ahAVggm6jh8qi1g/M9uMgKoIUhXlExsJ5MuQt7cd7h9
lLAOJ00SqJbMy2dNMP1i17FZAa7R6pv2zIb8WkDl05YV6Fuc2FFf9EsG9E+8cqAc/8/axp6MzG7q
3W2S+2VBWAN8py8VOclPW3Qvw3QaQ3pD8X/jvoO2HzWo8WiwpwVWbF6kKayN+9zLENTfwwjtafrl
JIUuKaXChn8+gpRO/PK9rGDdXMB/BjPl3pH4mez1QL6niahouk7cBWbuMlW5QJbl3NbmXeZlfG5Z
wWOF2k0ueRvW7KulegYbBLkeLQe40XAou1VPEyHWxLYtBw96J35MLF1U2xfbiOC/sLJPsp2R6gjq
IZgEgz4/vNbatqTiVrUOfs+RyG/dTS4JqX5z02lWPQu2gaJcyhDe6KjLDYaBxsyHkNTyrgU89lZE
5qCSh/UU3/JChS7mm6F4ipQFNE1psknuVcGNOXOPsOcvi8V2gD4/n0FpMmy0dirume7tBkZGdffe
DsNJAhjrRBmUiios1NF5F+XcQP9jzAGAWc3xYNCVVN/sgIAr3p4S6HjPzKud9WkzYK7G6sML6h1M
aHG/h0300isDaEnVBOR5BX/lkp1IXxmIN7M/3QUJwcmff7KsXq7DQytby3sChJKzL91rBaSE6Y7a
YvBYolwKZpqURWXtrpnGaYqnc49p83uZglzidT5uN83IWVKPyRRVsf4cD7KV02NslwzWbZ58aqU6
KSlHfRi3ungPaC231Ppxkhd+/Cef7s67TJfHz6+qpOEWvDXW/d5w4j7rwMimzsWcYqzER9Dx+166
TG4eADXCoL+oOy4q/A6pBNAeLh4URmGYc7ja/vrlzC5ghyCV3wm66T4pHq4w0/z7dZBGR5PKmQfU
jQm+tNNWd8n2ULzYkDVEtxWL41gmxKuIt0qm1H/Q5gAm0N6EnAKf7T+FcQHLp20B4xqjrH0fHb2J
D7qBoMy8LrbtXFbbnDolNWlxIe1Sayc20G3lpoCTunhYKcfQUDrOw8L+4Rbos31V2bYvuuly951S
qFF/Ym/FPs7eJKAHDMCOoWORSpab1NW6HkZtIK0KrZ38+sdJwgSyRndRHdwpyTukf/PM55P+3p6Y
hCrHudGhqsv+94n8fTx1nQToGWkpD7dZx8Do2UpKgg5BgKcpp4BRuXaPsK01h6HBJaGy4NuaJFWI
E6DAX8JhApDf/FC+q7dBsjzH8mQHwsQfi5D6F5cNAefaNhFYll8r45oBSJABaQcKnwzwb8DBc53m
cA+JhAMHc9hsHBpSdCR9nhmRtn2wydW1SQwFLK+DJ2SA/kmEOx6A2Upcd+jSs8YlPql3wTV8ZkwA
TToanFISl+d7ZvpGTC/KxLAhK0EKS2ngABIlug81oCmX0dzXzkyD0wjoF4iBK1jpxjOlRh2T0jQj
6xVzULL9trvX8qpt31SAyW/WySOkav+TsbQ7z0LRvujHMTXidv66Y55achbjkcK9dmY3SsIIO6on
Pg8q+7TWk/OmSNci8vbgNlPH4CO1tyiwDgvpYGRGY+BMCzNGeQnd4h8LMC6G9DarHHLbF60+OBXd
p91nikxZqcwmhAjLKQqHx6ZW4OONrz0taPPxwii1OCCUC0mbrDWCviAnswFYKdCAIdi7pWxqdC8w
VstMZz0riV4JptRj1oBsuUrlX5NSjTJLGbk0cnBi8Lb+dRtp95JUshwF27Yxyq/34zGplr4k2/3c
G6LG5LrQGgU1X8pXqQJqwBP+nEruBetbGDOBQ8lQOdXDkEWurySRVyB74WFki3VmSXTCdlEcgSa6
HMEKyYckRvenfOsPRT5wDnvhRjPqRGFkWzYfDKpuK6feQNLLp7CiO7kU9biGdf5dhGJ6rruoRS3R
3DeJcoWBliqSn/Mq4F89OrNZo8o23h+xH53v7fI8lFnV+cHiIWv3BwTYczBF5lvw+/rF7gK6dlXR
8o+V1kqoRv+TaYDLsTtXmkWmJRz/t/101mPeScG/ZFLzQDkOTbZZO3rpc4GIfPBVYRlXplPjyzYl
q1KNQlZwsEpweMbJXe0NDsAHvCenowTo2BE8aHgctQR+PI5VaKfL6BRlhSdbGWkPjk+kGUQ0q6zH
AiFVOTfhEhKkIdy5aCXG8E4a4XtG+CHpk1vqvKcp/COc5JVRMaQXpXHhf340iTPljeY6grbPS2V6
2tHHvADMve+Ud0fy8mZlajEa5X7dyB//NeU9+wtS/Eje4FIRuBjAVgaoFYXRLbWqvNHFLuT5/Gfn
S3nu9rdYp4sBJ3+Tdjf2EJE8f110HpKLmgOyrn1wQ7ivLbMMpHHXH4SJtuEGWKa3pCQHfs2eKutr
fSLOMkAr5WvI9olUaVxQNIDZ950jgMI1q++M53Wvn8XkBSXEg0X3j8OaqcqqYWrv7OcI46+8UVFY
96NXpJ/MaAIF4KlRfZKKtNYxLeYJV66nI9waPn5mqxKuGAw01HT9UbVXzCmZPgp5SvXbi1BzeOs9
jOxCiTt6MPw+BVkQy7WXSDMvvDe/BgqIt1dpTDx0dFXFFpxsdWC6oTHGcxI/FJ+eRQE66apnG5f9
b9k+gdIP5zbjhJOt8aaim+7ayfSVFALsnAAUS1O/9gramiexeMo9fz+iPPiAA+GNqSxA6U0Bb4Q/
qmjgydNqdDUYxTDJGhwRIF2SXelB5VzYrpRGiai3N1A0fVE9KwcuKVBOEgiADnkXA+89k4uOVeKH
Ss/Y9Jd+fYIWGtLVU4riqmemsbhR1SLHTMko0savSemf0WergGI2iQsTTJW9qMBnZEAYRiLzmX0K
CPSS4EVo2qIdE5KXhWI/AAr+jcTnvhFCqONb7FMfT2Pvu9TqfKF0xGbJA+6RxEC9XJsOBkEenkXC
jljRSYd3hXVs/7s/a/wd3hGPgdWXX+JWCeebk8iFUrSxk/7Q+1bSO9EcSnzAWxP59gHLbIukhrSn
aehl/Qr8e26mWMjhhLbtn5+zQggdQrV2oanbiKwEqcKeBTDgOfa2qsvXalFx4mAMHd1Bo7VaGDK8
vOrSJNgEgJ/8TPtcU9qzZzBpkGvvRGxPqVi2RrGTTMNVUO/6BGG/+//Do9roGpAxD1T/N1MngzKD
euHy8OW0l6p78XERL2J4KoU605jDNCPONEHDr9Q+nE+n0bsaZa0tlZMiPR6WUbn383OO3AGw6e7x
2dpQlp52wWKab0AaJzjsK6OI6x6eNeEZXfYZknd/VZiPICs05U6e8859CFhfJ1idRBlqezb/+q3G
U+/JNDSJntJ2Vpn0DZNZq/PcH2/s+z4zW7VVE+6aBeeJGlI1sEBzFU+mxAR2ZZklzcNMR64tBI0f
JbPN6F8/a4V3jArZsAzhKhmkmZ+Fc7n2c633PGvLKiqErHmdIusYSeTpjyeyMr6ExGJseFyp79P9
/a5DpRu4MZRjuGQbE3Z9sFMY1CfgvHMPNuApShSlVLlE10NI+8vr/tl3oBDfcixkY4gAWimeH389
IJ7PrBKoYI7PHq8McUj4grwJQ4mwr9afIIf3MbtCwCrH8JVgvTuBU0KZ5lHbvEO+gbNn/NIuKPMZ
jgFaovfmXZdnTtuPNUc52/sJ9kSWfxW9kJoqh2aRwxHptzak9yXq3XqdaopLeFYYVOJQOWFHv4dI
n/X6YFkpUEMr7LoytWLmD3hAa/Jsq+JzavLrYe7Su1NiCw2Sak/jnym8wIgJgUHrA576J4nsmD6Q
mPlFgan2SnDw0yU8oeGXOmCvczgJGqB8Iyk5IXOHM4ex3qYJzdE06t91b+hnAfRzGz9eh6594jNK
ovIPC0onRitEzs0eRMCnJX0MuwYjcU77GMmTKSSLI5ITFJuB3sHMNqyAMEUntz0oVu97sxpueYqx
pA39e0bMbG14RdlhmQL0DSHT+K50X0Y+H2S+dsFsYXUTTf5hPTZdTwcKlsn1zkJjKkk3Dz69xfEo
hCriC62rNoJEfR3w9wQ6O/tJNhaOgsIxfZTD51iQ5uleg4dCWgs8s4Gmi2Txc7O3jToyUvs66AuT
qOmGiAbvuKC951y/miS3xzq+NOMbHFk84IHmhxrR4Wn7SDC1nSCnCDW5wunhIT0eQnuNUda7HU2C
urqAQ8/tj5tN5KZGGQDy2dG8BY620kPJdcQkGlKM5bDcc0qpr2yYFD7CEeQKDQak7dRzQ9QsGlnZ
iZCwFjaBy+tHCRtCzOpdDYqtw3GyhUspWyINfuRT1/salVvvBu7Z/sGfPiD/XLVKb46tfd+kilXA
RIhSaRX1wAFP+F+1i7CW/lHYmEW7guCN5XG7S+8QzajieTjnieoE+SVVV6noWNP+HcAKXjAL0p+E
buO/ZUb0GnLahkgKLrQKLaKfJ0wrvokFoCtYF6HSCesbveVh4zXfsCH1KR4Fn/80kuGZigUfXjbU
8imsOahyK0K0CIIognoC2uuxVDmqeplja9jA55Wah0zIu0rQ9fXBOQJVxAeHoYxn6thl0Uxa5dib
R0ZFJ0kEQEf9vNMZOXYGQ/xsBPNcldZx98IsrMCuEq+jgnzQCbrCgV0Ox5+oJdNmNUOF4LlwpqCH
hPAnZD9/PYgSZ3HP54suJv0lOVPZap2+7DkeqqO0RxCSeORfvU/wuhzu7l8zEQ9zaYMw7bkiFl+Q
28Y2bWCLVpJHkp+HHxyzGr8N1bWzW8Z3L0hHf804JcbeRgwhvLyb4mavGFaZ/JHjcVzCmRzRfehS
ZNWD/khM3HX82enj9n2M5sXl8yPyooQYzol0icqTqLlVHoJvMZK8+MkaHWkeBkbctfLs4dw+L7HU
THnB2vK8NmcMfyrdWKrFNM+dXpqpsbrVVWYtl4MFcvo1arUSt3xicwjn06IMGaEiEWQwDQcbLHIm
NyVjxUIx/GWIDwdQJs20QVuuTQqrGD7vQR/JW8IMdopALywPdCKL2n+at78bxi0Zr15l7THnONFD
bgkp9GYVB8nE3IpZYdJwOgT1My17T4rhiKJ6oj6XnT41f+uaVWCDvPWMYXEzTZ72g7JsUmahjzLs
4P1KdxMo8rYmyei+C0NsrJ6Elz2wJ6YKmxSr7/5+9JY2VCIecrULfmzwx65XI5ZG23jjMa6bcZeH
RkPsIkicDwi85NLWDJH9jIdVihgFc8ac7rBhPojTiCsJXACy1Te7e5pADxoZvE3zCI255tjalRcp
yCrRwu5JLw2cmCz3mivx4XAh7fePQoeOPb7aNIaWa3465zWe2Tm45LS+ukCl1HwbY6cmw05TqrEF
2ZRdK1L9ONEdRmGxvV3WrIdPQGfvUw48wRjV7y9uuKcE9T63fKCMFn4EFy3j7jz9E3UztIhJllsf
iQsf5Tr2RDjmfUeuR2I31CxcifbY0zSCflY9xA4R2gLio6mVGH2BegtMkGmnG1XhIif/jVTtuM99
3eT25QVWtCyhlSE+QCSfSrhQuQvSAYMSqTk51YnIbszRnDssHdhJrcz4wVJT+vvI+L3tZu1P+ee2
4eoGDXPxyYlsJ6Uy0ce6nf2tPthPXNzJBZ/sJ/hsZs+djH1hlNkAFZxDTsqmqXShnPiyIyY0+zuU
LVBQOUNA91Y/34srssvqqHHY34cHXwDIpV+c/xs+xIdXhxdGkH6I2/3Il8gq64iUsfPHwitwdXIo
sNHO/1i8LJDEGQcji5Zel8WkBoFluQBUfqq8np+Ga1NioNFYdLvYB/ByUEO/XanPuKSnQFAPeeYj
D/+clslDYB7EtMsTOuM0GrmzMf1kOs1wwrii0lZtURObkATQQ2FFwZWKVTP2VGhxvqW8fpShYOyj
eZWuGjn3GuEJrRjH5k35tjzk+CZsJBx7dnBljGdNbCBgqBvy6Wfbwrzru+VhFpOkUh3WO8rT72YM
bUdsIwHCfH5ByA2SilJvpLE68b662kfq1HMR1MT2t6VSgOpYwEh+BpFoAzDmxY7IXvU+0qBhR5+J
jZsvIKw5rIGBteHcelE6lKrIXYPVHMoXkGfi2ZKTeun86nDiPdZ+VZrdNZosTKWuBx22c/JJPLsg
TQKCZMGFIzWAE/TuWxgKtMTor4zfCauQMunHLKppAdI9EHUf2qQp364DQpgKtJB1zQUfclQlmcT8
BcBqOSJzSbwiyQs1XEn/qpw7BnEKf98+RctQhS+HfZqxLE/TUVu/CGUdKWlXgQKdNoYwNfcyRkYI
7t+DPeYD9HIWQFS7fxz8cRRuJbXClteYQGfg49bHm/52KVAgEtHbZ6nWd6UlvVBYg7ec7k/3TLZv
btNP5eVHyGp7uXpJQQNO93hF81Zuoe2Ln3MQul5kNmJql08EDDF0X+xtBtwuWQzQzIEvdiT2kSbV
Ghre7B6yiZ/DtDe+YsM8hm5WLfgvTEI0dRgUFJB/pJf0Ll4vZ0nSy0UsYZc1iv+2ZZak5JA6IhDp
dxXZpjI12thENNreVnT3O5A0I7xBegAUR3yubJn/PVJ/yLB6lu9ISNYpkahOu5HRs7q/g1An3ds8
Qb0zXiaO6rslpwKADUS2vxFSqqiJUbJe9mUxSaklqFIqK53l9n7kYz8ODPu3q1XDJmqGAfeWAgx+
vy5ZGRwnsuy9svati633XFZaNKgU2F5AZ+GhVDfz6KmCUa988zMvsV25i9FhG0Rh0HauWEi+coAL
OnAqvgHnKd1PCG4BFHdiYqDVe9LfzJ8HMaoC+gkgkenVS7m7s6eCRayVMo0rNqdDWlcznnTfsfTL
X38MMLyhjMGsOteQYcm4/Bk1lfmlJTarP9zFKV/vJmK+gZ7v08K7lKHKKa3D00vphp1yeoC3K5dA
FjM+a+pus/SzQfYZzj0hU/49YzGG8HUDoPcHbX6rExUkg7L85OpykBnDYcv1WFk5op2E2xwN3m6g
lt2HrJJWseove3vnGeDkAGmg2uDmVeqsHSDyAZBBvKMh3MDI3NPyoVAozf2r0nfe6ooyKn42FaNj
CUN6XPydLdI4qhKqwrBrmGhntrIh2za34jd2wyJtKaTLrRcCwVthajI+u0UFqSf36u4UCBDyIc4/
axX4N8s1fDxnMaljn/r2LtvSQlOk27oeYZ2jfU5dpEIZoPMQmHpgKf1X/ftbv80Cyg3zxIr/ZTg2
013KiWLD6KAMnRFBh0PF1/WZekHjYhZxvMv4ygWrz/IY9ExVURE4+Pln1sncNoI9MIJTI/5+YKuf
ldC7zmFeZ0rM9hZqc0ck1CL61WS4T2H+jx2Fvk0MkhPqIQNnnX0v6Ms1a7v5R0tcSwXIwuCOmt+Q
MbKD0aODBe47OCcjlH1VRklCUIcf9x8jfGSgte2u+qu8OEURBubHR+94SMiP6xBg4n1rGEjwT4ez
NHx4bkAQjF+rcH6REJOmWBkWB/hkDWQsZAMy6CHcyOUHvqIYJ24+Upxt2hbwORKGRjd4HTmv2Mpw
pxts6+PBtkAq+rhoCo6W87SshsJHdjExU5Z/Q9DtJ0GTTJLDlBbm0qcvbbMxhE+I84Yikfx/8w//
gzrs4/f20ydLqE3URJG02pl6Q3oIXpfuxLetRrJOScJYJ2wv7qfWkyWYXJFEhO3HT95x0gSksle5
0j8iE5v5slsBx06GWjS0ZVcvQGp8dfWIGD5Nq/x+JEDga5KQoOqZ2QGXZpia8gxChSdrf6yRIacz
7fK6g02IFV8QquZknVkriClzdYXILNkBijCnslzlvOfn/ytHlOy9/ntr/n8ygSWLSQyrnhLvZk00
SaV12K6FCsugxplQYUsYyx4brjRaFWG3JvKeqlA1WNgTz3BmIM3NeY+OT9rsla2bITJGA45jxETU
OVm9D2vv7QcoMfMTvpbgds/WGn4APnFMpqZ0u7zsUqiiwhlgfAbbmLIRwPL1H+TMKUSOcAkwgBLl
2W2m1wzAW7sGBi4pi+igVmuhcMLZuPpuEnJt1T76J0MaUoEhHWgPOOF3M99RdoJ1YMh3Ahg66fjc
NNOKQNjKLX9kyhOfB8ZLFLAK8TsR7rMhPMx7gYiV+eWIJqL+Qe1szHkEmO0x5Zgj7I8DdT8QccC1
Fq+M03Zja+StAYugmB/XpsBzFHzmpJ+MaR4kIz5TRT+rmmJUL+5W5DnBJeKruIDulKfeyp0IFx6Q
fh51++xvCQ7WrgpFByHc11HfEZmV+du4g5353V5iQQE+S4wZO+2nI0zBZ/3WtKCXrJdJ4+YnT2pR
9p2Qc3q1qEr305L6yQfDpyPcJrNHxn1wnNCEt2w2e/Xmyqs+RrH/QfVXP313hi2MPaKXGPK48WuW
Y9VTf6uej+mAP9uj2Q3YnN9lo4RXWIY0u6xmAzOlaXNWtuYRTDK54NjGxADWFpUl1Cw3mBj2N01P
a/I1I/m0XOvVwTrKkWJz8L3rvcSMcI/eLzQOGBJh7hwY+hm7j6jiAjGtJOXxPWpn2C06d4Gr0Y6F
bPOgMfg/HZVsWmYjcMr6XKL+VyzGvzoSCSlXhv1miujpTOfQiz7Vzl5qXn1zqVVUhePcCNWBx+HY
UhJexGqvcIHMhzZxoOgw8G2DEqH/ZNL3iMvjGSz8+GOyMr5gbFuwuOWFPsin83TEe7WAfMg1RdRG
bvJlO/Re1MP4cZp5TL14OyxD5DeQWzgvo1marWeqzCJvzwrur3jPyJWYXLFGP9Ijt8+rNDiRFhW7
Et+jpBnygckprtt9EqtQJdn5sJSvBDZ3u4wChJ5Cw2iMJx3GWGGUwTEr5kyalwJhATHfXNQAMjcN
CwLD5ds7mlY1KwbWBLsozvm6I73MaSe3QFKf5PziT58b9McqD3W7YmHHuve6u1k3mZKdt0kg1C3R
suEWUlA6yWGsRwevFfI8Gr9v6FoiwRvKTlFhUj5oyAfq+nT2DQgVtWpFRnXzqL1/lWamJBiKUau6
3e4nCYkTnkmOHXZWReqV6vK5A4vkyYzfS7qzZGhebALvA/Wze0eUowrT6A/44c/gkExmPTrFMjjF
WHJNtp7Uy/Djqfz31s3qSCGzLGlfKUqrekwk32S7D3OqBgzgdRYEYv4UxHBu+kJPrf0XtnNVLn5v
TCBOhHdbFpYURq9NkVUBBld3Jh2xi/g+UMwhqKdoiD3Juq61aWkgmbHgI91vmZKgNyirr9J6kNBl
ajKKVoxi0uTAg2QxiUzhJcBO9kWU+nHCwZm0xgshkJiJf2ZmyQ+ltoIdQfwvy/6Zpy6k0lLseVZZ
IJhU3zO35zK+aUDMExXFc9DEc8uSN3XJHwgURxcm7ZSG/nIZoSCP4H0YOT9O8m5PhiV7WxstMKlE
N5mz5j+a3JbSA9jGjG3mvYsMt6H1Dsx8SOSAKvZB1rrd5ZkHYoyfx/Ft4ndbLpzOqBBmAhMMEINr
7joN4c+iaAiQ2CYV/4EP1+QiMCxEiNyfpZlgsoXigot4PzfLrbLt854x09beApCLF5G/vDLumg0/
Xnxs1l/ghV/g84p465WHIVKn1t5/4V61i9JfTxRGm22IHFiuIuR3WIA7zvV1z7jdapXyQEim2SOP
i6Q+hQ0wx6y4hbJxuOgBYEA2EfL3IZ9fllkfcSVh50k9tbioB0vYces0vbM8EQVW009GdZKfbFfj
fntHEp7yA6kacd9VNmE0E3OJ8EuF9tYu2M6lc1yXkR9CbW23xnMWxI5YQBQLy4qoMkvjoAgMZfd3
gaRgNzfAm/iQjQ23gS2WkmpLfinUa2IdH1C52+gBjK36eerZqYwJx96e1XKMrYrKwIVzDssSZxwB
5gszDyfjQKjrMdB9Lui2TGt3VNIjJDZoCiOL+HcyJ25hBA0MkFJasKTwacmxe6E4NqXCSH6sNEQs
Uf6BFVQbpQH0uZW9zJAYs3EL/Qas7QfO+wSnaaFZNIBDsoGM7VAgrEZuxcjBu1tko4y4MtW9yljr
+IPl/nbJpSozTf55fEgFcdVNbunok7H/q7oikffEhhe0B+Kqm0JNxNdBmtPKdViyxpgehhy12BO9
0V7Onm3YIP9BypQAjQ215sRalggbjJmrlVshg7PEYng7W3JjJVLAB+6cGlH1I8lgY56Z/3NMlirQ
VysyxOTGfjRL/9JwGJsLhR7Kg89I6/vjiow990L/vBqKl9hPmUO1HV28WAaGVsqxGFf6ws3gEfEQ
Rdw6SCHIEkVlkQyNNMNbzq/GnuIGSI7tt4OUihBLhwWCvcXU1y3mLh7+zrH8u2cTCbOUjVmXkaFl
bc6Cg9ANcxIfHN44PEmtTI+UKPoUtbLWvdqbFtcMo3nAThSQ36YknUsFcnq9LtxIeUzfeouTH/7q
mdjW4hGoaHstLJONI4wtjUba9WEpZiADFGnRl0KsuJ0Ec7EFiZzGBVFMj56jxLO8gTQ4S/GHVRBE
QtIvhaSLgVU13a0WkFLACrResM2xOZQ9uOk44/CHcesDXQNX/lJiFRTHk5K41rXtAM2DkZ7y+AiI
FuMJifwpU97OFjk/cubH67GMf9yl8YYuBu3Y7ZqVvLrvKO7p+pTQTYNmT6Op8wCUP+xm17GaMP4A
G2TDpFfI+SwH8VDPgFEVMx6DPKJXsNsh4CKjBK5dsRYUUQ0WMujE/TdBZPWRsBOU0SYO77DTIkBQ
yaRbEHdVTDw6lbJhBJAqqTk9kBIUJkjq5cWeRILWZfYR1pL7Bv58vixqblquBBhxQd+utzJKPC1Z
SbYvGN7mwcwaO9jZnYB4VlJGd9ZDQwKQ5/J7pB+/gCmFduLA8ezl1aamlmbFIpMyPqBPNHKDgsbB
VVYF5uuacaCBHg3Muu7xrXzdiUMYkJJH87XrppOsiS1zWzMs941bBis/Es+k7HhasHcNOMVKFULG
U9b1J2+ybBkCcOFEui57tnGxmsp+BI7trhyIl4Qbm0DWtxyZalIeKurUHBPvkNNa/qBnp91Qe/vU
mkgmzTee6DufRn3wvLKSIrDkgBLO1iKHk/qO7efV0xs/1NL6ORhtr35blu4G4eWV2oUMsUPYi7Eg
EUbJADZN0AmOMans6Q9WecB42rcLuBB6xtJT/OYeceizkWE6pLgaoZFDUcYz7D7eSHiK9MWnI7xK
jG+L/XGHZyvIt87xqW7DeOnTol0V0mekzVW3pdx2p3KbFY5EG/ylIZDuFWGfyqEGLNGxBLNOgDXv
9uEHDHiVil8Gtx8HaGXX1vPp4HTFQNpW+VyvtS/MVKG0+EjdiVpcaf9H9CFqftnSMQj6BFTVpExV
RjQEAu9NhzWnzbRsD0Px3p0pg9Er+nkZ8yDQ+NgA0hFU54SKiZf9/L+W4dOi/m1NUdaa2ZAEk3Bu
x5/Ilau7dQNb1B0BYuwXhcRo1+bO4jf/FSbKHTeCdlMfU0nhpPTL50j6pMc9M7FS0sbPs7NKwB6V
1BRY2GmgzBPsowziIRKbfknG/xvk17D8WBIqm+JbZvxHYe+afKIcQgpueu5sGaa6GS+nuajYsQJ5
gJ/Wh8xYZ+otSBj/PiWxe1TgWcXhW6cqrdJDjSWvJ8kJuRZwuvkOjOTLN5cx4BQ+M5FIslz0o1sw
XkkVMp96HcUxsE9wdSxTtrryr9VaQmK5i/dsVmnVPDwxMZRuJJ9Y314vP2A+28B0Rt4sMBYQzPws
plrGEexRMtfw584yRW0K1p0Hs5sOamKanLkd/6i0vPCvF0UNgFqo2HprPw9x5h9EHQCHl6YFaYB3
u8rimg41f+xWMuGjLzxTzscBdWb0aCEG8XlmGeFTnwO5xaDEhzBsddNpEq6/6qhGDu/mP1ALtgbZ
JNVcKWX9n1n7Pmt6kXfYP60D7tYoW98brfyQpWqkGwvpXve0Q9RJVXMLAioTBJFiQNzwZDtNTfF0
tAw/SNrBLOhTAryZXVD15WxTfBCyMTjGHigaywODPD7m4IwADcq575+QTInfPH8S8/AAo3rxgjuU
pHQuNQEuJ4m1DxRdv4vzkhWyRZboBgkruQ6lfovCk4pfnPYC+5pZnL5/f6+32Zqo4AauR0GoJ8Za
8VuhFu2q+KuXuQ/w09CKC6noL4UyXeff6Yv6j1YdOFWV6YZcoQEMxRkffvLwI5dHLBIwxxMaKsyg
+4m2Mdorh8IOiiYs1jHoCZ4qNBnF9n/jY7CZbhKMwnJwa/NwV0RY1ete2Kxb97r7Yp7bYZVW7mDW
d/WMWneOxAQzETUyjA10fWRe0/u0lboYSo7Tm7LvhgL8Epbq+c0LKJnH8LRlV+Po/SmA6igngzyN
xSZr9ynPzJHyS57ogCnosxgE3T3cRlgddRIwURvTnyjWRJT/HeLfec5BUiW/rYvlmWXu4nCkDrQU
FWw0p46FR5xdpl8OUD3EeVuzVbiL489NdRtu6iUid/qRxyvDt892F0CYbB3IXsywHhRCil6vDTTv
SfhD42IfWxuOfpNBFRp5z9LwERumPPuW4kprqoiKBevpc5KXusVyiYz9D5/gZ2wq/aXHCa01sWTv
kMa2QCxrTeUmkggX2gROljWXI1Zhq99tj0L6PNFW2oG9JgJWidu7opux1oNydWsejzDPkbFUsgeC
XJxLnDP4d6HvQFUK/pNwIJHAYevGuEdmIoCwJ8ROBQtznnbCsJn2p13XS9psD/xRj3NzBQRA3afb
kDf3CmgVQwECDybdlKvfU55rFeqYHtBd0AAvB2VJ9G3LbOPnozNF1yPgdVxvXaKuFdbOjDLNHTrf
4JYu7loYbPtI+FoSj6y6NgQ7B2f1CB2HgTVp55WL4hhEA7uz3TsDhylaUOjWves+AFsTIbgdS9Ze
3iQc+FLxqSWnpIzE1DVMqrmygSLfdCH8hUZOK/rQK8zaYwd5W+zfHBvC03sTOwnl1hLpFUzB14hL
JnEVwNWTm17UR78i4kP9KYPXDQ36vjs+TUhtklnVqdVH/AZZw/BlEOusFGomXQZrKXs06SXnIU/d
EL2Q/H/hVNhXr+gJMuUsNwydU9XcQJs50br2z1cLlKZMXiN0UEym1lafJBlJw9It7lqBee/ScIt/
hRJ4F9M+L7RTUJ5/iM7QePpbaMBPQ9fhRQodJNpdFSPH+nsOPOyLQHhOJtJA95BKN8fMb47JZ/Pr
NIuIe59hBjsx75gpH5qX72cBsPvf/u0OmCB/byY+ncA+vNIhh1mXQn07TSGTZD0YFx3SYCnbK5tj
Cf+qmh6hDuY09uxPSfqPRarqJj1XC39V1TS0qzAq0M3BZLQytXh5A8Plo9cAU28YH6FfVRDhem7F
fsp2cuxady7p4lssMe5mWrMlLBsun5pbbgCTE+g83JuC3hAyVDIq0A6Y/CldPd0TAu7CVQgdpICC
n2TnvYfpMlcwgQDfavN1BFiTAn8SI7Vwc0/Y21LbyETQIHRJ1qELAPcKLI51dwxd2OfsDVpQ464I
GpceMKIBWpHb6bBFfvsjo+R2bpR65icKw4hbHU0MJ8NNv9yXFSczSunUQNJwTkOpNoeHjh6kNP96
hNiLeljTtDKXWawEZM64yTHBpjHobcPNLyLVs8h1RrFGJYMVdjcc0pcVvwHu81MfA7Xzs9xD7XQb
ScYu0tCbpI+PoQIpOcUM+apoTxS/NFVnmhlX1C3PLEqaiMY0iQ7GnAuO1b5GRF6fw+Rr1zu6QfqR
r3E8gEsLzjtfWUj9H1BwuvJsDDYaKlcrsmT2n75WgHCL9ztLM62yh6klDshwd+xUxr5nj855xvPF
1L5a61/LcfVeSjlbwwpwBh4l33sDz1G/7gzg7AojvrFfS7DrKFa1bNuE29SdHvqGfEYu2YJ0Opq6
bWkGlR5SQ+UueUA0YsNUEtdC6+Mn4yt0dEtHsqWR77iDP+X5AWu8iNK2YCcoXm8OIvBPQkJShWo3
LM/IDcihgXElKxpmv+1FZW1nmWHZobasZl/BWEEpjLINhI9s+sRoPlJ+Hi/JRohsN1tCkXVC1CcR
GvRD55n9JwSI3kRHld75xEVmYObdhF7B0lmVvcvKL8peaf9uCQnKu7OKGHyHLWkxOo6MZBn9YA3E
gvQPCmUyG/JNp0JywcAF7qXzWnZrzDlGcy7x85T/Ajqz2c8O+apjZxAMqssa0bbAXyu23aSCBVDg
9GmzakGhrgITPRM2mBbmGfCRLCdtqPNp3MKXPkc0ZnQBEAtmPJTrq2XEE+tLvPIDxXAJztvvGxpv
pghh/F6DWi0Kor0q4MOWTnuxDjH4AyIApqESygUdOdKwirHgNJbCc9C7ZUIlLVtG+U2k5oI7uspT
YGKB7mDOl9jAj7YdZTFP7QtG+T3ujBGGjY0kjXVPgaHbIbVL8as9Apr4Yjlc7hcVuymcFDjsSIl8
1VJJSVpDzDY3jdZE1VLUDqWQ9L37bj6Z/xsjMui93p0ww7vp62nWZpuAtrKbCh5NHM0ET9zsD2Jq
iouamxwLIgFtBB043IPS5OY6FmCPOxmSwr7F+VyneK/voh78ucog8zQvawavx1v25QU96jugPLjO
QJNwvxKFPxzunEZPYtuOXTz7wqw6acO9C6zrr7801VqegymWEWQ3Lg2mrd4b+VHMcMYNwJMyKpUo
JoFfLNo5GWhUcdC8j3V8MD27WITeYxDrtKgQsthzbohqY52pcdn7gIOBau/K+O6AqwOOaPKhRnCC
Fy5VzxtklZkDTyONejTKHiQvwamUQ50tJd9SjwJEjug+Hej20S1azxmXPRhuLw/AAJDxjImRUGAb
H31IYCkBii3jIayvPUF+NHcsXuKpWL3X6M2klEt2q/Kz7r5QwRePsIyiAQTXhsDwkz73IYuAnyCP
0D4T2Rl1T8hLz+l+Lo3YGfXMNfZq91Jg2hgBO4sdMvoJxLug82Np7bVnZUJw6oH0SeC9VBqUH/md
TX46CRqSipQohvKJTZYf82fsjtrcjG61sfx4yko/gsbY7/skuRLWxe4tMEerAwwHHDwuK57cMvCH
L+l0eBNbsM51uCSErNPkxDJD9CIvNNyVQa3Cmf8xwxXvBHlih7MeCEkyzeiYM87tl8/eRHxVbtYy
yzE0hDd64DrOo1LI0dvr0TSGjW8chGThhxFp6zBKm5xAGQUk/7kOvMy+hnJA/Pw8Tz6evW8V+L30
d0VoK6L2dulxRRcY7uOjF7vJe/MraaPVbvcR/4WrQsxVgFMHkvp6r5PePdX0t1g4tLrI0yXHypDN
DhUCSdm0BbW0ESEZJpWqu9y2hQCxwHiA4bpnXik0TqsRjbYDkIdnT7+Y86kdydZHLFhD21LftIi6
kDfhlCbVPspvUC8zlg6AiZXAzaJcAgMArcNtuHDUV1Vp4mgHFh4nxdxJAREJEUcgdTlZ6IGFi36J
IatPUd05SoE7xd6XeDnbQrUetDKClTTnhnU/d4zGzxN5CXzNlAn0ydreht3qGfz6oTHacYZNGyJC
TFdrUbf6ykiIUk48MpnK+1grTv00SEw3PF8lbcbMf4AuPv16g8V3wI/OXtY+nIGmr3ZgmzwfQru3
AmtlFVvmLU9DW08IAWdDcWMyEH+vYTUL6tQar9Z+m/Hcg2wa+jgPT/xQPEOiGkX6L+IbR4DaMLuC
7W74qblGq1k4xto5If4UuH07OHx3mFhWjSQ9cGRXSGQO0F6G93R/sCES8jffBBqdADz+edkiEA5N
ecsOUt4VA5dL22Bv2exCyuE3eF4Ib2cpebPr+7CErqHghac6FV+JJHDLhygbYAkvPxPG1r+aAWEq
vCb27TPXfojyIWCjiHsuDA2vnISPthC1G41tWHcFdKsQuo34OWBCgzr15riDDNhCUvVzKTw+aMRY
rxO6uSTCkv44hO89XKt5FmgluGayF/eBP0Uw1TM9SOiesr7dHnizNC2tTQ5IZd1PM/xvR59vWStc
weNXInKT+uqCtQoyMAYYpwo1chTrrOwfCSATB7G7fVOk1RG0UfW9Dwb1cGyoGMbNc/gOCeSnFAxv
Y7RmPoEUee5FmRhdfgPvd1kEtB7k+liL9KAEDET8qvSkp5XyZ1zhLXBWnKK1TUrrrx9zVnN2CASY
KX+0BOlv+s9eoA7xdfTXV18Qmd9QocnWYOJRsiiyJoVw73HA2etwatzBDCeLRFusfgSt9O0+eU29
gNz2n5a4iAtOK8JlbFlRzgDvNyz25oWd4vdrg4pdJlmj5uxCHx5sgEpQczQuCzdIMp46SUVcOqA0
0sQh3sxTwLY8pLJhCFZrynEoQapvsY/7d12zRQ9cejKXaqe3JAOCabHeMhNG5GEgRiQW6howPpmR
GZ9dJElBsqbzsBQmOItUC/4y26JVdNi+PF5nvBOCAtsjiq9FkA9n769M0jgQQoz68O+agl7qja+Y
AHxiIXRrT2rr9q+CGCpzQxBBHZJiuw5jPH7bUkou1ea6mRZEJs9earn+52HrXQ/WolKOXxXe3+2k
XVQo/mo1Twxu3+0fNe7g0nqh6+qZ2B5isq7S1gORYs3jHt3mVwPobi+/PDSPCO5CEqWTLD/soc8M
oSrVqLq4GQDP8wQKFjF5bp4RQ9b1iSxtC9NqORjqJSWQD0APMzvpjyfVFZYXCjZlciqXsDrpnXx5
RvWc7M1efD3NqOmOanfGpZdfmjrSRTOiqDiT3atLvPe6MKLhy1MW79POpjMQUHlTDz/oWt/XJNI5
F/6f4lQ7qnPaXx3S7iMmsoB5VZ0ZAqkQed9BAgiDWIVT8RKx9kLj9oQ6vYMvZJzjCZ1U5CmFTgzH
WNLbjeUJo5EM3tQeTvpVkri4j/6XCsDsUG4sJKexSzLYxgCH+lSaNe6ghQehTEFKp2cHggcrVgiD
51CMkSM1dXjWW6wrS8V44SDvYQLrYFPn+phAM9kdY3LjgAQ2GF9VdAhSe8JEcbkS0W9HJK/Slk2H
XiXznDx7W0R5EuIcB0qNy2JOfrqSjn1zYBuOe4eF0Z46mM6Xg+voYrq7EdokFN/00urKmY+W1XSX
e0C0MTVCKACYzltxWmdTivxVwxF6QnxNawazvN96SsMFSvwzlGIGPRrLtksm/QJlU/wdGt5p912o
YG90mSa0YGWviuJ99/aZIEVjx36pIAzTdWUUBE5EISOBWJ7487Puaz5QjH500vdXi7WE8htW+HuF
fjTcx0wYtmAVelsDx0CzZRpCsVc2xsEs9henXaV4I/Zclp7CF10BHjLhZS+gYuHWblxktyiwWB/m
M4IdPm1+wFNXSwmXch/G6yimdNCHmeoxLBm0tqlZxGxp1cpquV8QNQJOqOmYpKZhnadygpsne9ry
PDLzzZeQwIFbnwCLBxihXHB0bQ4KzjUrV7o8/9lDSrFtWhmB3YwbZF3deaF3cmSK6IXf91xpibFv
NEStvHg4X/RnSalTthep57WDDEKXJk6S32porEp0JXHnPb4TnGFYocCUtnsooDx7SOWb1sZLKNDH
ZuSkJiq6ZwQGkttxgL7Mq8qtDaYdZLHHyyMdVIxhG1mPgLADWuubqGWeiEadUOym2MjeZ+Vz/24a
CK750cU1AHsxQRQABqap07Pz7UUUvoah6bvkN1cQP7yIxzg5/VqXF+4u7EHrzT4pYenno0y2akl4
5WB6ZcQ0AZXA475CTlG3KZ6irD+IxBz/yhd0EmY/J6rJCjI/cNPrB6DJCcsUUc28l3bsYhSJn/tp
wIhjWFf8y4iSCak+mJ7DjHXQIfNzUu547Mwdc5ljzKPXG9PeVCC9hYFipUpXNMRt1sBwyEsbh6lC
5O7+JNyyPww1mNn/uJjadDL7YVAvlfEHUeByG4cSNvOIezGznXReWoBO1SqSli++WO6wmcdRcz6P
7hDsFhPcqbEl5kzwOG1YWeoeTlHWj1q7PJJA3iOQ+6fHaKOFoBAet0/UMu4b5UjUyM09OCRdV5vi
MB52DlK+BJoWUxIxaBdl+o8+ODGLyw2SfUl+vdPljgzpJfS+6tqSC7AmrXhxQbmne7Udb/TSIPEv
rHBt0fbZ/7EPUHno3umiur4lPkJUmjCKnwh2qE9pczONhnzbPG1BDAaKKkWUXqN/FEAW3HLnPFcX
26VoBvyScP3E7ZD5auVRvSuEN0dd84A6BQWpW4WFiCegXbCgDN3mdnG6O82duj8aiLrH3NIr6UsP
lr+2AnkMcENBnc1ehUr/JxnKIDEUDetu3EyFFweBcn1u8L3JPBk9k/S1jxNALH1gpQs4lzyIkxZl
9QOjeauVJB7x8nqfVcUHh3ttxW1abQVnMkZhJXZRvDH34O6zykxteCAOVZeBJQ2eYr6buV/2Koo7
klWBvEUPl2LBzliSJ6diURnseAxTDzLlJWkIAUkMOaG9BnHq4RhKZSgIcy+XqBUBiwjbZ6wyn+Na
Q2ChhG66A9i7rDCU1UiVoagDb9Xp5zzeqH5vgm2jpRIfVM6IANMxZ8hf0x+jCuL2LL5KoOin3nCr
UxxoFjlOVhYHsRf1kg4q7nKChXPjhatppf6QqRYIG30N09muBdgaIwzOObrPTjXAMnPt1tCx7pao
OfovtBx8Fwt8r+7Toq1AcTa5er5cu9HxS+akL6jBbrPfbOCBvpE7tqy4lIaHdHgTwukTNHSVwe8C
2DtuRcLeRr07xY3J10nEdMmatMKNhOkl94Vn4GxzPXdV1ZCAA4PLPEYIvyw5wu17/lFGU4MBPEHc
qWGwn7ZP1jgf2kWwWQ1OrxdRkQsCCsoLH+SjsXn60+xcPBAw3SpuiKkdk4aj8+NJ9C8kzZhoAv+V
nkIu7zIb00W5+/15RaHQF3GbIgxhPVgqZcX0BgLzEpcvIeV/jDD6BMKoU93I2ZidCDZ80SndBciY
T5FJZ+ofzp+/+DugMenfWggXOGaVxq1VlCrGGVjljh8JD+hskgtjlCQua7rTIxd1gBpWfk9qykFM
/P1XNarifQW2e/bNtOjQRuG2hb423aWmoyyYOHMVe3PiZeWF9yQ/gacsexy5oKlLGPejzD4g16Zh
d4TgcrrfHpbjoeIW0xYslF5GH1+Rt7IL/d6vFrg0UtcplxthRIBkxViV/Yq31r36LkQjYAilPP0L
4GkJ+T1I1Hls7zpULAPTxcKH87mehyZN7KVy3nIh8X4ylyKnSy+PrhWgVwlS5KtrSlY2H3lpJxVB
7ppeFVfLO/Kg1hwlUFpyz5ZXo08eFptZhpjdMSNfylAE7Z0ah1ZCm0L8XvF8uQv+4rRMaP5OPR3f
ooPwP0thLF17EsMf4kiyi2A4wVnrQhvw56I/dj0+4AG9oeWPcLPZNxNbfXyTak6xijTu5l9wEhe0
JF8EVUguIZeJ3lwCbbdR/akeAz9Iq3zuOK9pHkLFSRL+qYHh1NfM4LB7FZH0kBUym4u31dOHm8J0
SiISPVx7R+SFou34NboCa3j+d5QUWz6WEJLbvAn9eQL0UsQzOPbVB16hWWAkRLdffxOHkdEV9BUp
fUSnhFJcDFBTlJ3HzXwl1foTwNvVb2xJD9r62E/Wde5P1jEve0i3B8+ESsgd8mdrt8H6VYV8qh+T
ezGZOihsu9+gyTmBZjW7WFwTc9Cawz2/Mgji+pEXmudo5M+kdmeapirOPyCI4Dqj2j91D/gfVoF4
AsDQbxksnHOnIcV8KvBI6Ng3Yp4qr+HrHBCanaEtF8lipPqVuFlQnYvikdc/QhdXSpKAF7bqZyQ6
rUkzVj/lGku8xDT96IhXT6pnl79yTzjCXi8caCsrrz+1Zxrffx5u3vLkFQWwPRdTiNeNn/9OXgcu
0bDoPhvbBbfY+OFCsk+5WV6ODnvbUzkEHqhmeURFbLdY7RjGjYH+cTuJzzpzINZJzmtWpSXkxcL8
1CtQ0OyxuxEMIqv5h1mbccxVitnWB5I12H+bNnFk3fgzqdRTbF4pdEmhYjkZCqphg1dMpYkRPIyl
LvfQCMuHNFZxF646BXlrSIR7LAgGWVGvhCufE/N5IT0vVMVR96iEe0Gxv4B0Zio13jZrQTPbf68S
yKmF/GT6oUEPAMbpYeGINNfTaLDRQMMUI/CS5SxhLzfLE6bprlSf6xMFvbV6s0tJXHV7dODyuHPB
BorjlqD7uEBPepQDOPk3yCwcyYaj5ZPm2P+zKKqhG0eVYtcQupTwzDMSlXwwkXsamGMzuWU4oh6t
UHSotfiPUx9Uwhgf8g2HxDuJ8znIk93PjJUeD2iDYlHFbgu2IDCy+ydiU5t6VIi6Vz4gN5AZBvV6
6BmaZSvBW5qvxlCs7iJVwyEBfAfILWAkbph2josyBbPxPhApxyGlIiuudNQq4pDsMMGDWExsmqcM
E0OaPis3d4GugqX0+wT1uFNdzJHcEVLeCB8uqgEB5BB5lIkl/HKmC8Xm0+SJrH3XSCWuJRASCdHy
3f+NqLd/KZS20T3LwUhIfc8RaX0m3fqIXWYH99GIESuzQyDjew9FVz1SgvccyhIWUB4XiV4YTUkI
eSC9V9wOUugqfoTTwmWu3RRDl0Oc+rL7EYAmTuA/AsapEloQRY67akJ9wlES3+Ua6qra8vODfo7g
//HdLgY7Yi71ui6U3sMS1A9YqHTIrJE6P4owqoqw0ZvAP+xN417+IVHYTPun2G2cppgGQ7UlsK68
MIX8olZwuUP95HQd//QScGRzrG+dBVecjW+3dyenOyiill4pPVY2Cv6hgzStp8NB18VLJS9Dfkzt
COAA0WMBGhWsO7DZdH++bnxuCaHKbksKZAvlIN/a0lJ9942dV4wWpC6RCromfDObuTKQZE7BvkQl
W+XYQSjvvamRfY1EpABMIEInwsNvW0WXhC65hHTyC1M2Vzt7+k/REcQBE7wMvv5y59gf9f0nwzei
7g4J36ppdrFKWgkXzGKnUjTmxgcyY5PlGxQqVRVcA0bXvwEZDdp5pS/Path7RyZ8HVlAvAR0rSPZ
EZopFNmOHnuzIdoW7MzxJn50ZVmuYeGFx6G75HvzW4hw1hXy9DX67wRakMtjCPyQ4JyeiIcjaPfB
xmLCYVuBYFY95T7k/yE6F86ndaKwmPzZiq96ATz6ldrF1tjQJa6Cgx0o+jXUjooVI5/UNQXZL72Y
DA1Xi1xetr0E8nI0brWDdpO/BQjhcpTXwdjGtsjXXQGPd50P1BhbQbDWS0OaTCiB9I5FUt+K0JSM
SXWRtY5KkQiRXGEpmS57zP4daRyBpfP+JZzormCPOlVj1GXqkrgYvCF4EIc/zbjijfeLmsvKwxCo
rFnjsRfWjvY1a9NjgxHAcUi2mxFZN5Jg1LacbcHoAC2QVyxyFa2wxAvSnF3caDxISyDQi7iINSBs
cgXP2oXQHOInFM+CxYRLNKFQsoD/DO+OInz5gRW40Wouwkrek7IkkDmmyo9JUtM8qZKeAcAkqEIi
TNUcVeqCHi2kD/G9opBWXQDd7M/0cWZyhsBvPmn3pdQ121jqfvJ9WxQ373cUdcV2l2HVl/Gva5Aq
UjKLmB6S086Mp3KfDMCJmVXp4dZY6/OZb8H5RuVH5qBQTEDEWQ5pzxyeMUa2lk+cgprdjQaCoe2I
ht8RoTbNHJH6x7HZKCd2jOsNI1hfG5Km+r8H7NabddcEGBrvKpJEfTQORGGo4BpJTpJ0jNUODlpV
3ldZCfdVn0aT+sDV5+UxjDIiD3Qc2MOMmVCG6bP8w2Y2zDWazcdC0HFXpxu1L+hT8gJNXJr/ANM4
suTCphBXhJuD4jMmKjyDLgzzsNMRO3/wN6pZXb2D63XWnUmpYB4eR1Tmrb0DnsMGhAJJbnLaDcbp
kDK8Wzj5lLjALJCErapS32LGFOe7fjORwgotfzgD3e1TBzNXDtM6mvhuTo3XJMTmJ+hn2+SnUS25
cPrP8zDkCsHyyUuAxPYEM7zenq4hhvSOKbT6BwITph2U7gS10c9yP/Wqt76+0OyQowBXUw7wtf2K
vtaB+FEXxJqc94UKRIxFThdmfQLPmblprqEgYA131JtrBo0fyp4SFOaTWvmAxI6ZfNEpLCJcdTd9
6wNKL2yxyQsMPG75i/8MisexsVAXOgG8ZCCtfqg4O247QS5VHSP5Vjl5i5FOMtvqIOSJcCD0ftUd
9FHPCn/9/e/Dmv50a40M2wDt5bVonzSskJECBmkIG66ryTAZn0RM3w6YuOI/T+biJjeVKrihpqiN
jD3hNC+ISn99WBU+qz0bWJQa/NXjkmQN13attJ8Kc0MReqjyTCiVMah/87uXKawhP6MUb4Puplkl
1/hbwbEf4u1JkvJZpbKO+F4bhvLWobXPVr3lgTQsx1e56Y8crwigi2ya2T9ydhyael62t3gcuY+z
gXGBsG7wQaJBSXYybN4QDWuEohR/JyJbOZitqYiaL2mmO1mPzHcLxVlc+SEHDWPlLyrrm2vyucWx
xfkXsZ1muvQoYkTCyElmuqhsMjf9yqnrd3qy1MTplhBn6VwZC6q521HKuUf39oz9rowx0gCTU0V/
ZgyS98ozK3ss9EZHd7eAeIht8qk/RFCzRUoELtv7XxGB/G/UKUTWF8EOHeT8Bhc4TQcIT6zddjYk
pPOZ2bdTwZZ1m1YjWg1I3GhjBWizkpQOpVlH7cNRUy+jZQlnf9rC4KB6eptyKFFyOIir+Aiq0Aan
qw5VNiWZ06Rt2Z85Hm4kKpekEzRXmibv7PCJwuIggtm24KpyJECjsXWJ8D9DUxIHwHoMxxZ9aNnI
xHQMMfC7pfmaAMGmTaNctaTkDL114bc18slbxioNkxEKUXkXKJbRQxLtHP9WhlcB+wWqOkEN5Z0i
lPM2ApUZiwJu5CvQ2A3m60K0xI5VNMmm0o/r5xm3nKOsEL8w+I00RHQ/pl11s7Ughz8WOtRSbVb5
p1jbSty0n7PQG7yL1odUBU3GxYA1/Ytd/ltQszRxhUm3ub2u25G489XviQsYb/AjAFvcnJkHb0/C
ZUvVvdBtKj8oWoirMV6qNLGZg4jjLtI1zDR8gWTBTa0zZJ6fK0oVhAwRdoC5bW47FpxmJIAe7WI+
3s5qMWj7Z+Wbak4064mXEhstolo1sjPYpIODyDjc6siQ+pjvB04/Dm9rvfe920EUimj6u7+Y1OXc
XdhPzkVaqlF8SEv08VkVoA3aOVJ3oquNUq/y64tnaY8tb5lfgZndpHyinLQDVR0wlyx5i7xkIbQp
eBGy3FUB0xI5XdSI4O1I8+7Jvv+dvr3SP90V1+LxiScR8ueGMYes6B17TiBFnyR45M46OmVTClmp
+d00yzK1nqTY0NCw+K/O2tHyUTVcwD3jNhpYLkBGtNWtA7gBBCSNESxiFDDnCXAUiQHf9Ljh4jws
Q8+ulv3PH+TCK73bdv7Hh35KYlo8vr5WWzV/U8DUniHciPm/r0a9o3GdTJrheusdFsVcfhZjIQBq
Q9ht9DH9ktG4oGk+GBniPvrLbIMROH8Gp2eyaDeOB/FeOmZheHyruELOwmFb1a9DgdAF/ED+kUw1
9LqWB+H01tJ2vHxhOJlqepWGMDJxM7zxhMG0xckB58AGLT+4d/UUhnNp5M6A/3dKjNCOPyPj9h7K
jZh5bLDfdcj9CvvvNxo7OBopa2HHF9RQDexooWGa6xim6Aj+cnYa8Ma+ju7AHBx0QC3hBAqcXBBo
ek97zPax0zgwUeoEtI0z2soaLs4ZUkdEAlEpDsxWNtxkQqQ1yJ7FlXvYmeIYnucsUNc+E2FIpWsm
56DdL1ZPHlGY2pmF+NSovljIrmPtOD26U7tY6lnF+L384fZ53IeMQYg7rtcVKtktC7fIvz1FDuRR
bMTAL4AQtr5jflDyqfbnBQB7Uqdka5yuUFfDawATrkIuNIB8/m14NCJwo+XooK/6iyqXSGNLpkAf
potV9jPy5HdydTkaSvHsaqF+mUhVv7ZqFm5MtyWVB9ZPlQ9N+xUTve68PH/RneZPbQj9PFqmN+Nj
vvQ5uMZEMxJeFkqsyTjC1tf82YsAkmZ2Fxy0QkIDH9/6VpbvEtrnxtn0EmZAnZqVvUrIIN2iHe1u
/786crmbjM8cQChWOGAMdJM3vhXPzhwG65zr2xAS8Xpxb3UfVXgM5aCefi7IDz6YP+a52VeoK/LT
yYkX5urcwrYKe55CJgu+ocEUk0dt5sbc7a5jzUs4pMv4xddPlIb6u//4k6FDUF/NKbTuabVHQzM0
5MGagSSySoaDQz4HMAHrlRXH6bxXqJ2gYk+bHGwsaS78ss5QKGaN/zKSfn580q8eIzAv/rvPuVfW
znhSYvqiry7yiMFbD2FInCqLdYEUBQsx1/v31MHzCyTQRZA1U4RlwGEZhF8Bqm0z1dEhAkCa0cMB
o4i++LENdFSPN8iGeqP0kWm85j4eXEx4xtXyftv6hqeF3quNJNqlCPLOSTCMyOS1ig9zXFwOume+
WlJLwzT8Ms9do3OjF+ijRz7OleUxH8eD9JdH0vNjGhSE16CVKoBCEY1CYZkSEC8wDW0XUWgLNkW8
pkAf/6R96kp2Re1KvaGKwL492BqF8jtC+jyb/4XZE3HP0yz4hQKh6ejzzkcCi7jLBsiL0CJCiC4/
JaLKgdIArD1npMt2SOlqXDC+5QiDLEiOs6DvdWvRJGXjnfb7rLT5sTSis01xihI1FAEl6OpWnBqU
OXPGmfbSi0ON1TR7FwzqaAS5lfqIrumji3lMpXI9gPVgkKH6W3WUZgBuKLishlAoo9foVbPdEuI7
5VDnzk9vPFMdjmOvCCABzkit9OzktRexHAp+fSMYhPf8iBdabCZOf7s7Tk6w8E32O4AClmQjMxEj
6KbRgG240Q/sLgMfIe8qYM9dPxBP+KS5Nlo8ru9Ay0bhxzps0oy2+Cg1mUhXo+pnV69Mo+Fc8sh/
fVAIqscNIUmNorH/u90UjOf2t84nCoooPZ33AhR7BHbHkUBq3Keodi2vd7WCRJpvTa2pxJWmZXeP
CisvYhnz2dtjCcixKDWpAG8x3hxeW0U1+j/BDXjWgvI5mbpaAnzU8M28yMu94Z0gjemeVO4qubVF
jfPoGfePCPoDyQP9zxQLb9ojsThwpoUVCdyjsTqWZZsAzNQga4J5l5jOlNEcabOCtWXDIhjN1bxn
1aof51GJWO0tZpLhfmDqlkSBIMbTWChOkbYjkMr2qU4TBOB1aVY6KIIHGRjzePB2HlbhEBWFeqo4
6N8uVtJjA2c4SuZO67q74T1As4TC+z/Ecxt4Cjgiin1ByUUdm4+VHXVEWXvz+j+3dlRVSaQ1MOJs
V7vg2WCabcLCU2Iq0e+Pj9LoqCiMnO8pQsFfeDcZBl51PGg5fQCl3CLVE2Ank8d8GKAAaiPuOwOq
qlS2/q5umgECGdG1xYBkB9J+ejS+c0o1+2uynUeCetYOikqXmaqa11Wjw3hL7DfG+lN5dWK2ZEqf
KB8cKPYLWSCArbPDhyoYkm655E09IPVomPpBZFqPMQQTFythmmIuzgoazbQLXrtr/D7Kl4eAO5+J
lxBaSlyoIxyLySf3VUjIQ86LEI9kvim/yRvkH9Sjgn5TNzIVK725kfq2rDz/k43fv7vfi+pZsZKw
Zfe4HRe/MZX16FDj3eUKxw+Mjz7zAiWSXZeEXydc+nJF2+LJ+XXVSnK/DQlAyCj3pDnJvAFg+9aX
9jw51qCgL56awEpe9tKxZwfyrdd/tj6qu382jZOK+3ALdO4N6C9fCFV558T5pSOHP4m72z28VJ+x
V4/XYkNH+iV3W8xDUTDA6Sow7ppfBuzSmYjpDS8kAW6lPDXceibf/hTJDPXJB2SinzU9TiWAqtAm
ff0MF4T8BIrLNgPf6cVk40magtp5ATZe8FpnWv42aFyHWVrqeTDKru2PiKKMtGaO3YUAxnBWJyFk
EFe+H3+aEbgtgUvaa4paIfozkJ7BSIxLNlczoxhekVceTPiBzDWJcprtahnDNldyChYvWjNd3IM8
knz3ZtxN3PQNZsvGCY29biN0zgPylZGMEteUCDajzPSezLuB+EEJPvfGGpGVHzSDYU3Yb3Vz0vwg
4mtRchXpkVzczCvNioqfK1b0GvU+jO4rlhONCnMQ/OLaAVHg7NXEyRq93exF5HHffYo7CDFGOZIC
rqGtZaCcNA3t8BqBkeWKjT6J22Wb2uD21cwBB/vEFYEliGKKa+TLshN+um8JjEFWLPSFSRwQUqzN
5vS5s7qVsUMfW+fY6a2wzPeFOkyQLtJZlATBmt2VRmfbA81aSNVIUnRVZY92iRv2BAf34CaWnLbl
nBK33k/RzwHHEpY/Rb6B1bKRjQqc8c+8bAmFs4Qz6mzmnpZB3k9zl85N5JDHf7RxjlGptEsFvhou
x4ZTf2RW1X+WBgsvSeZQ+d1rVpdyWUtbqh8Wc/PK/7axWlFp+p6+hTumJLGgczhbvGkUsAyKWUFm
2Nvrr0dmTv57wyeaIwFC0DKyhVE267Kz5a1WJqeetUegC2I2jvFCdrGR18xIOWLQjZGWKrNDUdQ0
5uuh4jkJpZitpiwVYDyyByNFRZYoj60zSHZUKhuIeFVFJrxy10E64kkJ1h6jahFcv04x9oWjgn9f
JOLfavYeuu9qvuZVix9dODHy54JOqnrGMZYoYYY8cAtJqFKDiA50KFgqXCIkoz6cO68C2FIlRKMj
JapWt9RtQjyrszS6jJVB+xQFCNx4rU5a1d4f3guHfJ+MBKwF8xuQ8ofG+WGYSdzLd6M0RdpWy9ZA
33UGTdn6+IuXx0zYT5nlosMwo+GiLlCXKACIphgScqnG6F5pDvwQLX8GJJGtwIJZGyBPgEYi7oi/
bIw492rvvNIt1mHk8TtGS4oUd1Fme8dlRazulz2PJsdQhaDdT/o81RDok2z7bxbbBF5cbZen7qfY
KtLLObIUFPfPmpgOjTJ+eIiW9b1xyRlCSJMGiX10S8eUSeUr2aqnX7yDTUW1AdOBJF7zZwORR0Pw
ei0IJulpIC92rvjxl62CP6Txn9MrSchw9F+DrRmdHEOB91rJOIwVUJhB1UoEpA1tZHJqe4BgAyQz
r8ktO7u99EcJiE3Y41X7poo23L2tgpGRxaxSoZZVC7vc2nwzO/Y/0PI71Pc3CwMCfJGG7p/yPeqU
xINQJYjXm6D808kJ9dRLkNIOJrP7y9EJ3uokKOowloe+B4WDCwFMDIpo5cbm4WkD6jJiwst0VF3Y
TO9QT8BwUBNhMQJ0ggpYjCm9yjBOsQM21M/bo9d8LKK57pXQNAbdf9B7eHN3L4JbkPmevAeFrruT
GO3AEzIjJ7CuHfNNgVzRGTIyFhjjbFxPHtFIDZz1AD0/k48R/3UKnufzFdHm/3YQ0Bd6sZQz0mtT
f1MLceFlqmWZW2levCAz1lQoa6+MSZQFs/At5cyM7Ibqxk2oWzRvnWMVgKMUrQYTlymij3qPDMVi
n8qy9NokyAioXGj9asG4BRXKrHjqIXo++0s2wZa18ztw9J2paYLjOcWE6tvzRa4E2raPUaMGOsdv
bnyDCq78yyUvOigM+yFYULL7q+Ri3xqdBogT3/LiXdTxhnnmCTE+tgadThGWVW5b0qulEv8jKc5f
FSXQ8jqyprfzB0Ar6ZEvgzxkukUvrn1g5tVIGxWnoxaV/7j85ZwVqLPXqxGE3cccq4pGe1uD4ysb
6twqET9txoaXgA3BDMwiKQ0MT7fGeBrxa8mqYV7I59SgXnJO/bNBLIPlPsd/JoTCKxfgA8BEbt3h
Tp2IGMidK8yacj7PEYJrwee64DlC/7B2jo88J1nQsnBHK2TsEfdv6yyr38xnWPsCxx5CUtUkKuAM
SwwJX+H9ykhyneXHGld3AkAdwlpwYKI6UcOy0DbOzOuY170db0Jt1qtWS017J55EBQIMJbP7xzTY
EoJCVnqy9wDwv7ZAoelDYpT8fQhdBJrDeeugRnBVac3aF9ZYx9kVvK1TkNgFyF0s+CuTYwZXl4Iq
pFhq0KWkQMEqmTprHR53HlU/WBp/eFsQn30Em6f3FK6DhPwQ2YnqmR3yyH/TGw/fRed1/YphDf0f
XB6ibM5AkAYO1c7dTGCMKj7qg93BdC8CzIXM1VhHWtgnti+BQuyo8X817yt9UoCT965eoObBI2/U
n2JNuICjxc8ggtWYxNteyWg3qGpaAe90jZV7CQE1NC6FHSckY78TwH4NUkE7i0DDqZduvZfAn152
s7aLG4/tgVYsv8ORxKawvpAJsX62ge5SpZGA71m67fdjc+AO7+dU2n+Df7bbKWUAeclJGWBfabxj
H8V7OQ9Ibq9w7dCHfaK4BuE2MNTvANBUFXzUSGG19t9UxkAEMeK6a5/cX7JgpMOSQFXKVCF/CDZ4
HNVfnZRjfSRfTceXQHbBi63PkF3/Oaqo6Klz8+I8X4/Dk4tWKhajHIAYboSGf8x47mA3fmiMW2D3
C/oAOCoXRw7NF6sAML/ivZl3ehHFekruR/3Wx9oKzI78XGilTu74kt4E0VZ0INlpHv5tuW3fna7O
uuXngsaBAMC8A4gtQMlqcq12d/LMv/zst0Pru9Sg77Ps+2HHUbKS3QsaW8L+C352PGkjbAy+4TDz
8XinC/awcGJu/xHNn1YHciViCVwpE6aUPc9riJOe8Qrp9luUbRCAVvN4dIf1z+55sLDqJEU92ixM
z67I8AxM7KyIonZuT2DZBSQdftEtDtUWCupQxKG49+fLFHzPFV9AHMW5FvjTNDEueE5n8NgPwLBi
X8nmk9s3HxZ9iMhU2YollBzq2RoQrQAxlVMUN2ftu4Qe10lWd8a0R2Rq67JGxBGnF8nQRyhxVKy4
m2NCAM0J0vP78EfPPaKU64ZZpPtxUsQ9hI9vHvodWQOb63pxoMTRdnn23tUrocomPIhvURsyZmK2
p+A919mUWEGj1GrtekvKlpEe+Bf7jYhjD2lD3YRjTfzrfzyAlHCbaOs7g97wLr8dv/22/rHtDwP4
X2TzFsUsmj3r5relZJAR3GFigmxHA0ls2xrMhKvRkiM1e3CXRtDNDO4zuHEtTaF9/jXU5CY6Uh1x
Kcd+25Txo28k9cY2CFL+F5Mx5wfchabeA6a5Jf6sIJKj2Bv1Y6XnOcIuoDVJBe+6VUhMfNRg1g7d
ilaId8HFLxFhh8Uw+IgkNyF7EvUesf7rdk9F7UbKkmgfuoHoXUC0ZpJ6a/IQh6XBFvsHziXhZanU
rS/f9B6lL4lbePJppb6b2KwiUevGxfgWjcK8ZW8CcD/1JakZbYKR4+/KTBUZ9WeCPRH5xRvnJy8O
mphz+YmemVrCTFgP5G+ZRak8+Zk9rBluGkjhRu25j+3Z61RF6Zg/N/93e8Oh6cjHYu2o4Fei4S3b
q2ekjTLwpWrOHSJP8F/NUnAJu0E0sNqtohQoASYI43/H6oci5ybNGzc5rPyun/KXbhGWnziN2121
2gM9rMjRyC8WuF07rmgpEyZCyJAEdCOAjquZ11KjW09qx5/y67ieRkWHdh7XuhyONLPEwOQj0w2z
+5+0+rGFY4ieRX5WMUnZN7bU347OpEki77rkyh/Nx0+aH2BTpF0w1RmEn3fI7DKmdEmuHpeqDLGt
7nfSibI5bU2ay0SzCmmM4LHJIsS0vYIoH6GBc44rX2Wf/z5lO5Hhhyz3eucdqiQBpDR/sbmSRcDT
HOZwrXQ8NTgC7IlaFqsCEVMtAEVOX7oU5AS52N85PYUSFGs49fXCSQqBcOX3Fz5QA9TNHQBk6WUE
DB5+JQAz2b2JiPKDSGke2KyLnv8UyQa00648rZsW+6lvY0rB+wvcFR8uNsEYzL1ORjWU37bL/naI
YzAfhnxg2g7h5cu7pAxTWb+wr6TeZVdrBf0obTf6qciLMLKxL3wnRyLuBV7kIyg9e2icRyce4EGW
Czsr10WGE+XDD5tnbVJvCltPCCqAOLxGmhkZBDCo1w79K7/PCDPb6Y0RsJNZZ5IMMdCdPBikEocO
DcukpXN8xBiHj5ePp279hj9p1tBuZ2k5FAL7IVa1tvamzO5f7i1Isl1FcGuZQggj3NKD7eE5Kb1Z
BGeEedLyTbIXy8eyVJXGW8XnTRQeQ234TtU+gipxkpls6LjY6oQx2pqzhDAkWStHvJY+i8/2MsSC
QULT0W7cJhjZ5LIDtuZjRwsRxjage3RyrCHVEv/VArf1lhnyV1WavKkyPjhXBPZrMWr+ahfBuCce
5wOpoMs9uAMzlOyU6MFIq9zk9jYAZEXaBAUjqF0bW0ly7Sn2goW9HOpyVh7OxCK1hTMEsDANrrId
E1DBzQqnoGGFxdO7c6h8hYB+jV6ahXReanU3v6RBvc5iYxxAXI3/p3j7DciivmiNOjxW7V6GWCIc
dBnuDH8a6lqD5axx0IDqhgkowrrRp0osMq9sLpvBGSb2X9c1z4Bi+LoXfj0XpbQWufMGGCDm7JWg
ysgHoF4yqH41288CS9wkiiMyZpIr+If7IieEowwUqLkvcKGLORulMM56tle4ltU6I9M00Cm50pxO
wDb6ZfLVE3t5tLzBHwy0iMX3BDo2ZPlxhzIo1H9XVp19cAdugqq44dik5mdogYulERRb2hD4edeA
2MC6mESE1U67rw7RMQ5rz2JXYEV3XNdoAOJ2QeKuvDT2ObkVVpA2dycuJ3wTTz/7MtyYsOtiJGWw
6IKSaLKC0JBV2znGVD6QZ1R6ZW3h8Sp7QptPbQoU0y4YM0HdUC/iYrdnnRNv9kOwTRBEfDDOxEwF
RSHfZd5IPLVGZEHFzusG2+ARvdHPce7s9edUWxhfF8+0W2KbsOBYjuoTU5GF5t9/DRlU/ZQkuplY
8aJIJD8mc8yTL9+zJSZUI8aD1O5sQgLyItFwr7XE6LlGeK3nIYUFkce1i2nu537ryz7nIqK7wx2x
Z3waQ+EWmexBIf08Y5klvqE+gk04MCb8LwqkXf4Z2VqyYrlBInd9UkTieYgNOe044Cumf4AW7R26
PTSBnpmqFsLNmv1CW4rV2qa/vQ2O8vT86yMfkoxe8L978Y+K9MIDwxZLtvhoZ8rhLPBUrfsdoivb
cmN6JwyEwGwTiz249oaEkiRUV2ngYqVAQVI9Q1GeHLo2qK9SX1gVfhsA2uNPT88BFHlmB7NcfPPM
H3wvO4GC91u2tRU8hVHiati+gXtaJO1jIoW2ycoabDJo4XqmkwxsH2jXOt1OvzqBs92geBX+44WB
i30+g0ASTyy8pjQvtQKl6uw0akJVvDt7kdvBdPXgGoEeRIOvzcT7JZZAqFPVTOAJtAoPO8rr/UpK
7kNPXgZKVWzrOfO1GMEnqUqGcno9lfLP67Rt2ZTyc56cPAz0H2nxesD0k9PW0I01jIGrXIu2aKMi
SeJQTx8aT1ORyfUljkIBLjurbe8msJOUBK+JCxF4O76ebHRuxb3SCoK6+qOfZd7mx3nzUAJt13Eq
EtSw+RNDNzkqqZYLGw9UGJSkzwqaywvkqTqI+YA3gowdDI/bj3kAuz+Pmg7bJmG4JAkPMkyIwdtu
43rmOVD76A0m2/nQieei+T/nHl/EFuX3djR5odiKM67yRj93Oncwi5f6lyp+NhubthQVoQpJNglc
dfTtD3/dlArmLyAs6oTuXRuq1L20n4E0LKp5z7aAlFRw6OJACkn3kVTqzzoP2NmB0vYOB8dlcJNj
flijpRWC12kdR0jYfscsLcZIaHt0K/uphhvYatA6MAvXi5646n0iSK+4MXG4WWbspjDl/nGVm6SP
bH8uYGN8HiWrdtzwaNwBCsDGJByK5QmAKhxR+yTLniLOb/wajw6mora8DRiq4DIbPy39JfR/hEMU
H1nR8jgV8m1LWnrPXeozIInEYGnjYH+bjKMnRCzr2xcYLLq/dqzlaqp9bIh2Gt6nbdZ7knIugVZG
/re65tiW/aKoIsvZFdubxoOGJlcRAVFB8OS8tKNVBJUQ/0qdfCBudPH37jJw+kTaigMvorPuLyqZ
x8rErXD2JHPL4Xq+NCKuQYcTwL5BiC1+FwAA1uD+re/FVpCgSBuZG8mGwwGMugrBij5UPbRLQ81W
yWuLn75PxAWG0ASJff5vvO+EUuK6CNCOMZWoL29uCa/QiOMS/hg4sySw4gGL9SQOhwL7j6U2zubg
Kqmd511k3RISUk8pFtZ2CydtAyYd1eku+1hutk1ioaziA71speIuYtIlcU8boBeI4bI9gJJE3DrD
JPeOp6RskvCdMl8C4Ce1+jQNaaWHme6pvlZBuiPwVtAA19W/2qmT6ofKtBPUiDR0oSzWuQMX0kyh
GH2VRCiRARShRKa+VhB66NivrAkqmVfYFCFH5OE0qzZReRivVFPCskxQp+JZ5gCNWpEBUdF3TAIL
UwRHnbaTo9POlhjZeBr4yBxKmwi2Xwqfn8SG4GceMVGFOfinmVQ1Z6iFoGXPwkmv5RcTbkHdkkUb
mbV9NJTPiuDf8+A6RLaqmpCeEQuBGCTjgo1o/d2lOmB+7LvO0zJMckpc7O0gGHIpML12FUOWlUH4
IK6bbrF+EYQzclJ6ESyDmYcIW298PNgm6cdopsfgXhdAK6B20v9BFIgV7GOn2/qQ31mdYL6lSC8N
6DKvwuF9yCaj4d+vC+Lhy15ndgcDudah5XdaRtKFl2xHtw34Dejt38vRFoaU297IkGzE+Hap5Hs0
pJ/weiTBQAPV7ranqAm3vX1rBuXwefT5+xs5UGoqwulL/xeULYpkOAgCJTPO0h13sMNPQmJc/YKp
GfX024gh3NHzTGws1FMjfsyecbxUAYivK1xLVREEVuAzB31+LIKz6RcnGWdxZba/tYid78qS7I2t
/qAfBSnNzcSSjEQPpOGrS83JNv6rvVIsZUAusmRGE43u9mhUU8F4Iv7w8Q+GG1E8v2ZdnjO08J5g
4cCFmtbNEh3K6IniZSw/8S90UZXYvTU5BGzR9L9rK3chCBsU9bLUmMf4CUlmnDu92NUBmlYEUwY8
9SwJ3GHrN1qoT2jZOl5lX4uQ/l1xjAoCygmerFrwFsYcozVEyy4cIHOpFVcPet/Bd+aPMfWFVp8Y
6Jxj9ZfPQILxuF4OEX1o7Hx2MlRzZGgIYZD0lLiovQVg87vKq23w26FiL747Zte37VwL2KjA7ezs
YgoJkj2Yf5NqeQlcL+tno9kaTCtF9RqYoa1Y53PB0Kor0rCwdCUr0yVcvInMdfoxDkcWQsAOcerS
7jRGLsMZWQdI/6zMTDwOXEE59UqXpoyhD9ztOMfSJ0dkgMdLgbzqw5Wa0Up4or3Mx5gCCZDD4gT8
9NEKrfHursXvuyQ9XosgK3BMz7PQ8t1WF2u/aTok+UrNHzF904x0pkacQtpwyoAM2sxppk6fy6Hs
/PLDdWf3CQXfvhTrxZi5lEBJeA4A9G2FBpep0EULG12Kf2rc62pyMkm9a/JWpsV+j3dSFenxe52u
aprJKj4DPkPb/AGmot5mUONlUNI1E9jXz7XhJAc1WVLe3pISfmkHkViStDnJYo4RH5I8uEwk59ct
3fkAet7cMCWAR8rySa3surnZ8gGysK9fej7gJMtHlISd8i6o0v6tYv5cpysGevw/JrpcSvCHLRZi
Ep5MCHcrP3udU1R4gNYgh42UVBYapsxcwca6HthQiAb7I2paYCPIGRy0WunlrUwYuMfD0bgdbJE5
hU/A+4dCaHCJOv6rajLZ4P7U4a9y+HzIGmiKBcvis4NpCTeWl7EybV9B+Zqa50j8lv76PlYDDI43
oKojMFlYTzcQsZbsDyJDofQv+Q3aQlBwqe9mjhhYEl/KjryoUi1AXlQWE7dkCocNAdqLJJOsnAtc
xeE1Tmu/EklKgQeshOxuX7bolpmrBaHTbxhPRDZuDIahcOINHOoofK0WvRhuZfvKUwUpUv8WzDK9
dCbydPlJcG+I6YDU7VJGxCrXyROT6z8iK6NbWAOi3oRhf+i1kwZgfNyAeeD4DES4wVxXi1xe6UDC
zVe0xkKRHm/JZj+3Bf95Lw4Sejz23v6tgPhGwTgBUC8nMyVyHB29L7aAiAEj3h/1Ol+hp+3falas
LMstRtEJwE7BfDQrgKSKCg8dCZoUJDOgavxeAKdBdF16x7Pf38Fr5qADEpIWudtIEXjjHYJF0NVx
oXMzzcJNvG/xyTLzLFkHHT91gueaFP9qDT84lcE7PTMzkSJ9JVOvuw7moE7N/qvdCvNbgFpKW4OM
9y5U2o6tHS7by/C1Jca/fv2BGDd3zm8vpODgXAs8KO39lrP7Zbh1COJBcX1iahqVbDtIxws40YNC
yHMchdKGbx/FYYwzptiLrTlB3FmoWg6PuE+fDp9APgXXLJVsx3jfLIl1zEDdV7J5jWJGVeHGN+RH
HPaf+clSPYaIiCmbksXtSKKAuVwGILQy2uI9U69U2JVcmTTBrVEBJrX7OxK21JLGZXhUP65bt6x1
vfVkqUbLsdi7JGdiQ29gqKH+E62BF8g2ReCi9ZJExfi7InPiFL4mZ1Vs1A2ZpuzS0zJhNRskC4T2
ufLNJ/4RVaP6wufoxflNn/PM3eAv2H8XSOP707xeuSzPlC7fmENjCY1CYzPCiGcxtiujbsvTAoZg
7Mn0em60/TTHjpXn2licZeZkhpM70Y7xx3oAf4YBpIldG0FURL9oyo+cKBVEQ8VCafsr4tljERjp
aC8b6Gm8VQRBauK9hbJNODygVAXbGE2xfPYlabi0NFmk+oFYOxxzSrblymMTMHB/QSv+w7yp2erS
B27pi27jd52E4bciNFQY0z18WgbqLtk4R5UE6Xc6QPspZfTyjP6v4NpUFXNa+TppVWx4yTjoVQfY
jCUXiITOTQ7fOr/5iSmy0NYmWjv4c+wGIk1A/CcfOFWNSU2v0dWipHMHhf9izCcqf51sI9GFvY+k
rRlSMYfpNrntgw269tPntB++7xHKC8VTvL++fnPb8bkJx89RIS/VuJgdwYXIomO8Mlf3jB7ua7QV
qp6hpeKYAn+v9HhB+0058ho3Cfqy8s4NdyC2K1E0V3af7QcNQ1n1ms/qXzSJPtAjy197+C10o8CB
UqUpvPjpzXRw2CfOmwi/qZmrftXpjn3x8sqIc/QQ3zzprxbQmviSVYWz/dlGcSMSR36B+7GOLz6g
IU9yo/qIodJqM37IolD9S94jbRDkQUnsJr15WvicsRVGCJoTQHRDlbjDM/yrLS0OWohVNqJywLJR
ET3675P5fRpkYvGWkTUe0IWW+0GUcJ/hPmk+5ZKfdNffcO8qKUJMZiWPh/t+/xEt6EFLCvgc9UnW
omMrWUbBkpEV6Iyc9Ru3Qy7pANIGRCkkzXo/G7c+cDdHTC8FfClnvMtiPLCG2SYHGZMg2lvlNY2t
tt0ExoYoEHBRurZpyb8yhf3R6ZlW1piERiXbp6V/4sVdJ2+GCciV+FbrhQ1J4jm/1tOt8ZxNl8tG
W1tvjZOPLG0cI82aNP0zq4UKIxC7XmfNK7qv3E+VQdaHKSsZYhs6gC3mel0jQg4ZWrut4/68NW/D
lzq/fxoMFykI87jYNgtZSM6/EQ99aG5ONyN+UzdQ5Ypb1eT+VUF+zhFLh8VOU+KwE5YdJCLIorDI
+oQasTWS0nFJmAWRhxMckYe5DgKwE/OKhKJV4/sLNaDIg9A6awJjzCk/ZjJ0TVSD5UJHawSW8NAr
+fj+Q1L0pfO+jmH06PrZAWWwBW5zaNQaYTXv4MTJWAVSDtCdffzVz+cp0Z6pGqF7RQkrQHQG79Hn
N3hw4tZoVGtIYgrITWK5AFCvzJrBB/Skufys7XDQY7K7cQIPRE0SBLgs0vyFgExoTavAEUP+BR69
mxhHZEsNosDJREhXxXFU+b7euwk6Z8/nHlT5V9pFv0T/BYRjMucCafC8Kk6UrYwGw/m3eiM5470f
sPZehVsHoeYAK2fiP2DEtUMKnNTYCu+amYk2s/MQVq6gxWaWolRLItjXegJoEsAckjv4e6K9wNP2
OY6awOwIWIZpwKrP71u0LdIhmNLpbGmF+9bOr1VNUI+0BSWJRxkHL8Ut6kuHcwMGUpMuhnAHkBG2
U60h8sK77K9zoQp2bx8apxj/lRNnbD5Fp+niB/e3PwgBIPQW6xSu3rzZBFZmlULq1qLiiq//wZCj
jrHgzEePzluXV2hjp5cZq2+XV8oC2ua5hgMRKnWoUCjXH0xEd2fnxdpdLTwGrsB6JgtgkdrgquHu
1JMLWd5l77W60ab8jck+hUL9E/kd8DUHTwFykBKVzsTfkZdFFN7Zz40obcHWSCOZ3lMEGeymeQti
VOVGg+UbRQi1htCaxyYdmUvX7xFfXygw1YCcptQqg+M7stKMjAsKt/ZfaJjjpPTGFdNg+X9YMKFx
ihpjh/Zl01abxn9UgjEhpZtik4VIotz2Uzeh5uwMEwHwhrHq+OySa7m0JzD7lLZr3bNd6uunMTRY
RWSeQzSPGnyQm/cD6nch2c9e0Vd55pTfsC3F3Z8I9vC85EaeEXNCaX/zPeelIhT8haO2y7WVPH+f
5lklaD/OhvxHLmTVk2HIxmO6yvZglVS5siVQgV+jBK+9P9lY9SQ8552V9o3o0iyZW35H8I6w1vkb
VXg9KrcGFICt+gzqBzdARCBvEfRJ0GN0EB6Gixys2iAGGaYUF/LisyKM2ExZAj4wqdgUbBDgp1QS
rTQTAW6kosnZ3Fr4xhqSrAkJr1CF3ys+vHuHNowTbDuVf3PTXPy0MF+t+56tLgPxtOQUU56p95oX
T0dtQRb3IJhiA24/I4EEUQyMsQq7gljdYhInoZkXaRrIqmwoH5xEps40kM95ZtuXPjSPR+Suqf5H
21ew4UDw6cQkhY311Gi/2wiwcNA4fFgwb6hBr1ingSKvuC8TqhuhEfyqIHfE3ifFF8c9YQmYx75N
PcnPAoOfsSMoExPY942wQWtCoSHQWZkJ5vcj0zTtmwp069EYqam9VRZSsfcEwZXE2aMy+Qtu1ZYt
tB9WzGL0oG7rYBVqmhFRzWc8Axcu8RLTwGk2lZBZyGODEdT9f5alqzPk60wW2otn9YgggCkkQLSM
j6t/QOVqKuRGZPBCq3SrAtmQ2MgB9aF58o93F7JDO/xNQ8o2oj1PNSExCxU3awrREiMAvUK4vwDc
4L7hf7zew6zY8ewj/GaVuiy+ElKIfAGwVvzVmsGT3nRrZtPDlIh1hWEb4/w0usHveY4nzCGvWpWq
9q3VUmi0vVz9uxiomgvjkZxjfH1YK2i171oN18Yj89wamc1bMofBPPbFekgApGS1vbs6daNM8bva
DHpAuI7e+IM19Nu2QLqDtoQJGv/nyR/mKMMsId0yGvW2+K4LND3vltkiEAS0cg/f6iz5fdqdUi/F
4EAfEQqIVo5vKq3G6ziuhdrgPFY8skXABoppoP2QEBlQWkjGIASHFAKBYB3Pe9K9ZRBsCC15fojG
kyIe6tRZCT1grqWhNTtwNjP7ymR/6fibSjkRAo60Dcs61ZLNkqnbJhIXUwxmUNralK61tpQCfb6c
QVkiHBnMSuhgT7aXwMJ1IIOKtiD8osphUJd3cmcTPF/WYDiikGF/Eg8iB6K1Xor3G8sQLU3xkL+r
qc2Pr7G3I8iAAwBmpcLqp5/nj9bndeeNCD0lihLc9kODf9jqaKI8wxgX2idnctcRSiIsJ5wAn99K
bHzsD2gTEvAEJsgBcsQyI1qAVmn+S3e8ctbU6dmWvqx2PIt2sIUk3s0K61hzVHJlMUGWfajEem2V
3BE1/d6r+wE5jvplL7dqvwnUTpGmrIhjxRS35xhxh5mKJuqF6RrWp4p7VZgYlNIWrKOcN9oZ/plr
pJDP67c30/DyDfL046PX2cXuiy5wyN4ovbxOruiIvgH91NLRGwVeDQFAjgN6ipiLQBAWmrfsxyCD
mhOH6AZp06MBFez8hsWmWg1iVz8/dPSosloZT0zWKeWg4ZVCjZca4MGHs54NqyIayOh2yyROZ3Vw
28HeuETWqlxr4Ur2fbMiDGe83p4IUNXF3DDEEqd0mkLOtxEMLlqESODcm3C2qad4/CRM0ivp/NI6
+DCjhMZW27liBqGCdf7JlYOei72Y6+qCJ/ZgCOpNIwkVLPPyw+Qz6MB3IF2oWHiR3L7n+DeAweW/
RJkdP/+D1JgtG5aCIKTPRQ1juuuU3WBEGVUYH8lncZBGa34OuzzuhGUSgUWGV00rERY/Q8cGiWGS
zu4fYYjJyUMg8SJkcHUtSltffCOGeIYnUvQi9vyybVxHHyo1MbFEti1sMPf1s3qncMqycO5hHLkb
dMH9IJw5yC2ntOdlFkcekcd+aw6DSLsjCcXWi8xRWN2aTq0EqqA+pKAQGe5yzXcWQ329gDktqhrh
lyqrDbYEKIhlYP1f5WVObfFYce98AqWjyaCYrQtobV1gfzTYQD+CyajCkUaGpQgVpXa24wn1x8dE
hJK4dgrSWqBtnrq1Dt4Gtj8n2+aj/qHpMEKO5A04/erIv7XyzTx8Lf40/wozW2kuMLcDvGbAoDUP
C6EyTVoyr24yoamlKROUxAdUfdql8Oty2sd0DAwFsDMjH7UAnJ/wAAUdZ8e6CvJJ6uHkW2ktsjk4
J7mSF0EAzBTrm9I81jJle8nJzOVGalqhShYX1qm1G5rz/hJclpaA1//vEx1lQDXb9vZ8NnIHb708
+VypKeRejn4nxfpuDktEh0jumyshaJlc0XY4diQLxOAHwl8xLRbLmlQwxlHhALMF4Ev5KYCDsU1v
ezEZ8cqY+XGv+0GVGd9tCO1JmeLaGhAGci+iNmZXZCmmaW1s8FxwwQBkIOzaaoZHgaUS2gIEFnTd
OHVBpTXCL6i1O+ofr38u5b27zcx1OrkPRIxIywQtst7jAp1xitHG6ZT2H5BHQSGyNPyI8Szp0GcY
Pqc99K95110F1cEkG2RL4aCdQ8R/0222hNvuB/T+erK3gt3FZ8YhBdyEx3ODeJV29RVLCAny68zj
I7vhTRdOXGrT/4TIzZUEZmgkPtbWEPzCA7sh4JLdvCm5QV1/w4ApxG2rFR3BfCmvXFc8MFxth69V
FJ1Gkp3/3bsrgCa8qFsbQ3td3xAWmIBOb24QF/QzRqd3rm6YdlqbC4aX42KyIVSTkRW7PClBqTgO
AJBa/FpDnDj2wXK6adCEZXU1/gh4rXjj18sgp5UIyz88xXVbYU7Yah7MJcd9UImMj+cIFfZgd/CJ
2VjsBaj6gTN3LGj70GHIfab0xbRco/fy9bMAkj8y1ukovb8Am4MUHGZVPweWs2d7IcqwBX/upOnV
VqPSeNSCho+JwTVuvOVXfOBBwOim0lSZ8+8rBuc0zYSRYx9faigAejibQoN1HoU5sjdI/seuLh3m
YQpHipMOFFT5Z84cxffgI50SrBdqu02rJY7qxErYL3/XXwWrZz3Vzc484LnRjUnppgbO5Jo0L/vx
bfNLlko2f9I1sPEYfdfdZzCf9dSg/uxl7dgsbnrWq3Njx0iN2MWijy4icLWRt29IQgQj4qRoC6Bo
pl+9h9Ti1FN5vyGIZZ+SaBHd50IAJvSe7JmNU4iLVfFaRF8j/xpf7SsnW5mjvacTKTkE0UgGBEGv
Ae/9wO88fn5dwIFxgoIR6LX7Zts6UUeMZJkVNoIe4pY98RRSolkXIMH48xoEKi3ME3MjDrUEc3BD
8JgZs22P/3kX9Deh3zdw3duUxiM0DoMve6Y1IMptGuN2l8jUNKKe6bGeILv6jmu9FCcKlQPggOW1
ZkvgBQvAKcbyEiGjt31avdiPwSfUzu+8xHxYrXb/okvBjqsrUJhvYV7QOkPp+1X/82pVpnX+TzFy
pQbnCnSgPkFj/zXrY+2oWjPzM0wObZHD55Ga9/D2eP7mZbe7LjFerk2wqA7aiVOSwCKzIGbRordh
83wajVuxNP/YCIi4H30yCWIDS8/y4lcrVIv9SpCt9Aj5GYdhUbNr/5Fvi9NIEjmp16e//cA5g1o+
HGm77265p4tdXpvSaj3tAk/pCr6l5a4esYxKR8DzBhaqTPcUBsPhuP/sY4SqctB+uvZNNPOdSb9r
qL8npgnX9YyNLWoGtvjU23CytunNqI6ukjQ4CJXul8VOFanNN8oJW8yW4tBAiaIXstlKw3E0dLOA
SOWtnnzIN4IDZwjBdvcxral+k4ZXKmZHwJyWTkFQl0mjigm4uCPojXrj/kUxo3hbdWiPo8LFJFI8
MlUxLbeMAblumd0APJ1HKTgaqfiUEl0z3rr1hswA9+hPuto7NgOYV0rp4575V5DEzhpEquq5sJED
wsjOOikr58ZL5g3oB8OVHWYp/Vu2fJd6ei3UEK3F3I8ulpms3Gu8aYTrSdjgfexbr4+82lBaD5aV
tatSf21cTM44LRrwKbW496lptV+uahHk2HWx7h9MN4I4LkNUdcPdVRpU9H/4nmb9p5PYu4WWKcPk
v7t/66BCOL7jjVcyR2aiVLhViIAVsSvqT4na/JD879/XPKypMLR7qAMtzrR+cVFfPvdnmdwfkbBH
CtyJT5H9sg9hQY6FLz10D4EANs3HFZDjiP8UGUbCpOuZwTyjqJLYfpMGYb6fYPRYWsBbimKuYAFi
P80Te0EZ6X4nAZsJgVjMmlVL2qa+b3/igt44CMmzbrAkShYd76WyjQHH74rN+n3A/ujtmy2Eg1rS
omv9PiaSd18UgOgV8b4N8W9YE0vIBRcekbXuhuCiucm/rV+UtY053XzDAWK5wQsjVkFWL4Qf9k6Y
4fTYuJovS2LR79ZGvnk4x6kRI0AmuWwHy730ZFt5QLNEA4OwTQjB6OPnKod72eNSMBJT0Co4oaz1
7+CwZzTQd/FqxqoA30OMkTctT37p/Yqp1V+MUb14EGxc8DDuZjAmcZRDF9obkEFvwWP37Fh6UVQa
abXUUov42m+c32wax+QOUGPQletmHsRpexIAr0hnARCIvuvC8OhvlA9eQi+pK2egJfW5kAUAtoPZ
lPRVp8hS9zLo0vVW8IxL0LCMdag2aWsqZBFAoG6Itr7zNHX7/IoJLI+FvRv2/HpehwrNFesZgVeg
pa+VjJOGubVCWodMuZ94MY3NaeF+21blqtxyPZA2aJGb+gjtydX2oJFt/ShBcgIjeNapNya6EMt8
espxoB72C8GimP2HnVIRXkgIR3RcX/DF6yFMOpPxb2SO8q/cKDIe4CuIHCpjaZIep3kAk07XD4lB
CjK0zPh1ftSHc9l7JOhrx7SNj1j93uOm1oN8x+gDNpQ9DThEMWcWp1zMWTHZm3Wn+cEQPDt6uVTA
CpUezFjnh5TTMphKps3YOhg2X3dkMUA1GG4AthgudvLdxjVmrVUjPOsuWOwGdxhm5zIe4xJWhZcF
5zeBOGfA+EU4jtJ+onup06uFb6+2od28qoOcS7As7a6ZG3lkhu5sy2aLmBt7ZY/gFYzAoZSVE98F
If5q++S8k7L3iJyN4CQuUcCEISntDkC5SkMKTxinoNXjNN2s4oMfB014jcxHSTtozXeBlACDjyr8
CBM8gtRjM+m3iDgBSA5k/wJsvR+yztC/3SmpGnGbJc5Ou1ME3B3xV+WoDvYsnvDWiIK43ti3GJtU
GpsSrbBqcRRniLXm6IGkVgxC+wy3fZur4ONMtIqtBaLaQWxchDLvKV8qhvNuRn/gSIlECWsU28ZZ
2qS6ryOLd/uSncgoW8fyfId2Z5cSzizQLuwO9aqclablxDyU2pXfJZTlutr8YZjNScH2ja6IqAQk
mcTTbeEsYX+3JjYodyxZZEsbXUYcIsyScAXM3OxPzoXCzoJm6haqdwFk0E/dTMDaGZGru0PI2HhQ
jjAT5j9XiGjR94LWZHkCj/h2Mb5E4vII1LR/2qfUSCEEXwKmhWl2GgdMV6QdM/+Lj5LhKOUoil9v
KFDl1rALcvM5VLVlhmGicCOYv0iXwsJazc1F6KFYofOAWdnTHGd/ahpa1uaGR1LhEZRzf/sTiTh9
UXwTogxfb4hvZLbuNGLFMQBQKKJG9bsR/stIZSip+HR4mFbN8vz9TK3oiNpHBYJFn1bRSUfEP/Qh
zM9Rv1kzYcncSJipPjgWHnLxqvtGalu5LvGjg5bvTgJSd5OUIoenrUFcGwDeRJhEmOpnQxTzR3D3
Wc0B15ROU0dRqrpgCc7KItajxJEEu5rQ1Y1rPqtpsPRNxIAu23gvxFHKOhIow5CU0HQaImL7aKzr
O2xebYQ+g9Y0uvVW9thRTM1MHeyp5TKlPEr81O8nnd8j5ky+jP/0yfHjJ9+1JFN+J2yS3Q5i/+Pj
mwvDi6A+x3JBVgQeJ/f/fWesAnksjKf5MNRZOg5VHs0x+D46FP4mqUuuS9lBbVh1fAE996e3rqhr
kbkNomam9ILgll/OxgdR67YDhO/aeT+AOX8KrlsvRClNndLkZQVxMTx3enOSHe8LqQUde2ZH8NPo
IiGWt3Z4ffhl8ljEr8/ToFtOWNf6OLxtgmzkULYlYROcMA2e28GBKBCpEeFH+Nw3lFFVt+U+OoGK
JouB1MqhJRihDomBONqlzuzxyqP0TgmGd8TmPTyPVk5pVCqTOGmRgYH++zqdz1kKRdWh/AG2Hod9
tan8Y9OjeJqnBZJgXCDwcbAMwZpvqGsUVLIZ9VzByN0M0pcSZDzQgqj0qF0gjjX0TFn92ouyoI72
P4OTpH/0Sw6tkVoByber1Q63lhenAQSPvxq+Na04g7XjCx+d9mtRjkeMPSb+GksJu2uIrly3yL6Q
bLEjuDjd8AhvaqWEBCcnluY1O5yWYbkGR9KtmaoNiLI/ap/op2gGwX2o29lSqsnsjFabiwyEzZ7I
0Xmj2BZKsdTYFC8dyq0dtfErUkRACJn7QvKjzPSGUGfmPva6kl9Zfv+neQdgqCZs6WPDCgJ272L/
iCPcJae+JyfPwU6/jOd88cAL6YFLe1T16gSNZoij6i++VHOmQvi/RbXchb4oMuSzQeyT8b8snS/I
vU5J6ja5zgaG7kBPvijT/Avv96dgE/fu5C20C+ikGQyBxLuhmHJAa6AkJ8Iwfs0t3LApsnV8hx+e
cxf3mE/3Spc7cXPMu4+FrD+yGobV2lLVK2ZWbqyAoR/Xk+v46ek1hcwXnVKmX6p9gSONqfliE8US
2x3zVXRmlDcd/NoEpP9/ml9+dfSYfS8Gqjwf75uzkLprfYbkI+YJv7sV4+9r8X67kWYr+ltgfNIk
iFIswd4nlPC+0k6rAzKPIRODlRA7cz7cSN2c6D3y7t9EtZ9oMF3M+F2eV+fJVK+jEf1ILSAnIdFb
NQ/5MD3uYnXcXN+mE21TBGh2vjLv15v0N5ylYZjuTcHzOUTlNmzkXg15QJV/g80dbCO3V/xNraHR
3S8dAF8Bv3XoCjoh+FYGV9fwQWy/qgWDhlUj0SfRE7qjVJJcQKYlgfFRM/QH/c0qyAkiFdHDSCJ2
n7Z9wl489TvuZNp1iSx97/uzL1BiS8PU86yiMsZRnnYvQxM9+BJJTmjOvPtn7qoCz84HVFvBI80y
54td31Q7B6Jcj26Usd1paAo7VW+xEt2ER4H3XzPJdRLFst+fgKAZ7juCaFDw6HogroU/13al0f1m
aUVu7s663iwJ+jC6ja5WvufkGII59Dx9qvocj1FwqkzmEt+ao3GnqpGhSVHBOKDv1TkZ1bciCX0A
w180us4b9kbTTdBx12Me5fDrbtXwxqqKVX5yRe2esHfAc7cTc6OUMVXMdvB1bNuhFg8oO6Y7OGRb
Gjvxlp8ATdFD4X3eWpRtRLe/xZqzjoNYDGTLtbPmmwule+j+WkfqVLBLD/s/E3pZDE5IU3tm5dxF
7QN4ELXFkyipK0lpGryj5b0I8naXa6K/gAve9NNiCMk+mp+uUnjUB2MuVIRfVEBYg0oRfOt9UaPR
y+PglKjWSB1oFzdDDUvO3zeIcJa+fhs4AXxC7+guug0vdZcGB5sX2lENC4FMxtHD5YQnJS0HiA/Y
zVPvm4LdnLL+L62zCHzg4Cyyitzm7/+H75Pm/SsDEYt8ProPKoOdocstfMGq4VTH3Xabh+EAlarO
KIFabHeGDcA+ZlnUgAmK5DwqCIHrVVWNEyyKm5MDe9japngPkgO6foyWRsw7xCP/WGjfCMYUI2Kp
KD/YtqEzbosumTp1ErwSPaPWyk+GiQ5eBvIJo5XmQ9d+UBedlYEsGfelbfOifS1rPR2JIv+7TI6Q
iuQkVianrxxr4KasQXOb//sGbbEvPinVR1o2abfnw68DcI1I/mKBtdu1wAIV2Dc9q232X0uxfpyM
wo1U+usFweFORw5SdXRSo68mw7DFx6qJxzks/kz9lpvOMnQ9Iv4EyRLIXpSgL+eqPv2WuHSeENDd
gFQEeje9vYUJkX3Em9xmLQfD7Q38LKWq5ayngNsnqNHPJXrWoKqqZO2Fp5f2Ad2YNafb2ZPM+c1Q
6sFwYUhowWoTnMlXOMJr59TFk+AY8eQbnUJesDSEj5+30p5pcoSbm8/dnBO9480W4JqwgtoYU0y4
h67VXN0eNSj1kciYtUnsnEL2A9qqwLFGWBe+DJcEVKglR5P93N/xk+7kenrvhn4nXYTilKrXTI0D
FbmvqPMnDsqGE8cG2HS1pMbFWbCa9rdgEfktGGsenWoTGqblv4gVu43d6dRz5VXx0GyZTUE0/xM4
L8GgC9R2Cc2HjoFWTl2/N1VApU/3q2Sfu2H2C/9QvoRdwAWvjquP47qUCVlwr+0xTbSbblz0hf0M
dTii840lFjktgIoUQGmZZwZiBFpj3ycMcsOx6sDi8COE9vtXfpBLwsoVxroa/vJkYY4jtmzfTJ04
8zz/SSzo2HkKfvRMy4kIS0BAll/3/1DMnbJXTJnPs9tK1gULH1aCDPhz/UtnJ/0TZRtN0baAHE/d
x2L6puxJU5VGCmCJGx/JPH2ikodlJG/fENdix3Kk23ypmIEvp2HXCEzqBE/Ssg3ZrOvySXzV2h/5
0omrq/tCy2KFtmGlvFUvMOze8fMA62HWTotk0BKq+ad8bYiGepz43ZxwOBZARgWL/7kGds7fA3Ub
YshTq8P1Z+rYDH76grBn0RJpymhMdHd7dLW8osiKuaBy/gmREAXOFUpUjBdR9v9JB01Mw+9BYfzl
46+irQsCtO3rhV+kSCGWzG/8rqILzxXBHnJ8ysux0KD4K52orKMegdUkvTTdp9p7ATJz/eR+9eNh
UjpXNyDuL7APZM2TkUC/AY+hUsYTNJR9/9IAyWB045+p2cwp6SFYTDmMKIDREJpt0atCIhMeEs3/
iHguSvaKZi5azS5ON/4/gWfeonUJI5W70cjbhZAs1C85XVi1YetjtncIomxvTcJqIUHwPt4lawoG
fUPNv6fuvyAvpUhWWaH+cf0sq8HDK7Zgwp1waxZdb8coK8E1bAECw+1PdZB1wIO/LPG2oajm0iz/
ZnAksqJo6ntxUNDBVyeq8JoDU8o1y7vmi1BYb2m6+YLyY2rIHmagMNEgynYFMLWIEcNnaBJqi4r2
DHmestUzbCqA+uGIFT6nh80ygktRojvZlDDDxPLnYUyfBcyRBnnHTHoJsRqw5ULl0xV5Nf4/E9SW
XrPkkdGQWHbsxkxq/Hqyzwb0wYvLt1tq2dZvx5mgKDAwZG6x5SA4SGdxhvpO1WRZUnZMSCdn+oWg
DliyB45U/fNtqUDJEIllJblU6wI978wR9YrIqaZIiPIEcoO2uAFkcTXTa8HpJOLwSmZkmCmG3MK1
x5FM9gHuW0BmW6wGejZxk+cINwThA21uHEztF6tGwJAnXJ/2yymxpxA8/4PS3MQPYZKni6NKtnX9
SoeZzqKqhjH132Kcy2YYp8IQc7q7pBDzRS23HTjD6s3ufupS4Kvgla35Z909FCwohCL2LjTwysVk
Vg3Y7rRpPWDz8K59f5pd94wp2mbtGW1v1bWlgX/+gHyGu2VMa9W51L0yq4vDSD8lnqqvrMpo3vB+
ddvrr1Z/9fWuwkAKmr9sTw1zkb/rtNokOw4HNqeaqXe89wCIgYjJfSKjje2HUOu/M/4e9ImO6ERZ
KC54Qp94Ckkju6Nf6/XXTgee6ApixWqkWh2rYpUSwRepW0S7PeMP2HQrZ/Dynh5Aq3GbUyBw9++c
VAWcUQWZFG2c5HwIkdyZNLFETl008b629FAWWyV74PgfTUDdKO9qteiyT9owQZr+sIzB9micmoe4
l2SXc+rnGiFraHVtXRpuk60WnHGQE+9XMoIk2xQm2Dkq1itQJG9UemS4t78WmhZqniHbThmWOhHq
QzV/PSat1CbdpkLBJBPHP73AiBF7zKWiv4gR5N0hfdkYmzRoTxtSPdl+OLAnNZ3lupoKf6iLCTsM
y02dJkLQZlKkhdULCw2y5gZ8krpjHF6wDFMutdAESe8sYw5p0I9LQKXPRXLzp7NUrkrsQ2nX1EOe
JvE0fag2ugxpkJUOsY0w/Jqq8epKZP+tiRTf8xoiSRP68if+PQyy4G/RfYrQlNKhKr84ipvTotjb
aKjsR9qkp4jnAP9uKlPaGWGUti1CdLMyKbblOgKJi6fNEBFz5TyK7VGwGNl1cQ83UByWUEhyVXLa
1uhI7M7/rhoNZJ22Z3zNcYpOwDAWyDd9BnIX5rkZOoNAfD9z4aOO5zzdwm+q0QwYA78uLXTL7zMS
psR4Zihz1RrLd8HCu6a2Nwp8ydWYQ19MoCX7BgZmbsIh2u/xoLhkKrDNxj8h/N84D2b6+l+Dla0q
KhSm2JPff69g65bJtmLv8/58SI/4dzCOXfyT8vHzuv4PEpihGkRasLn7EcBQjIs78I+x8oQrnnA2
zXtiJeuBQMTF07+h5RivRIJOOHlDfr6VGPaQpiBaKYhiycU0aVPhvpXtjX7Y75IF6+iZy8/70zrF
gP7LvS/zdWDrZXKRGDDLGxSXafgwFhUlXfpg1cdWjVpLCS5gbxLzdcU0R/7q5fhPRS702sc25+cJ
9OCMvXdeeqRYgRRAaDCAs+GMqbEWEq0MURbX7FuC20M8hRnbNw6uGmrJ65jxUodzwPu6l/eJNG1N
oLq4FbOpIS7+9AE7K9HWJpGkNhZxeHY9LlCpq7eAUFGIKotSb1TMFatkH5GztfUa4kbszCNkWj/c
LalQSd5W2NFaLf++Ep/dx2qm988C3e02561jKOgAbOO2rzTsnIutqKjIl4pBZBbUtGp6zTo2h5B7
nVZKjymCsumvsOnN7PwzYwPZlBmBMM/H1kg48GrEBfwoF664IPXo6RRo2H4oCAVWBWFJCMnJFcy8
q6E4IVt/1oLMKucief3cODf4q2zcMWxpVWMtH2HBDmTKxOBoQ90xWw92UADkFxnM1gehp5G7ivxv
hwNc5EVEl//lAKGagoDHLHWVe6z+QmNGqJNEsHlP0kTJZb0jE8KOvm/H2Gx82MFiAAESPDAHcQCL
OKKh6g1oPybnIIFO3kOihWj0VKrzKaMPCMwRbyyGzuThqvC4p6OZ++ToDuoHVgXXvrJJJKcNJ4Ob
y4KKwndO7TLm3G6TPjp3Wz0wiPsuFbvuTiLjkfKO2x+7NAeixf5KD920OdMfYl/0jfZLve2Ew0Cv
sJEOknNhXMDGwTOWEw7FP7aIkLZsKhwjmxtRn0v+WMLA4Fi+ml+Q1QgIgs/TLEMNt9yqQxyE8lK4
Gu8W6TyZeQ0p1/adC9zHmDnN39ObrZfCl5fPgq+1QjPi40Py83jJZZEM3GMBLmQWDp184JhJXOt0
qB3fPXP8+faUUPjZWt15NpgpAvPuT1T8TzSo9EUTixKJZQ+Es8z7GAsXju2/u8eHE4JuGDpDayDu
yUlWfIoHtlTpngM8sRBC25dktfSFfd+cSpkL2kLtxj2jvxG+9or59fsTfpaXqQ1k3tnyf9d9nHWb
CCtUL2s49MIwwnFo1FJ3GTc2k6oVh2RhR+gi13EKxSRJTgOSv9C8PUSYZ3ikbbMXdYCwv9JPh24q
cHtPpBPQMSDm7wgoD7O+7FM16LaLdmv4f0W86E/SFBBWLzWHOlXwba1BuUv39lhLZBxPfYe2FW/F
fNi3frHnOoxgJB3kjSCp85cJ5fdKgD9Efl7nBmEXTDJZPn6GEp6TI00HXpF7Im+VKFzfgkk/lc+Q
rIYwDpTYyq/n5Lvvb8lGmVLqCNV+GYQyp+Zf9wj0zsbrXcW8/pav+qCOlTzpKxqt2Csxa2Lqm9J4
0yAVid0H85Y9n+gS5loN2/C3alhuy06YHZunMAsw3z1McG0MkPjJW9VoY/jmeajkbTMFTq+cSt4K
PJvzLv5K+lUBzCKiS8anQBHiYnVnPMPxnLrWZMiYJdtosB7CiTMuEWNxlSvgrcWzkvBahYjZh5AA
dJJJrJSFD2Yh16SBSlSCL3jGDbP/PdwvrbHbF4MkX7TZk+O5ULh6cJuQ65G3o51eMFchu4Mrv/bX
NS9/kbHt469koVRODn80dfGS8t4eVDUqZqzSPITAfIROK+2HOKYO4IiSuwlImDORSAurRortbZL4
sQDCJZeA3C3HyIV/hA8Q8DgTFsa8Z+gROfa9y5BJxCceTHwdviFJGYDnFCBp6Vgf8bz36lIrl51m
tUk6DD5wyMSYXJO+/9oHutfJRfw74FcRVwdfLdX+iu5S1WqGhRrGZT2/GbAnRIjdYhIL+Q6WGIOC
9kAwdpYjN0y89XZXeNhbV+X3JtQqJLjhbzGW1iqLxc8XaD+4E1Wjr2bf/nsX/46oqIFfhIyJz8lw
YdqQ6J9k7sk3XfVz7bZG1tChUhr2pSMgq0ax3JYmKrBRjdwgM0YgRtk4mWpXj8cr5/tyAPdCk1+v
ZsfXKtm+twnFgrYV5/x7D968X+t54z+d68WQo550yrDGtq9YktfWpzkHy5u9VLD8xgYIRitNP5HA
cd7axbzp+31uiwJMRkHc6mOSxYgK23jX3+5V8ZSISPjdczXs4lC9T2Ws3ynC9UN4D8ksDWRDSRIx
BqWWeDugYsMgxUssvWjGxxCGESwpnSmMi1gLB10LSmBIvnKPKCGU2+ynISAM7xJGflpmH72q4b/L
A/3iDuSaisjSMULoUcWErk0E92ZzNDH6eInIz1bi5xAx7/jXmD6sUkynWSEBAz6XCjdN6qpSmDgO
naAu3hBSxKZP9LE5t+k3E+iRdstP6OXWLuLpYKFPOe/SuonE8ag+APxTEuLkos4Lc28AmWphxukv
kB/u4xScv6e3mvErmuuTnmVdpSHWt+MR3fS9Ors4TvpYyQnu3yVUcgi/EJp138WFe1M5bjsEF1e5
MTH80Nm+4pXSYq4u7c1tl3MvMSLRXhGEsk9t3eWS67+z45Lami5MIveNqRshB4lIqfWFB8iBeTW3
ELqmGUUnSW0c+wr9m/DybcYG/wJ7g3O5xOf7rqJWi/MescaCzqnC+/Xn6dNhHy0dwXpKExy0iTPx
HWftRc8mtpu/tw5vbIZ7CwGQc3GKpNwhbAqjBCmdFo/gkIFk/wDH9GT0RRuWpOndDz6v9mKpRWMj
PlLsIygHuMgjZaudJ5yOVC9rkaRE079Vpi6mbz+iZx2J70qZ/Kdsdv9KxeC26LZEjNIReoi4TCG0
vup5QNbgpFZkWf+FtYmQKdlwE/ZejZve9qKdbELeSebM0dg0GbjKNE1vhK6W/B/n8hhMrAiLNHbm
jB45VXOKwcK6002YFJsHRmPoXoUPz2rMeOkHWOCK2MWnWYlYk3uWpmRCVXfkjb/Eo198n1XffVRO
PHLLvy+cDmAMzogci27rtzNIym5I+GvonHh1OOMzrXJYSumkHU4XFyeN9XmeOnFsGogt3XuqQC0p
stxlIO9RB3mUAhvvjuTnK5XMvWq73sGjgPciJx81vSw+mVbsqANOQyAR2zTrBb7unvhDo/gsFBe3
0DnDTa7wWrjDqXto68yQS/rKjEVLnKbv6wRb9OrZe2kpeWDOrG2aXJdSb+278BVnoPJ2b1zzrZh5
ZJMdszbQb0L7XoE92hvfazq8KIaqNQP/yKyO6GmCWHgY3u3Exu3TTWz3r3LxxZq0WVhU29X2ekD5
W2y8UXTIjJAtYLlF2dCwbQ6OHNIh3AbPAMvDAM7xKorr9TEhDZBKkXbMEhyOvjAbElQ8qAQSIJSL
G06bsE5cxysnj6dXBUEjsyg3FUXH1UCK6bd8JvAsUZAxgAJNt4zMTdYj0YMPM79tklun29y1bh3S
QPqbUHFVSd+kxJ8p1f1DBJglK8bu13xMvWrY+/CV4ErmghIVJ6cyaO4YvVSZG+WLfUuSp4Ekh0up
5Px+nrvPxITNPiAkAjRtWUTSLK3aOpm5MFPR0G5w8fPM6c1iUkLOTTw95kUqvENfvSsw/B1t4Wpc
kLVUl/9Q8dlXTtq3+JZW+lMqA+DEVjs4/PQVrVfEj/9nzmIul/H1jNkOUcbfoldit8z3fE6XLsA0
RB1pb8u9GmTObJ8ozR+m0sPLbDFh2eh9E8YgyEr5jxQjEdtchTFX8znJgKIRJZ1QoeL4gApNvXOG
9dqhUfACq3htf/xwmGA8UxUfg9to/7XNwzPj8AYPfmBS9VjLWFkvJzYA49ixoDX/yn94d9PO4lIX
790KRwIRCHLkbswv4w8rbZuSpyePNaeMyRMTqfGEGpUrRolkieGZuMBgKH81qhJZdA7D/I/axOTG
Vt72nRLoO1Kb7oDqmw2YF+VlB3DZqHEKc6EVD+jD8v48S7dzd+HVuhuch3kH8VoWN3y/AOCn/WUg
GuhNjl0lGGunJe24yCN4G5kAFUkv7JOUWwfpIzvo2U5oZE3LYw9uLB5vBvlKTsYFS6QEmf51pNzm
npNk0MMPSFrp/IpEmaT8WctqwxVJuOhThIpWz0Iwyy0RJfIwNqCZPemWRhmtCxnOBJkfHMtwOVJ/
ktmIOf8VoSAVWhyvl1LdgLJpl09AVGaRlTvWWA/2GuipZhEnxGyZFNIL8CpDuqqOyqvoglDeUYhj
FhHetjN+nJSZeCvV5EHnG2oOuhJSdORbBypiuQRVM7pbrAMrqtJAeojGIzDVPXFhMFcc1uXY8nML
e6gRsxWkwBz7VAXncexov46rYGfkItkfUOwWYRE7fCTDkIF9MKg+6jE5eXssO/LN+EWiD0suJt90
+j/f1ePYk7u6jFJrC4xHTv3NtmO3zfHeLC3f94J890wgTDkymkUHsDMukU3LdS/NGWHX9089Jd9z
GR5AUjlOBTTKZnUWgzLDrp8oTYqWXGg4DFTrP3A0dzQ+S6yC6v9sIgsmirr+CB1UYcaS8p5HvzSg
bFxhEuYHQkMaQSI7hSC9NiCu05nLgMENfXH0fAKijsVzNqxt8F6SmmuzrhiQKTT3SOTlZSSDbwbZ
4GbAN+CVxFw7kEUoLhtZDi8EZuqWGqZvqcV220YdBelsl0HECtgJrjuFnk4D9Q9SehjRqNslx2zn
Due0bDoMu9HZWzoayaxAiyW2/qoWqrQF8uVh/5rK4EYcNFMZKMHFKOzMmBV1/PwQ9nH0GT30mQVu
tlUU4IlA0PJVDe4dpJcyPftK2dnrtmxoGFmXre5knszMhuqm069K5t/fsp3XapckAmthwZ33vSAR
5xuXpm6jU6jBFqMAViaDq4z7ss0sbjp6PSd4OGq5fwxqnjY7jL6FzChk7RTo7x9jv6jdEGufT54W
ECGzN4MEM3o09G6qeAPdIJdBbM02olNjDpz8vjgGsy5p4eX5CxhGgpP32LFXbi2VGewQQMS8Hssk
vpsoI8LRuetcaYqyHRhVLgqVFEYX576i7CI3ZhTHWl4wyyTAquvJ0DVHwIPlOXsmdpogpeayoTD1
86ivQHwPw8s8t6pqiq+6ElsQs03eg6SxUn3Aa3z1JfTroLkPAstuFz4+JxohJz1sw0rhexo0ByzA
rPEMEsm1SUqeI4Wct03E1b0kbQ8mFbv16ldzwaA7NUlxx43LtkWZ9iAXawamqo8I5uu8EWnV/HiJ
N0UVDEBlSAggcDZDE9QPGdrxWUvwwwmcfBCx0VFZb7YZWbuqjGH5mgSNqz4b+wE5RJV6X3jH1Alg
zGcQUwUZs9Sn6VpUuVp8bUr/8ZbQh1jpU6IjMEZ9Vy73gJJdokL/+mxu8AeQoXpPxNW+L9SvGEIX
dKCT5gXCgN+pZMdm5RGPy0LZnvRddfDc1b+X6MAle4gg/ROO60nM0gk6ycIpjpq69hJBX+ZgFuY8
ryLr1txgtcvLkoPW8Czb0VLY562n8ZltPmye/nSSuWT8AqVKoamtV5QX5Pu00kbhRlozZaH4vtjD
ncyDsf6leGjTLc1fobJYI8s52XMOy06opJFPuTKV88rW9CKOxyOfD22P7cdU5JDxEkrY8kIPqDyc
C5Q4bJk0UI1LMzelGqG0vJXStfZmvZx3UXBbXUWNFUe1L0uVbbO6CXW5PQH4t40aTFfEPvfmXRNB
MWMks0lWDoWdyhxhlHs1VsU+UnNGf9Q5ztaT02T2K6p/4dHgx/20ka1QbQQd+7DJUd+IC3NonGPm
XBlDOBQLvIiBa98QT/OMisCop2K76VF6aHHG96sSReYp222qKyluP1JhLg9XHoS8Nspl1bquptkS
DLnkVtzoPWFDlz8Qh3HM7/M9NedoxA1CBNatkWBLdmEs6oey2UwLPdjSnM/SFWJoo511Lb5Ju9bF
gSOCUu8Rs1lXqlHZuGretd1qR+1BLrFPXbb7mubRrNsHXgE24tWYxKiQe1YN/1Bn99lbQ9Or56T2
gJJGQMXUu7LUBAkXs83YY4slyTAfoD1ZZdIMtE6ZHoToqSzHCZ8yCDKxXsZl07fvblMbp1y7omOh
gdo1lGnGEmiBBcFTZ0v8KNAydBrZe/akCMR2DNTzh27pijicjx11DuY6KtmWLdJoNORKeWUlSIVN
ZIiCZaytJe7mtSaJv//uEXUG1ZyL8VVAvF51pylwibW9ZaO37KC8Rls1Ywqm6pJ79MIkdBa2Ee0B
yd4Rxd8bIaL5w0G9EJNmcfZXiOhHkzMozCJVLr9ahZAXkHGMLI/i41W/UhCEmBhZLR46L2mEsaKE
hfPlRuPt1a3msy0RdDch7NtyEJb+QVBBFvBKrAZiX73pzWV/CFc7teeT1IL7Ov98TQ3eCGWVm+1+
4SDTlf353LmjFOb6j1xq1cFqRoR0AeaA1QwmZkHOux9njMks5XeuN2H1VHnWys7N+L+5y1/eEs09
LUUohLCSKfphcEwYzI3D576SJC6XV63vEGrX32+LUjeTAJk3zSiciWhBmTxtZwE8NUkHt5f23xtH
EUbd/yTVBuT43+pyG14BI8Rx/CbNDrXxr+w9dRVsSHhbfkmIVSA89JAX1wkPAuI8xf2yGP7PzBqC
HqmBrNaiUy0pUWbl8sBUy8eGrhZRbQuGF/3UA6MOBitQYAuqesTnW6++hmOV73CH74tzys8EyCCk
9gP3zqni3INqZGGg3ZoxWDGUirvIiLU1AAvdtbdLXDc+tFY96TXmwLvELrdfd6daM9G63ZpNxOi2
SAfKTKlLebH+92yCWa0wciywsNEkiboCKyI0fjCpZ7IB6zYdEVswoW26OodAawtsWxt4rwyBSgve
9U+2nxMeZ7xzHcdQHTFZYl1Rw1O89k9hsllVYm6sLGB6Sb0ob7bbnJruXHlQSI5p8HV5Cs+YlV4X
CQ+9E4yzPGxSF5uuwjRdxRrgyCCBXnPB0Y5IWQSGeV7k4wYuoaMmfEHKbZupvdcVKcVhqJzRSVYp
PUJ32bzPT5l7sgvIv2V0TI5uveLPjgqAWkuGONHoQl6QAGt3W4T0k2YShwxCoXrS/b6vJrYA2Z2P
XJGIIXo5YOPFyMSnYarCZFUYePAMIdAj4UcwXQBOa2d8KmR39rug1dI67mJy7wKrQUSdjVTGY5Kq
Om8ZAHr7NDxK6NI5GjHqhiZEH2N6QqZUVKYMB4anAME8FGyAgje8+M74U3n87En3T44yMBLFM63I
WYzsME5a0AlIvgk8z/yKvsHdS5sn85przNOcm64QCq0RZ9QTLZtChZ+EHNoesxIbW4InyWTkGcVY
lwkavyPP8aL5p/f7orlJLej0gQ1JsT1025ixHva0UAvSEHQQqBfhqDEPTwZitps9j/FxUvi4jUPe
IqQtQiPPaqzk8vsvgURVFDzvKWDqsOpQrg6e2RQ9hWWWbohZot620dnDB8UJnxybA8LZ2LHm70jc
e8FXDrA1K/KwVK5B/nPt2LH4cTzEPAXRrn9VBL+Q2rQedEyOfSk1HwZ6PPErEjLUjtWfLtL+2fEL
0dEZnbMw7oY0vkuDZMGtCBdBJpBTSqFjs8j7ZiooAd/wT27+4tBfLMtRic3REvjS8zi/KXTl5z/0
/r8vU8SFg7WBdnxwmadrZYdNGaJ1VD2uOyncovUz0F+HLfi7RpKAbbZYRQi2t5wwp+C7UhbAUX7R
i2pnwLIPtG1w9D/2NpwXdO1x7xxrzLZzDDTjfT/L8ODx4nmU+nyT7ENJMtRWQ7S4W0xX6v1EIbV/
4X6sb1XEZnXTr1ekjBIPDqjqBxsTuwkWy/Au/ga/GdgxK43djnb/1sGgQPeiHRLJsajmKAGzfdhc
zGDxcNOOaZ3kQQIjW6p5TCf7BRQ0bdSGHS8K7sNAv7+y3RyghNo/bByksbRZJhXS+5I9rks8zA7D
xQNk9tliPiuRgy5pHyVjrWgj8qVNHvHm7y3Lt4fXrilh2nUmeNjmYinjiNH+mjnke+ZFqSLk8gzw
GWyqPzv1//A2nvQk7Dk9ul81OUa8KecHkpEaJrvXPWKZlNVFmmQiPs0RPKg40xJi6KxPeKNzs2fe
yc5nI57qqeQXdHLz89m3WKNFQb9OFZeARaI/2hJT8UbawVh71Dyp+uy0bh8sbg8+4eQDTgBzQCOv
kO3UDo07bGtFZpSUAurUmjpEn0rEj/SZTWCMlG8mabLxCUV15zg3SMeSQcXA0u8Zl8LaZnCv+bnq
ETq+wtW4q9c6GFREWUJ4HHmz+TaTSU1fXlo6iwJ+aKSDz7KYb9zMi65mME48o6hBvJp9Qjf4TEEo
4xjGRI4l8EVZPwC3QaI7xRcZIKy5/ImYUo4am9S2cX7RBUjrkP+N17KNURpSXsfWlZPKIyipgDpr
RbEMFlY4QN5XLmIOYu+XSLH2cS2C52p9B7NZ+lY8kFUVTykXlUAMozORG+9UZ9sQ3mBzpVQE2N1t
aXtYsbPBs19s2bJSgrg/wROdnFeRUVxLZu+/Ng3QLNL7eoiXlgPjGuYOUUkcxGp6Xadjxxc38cA1
t2CdGunpv3cHbbX5ETTEYRv8Ckc9gQqGtzvy6h0tQs0ETavKmhL2Ko7kCU02Mblsl5sqqNPF4iX6
C+p5q2o7gcZbG4wfJEXJOn3Bct/ladl+KAMlKIEsikMXj8QxaV9olSm6h4WpH8/gndbfI5JDMVtA
rP8tToKgvdBhD4lpyqH9sGuY8yn1FH6OVvOv0BXpb1fJckF6iP9yvK4SD+d2FXfZgf4ajFfNhQor
vmsqZAKIglffY+oVJM2DXK5D30x+bmY1ZIC50iw78ZesC+H6l+1n34sevbUCtWr/FJpQ9l/FM0B9
A6wpcs1paIfQV6TG+uRtdBdgVyD5zXewP2RsE4rBSmoI0zxtiD3YX6YLVdcqRthbP8jzIHkTcDi9
s0p59IoEOOpUUrPc1m31sRsgw+7YU7HiZS6BIt65PDMXVfBrXgnKnC5+27x1yM/9wTaagdWEFOBq
Yf8tYjPD0dWEN7ZJIycZsN5D1kfW0t6dYEQLBljePTioVsXCuSLTEASEbH1wsqLPZeNPQ8SBHfOq
s1laca8ufvxQmWTaiSniHSanz7dLPrQx3cF5iRCuqHHgXS8MpVFBQPNKz//TwDAW3SOK3GegZy0v
CFy0cwpVT9l25azfP9gK2mnxG/0Ajq3Cvij++lPVOSVwgTDj4T0nk+FTO+OZfu5KiNY/LzDx36I/
eoefW0zwEzUWGHzcBoli833ljs8Xdp0snv0tjKf+n6hIa35eWe7c2n3YnYuXS2VqSHem5r3TSony
BMKVPv0Br8SdeA6JvW2/6jPbunDiA7G/33TfVq5OIijkn6fRRY4WoofYvEK1T15oKDZlKpPn7LIX
80vLJTvhglZbMDLfX65jl97wydd1iip1DuVi8gB9DdHBjLejeac4hecQXfyPAN9dnSAs9H8EQDV9
mQ5ey2HM29mOhoqg2gL3oqBDZUf8DefYeb25Xtzli6VhtSUF6W1Fs55O3paXSRfI2+XPZXP2wLri
C8fsPYKokO+bilqoCXlpBuWe7PlYHI3s3yBCLoYg/HrFndjARyJsfeIYf6JPiNbHKE8hVIpy5E6S
U7hXKrCrALU+flwflHz+FRp5SVZmbMWnarGdLVP0yVWUYJLXdxnAgDINBIxe6x+faekH3JjkCx7T
52HtAo/uBus0hIsT2F/pwkH/CiQiUgKCvhsgo8+xO2WiR9NaQJSjeFvqnxCg5kj8NyZ5P902XCM/
7rzAdoNG9Y1J3PJpsnvKB3Y2MubUKhIEHHbdAfZ0rpA0viIXyDHxMvZA6ZRzPfuK0yp3f+QJ4Sii
qHc90ue7BHCPZmGP+9JX0+/Ncmcr8mS9dIvWBMy5BLIJbP5ZoBsEBLWCmGVbaUFeYrmIUohqbs3p
8gu8rZd6PmcBJJ9/l74Jm7HuzOGdOYMf4ksSCTy2jvlvmWAV4rm5tPjEeperQupxhNMv48cKvPQj
NHVAZTx54apRT0VvV0xf5Kj4ePYvBoNLt5U2vTej/yvu2xqoxmCPSW+npkKLmXwKCF3TXOw2c2WV
0jp3nBg7+7RDtlRwJmy12ohugUvcr+xg7r1rAUd6zMq7s8y7jTE8XAkCarByijIiYfFjw2RbkQg5
EZVO5+h2cHx8oA5uZltWtUq7/+itLlSmhak1yj+aqmD62v91ZL60E/gYA3CSVtmNQGeOypxZ0yzx
P/5RRIqMQqZVPTH1NnPpQebqxtJKk8YMTjPuIo8yLaTsw56caRqriQjClGTbd8DvGxey+8Up+5O4
vmP6HXt820rtlB7ujNLoQzASnTBoem9nN4ZCUL7YOlR56ChHcbpOCpAf+aM12cHny6i6kJdFSBKj
sjy0lhctQmbqvUPpJe5h3ClA9AwcarkUrBbuECZCVix7ZZoAcb6MNsr0eljLwSHj7xcsEQCBUKc7
4Thl13qKrRt3JEVf72wQ7KTNW3nBifac7dUpTsbfEjXPjkdiAG+JDJO+xcM90ZDx1sML5Rq+ykKD
ZCoeKyNLHVPfrnv5qkInvdn4ycEqhzE25UR6zvSyKlxv5wAfPXQiO0a7tabvprTdCfLbVsEeTXXY
PV5WYcxBrNGVjT/zHOv/NwtaVE1KYnHybKT5LqBvZ+kHhdP7uIrHgx7ca6O9RUP1i7E8ib7rvFVO
TqqFRDKUI2vDwsAwjXgYRLhppcrK/lWFqb/Z2P3TDaItuWacm9/GHTbSXXMbpXkd7Or5BHafPd6J
fVJgSdvhVmQjfMA7CYH8K5t4BvEH6elV0zI9mqxiLvPX+6ElsZDaCdB9Zn9AVS0aaGcVyOrAoopB
bW6TjKhlezTynxUs7+7SCPmwspUNnDHOomUPNnqDtoa3hIv/jsuB14n9EBMDSb1ZM4ebvmpvgHTU
sBi35aidEF8nw160yx3hYNZ5vVptU6j/r8AsYjKdv9wudLpMJ4n6MqsGYc+/1IRruGFkEfwuw36T
Q4Sp8H+PmQ1LYcb33cj37itCf8EDbeDKkLRzWDI71Om0d4B7CksF+jAxMAHC4ic7KzSm7Mqx/UwR
gr7nS2GLbD5TUbUPOc5kZO7FfA3A7AWjx74D65HgjmL1J04WAWD8Ut0UnqVt57bVxex5RH3pmsPR
9xiDAyGDm+dCGTKpdhzIC+RFQbdMYdi2w2YdXvZAU1Tbm7m4Xgp/n6c/AaWNFrUdpKsotEMsBFGO
3vVSTtzLlF3Rm6wh2wncZzwyvWL+PBpCzXgJPlECkXTc1JAkjJXd6iuNr0po6aRciwbr/VRxAXEa
9LFkNAe/FzUVWA+x730sk4LewEsJQJqI8kVFXRTH6B9FX3kmzIy4T12CVaBKqNh3IAjFvN8BEgIY
BgleuuJSzsZtTUkvxeZdR6ubLoYbHdUOkRuW/xQmtr5B+Fh3hrQC8ALW3OBEIgY3MC9HQucE/o5I
8MRo69DEsrGU2eVPwzqUjfiq62FZxEvY8eIWHRcyt+tMyDiRQsxHmcrLtav+CfrfhVOXU8M/Zba+
ZyymFtB5xRjxTfDLRGg4UVwh8lQDoXMB/+XexXJxWiWnwDqxYk+6X4q7yR8kVGbjS8t2mU+NL6u6
EsY7sP2YJjmWFvFSGOy1IFyslq5/69HOoQy/C+X1YTPeavEdzVKt1BjRw/tZoJn3NIH4V7R801qi
rICpfITA1VYb3ljAggpJwvTg+8M3G56niqaHVPtmKEv4ocwBLqqFCwOReF2U9GlBhm5a9N+ZfCNI
pubfjOel4+jPI9NUTa5rGXQBAFZ1Z7zZ4qEyLvklCKvwqEpLR7lfgye3Abt6C6ebRyKEMcc+a0V3
sPFLuMK3+rmZCrxmymwpdA4eM6Ak6JzoML3fbpT+VNgvo+6sSGYFK24TpsESG6rQwIlmkzB50tGZ
DEVzYAfizl6HXR6dLd4I4sJ7Sd96TKac4MoS/BI2PJRYGGMWBadMcpC9rKianvGKlxdyPDMKIsZr
CTsYo2QMrxwx1lFSocGLRTyXvOvlGcmR6ZXmf9b9VU/ddpXExw4noC4xudjFBYX1DD5bCYGaineq
kkDsK+zBsXzjdotUGWYGjBtxwCPgBnmoNBZz/C/9M9CzCFqmmVDSwBtvma9dzb3ezlc8kUzR8I1C
eQB/yqwmWf3sZzYa+KhOm/oPfF1uVyCyWTff3HKWzS3RthE7YdS5S+PkARnE3y3dEWBvACXxAaof
TWmXcLLSN6f+C6zfI1hLxOLyZNV7/CEGdZ6fXDrf6B0SDjccRTW27Viz9xgoGNtaH+7+UW5TUfIa
l37AZunPeZY92nWRYKBGeyG4W927JOogjwc3aC0Ysu/NMXso5NLOHuobNJvsSrJbJ8jvhpaX/UJT
m77UWNopGdrj0Hi5wwD/5P+qyASvTuOthBKytHs35V5zRHjg7Hi2sKc7NdY6NiYORSHeOOiau4vX
aj9nfig11XwJaVLa2RCxfmnjR6cwwtXixqk+y6IwenG7FmNDBSvrqjndBjTmghxgHLcd7JuaE1jr
Ubyire5PvKrovSImrLVZPfSj1GlO+eHhYeA0DKKKQL32DZ3EQ9hFoxDpwpyVAk8OFyPyqJpTta4I
8r0n9gGjyETK/jCBk9olKKJQdgNFXtx+PtBl60n89MICSnnfhPtsgwWpIFmQuDOJ4mPWiL6GMpYy
cqyIFa4WeOrS9E1l8Dm5XRLz54dmT06zjx6gsy5y8Dx21l7mxum3Pz8g067TtF8RIetjzykUpo1v
owKJdQzOYy4e5hjKaYSON9hFr1LZ/nya5i0QfvNEHtTva1FY/+dpawM4J1RBJyv5iB92cEZwnRiL
w0NPmRZJtLf9Xm+L01j0vE52ZylByldHm0Ac6syFa3xQXJh9pq/N1LC5TI8f3Ihgi862h7c8TlqM
y30fUOWIw5EHRmLDNDcJe6JJksH4p4ZpbyLLMnMMgZs10QUBeA3msewTbvjZcqgn+n7O9XqeuzgT
j5w8fbtV84XtaqbTWPsMRAsd+miQZLTMSOyu6yWZX8BxZI8ukWyXhcxb9PHgSPMCN2YxCMomH5tL
sSy7LUgM7Rvwkpz8bPZ7hu/Ucw69NH3Y2bB02uENuOBEQCA+ubEjRUeMW+c/sn4b6pNlkgOPWGwz
Q5fVxQXnG602ywI5ESbFnDF/fv7fe8okNFcD77NAMlbsKcZhp+ySMrQSYS848nb+lvZ7gBQuVZlN
A+K8GaLU3vZp3vkXP3vAczah/tHTESlZ0b2dC4Li5I3hw5odhSPU4dF1AhMS7PMcmGznnC6ClAUy
EX595VzOxc2H67DlDZWbCo9xrsGpTewuUXbbGKuu55bH2LwRqkhOwyrVFYPQp7n0IaK/AGfAiUwI
lEgfP/5ASQP8ELmLC4glsMr7XkNzsiFvtCKXIEY7bhVamAzkuG3M+vs5NoADuGUpjfR8ikEXIBKL
5I2AN2yZyDxxuL90bWuMXnOktvLiXEMTWSWOBbeBrLOeL1za1GgPGRUSb7MTAiTyz6hH8u8ljGuk
WjJKtCs5SZNyCRFWS9j8ihvEoKTMa0g3sZBiVlGutNjwemHC+WP7R7Ij4F9b/FJeSk2DvYaaoRWY
BQJl8gF3V2TUPz41sE58TSMwbp5AYHLef04gdvgPXB1tA5ChkNRopJ/pDIHiXUJtvXYdnBzp9si+
knAiJAVtkxjLr+f7Zu5bIdF+Zoz+2Alykd6MJIWAfa5EW+OtmGmGTXmNSuibyONH4XSVt10DlwrY
rN1rOmNyucN6k0Z4AnMv9E9YxpTfyUXMSEfy0X+/6p9P509xOTENSXirgBdVLtr6Oz0Y7fnOXBFP
kYcIpxh0FAEb+uTZuJcZd5IbjKtQIgOodKzVTsVSPAjJvW62mwkX7Z12QPGw28GssIjH6hssbhRK
ogsYeaihTUS/hhl9gry8xp4ru0gPyYEWFRkhXNq+glBEJ0oJTqb6srf3/rTXGb+UCaLbKOpJYGIl
/mf54bL5kOx9/3aPo1xCgWSGj73Bw6UURlTX4k/7/+ZmTUEANUAA62vbbAC8u08ORicqKw3+E5ag
gNcERqU8YQbCLqo9efmf76CCNktzrO8R+JA3KiO82T/U+2n9SzyDsnDE4WsPHBnYaxpZ7s1riVF5
x9YVYqc/eusNNDMtrPO9DM+ZyFnN6dj/Dfc3CE/k+1EaxfcyFWAJGzaGxQRVlYm0sQQOPwXXiVGW
njUtGWkZfDjIMPz/xSBd3lPf/46OPTr+p+6xGBnC5dZZDd87xTlVe3CKCvvEw27t13QYlM/NNcM3
YuwkYJ0vuGWv6saEHoij+zlVS4B7bIl5BLeUxwq8B+X3VRCtUeVJ4Y4l37a20bAWQBrr1C8S7wDR
1sp4wWDfQdCybr0+79QS1qJmTWAFZeAPoFdygGCZg9Ppq3mBB4NKNKVZzehwk1zh1l0JucqPyxZw
toMe/bdSd4GBs8QzvgdX70ps5hsfUYZZxl9fadZnHdPh2Y2ybAUg+JRPLk5oYrcUHu3wUyDIwbc7
GAQVleqjdD9xcggD8ExRw9Y1KY/pkv+/E6lmal5vh9WkPbtwgyQbqlsd/3+2siGgxgGqZeGOLLwE
OZ8CuFKti8fs9/WJIL3ilzIbchEUJvOA4dpLnMWP7Nezr3DxKshMOX0PERb5FBS1nB6dssjVZ42w
eGWngx0U6opzAC+u2N8qkyZWP41CIzKX/wruK9mmU8y8/09rWOV2Cv7Xxfoy0RG9oFpfVFkpz7hG
yGi3A13965qNM2DD4+Sr2Iz4eOEY9/KIJHGwExJZsXhIB12q4HJvIZXvr7HqQBEG9Mfox7/cmIvA
cmYSYQI927LSo/EghXoojc3BQWOqZX/HSLq6PVUShSFxW2TvgsSGPcQRrAXFMZfaPZOER0EWhxNP
d0w3R6nqeSuXpBiNo1hIAAwH4ap9q5R26UesWNzAtMsms+/kZ5W7LsvFNkBAxiYXPIey746axjJX
OqWLA95Bdeh8z1yNvFXq0qFV4GOqE/gc5qJTjJl0ifm+6hCyY/EjLRVumyu3WWaUTJJyX151gh03
0CDVJdxWW+BBzbYEMX7hl2TCztmwCFufO5UNMJJGd5RxT0Xvz15IDeOVXeQZkCb5wg+dIpDK0I6J
HQerTVu582F2y9tTe0jYgyAvQy0TlnbVkosTJB2DGQf2WyOILXcW7ZU8GNpZ19LfDJg3/Q9e96Ea
sYWjwCDx9aOYyY78FUqr7ko8yieGCMwdl2ystV9AoVEzO2ggbwnV9fHBsbaXBXCgCXOzp8WKyY0v
oDx2Y+CpiZsImZKtIErGyprLndXI5KlPVhIwYkyf/MSTvZzKkF5Fi7IHOt8n7HiK5++ZAQ65dVFD
XaYp69xda3UCbBC/JW4zOViLK9Zf/kL1bz+neJmQf0BfSh+M0G+rDoYYLZoy2ZB7e6cjK6cOOuVM
GpW7/X8SfUw/dij/pEpL0mvRloj2Key8Iu3yByPJ2epSkm7hS7Ax/ZXkxuYChqlFEItgUqWCv/i5
I5sk09E2m2ORXiHqKAFjFeKOZTxfmXoj1JssWhsrNOsW81dkYazFtA5nyH2nD3tD5oosFp5jF31n
L9Kq89iVQYCLaDNwYZdzyB/BcQ1no6npoVwQV5FrQY5U2tohVsaMrhuS59bl5ufu4f6gH9TLAicc
EinY869LemD6a8FxEwHlqBa+GkwUVygky6i1NwsU0rE6XH/LPY2dAhYBYxvx7ReZmM4S6WRyxdLa
1TlXnxW7Pf5dlhKe8oqyIxiPEjZRoJm3IjzBt5gUwgjYLMCLySvw6PKPusiegZKAH5tZaWgamNfN
uBIeYtnrNUKp+i79UzLfE+wp2fDAUzmsZKfGO3Kmv2Eh5fWv15RHjW0EyDSm9VM65YpGPdSkBw/+
+8afNiYVBxO40cyxWdwuluFtwBS7WLs1k2xb9GmRTiCafkgTpdr7nNCLGZnr9GcMZC9Ped5sUX+o
wCfphaswppaiNxcSsJSMdFH7M9hcfGshDdN/cRBQcYjPdBIRY94K3ieEBa0dUTJMQcpGjbF+oMib
nLSWdJgqFeVLlmXMp4j/6vVAda+pewIk+ay7EMlIvrdZNAeWAUy+y2r2n5RoGW0unjlW/XWxhFvJ
H4kzLJuQmaXTcDNPuoFEM8aauOnuR/MqM2YFjSIjy2IBbydA0dJZz/nk+rSLRdU4MXvrXSvftGvr
BBo+wyLTHo5QIhkjKT+K7GnXnPNP6H3k5B/SL9R+yNJyvGkJtK07V6pyMKLqDkdQYc39Vw1ue8uE
bGQCRixxDOMA83SCeQib7cNWSAlC4mlDjzy7ZDrsSEzgNWZTBfu/dHiRlHYJyMmh65tHDKNaM8Gr
18j263CgFhOcARBaD8YOUOOHmyMbOkh59GuVuKmsZzIMmjwysU2keEuQXVLlEvlRtTGyVVc6ZoxE
PjROzbZWSmfxtRxGwXPZgDj30F5l1ljTBPRlnUTQ4VOSKbmTqigPfxmMG1eKUnbbYoMZQzYvh+nw
bn6X0dE8n81ta8lfVkNjFlzqEGeNvV6+D4tczTXAhtXYK9sz3CzlhJ0+Fnv5gC7NruFApg0vNrSO
V7d+zHIEkgb4DwnNWbJIO46V6VsrYBx+swFJ1zz6Zt/guw7g2pxiN8CceZMTem9VXMPrs1hZuEoo
hNKW7vIBSii4L1vQEaqBqiUnKpJm5LtHN8GqpXVv1yRsUEW6N6Jaqy8Vz1hFQ3yhidaLggumvoky
1kiluGkgx/bxQ0hNhoPGMxB4tlnYnnrSRaM80p0MzyFCO/xRA/5IGJiLoIxUlPVKwB/3LXU0SXko
wrC0c+Uuc2GS1FLIZI6PiDTrtFjVYdklYFfxgMKxVfp/QIQZN6GVNiY++7XosIJTQhCySDTIqNuQ
gk8dU6DL1nNCMlL5YpwsXSClW9KrQvxzwopaMpB3d0JZZIaEvIh38jc4zPCUPTbFihfTzxgeqk+r
+ZP2DmroMBTXDeXgiAogbW2kYplo7Baqk0cgourk+6GGr29crPk7aZ4Rws/nvmLYkMTAeAoaY9jN
aZdgMrLEhHgdHCSi0jQ2lG6mx+4RZ3dZtoQyxZWhLjc2TP8Bo6YEbRZqgXncI8NQKml6HBBAbEZa
4twgeX6LUbV5mwkPFV0d0ZjvJnIpyxJX8QkQ6lRh5Oabzcl9s5rfRXyWMS2u29j0fI8aJJA0wYOP
FbXTxFc/8rz/FuN9a7ziJ+k2y5yvPVYmXXdLYyJlYX4guNoJm8uceMYyBX3x64RN70hYXaYyQv4B
z7QS4e65onnDtTD18PlUqH4n8et/hl32P//dX37VQS/guhXEqrS3e8Z2+uYD/r6elU+V3pXzN9Jg
lhbLbqIntQKAUbfZ3X6+m3vkBkWILCPoBD4ija3APpCANCMG7zhbkyRkLKvxXnp1dkuXchp4a1rS
KMd9rnXR3Wt3f1x4OVfMhnXobYOrLfgn32upp7oRsOD0u4w6K67Od8zyj4GPzbT1wI3SR2ZL8qhs
fpi4ctiqM1EQzd9BK+KQotb+wVdGplkyMQ9Btvw2Rtej7UTQKcXWv/YJwr947Lzc/SXkSU+lcTqw
NhhHmfKV7rSlvbzBnbEe2wNtyed70+LccjnYVgd/BwE9xjNtHjzcVtP76GqRYgBWwKt2xE93VU1v
CoWXj75rCqq8N21ly5KtEhHvATSuODTq8usBz/FEJ7X9qxU24Pzlxiq+Q09Dpr68bmq4DbFKbpJJ
avW2e631vYVvg+jWxEx+CDZTVLZc9yLftGQ6yCbllaCAyiotlPOFaumI7BXDgM7tlOVXIpYbM78M
nmwHZbIWiZ/WoiPwpt6ovRC97caGWdiJOFxaEPJvHomW9tdj14MPkIaL/ZtwxWPk+yPIVlHVkaNy
lobIo2E/fg+JmV2tp1ELZtIaN9ZPNbRoC1yDlQ6w2VUeiQoxUvkcD328jvRUhSswyQ9nn/AMAu+J
r+nuo3Txtid+W9EqP3vzmALanmTWzFAEiWXfIClHEE8aSb5wGSzc94Pq8MPJ/kzTYy7yWFCaLhLO
SHDuxv33BgTsv3r/fQMGc7qLIXx5pjNmKXFXRG7L3ER+jxAL+L/VWdMUoN7677ptt7nl8qnnCTGR
BYNpY4lQmIkKN/i3w/dFNkqDPLxFsIAymNIWWAIEx7lGTWFkGIQf3Aab7Pz9IpOrqbdgjrAEt9nP
p2fDqFY0R+wGxqp6P/lWyupZEUi+p7mht8EEiUqa0ycPbuKcwDh60lJ4srWif2g16a7mZvxzX6iu
mNRvJ7r9mSJvvF23ijmTvg0fy1ekb2BCECvR7SP4UAcpJLsm17qaM2J+0ODEta2KtXfgiSOCuVhQ
QGh21Cxa85lzbIjXHCCFGtHfo9wcJZ4XxoMRhfNl4iN9Qo8SYrK+iqMsSnVZ579UfwCWuijAFWFK
QuZXPkJRHfjUCWZ7vl08HuRT7mtlazV6NIZlX5QVSL16iarr6kmJs+Heulxy5DdEPlau/g1Ir/V8
lD5orusegTD41CsyDPKM4Q8B2hkvkAjtHqItFZ8GvvwhFJofgfEz+5tjzVx2O4J8z/T2eT0uC6mr
bZL8BPjpqxX/2lhoTCmGV/AxK+4dSOXMr5+3UZWyZ6Ktt6RGWKObp2Fe3c3Cyg1scJ6930qKdWZP
kPB89ZLTJh5PibcAAOMrJp0lSi60kaxe4dFu5reYgM3qk+aB+WAZHx3vrxsnhFZxLgoMSpKPx0HT
mRUUXVWIn3IJmdXSxsBUVpHmPN+L1Rv/Otal7+gyvCchq64R9lUdmyy43nYN7kLO+s2aKpSOSPnu
O5EMumUuiS7nGbjGkyZQI0lCTxECC56UefIh4XVm7XqjS7nPfz7D4kuZsXq1OYq3/DP8u4r2ust2
Oyt4/4VRTZeQ4n2E6OuESXSGdrJ+wR6YfolnaLOPPd7Q1eP+XKuo1wnge4czYatvOp6qQPbe/AYD
DsgTY1Z1c/JNC0TcWNhNg6QOCJ/gneKp4cMlmPMEERQzI09vLwB5mlKAPIciVJJKiSySfx4+2dZN
Zpw8eqZsPOQ7qVO9D/b6G1U46AnDUDX9mlmAEzgEsdzUfySWc6rGYgT5+1wRS4dQbG0ApSzpqC0m
n7LQg0Wk3oP4CTF4K1Gys5Yvu9ljNFuPp4EuEInlQkr1qx9TKriPIg5MK7iVytXYqtXxF1XltFDv
3e+nuln5gln0xYbcQmA83ORroQNEqzLC/fSj8aYD3LrzNWyMKrvQ26UUn2a92ZxDYBauuus+R/FH
uY+ydBZtQ9PFnrL6RztWeLfwHx3haeHDfxrydN5abkTkOR83a/cTvPGsThh1uksrEfX0642UCCdN
f0sjGAbY7c0ztnDlBRefiwYxy9vNuHZrYa3U1HqxaKHyGto/eiM8PDzSXHDoV+Gl0ExN1d9Lhzer
Ss3MFLDf/TGQ+k3rR8tNQjazEmNmBfWycnINkqQD7KXvXuQP6J2vvGmlpbNNu4wiEGQkX0u9xm/6
UaekgtV73iyrKX19SjGj/pNkBK2A9OZ0W7HM/0zgE6CSoll87jFXTZBZbIh2GggB5dx0ofF3BLIf
0Kx0qVax5fWMWL+5peKdWLXyKLtPIV0fm5IkK4HKhIr4Bsea4Jnd8TnwBwpkdAVBplWC96cVxiD/
haf7BAmO/gWepSSdVn4vyUgCcnsflar83tCkPza1ujR2nNxUKXF3bZCMK16qY9cmWxYWloW/3sVW
z0tPUFtYg/IyJXnZY6Q0YzZgVXgA5wctNAPRQ9HWIpSe1frihxBt0lASyjNsgHj0dgzmegxkvxdz
4Mc9xAY0afKg6/78e0iizH2LvoSO1Z+rIdvKZ/f5iEUzWvKnF5FSYmrqiXTJbTFaJ6LnHWmrrx2F
tO4RXC5BSudkR+sZTyOZh2VevnJpsSLh9ZUUxuuZcvwLU59Uqmr4zgN0GMOeVgnwCLGBnzVQwZSD
a3K9pzfWsvdh02G2Sr5hd55HbMl3wooTb+IIWpijwcPma1gldh3Z1j6aFk97wwjdIPtHqnGTI7T+
/bMRfFyxEcvlHfmyJfi+K9J28z6YPMEqhTMbpklh6OFYvPM2zZ1pnlIdhVa8h7//Q2dZiTHQZOzt
J3QJsJi1uYs75qy+SBCSl6nMld7uCZOZHX3eu3TsKClIC5cE3P44V30qZMKsnmeQkGTsyFM4Dfe8
qSctFDxwWh3zWRk/VeegW7dSshdJg8kjKgMLBDNqVoa1tVPBv+gwe0f4CFRvQWdUIXQ1U7+CYajH
5GEYqHxSh66UAjl3bdVyAi8OlMIAI0wILts+O/kr107qoMwtnWA0SSK7RxCAiu0xpTx9ZnLwGBTY
pDwVjoRnmSBI9kbVQNfWWIMRsepbiYP2KAFnpoAa0Jg8KuxfYNNW+EHDsIWbh1jHgnmRQ2XfcsQw
qFat2zYTLJegsuXs4k6zCniNyoqeqMY05sCzzJuYaVfCwByi9dxXiBYPOSL1qh/BAB0qLBnPSBTy
DkSsRH/mpGw7J+kRVlPsgXxua5wKBewZCkdNTRj+EJJ+HaC4Ep2NqfC9HRO3351ZeuefcK6qBlsr
pE0tD41PU68+LquErRFR4I78636IlJ2p10MMPcxhpd3RQFbfaL+kUJlACejqWNo3kCFy8/l3A03r
BIps6WjQu8MzwFvFOxZqD1M6uSMy/jlxcBTbh8wch0QSkpMW9gHM2RrW1Auu+mWAT8dZ/Xz7swpu
nKL5QfDWDphS4IL6pMmmjsJV7Nl9fem2QxylDGgUDT4Q0bpTl5e5K+3dZMW1L53StdOIWkD+mN4Q
izL9Je3skYl5NNmBkao/r8gRovtwcXqb19z+o32w0gOFt71W/Q7UTrezJfS38y+PhUuEJYh2JXEg
dP9oAidV5ZX459jNgoia69qcQnVkkIL1yp1+MREoDr7+n+AIwHYEfta63LQS4LMpzinucy1RAVQ3
BF9bSxRYh7jvSE4klaS2sXwWVOgQaOgch7MMjixgxkKvNEaZ9fUTmXJji+5TskgF+1Vx+Iz5t1Rt
wXwxYJc9dEe5lCG4c5XOLLoPxa+0dNZH0IKmgEdVAzWNbK/11lwdgkv0gqUh3fDJWo+Ya04TEr8W
UObWZTFYT3JNCsz4Fo83Sg2RMyXlgAhDgYQG22sdOeitg61yKD8bZE76fV9oTktd2/5feToSJIsn
njmshnMyk8QI2pyrAq6JIbwPY87TcIrVv9eoZPUJpbV+YzmoWikMqv/8jn/dJFCxNX1Pw9SXdURX
yNXujTYeHZcTzAZkuIP53yrinOsupqo/2MpNgS5sXU5Ex+Aindyg6DTlklCbo+1KckHhf8IoAMIn
Bg65lAfGDm9OiIiaUvqKUumlzo//81kgABc2YZOfhFtKmZmre60CCyK5fyHlI6CHnB5o3wVibtrT
eVaOl66x4AzVjChhrSMNkjZnKLQA99BwGLMLPt5ZqCf9uluoBMp58VAKOQQM4t/54RoDP/1a8n0z
nyH8Of3uqXQtLk8TmgP8vSgtDsTSQavJO6QYGoFpngZuo/Qc3v1OYsErYDJg17F/6UGFRTBpg+qt
OxKsMs2AFZFrKhLW3affNFrHY33+pPyPzERbyGGUabduIfvusmJJrlPexS3Bs5UAJEC9lzju2B/k
bvHF5pvx03LcCGVUlRv7uKXdsn2c1M10harjJ5Ganzh9R9RTsRhdP/sq+r0VpUxGN14OnkelnszI
/MWvRYemd3TGlU9LfoNyX3pMLSrLW5vJKI29KNDqkfNZcQcTdo2b90dh3i4RzYlMM0I59PgrnxiZ
CE1L0mlKvAAD3sNNfVSXFe1k9Rn7d/Jezi8T0Bu5w9Nesutqd/2qMYHqZerdkBFpZmn/ttJ0E/eq
g+I1m83SvF8M2L13yrS+VHlnBQxV8EYb3674hc80LcDTUtHYTGwHLhLAo9ONJXyQB7sYYyDOx9RC
0aBEEGxcAURb8Uk8aPiZAMJs410x5iTkU/tzDSIa7Yx0OnFBKjCZNfL0SQKfSyT5ssrypOOvC0Vn
5BWtdXiROBJYCOufkg/89Dc92wfD5fcB46C+F9YjB9y8ar0S178hdLxuKTfpXRg1xxELg1126TQ4
cXXw9WFNDfMcHFiCihxTLtKB6OWq/djdi0xBGUwHj4PwpVZZXTSLt/5lI6iq5KUYBhHyBFgwwjpj
tl7nGcD9m7L83dDExkPMYbBVqwFZmSWqCcQQ6IRW6q/Itq/fCbDgb9pXLVc29iz0yDuvbLjr//Dz
M1J7fbMZuaYTzXLoH7IMBY8kbVi4J7SnTLQqIdHGFqQ8pR/j6+90yo2YcrZ+n5LW3rJhGW3iUPqQ
TyQ5d1W0wmwTFUahM8Plsyz2WruT/mT882shvvUMSdOsylhxYZjOW5PipDs+Nz9+acVSB33xNXD5
3JSuJxQ7lzlp3kp7pcVx8g2/FBtnGejbAWP/Z8ccEpn+0bBQaRmtZo4sFAB4sz1+w++Vc66kt9If
Bry/BTQ/FGsOCC1t9PVlB1P8bEqMYFjIgUTTw8FKdTs+HBwlH4m4YkdOL4E+oSK0ljsKDd1kLaUg
KBgs8hPYYFDoSw9E3qOWMKlWlZXI3jAANuPvSSgOa0bQpf9rtXLCH4fXyF/+dLzm8UPd6+WLhMuO
h0XMa4Xq14LdKp/7vjMu/ZsmF6UTCSHEsZW/qPPgayMfykvGwCLPX1oSnrXGsxUJk62L6Fihulb+
ORb/gZ1iGNRkK/nur++cVC02oM7XXsrxsZc+7P3HdAU20XOLQoB6b2MPtL4zob2RoxS40kglDlv4
Het32lszO22L4XGKLAlyJOQYevQc5cfgDJdMdIJdAfNS+6/rZR5KxCgNUVhDvrsEEdYyW5Jqy5AP
pYFOI4CMvdZWHBq4VaHR+Lr+Mew2FcvXpAWnoLfWV9fgY6BH6xZWb6wGW0h597uoUJySA5HtlCnC
T+R9I9IT7NhVG/PVGPsEXfEr308SDY33lhC+K5xr8Jjt0UPMl7WwcCPp2kXkceuQImvlWFOMTJqO
I7+7ME53QUEXSPsV0U/02702uHHfw7ZojLPW7M5DFmTy46aZKsK6S3+5iT3izCEWdbBrwKu+iFbb
fJO/P2FDy1gXkcQbPKo7siw9rX4IVvDd7Io0uGjQl/fa+Vyxin7m/bh//Jvicb19ZbIkRf1OMUl6
liUgx+y4P6pvYYV5tqnnUKlpIx2VboX9O4oZRRrYQ8coT1/VfzLNOOBH1wmZab4y42Kkti/vWbp4
X8zjc3XqrnqPV4aDTx2lAyuDsxCV+xDUThYx2qy32RHmnVFlGSf9ZZyHUuP+/Z0dB+Y8uCv8lG7M
o3C2dI0w82ZTWH1SX/vx1Ql7hhqgnKyBr0R59KE3YMVaX4G1VvOEEyee8kqwamy4Zw3mOOPjrTBP
ptDF8yxmtdOCku+rAmeKhKzLNRmMkMaTnw+hHGJmBVahvczTzseTem70oI+oSPYbXQwL6rcBzXEK
kWuKLgCST3C7OhiefvWX+eeQ0tiCzNcNHSTL2pkEcRDtxGvJMiHcPvHg1kijrbuiokiTiMaP4bMd
71VV4qdbro+K8yPIY3i2+o2bSmNK+7gvshAbAeZhnW5sqvyibzl2bmHrkTxp+aYx9a0odBW/unrv
+cTqnVyOzGQxerUoz8NYqmxC8D70kZjJbCeJrnEgvIPJCLaEueyVVlBU7t+Kly2C5Cp07AcR2dfs
aIhqzFCN4jZyjWxita7lgSKgUMV8KviqLvTDko+P3agvgDdiQyWguSzn8/dc9eKs3rmmDzWpAWJL
prncFNL1SaVKpmWeGIyf/d1hny7Hojcni5K/LACkfIRKUmi/GDJwkQlHKDwi4979mKp+bA80tR/C
cMNA+oUtdHsGuw9BbSC4xhkm+ZWMa+rY3wPxDBjFluLIIf+FEGNAAq3viQiLtdT2BuS5QjaXIX1Z
kkq6Fxp/Va7fNkEliUGqh4LdkbfzrnQOYNel+7FEk54FhNQuYtxkmGQ/wQZN2b/QcBG4PMI77vDd
9sxbo6+5+37zXlamXIItefBjGfOagBxvAJQxoot5GlBRttAyvUaEz2m4iDyIfsPreImc9wqGy+nh
3+lUwOpsaUVhpAjNPIoozJ1KoEBt3OQ9G24xQqwFr686AlsxE6wX6QkxxVGnjNvexWMz1KTRwWNg
tnJgaQQe84lPM8f3RDYeSHX5LpEIF+x1eu3I2/91DZH4C/sDOgoEbDfcdWIUS1LXOOXpkCelrW0M
fEUn4u21TLto8XijFCpc46L63JWE4hansNCKiPYF371bRe2jaarrq0OKManbzkbARgXcncPzV3qE
DQiz/BGxCZIDM2IeiAWEgNqDluXhv16L6V4Fkkur1WhEsQaDhGQKBfeIFq+Rg0EyEu7pXxYOofqs
Mde0NZtOukB/zF5F9ncBOS5lZc6rRX4Uagf0IjonBczWVkbbHKGh617MXOSp/B2L+9IaWEhsZGjo
tGEt8OpZAMzCJJnmbQvXFjgQ1elbOefRzhkQNWbnCDsIcE2OAtjEKGOd440RFBdeaGwkQ0yYeX2V
LVSghCstyk2z7c5fE2IwzuE4ZmmB9FoYhJkNV0lzBQVHnycd3vcgm/UzGkNWeb316zmlXuEEQshF
cG7BQD3rqqb10bmb0W4Y2KNgxb/AUwj+uJSVC3Q307xZHPW80O3rn/foLYiLcATA+709YDzqHDnC
/X/lwxC3th3zmVXw9Ef2Da+LusnaVOu+0oIOJtYnCp4U3bjx9Rm7BSwUK1xT2cSA67VjTrWop2Lu
xPw0aSN9Elh93wvloB94GQC6uwRl2Hx62n8RDwnHmByYP0JwS3gksciH8u0ns/JIpav4UPrNto03
IS5Taqh8rezr8ktKWx//JJh76CN509vrauaMr0D0u0Uq6csppYe/2YvRebckEATGLCMkshbmOlQo
lU7gMPST25qXmbz5bTJzUq95GISHJ05m8eO68VQDO1fgVw/9WVE78dxiCc0rV2jmohpTvDZXjsM/
8Po7EQKAO5xCHYxEAHvjmdkInPn3WNXbkkzhSDRZmA60DGuB9s3k2mSkXZM/xQMrQGwWOERYqYkV
DJYMDxRfF3eRfXEVodhazB+1ltHrP0r7y/01t0Q2dci6fIkkqf+F6KwkWMHALTZIsfpF+VtLyWoe
17wPd2KQt399E63wdjRt0yLkUhwzDa2Mt63nN1ZGocRZUIjqmyYSsAoNyDY4iODBOvsMXjWwPv9V
LXrUYTMGdcur3IKxcymru7HjarV0eSk1o2ODgmvnNic2wGWV0kYTswYVSzuv/HidaTySjzYduJPX
UR2pFjOsUx6OP/VVfk19HZ1MfP65mlqkeyw5i8PljzBWXMqM9rDZ9SW9y/RaWccqELm3uXq+0J5V
kOeNGDxygLXdK5MfmC4rpk8yHSZlGG79EMmAtzWmjggxuTPNrwxoJFbcmF2fq2OC8H9Yp8V7gSvU
7iacejlFaKZQN2/j274rBopskfgMsXUGJcfRxUmTD6Fm32rIvrEQ4ATXEM6Gt9fPXppfsRfrvWPO
S91E1eERor68qU4iHLRICtmdFyTt5d7MUMwbTHpjxGS4MjCKPvfiGJCbRd0VtEseYPbGEZLSGo2r
jR9AavAr40kaNUqPwtXm7Uys2e1xHEAEKA0NpOkYq6/RPIORJwF2CLYM4bm4CKfTDhyFcgsCZnUs
SfS+Be3e2f6syvulWzog1v/s0p6ayErwSBFg/cMao/LdI2G5gQc0Feht4vgaFBQro7UlJMNjqU6R
diRYzif/fyg+TqDS67vSjEq9XSqNF6a7FMetmD5OvxNr1BJ47DpW8s1KGGOz8XG3fmTuVrKbZGF7
kT8MRJDBr9po32Knl9t5Com3g2P8uT/x7ZLAnM6XdbK/bdPMHBlt7jke/7NLw+DKA1u0Bxntn4wo
UczX7nv95muL1uAsfjOl9YvumfBa5SPP2HUIU0Kyl0rbwUB1lO9AR5kfYlLox30fGQE0x2VqcuUC
zVUze/oR2bORIzUoIRNennh8AyTGIeCS94a8T7vbRIWdWaquUnE84ov9LkZogan9xjnJm+m9/UJg
E8A7UA2BKUWhC6rRjzPSnlneo+rR1wb6SdQoY8XRWYNTNK10O/V1rgoSHQPJa6ZhFo4znXkfgq4Q
Lec0eKQH4nXoQGwH02PrFKDnPty/PJXo4RN0B6gFH59WV5eEiAn3dNLowAlQsbUhTW0wtp7qIMXI
VjafRd+RaAN0x2+eBCj7qtYxk8huBvuknaiY+Yj1YDtd8ZGdwVUsMzdgItd2epaSCprVpRdns3cb
lyRISghIYosv8qwF4NvjzPDnteopdYHp/pG9xyVCS6xk/gAleJf2OrKZbU7QJszv/7cHIAy3YfQ5
6wo395++YeRo+QpCkqi+NUHQscLHnUfGnayxx5OtBHQhr1Q/WYkAWpgekUoPXH2x/dhDnjhBgYRu
9gHpoHCDapqDnv8tf/X/yTjwq82+T/uqFcdRXt4QPKTcTG7cS0/B96cNtIYh8Lojr+pbIZUThLzM
iWl8re148rTwtCpnM0Ls99Yew8I0WcLWBLwPTZpGPM87vn27eF1Gg2eoHoXmXXZC03BCPJDGusFZ
7hN+xMsP1w9Xvs5ErfHQ1P/ePpWt2Y7x5pbXz4IaHyocmM1q1ekexFEKBsliPyPeW7DoYZLcj4Tx
+nJUSQazjGfo1Vqwo2ZHJ4oPOwZTQJVs4wbjYLcDOjymVMsuEnr5FseGUV5PrWI5qubQJwirjFhe
lmf4v2nNvkQbi672ixo5EKJ6zLiRGWTMtiB2/z7h1IxOBBwl5XHY3bis1XsNk2eGG4eU9I5kQnjy
ILKa/yYzJOm0mk8q7z+DT/b+S9KLYJoWMmZUbFC1ZbcFSaiWZIxxh/bCYtta5YgWj77vfb9k0VQK
eOR44kr0/QNVNoSrv/ZsFHO8P2G4JsAqUzrB4LFLaau07zGawkaIIwc1STVfgiekDckLZ6p8HhwF
Xm9gf38S8raAPR+EBcE1eSDi+1c0kxHoLtEZDN0+xst5r6KaOCNXN6FQowwhrnMpV/AzsYCyJK2Z
vCdykHVp1ECAyfRlc53aBCtKyDFYGCAIyjXRe8+/46pBwZJVbLnjHClULbxU8nLLukYT0kdE5XAp
qiXixDp6CbsAyIex5lQY0txSsMQBVeGET/MYJlve7pnOaFxNMWcgr0wU30XS6lBRzclBobSJKnTs
ETU2PHXdJTQ7qSKQIlz1Kzefon/bcO5JSlwnef4p2NQcRDgCs79NrHn6GEuZybYWZs3WC6YP96en
dJnY3Dhdbp3b6+NbQnNvuciGI+JVnpDofpgtxWJ01+eePDkuQReN5mlNDDXPVmoZD9LWhnA7ng6n
Uw5D/IGgZx7ifJuJLb/4qnh8gKSIXCJN37k819H4DUxeODyPSHO8cWYM8D/I+51CRhMcg0c7As3l
pXuf7YjZKZb/MNhrvbhzADx4pBmvf0Rwk1WJEQOcPNhAYdWETLlwRmlsdtfaG+Y9w2J40NosfZtn
Vqyyokg2KgI66UzH/9jrI0vQ5zCFa2xqBsa2G1RAGeVSX0qcu2AKR4m3lo0Pm6J7QuAcROQQxZMO
gUp/6TZgJcuQpDuhIOZms1EiZwZnmX7XJcto8SlCclLKSwbvq/2/YpkO7esDqGm9+aYncHbbxmh8
STukWtf3Rk+VyAjVqbfgNq1zVnvCYWRUPO7qvr0If96AGmfocGuMai0/PMLnM84o7tWycyh+Za82
o3DhmuCsCav1mrGu/DzFPpSUxbKky0056WqsQpHD5A6DT3YdmLpseyKQpBQszsTBinhtlnomoc8l
nlkD8xWeerhPPf9eu/80qCRuQPU/R0FSfrJfTVqtkJ82b2PwqMy6YYAgfzKETaQIP44LQp8ozN+5
X6lty3H9wPA/DAT6z8gmspW1lx+6p0dvEYW4odDWgoQCbE+8d7n8n//f/aigrrD87PRGFcPr39Jk
1KqlD3DtsZQ9hSpfwxsg0l/Zq+zBA65e2v03DG4dWKLQ/I5PP/Gm+auslgvaVG/OTCWckV70FaTZ
kqY2MID1/mFDSRobvkL3vZftbtTkMh0toHs2YKtbBZ90T8djUuz4c6AZjytVZeFrvhxl5HpxzzLS
y5eiZFhUUXg1cmBLmttr1w859UrMi6XuhrYuViFaqBTTLYria9+4f20/XGwSCuPkr/GBRu3j6uQE
/cEjWWzLOmYECG2YFzk07iqxkzKNeizTUNW3UKv7DRmqhljlQeEgs6+KOTrJMTWAMXSEGFadtSDt
HyQ722qLFPNxA0AKEx3Ckq00KQQ3YeSom+Gv+IJ3xN9lp3MvBW5yNyFTzhjwPw7TIQ1JLbXlrtAf
mB0T6580it4EeEqfdS/ZAGh1zTQjj6+5qzBSVyVWfXVk7sdjKG1X2hAL7J2zvkdr+sVjmsuzaU/g
WptZdb/yerhfxNoOasiuZi8pyVJiQiA56LNuI0/hS5wQOpaki4NlXwZcOdBN8VzUm9EVYvNSZ58H
ize1H6wGsKwKcqdL4luSQm7+Fw3Af/JkVz85xiyQXoeh3okZqiKHdrcDCf1d989RTIK6Uz6iKKKi
4doHDaKA9BIQvswryYxjPtD6lryAW4+fJKxg12gsQuXGBBxYsvjAZz1y0VZbUX3tScL+YPTt7c5e
Ifvt503Tp7Xn6eA1IvV07Xf2T8+Vuytpp0U5LkCEP/MKbCP6NM2rv3Cff9TW+/ffPmEZgNz5gwG7
EQ3uhEmkI6Gqi79tgC2iIV8KV/t+tjByY1tVF1ze0Qp2bYGZNa3K5QHyTOWaxS24aXoxsHTOokPX
LYK+tLYbJ/WVTmd3VpnGOvbYGxXhMICDr0ftJXIv/L6JcT6KStaEZRid0i0+mAAjcj9slbIN2fUH
xdqgrMpDJi7haXGIUmcArKuaEVdYGRW3OKKaJhv/68owfQLrka0tkx+0v3Ms8XY/zQ+5dxVsZ+y1
0wfjd+9vMzmzLBvf4JhiPSWoz6XuFFKPOIjLxE4VCYZ+Od+hM4jUmF81nu1C7mRvS2Bco41/ZdHA
/0bLDoLWXFGHAiV7WZ6Du5zZRBbRXgZniAlxfOatOCo7QGsmjV2Q67bB8mjrs8YPCt7OLleR03/4
o2hYIcW5asRpCUxMshxHlWAk0jDJ/7UglmGxO17OSXpGYyED6BEXGglw9M4qTc/shAc92I5MmzyS
bu2AzBzw3391CQdJaOtaNDoxIyx0NSnIXRl0L05utcYJLQqVFuGOInZv4bJVSAwo5s5VZ0Cdb3sq
IsyBIxhSlQYgXIwwVykI4HUNJ7MGRjI+JOv2wXPo5vHNRTprUUHJDUPSChMU6JTlKs6hphzymVLg
5TWiaFJf2neVB3ili2PixtntyhiFewqToUtQ84/iOe5VGSyeMh9Z5Rt3zt2wvlIYPkzczabVDiID
AK+56Hin6bbF3ZcQiw0YFKtuVPbN/rKI9yvkc2TZIKiGKvFcIxjJOpGQTHMN7Wjt5ALHwsO2tNhR
j++FGG7FXlHQJ+r85YCCnSPC2Fd4E7hDIagsf+XXhJmcIxRX5tP4W9EkjYN8pQeonucAdDPOOGon
TlpeEBucext4D3+xigJwPMqZ4J8PVgi/y+oC/OV5kl79DZljTvC59PAfH8n0DF9La9F9Qhtnxhh0
j11mv33zESIcvCQdD297g5KMfvZ1np6rkeXrWwriYs+P9JPoEQKKrbM9t09NShOA/O2gODMbhr78
magYvhCHYjdRRKBoURdIksxFCLHTypQKSRPLkweUeA8MqIzG8pHU+G6CPVevxOqDFeESp5wZcdFS
um2A6l14I03FrrN55UnYaUVk7AA6M6xp5GSykb4H51gFna+B5Cw/HJOVb4+y2DS7gkbil98aGxLF
XrhcWalWrFvhbI8UzBzG4mMxuAAbpMxEAk+i33NxCN4l7RJptEDaKYDx6ddUV0s744SCXl2nGTAz
b50pX7QNxAhdtWV6CkFnU3w+lBPAyUHtpmvZL/EFdkb6lXcJkZ4mFX+qz9oXXsRvPWJdW+u6PWVA
ht33ADHNrI1VflkK5frkD1aXlJB4JfEH0A30Ezta2XRSUpuB08V57HZkYQoKBHWYMpogqvOeql4w
ulHDQVeksItLZfrpxeZcvbMWoqpJkQcSMfeYRTqJ+G8Uboyy9XqxwlR/R7B/MhRXs4MNVnASeBtd
2gMHSLKpRxzT6oV9kFVyaoXddsRe1N9GAv3iEwzS1DobVuikmxn3keeQlVdU25HI0g64ef6hcOKX
XLnLOOJdoSa7SQqm+Dz7pjEdlr3Js/Y7G+7ib6+YCnS6A+cx1/yzXuqnmIOy48QySVqJg7elSEA7
qrXmbJYJeZFXOmdnJEHYrHhseTGfsRDpAllLRzYWjOQQLX9BDdEOyjvEszYaHPE47F/wW3vghxY4
A60d1U53q7K+mQL7DH5hvkGwT+Wo5OBJO2FqnD2w7xEBpMXRoTF0ozEAEVDJ+KbXnZP8e4/emgql
b9TTildUtQ5EXJorcMS5boa5jtRNphO19ampINvA9vJnqTMYmKULxPJsyPpdI41mI1DmS04B1xHF
FoeMLJYrkUei1LGzSt/L4Ub2WKBFpN8sD7/nLYQGQUCrowbTpFdl53r5P26JRZUj4ZT40VDYbH3K
TMUwRR+0zxGrKDS/hye1dmPaPNGvRGO01Nrm+4YCS5ZLdCzkG9VTNQEOR46JgsShN14sRkNM/GGq
GlHZtstY2+tVwh7x45Obrq/f0gGnPCQdaHPAzGfWO3TsbkyWiy+Zq17xwHTlw+XPSKC3B6QmAB4A
Dr/PlxWQGK7hpYGAtk1DaL5J1Q9IGlN1qrNo4TODTckKSiLkvi7ORvD8VJmgzyqpI1ZdDCY3sVM7
UCqdEYkOSa0MQjr+MjkFM5/eeSIK/ARFvrU47yXXabA4+4aoXzUhPe9YN7q+vh7Hs5KVnLgcKF9l
YDFfbWZpaOaVjy9ItdgPMnz1keFCCxDybdCv6mr/uYuEYGSLCQ1XWKif4L4Rby4+tdNHbn9Pugtt
ohGgFktG1jnej0abgICedgF1rrJY0omgK5Z7Y9NHGcUnAVxyNZRhq2UoV4M9JowptlMKpZclYMBT
1S+MahJYh9Bt6rsdgVubGL0FNvvxOdpgW/LjBuvGy6FV4eOFReHpT/VB3IJVpIESkKPhgr65DB5o
qcHiP/px8WXc1laEZMqa/F/N9mjeL3FG5kPDhPcwNm+C2ZOhaky1AyeVzn5ZOHwN7aRddayqG9+f
6ANoGgLPdzpEl4fZpqZnaksizJU8piDZBnk/1jOjUPfkz5xooGJnE5GF8odKQAwXS8joAL7nE0aq
sNtL477g1DHoPQ1YhuuNSglNXipSh/v67j46c1Bbz8ZBUZETaiDeoBoLpE/2dw0iMOJaM7OMYsIq
HC9g+QxXsih1ehhJfoqK5LzkkOaAOoTbchafi9cVCUAi/FwxSGY9ud+ynTdGGP8+Erc2rl51DAT7
CuXQCM7DxrcjX6ikCYYh54Bj9+n03EM7FI7Xo6nP81ra3f+LTFWiEKtnDpJkP4Tho9sf5ay31Mqj
g33ki3fGxo4Hli9o46qECwGlnFGpvvgX8Lg0wf4rEekGQz0W+PJr1LbrRn2coAFhu8hfRNhAHilB
sS6BZ8cReULWDalhCR9EuipQyQdzx+7X5w+790qJ603cP0smv+ftz987IeEmSs82PZHWSjJ/C3EX
7RWOZ8xz5ni3UpPU6RxC4dpw0M9VIt4wlgVAallifoWFeljbOuLQqxZVub2qVB21f3Hgjy2/3i2h
PQ3A/Iy5UNaQav2mVf0yfowX52Vx/O/47w9hFAPyGNl4DyeFlJzlIhvBEhHtg2+78p/UoG+MQ81/
Bq2VABMedNF6SVUNmByjP3bMpKMV+rOJ3pgLsfUbuH/O67uW2KcOoXr7DlpkoVAz3jT/CmWgSJ5V
3gErovGqE0T1bzc1E9CmGgeAk49sA+Z2WrK7OKyWKPx7hY5eVATDNxlNNji0/KpL5rrxrWv81Hbm
p4+lJhfUeu6ve/9aBnL2LSXk6PmyjVVcLEJj41WtgFqNj0i5h+CBd/z3NBec5s95li0Gp+ph2DI0
o5O6CZfp27dyxfG8qQvpL42vNzLUyaamjIsPeTQMCqFFEJWYzDhJoaqMCqs0geoPqTKVI03qZTVG
wdYlLJ258iHHzDzmEysVq5ar1WHHKoAcowR4DN5Q/syzD0LEC371oBHa58CSRtT3/q+dGc2um5Av
VjsYs38B3FToXeGXwzSGCGe3BxIp0gZueNtkQRxilnud9x6H0jSxte0I8gEWxbwalnbftsG5TzGi
1VsGsUCaK1aHposWBiZBkJOl8Y1qp/3+tTXB06gRyPpv+w/ED6OnViQVHNbcKDApgps9kWaJK4uR
3sdUyafVqsSgd1CNay5i9P/lYnll447X8YvHShWJaXMXOY6GAqDwIDClXa5Hm89vYcSv0+GnGkuS
WVUiYG6d3a+COMrh2duEgAPSeskclIiKDTqWjapk4Zk6tA9SuQMzZSVl6d9RZv5aqmkDoSKGuWxL
SeAGx2p44uoIekfD+88mT6N6N9AeCBy6WVONDpTXZvqt29GFA+Vi3sa6Gs2Zx1hCmbmESvbKEeb0
6rSBdYUmpwQRnOVGsEMqVV2Jp9bk5hMsGrHJzh6/otDWjIxyjBMSZVpk3Ed2nsIjRD73S+6zMzLn
J5Z5vo2FplF45lXuUg+uSAyjGzUFeQpKpSopygPTYkTrprsttWGHBVLWrAxxFr4V9NfCYHfC04FM
NZQ2ZclkKMaVP2itcJ7m57yXDTR6FvfbdLT7PzPukzYlSOqZEHJb+cmFogrxHbjGBdm8FummpKnk
6xf+abZKcf7kxxolPcF1ShR6ATPqRlS8K3tL0510TasWS6yj17i76AvFADE58Y/RmlMiOvEnML76
bqImOZsQFAz7N9rc38uXDkwD5XaCHcX05JcgiwHQVvYtwPZT1v3+SLQRcDg2qifQstBkkROFLWP5
k4dSJ1K1AnS0cN+692XodEammkKYjjSTNkAcJZS6V5NEMmMfEli91n8XlxCbGYK7sKwlk/YQ/cC6
OSmomUPeiaAXdo8Oz476SZLMCcKSYkh7VRJA4qI2JY4M/3imxwc7iNN2XOfSRjOgLWMAphyaUeaS
7vmkGVCRMMAuF0w4sQckUF4ldgP03rrl88wOK3fPwHjP4e7CIqU6gqC0b5QH8eTdjIG8QjKeTp0P
aIOK02oINEhqEJmqxtbTfIDfdwt4iFTEt9R65Y8svPnuanQyCKt3fsEENFYLL4DGhElnO0Rl8ZLl
mXDnuSq0WPCbpjOFg1/QhXDSYmXjBjRnuF/Hz9Mc4YLxHTMqgCYo6equSECU+k++lM3EGNXm2eEF
C/qz6iCYQe5dO39Lpt9st+Q3DouTusFlJPYIRcmYmYTsnl+1yBZxRx116kuTTwZjRsqElVExM5v+
3srb+RQJXWO5WRn6uGY77bke5a9NerftTYybyZJntYxpc3m3eCSDOFDPDmxCBh/Kg7/j4+foFuin
mWs6SVUmwHmvHcvtsnaE9Ee/Rb74/bEUT2X5+3yC0qDz1pg19uOTvckaKzgv7Owgzx08NFIPvSoM
EXFHKFA5/0X383sl0mL+Nw4Pz/aKod53PIp7GhVgYKju3oPx2fyOpodn6nGNTkDG/28AgeMkdYvy
seV/MiWRCThOCPAadKaNsCB5LGsywpzTqAZMUjulpE60AF0LUDmwbs/G45JoGUKNvz1JDX+3orPl
bqNCvvYGPxy1xls1124wIIVg2kykBTpaFOZ+UPmW6xdm+xbO1kE92NtV6bysvjudOwzRltVQruro
HZDG0E+V4mQenMttMX8FroE5UmdnJFdiF4B0SNW6lezpV1wW0kOeul8OJ0bjrH3d5eHPm5X3uFE8
ui0ayOI8UUvPgUJdAD4EuzKHMQD1TQgCavNBj5vQlSo1wSbcRmSkka6/70V5/Q0a/0gl31Pjw0ee
raLRko8HEhyNxaqisBFy4gKMF4ZqdhuU34r3HeoMM2GNVM6+9rGb1cUKzs3k1rXGuW5bIYibAcXm
4V/63nusRP9IEBqZClumx3vcZZCwQVP4Lyr8e612LVbSv7V/iDPEaaTOkirDOl2it97zU7NLiDnw
f/RtJ+4NXQjk+CosOQQAnNdSsbLmQmkwyWpCj4th5nrOXfbIAI3jbYp4FjeOHb14VbY66JI4N4uZ
2uL0tIVOWQYM2sGNnUxgweDppE1hZWX3wMrPNWFm7ixZTnah4xlH6pjhrT/NIoxM36FFkuL3OGrU
tSrgey6UkabBAXreE2kQj3pMclOlAN7vrLCGy8XvpmkZDvBuOmxsPdZtC+xRjXQ4vx+toZh2ELQI
HWscq3YJaEVnhL4zZTIwyoRi7bmd5qsF8/LXu+X/EPRXnjrLbJzmdzEMB+C69UYL0AbW8IE+Po65
1df4SfZHgxOzhfqMY35NzMEQxxEeANaxwhHsk1F/z1bP5lFljRinysah+atkC1vBu3iSIVhwYvaM
DCW9XaDgaDbci2uFp+dZkKtON7bR0VCqLIYzChaSPrPn/e0KemBt9Unr61noSw4HQbw9jYbR3qmT
rzfJvxUM+aSmrRIriS1gz1P2O9RUszdwcubcgHfY+7TrZnLdUzzSPjJPv7LF15Bcc7KAbzDRJhSV
ZVv9GBUUP7Ktbjx+IqBKtRC5E0mwJkJkpABcC4cUYUN9osmA9CLfl1xS302izDmQGIzcblOnOgOC
2XdN61btzY/JNGIHjjJcxJKSwDuiKOq5DoMXLOn1XQCDAx06AF5ZyJlDrU2q1GQMPMxkeFGPziPZ
1CZQEDDy6SJGbBovK2oPVi0fMls5YZqyYtuCg0VppcpHQjOKgoxzG9e+hJADhwM0V7zpqi1b5vcn
ANyu/K38vtSHx/AyRUvLMywXSucKg9cV16k9I+k2n1A1RyDEggGbNkefBoQMXqaKmeG0HHjLvBrf
kBHKlznDefmMn8/4S4Etc2F7Wuec9QjtadSR/31y876eG/DOoGAlaaRG7HdMR+7sfvOGCvU4ztrR
NUFuQJCrlInhjWKFHj4IU/EEPYZhcyUsTSsVUX3t1Pw1P+0pWWASBeBQlv7GkrLgUm3FdZNZWEd7
amc8C6B7ndamYfDiCoOanQ1Zcn/21PHg7X2xzIyL+yQau5YspnglM+Pr9NRmRpk6D1EakI+dYs5Z
+M27DjNCNetbNPMf3AlM0qtP4nCDqmf8HszqhBvBcKR84G8JdPd1KMMAixWA0c/k+UM+/OyOFwbz
rVUmSzEcGZlXM83yHumgjIi48uksIt0XI8Qk0aaGESnEMInDV5UbTeidi99mQ+61+99LGgoLLcKf
gr/ku5DDmlNMrIGDEe48nOHhV+eHrR/+YEb7cnSPLfAKOxXR94ussXldFgYHgnrG22cP/tes4HM1
RrXSknQLZJquIhy+j3W5hhGiIAeXkzLGsXRU8WBGGhyxk9d3yAgYAm28ItJ5KRUN1ZuPEYb+zY5v
0s84rUshMXwYMKPq2fstb2OeHYKAP9UaUai2/ecgHsK+AnWcmqSeoIT+VRTYRardXcH7R5GHlXMc
BtuoC+MJRgbGc3lsbybr7s9GkCL0HI2yT7hBxCnn0Zpv4zGjzBI9jgiEhYyjF35+UJ340aZyO08r
7zZrrQZTd6+I84mF9QGIPL01e0lPmNfIBd18dQQbWQCkdOVruf8bwtB7PkUpFJEKw+snFZ+wAf5E
yuoZxC7AeoozM6vRDEZGF1kWkWp1Z7NPlE5lYw/p25+LSZYGBy598FWnVSZICilZ0rq8Mx88GQwA
us8WMEttQoaMYOHuBq87Emy7LZ9ueOYJNGeWvLjYM0K4fwoC4296tZDLfKBKcPSmuiZs2kzGjsyZ
M137oVoaHFqjl7Yxn79rNOO6KaTjQvue5t3ocfrVBzzbDNhZfZSHAQ4vVtWtcP/zJPcneTXhWQEJ
UH9Sfob57ak5Xt8IzZO4mgbS4NPbLNm8nJoCcmntidr69tm+X5RGoRLQOEp+/sMpyMAiTwV5VyWw
nQAieH/Sucu3kUzFEqAo8OYnDqOMoYA0H1s+MfWvKbxUd67UiPLjRbWnl+Kq5vx6RJYuELi2qcnE
MgourBOwcQfwWc0Vq5ZAqVX40dXbHoDTlmsFTsCzimuuMQcc2fH1BBrXg+iPHp2AlcbzWV59W89t
B/aJ7CrDkDST1d8vDsADsyIl/o9lrwVDp6yqimnes6wvD7r9fg1bL8UB1M5QnHvNA8C95TmDHybh
720FzenQbVElpb37mfwN/iiFUCsU5d3xjqZ6uQYMlp775JyaH8nIlgRkvx65SeS5LP/8PxCdL8bw
chV9kbJyCJwHa6781GK/Gd3kjhflLnvERrrh5Zp4OOA/CCI/LQC9izHtqkRdn3LA3q3Y4raLUst+
X1h9lC94PX5wy5YXhxOulr+HImJjZovl/jbMUYXShi7LuH8GjbSLExVewJlx5l9iK7XEqKzqRN+H
2QN3SJnhp3BCEH4Tc5y81QogauRZJoPeGC/EYlh/g/6nVE1mN1D5DKeSX8f2K2oNlaoYmmhxcpcT
x6CnMnZbdqw8Gf1pbym+X74u3TjEHBHgcBjewY6jJN4ce9iC+ZSPRbLP9MnrmBwRMDPCw/35jjYQ
UsYu76/bB5uaO4SYy7e2DdgDr+IeZOb0hTVVfpbSi0l/3JYph5EJQNDVsoIC5e+6IXOl+E4NGRFC
Pk5vaCAUiihikdcWDlAEsQgXezgA3rkmdx9CdJJNVdCHVXVK7la2K5ARSmzh0kNjRCAxwIH10RAz
DZDocV3xY2Zx0bvbvuVtyz7PboU5rRlheDQJmKWsRCa30n9hjDJ4M2N1TDVnvZnuEF0FFzF0ntFm
OpVC68OYc1MlCwl5WR2QO5NN1bGkTDxOEIepoA/NFhVrT2ZXMUIK9g4QNMHjTE4OHOlrJ536gT4W
NaG+OmFmRuPaub1wyxSlwCeVJFpGGR0zRGggDOwDknEA2AWdJZj1uIY4pw21nEtVOv6CHWO9kNjw
Pmiz3EKmhM3YOCfnSRwsujwS1Nz9RfMTAt2HFfB+8w2bRgZW7icdGDB3xQUhfMeq6n9qVOqyPYhe
W+fAZzakokC7WmqXN9t99fwCAkCp7G0ToyXVSGo/SLFGDXukQ81mlr3Y/MWzTt8QBHCxrBi46iVE
vdBSVytfmh7HYe/2YJCEYwV6Z1F5PgEQv6K891Fa1MP5MXzNOsbRs9sQHo+4Uvepp/JCXdvi7bwC
17HJf5RK9BvJI343Jqm1Ikau9fccjyQhK1qryDo4uDv8XrAt1ptuhY86ffHszEw0Eecklgu6Pe07
Iupo52L4vm591txXB3GM71jwldpWm6UxvrUMxXgZn8vnzl2pWbf9i2LskE6U9AaH60lVhuswIpOa
lx1qfgzeSfn8gTc8RPwhK59RdFoyZ11+QliQgFthZ5VzHDOzmx4Ao/G0OAthFkiSU9v/IWjRH98+
zoj8RLJ6m1u9pbcpcbYiLyXiTeQyvqTJVUnwXv+KD3EGLUx7RsK9vI9b+4jaL1Hji4cMlxw14yBR
7W3OPakaYKaFoie2elva2qK6HVgRmfFx8zvhwnlyftMGPs+6cL+UgAmK01ex+diZmblVkpX1Stzj
4wd0zi9md61GbCT4efP/4XIc/AMAPmzyeMLNFRvJFE9egxg7gX6P2ic7CYwjBypuK9YSKm80VLXf
85KVQdDse73fT0FsrznNuUBOUH0pbqqoFyn80ymDENWDCFSQYDU9r1Z4FXivLdglbpiQv23M7A9K
Fcwm1SSkP2NPeFCYAVd2tUvngXEqazLUVYbM71sDcyFwjkcnYyd8eUvhQQgOagKAq/tIlfQXRQbe
pgeyL8Fd5GipQTodqiMLSw5+CUBn1O+4bKWR2arp2YdLME4M1XiTZqNajNIKZvPWUuH3CXK5Vodb
XN0lZxXtu13GZDXPAiGBazgplAYNm9ZhnG/N7wp0WJvyJ3PuDs1fqAgNcwibbYjv1IuJfD0Rx78z
xtIvFc6yy+JwBUZ7OWlxTwnUOmVStze5ARkkNhpwvwCNH6SlfIHCdCW7kMA1qw6bXx2wRwwLYV9p
Pxs42H7rgx4E1LbchEIe3BvOf6bFkIPK7COnjQatKDkZBPB/pUwP4Mt7SdhKvDV8BmfPzxj/+6ud
DBT99thh1bbmK0xg97ZloPgBQCvL+iu6XWsGIo2vIykxdvKyUaOD7NmKJgdO+kv3k5pqYRPJKTFB
WXB//K1OzrIlDrlo/vBVSCZOWqlgHyvCC9ht4vMTlZ/X18kVmPhbeVM5Qdg+bK/E/ulujT5CBChm
FKKYi1gixvfeLDLeH3H8/fYuXmtXdrpNWLCNvtRN+dT/6solBfpG3yi+1CU7TUnxNy4Tx9dUHSRt
Ukd5vFCHvQ3yRmhl/I9hy6dNvvc640vjQ7bmnDzgQkDHuGOzk+fE70OtHg1TG+o6U/9+I1sq7R8Y
XT98sQMsHDMqN0Roto3EieUrd7ZciQo7/Ss4HNUtBIvpXejFQSA3S/rHYY+QhIy/7VaPcS8Hebut
Lq1faSgII6pywtQd9tF4MeJZWbSQOt3Gcuq6ziTl+cDQga1j1Y31ACrPv4vDUrk5yJqOzAC1LQ7Z
zVTkx32vpoNS3p0wW68EMUFCoORtnkcazj/r+BZPDaSMyW6A1pCnR1P0t/eJV3OnYY/Z1nXHhphg
oOUAudogQHFk6sbokG0stCQMJfHlNC4fjVAq/pbrBI8xvMwhXg/saRRNg45Ds7np2u4OHc8loSg3
y1S4jmjeA8wc1LX9jAFRUsr79dYYunFtQzmLSLhl2Iq/lpgojw92UlvDvImlHojLdjKJv3M+RJHi
IPP7U42HU6xufzuHS3VwIBtoa+6mqY3cXwnsYawDWFLgNeIjpK1NX/ZC95l19Mulzyyk5tHyU4tw
NHImCSodznLzm3hK2BpDfhqiSvE/17QPacyTucjVGSRNl4mY9mO8M67RGVfhWeoSGNJ2pM9iihfO
MovPBOYHqTjMqtVazwllWcaHK8sidgKQA9xA6A/yY5s3IQy76UK2HIJl7b7YXGSbD+0zpYl91O+M
pBIgk2uK6Ejzmp6YhzItfWoHszBSJEhiDIN6Cb61mmBGlDVUQo15Qlt0TGCdGoXV+Y3E2eo116L0
jYzEXPNcOX5Vh2F063I2m1Rmfz2lBlyAVe6lysryPxdqRFUiTMTjGDcrcT0IuIDnIw05YnlplQYT
92YcmVUWOPaIg9M+ErDrmHZo1WPqaXP4gkN3JWCcOdsmIafI+ExUqlRznk8jUQZlsghBpmgJX8pg
9pcCtk8vsnq11kZmnBLYlu/gQV8JUEFM3M5k85qrkRHq2OizSSqY1EnklbwRXGepMaG4YuHjB2H4
/nrB9OVneJU9BkXOemX6GqJwnbnoeDbPQBiRhaEutVer9iZJ0JhImD5x298ZJoKnRZ6+dIIqtwBV
6O1jq4GYweMgk6nqIRsb/lBq5gwW9yNF1pNOEkh0Pbxca5CwZx87bkQ+x9umDQ7MdLuxkfHmijCN
LYKHgmC4lzWviU8hxT/vyWYRSYmMtwQ18mXaM0DoEono6Zo2P9LhZPHjypvvkRcMwinaupjalkNd
H0svm8QpgNtmfQVfDJua/wNIC+BeJ4fk8CEfzQ8dHvPYLdNJiHZMeta8zrOC4F8mqCQ71wQuvHP0
bmxJE7BL7Mzk/ecnG9Upv3FHgfvtqBB6thn8vANBJCRCBUAkjOxVAa8lYQDYq7Tz+QFikyFTrGVk
TdAG+rJx9UaPd5pekXCxMV+4RFPUSi3O1cJU6svXIOXaw2wlCbajc6fvOYubJvkryoSQlS4C+O/r
vDn3PMbHLLdug3wSIfoWrpIqlQHvi2BWkkG7PCa7dlBQhje1qReDt4MevtIJXZqSSBwj5xSK7EGL
VhwMf4hAENV8CbxBxDoBWFOfJFmSkDJ5AvLqomSB0nc8GVWU/0MWj6/2i35UkWOpEqAHbq4h9GOX
9rm1TRc5xLEUe6o8vf0CjgvQ521no7r1Pr7g5R4vRcAGwPOHWC6Gq0sUJHXiKNEw3AofB4gRMLso
uECRcMx1Rjl8h7BX+QMgoA63ZEWDruOpchBo2EaK8D8a0Z+lrU+QFOzHfC+975wjrrupj41hprHo
UgpajeEkWc3poNNVamgLbJJnakBWeaDxONEqbBwmN4uKVwCx/ThcXO4IoEVhHvB+HKHrgudhJ+va
KRlIdIBTu8saq21dVCwgIhTlhC/pycVS4wQCcCBUtXumSgb5QEtGHPKryhw2uHRyheuYxqxmtAm4
ImxT6kX0LzEvnJ2/IoAaLA0lifvbvnmwDvfPC8/EtSnzX+yRjrjUd06vMkeaJvvnB92A9dmv7x31
8spvwJCsuQYQ9kg8e0pstCBT/fPzLPH0f/I3Mn0TV30SwxdqbTk/QyfwX2qqHywvGrx/VDQDAVA+
jsNUK3gRXevzXLHTt9a14HqIDVmWolAq88JOpgfjkYWLCLhfB/IHZ6PJ7QMtrXotrpb2ucZ21Y60
VtZJSYSxTRsvDzHpUEiR+nPaYe5CD/1StOgT9dlB0qzYKPgOm/EfId7wEUJJyizOZC1hIBdxkbPf
yOpPSqX0QWwgkr399RyCUd47cFtjeTzWs0qDMJ+yNJVkkrJekFVFA/hJ++GLyyr6wSmCpP5zHBv7
VBFbLlVzsJ1vJQ8boIH9ZAYH6xmWEcIlnMdmwcV017/UqPOARxbmPicfhntgK+ygEQ6R9r53ST+m
fPF8CZSCI59kwtt2qbKbl//YopwSBKycjSXz/mmn1MZKx+/veyZumR/Po/BEfW16Dg/B726FXmGP
fJbNpwckRCsUTbxofm0kyphXpyjIytFD2bWPyU5daNb6q2GhVH1+F7XCttmkOOprQ61wV5smSgr/
8DIUQZQi3X+bQ2cG+BNX6h8ojVM1E+lYuHQBxFBo2aUaG7MuLDWmsm9+FQm2bV9vRAtJrpqEnksI
TYriGBY57DLcD35qikaKUPnwoMVQygF7s6kBHwdjT2Txz8JZLnQZcMpiBdQ3hhdNwGvVmRmJBfue
EP6OYIgv616bkapIc+ViHSqNcQLI8PPZ86enfHesaw9BlBS3lvlnYlSCOItGt7Vg9TfyTABlaDt8
2IeaF9Vv65ewwcdTGoWd46bdX6L7HgVGJRoXSJ+g3KaRF9JsTq8OBwcAI5yfoGJ3Egf6MPB2pkPG
qxAIZ/AtPaJOBjhM6GAVrUgwmM2eK/XWcSBg2e9G74R/AfwciK8oFulQD/zzYqUTAeD75Pv2mWMx
zy6UnOAmT4yN8tXomzZZ6Oembnp3/OxyMtlqi+aPvefOv7e2KRaVqoUImv12ptIBxAHIKhw+cmNc
CJ5maHT6NkAT9/uTdWyRb7/8gbVVGkJ2d0tn3+T+3/y5CfyVo4QTMh4WJ642zq7jFvkO7NBnsB/7
jklL8YAg1WBYbL1KQXQVXvwgKSkRv5qffVa4CTNBeCFS9PhAvFhs4ckcyETOr0lsZbgYhKhtune4
IsRvVsDG3bMJPSTTrWYdshwFzdqrBX2gGSQpSVFh0gbdhwBGDLbO7bl/aqJpM037fz973tq3Dba8
YsLDG5G/trhAjhtu5mxZ7vnxvIsxw96MEdSNJp3uY4b80xyq+oZkYoLcL1O1M2g+GFovaBafMukY
2k+AvehrfUtnI4b1c6VO4zSC5pVsUynuxkTKwn8YUK9LQU8sIhTwxxYDOgmJdWamBvUTXjDLKQbO
uoRG3gv5t3bdfzEW5Ht4N7DB+p8qQBckngxdO9moqUP6SBXAqyG5gw2aJ+1iYxmZz0BXUEd7Stri
oouOWSPsFbxRrB7k1HschI/x6wigq7aSBH/O8jd7b33U3+9bTYIEES87KS87Q4szOqp5BsMQk35Y
K2rI2CpsDL44uIdz4zTxvreHU7l8GrPlmVy26AWh5YqqgHarANW7PsQxqzikP0F4x/yVpAkrlgEO
n+/dQ1Zd8I+xhj3g+ALjcKXBXSI2fNqKNKAqXClDn4py5IQXXX4rLA17xQ9pc/LPBxzAfzyTTqhg
N88xVoZ909TcvOSNfBEmxjN3GDkhGnxJFUmprApIa/qDNjnLP7BAgDXjeGqJaKulf6gN30NbLmfB
laP6ashILx9/877fPEgI9hmrDCCLE6g81BoFtzyWVeFn2t1r3YGDJa6pr24deh6vvxjAv+qOIp2U
Hon6OwjY7gZNEqvJLRzuK49ombj12XVYNgTy/++ai2tPvD7YuZO2beT7BbvVbHvjIbV5iPdrq1Lx
64naoZLzNsl7GZ+15/C8TwIHIkJLb+n/sy6LRE2wQjFqA6b4Fp5hwU5TbRR+RiQM7y6/ZUDXB9sR
/YF7a0rF4ymRs6lfLY57k4MqtUec3EPDUmhtQUnMPcVrH78YPY6gFBIQqPAW9Sr9QIB/y6ZeNt79
rUsOdUz91jTnQtm7v9SvzEEYX1wXPO6l1dkmBCTonafm9+JpJp4xPiR0bBHaoNSvv8t2DlV5VgbR
VbdZzvZRC5Q1WLcrrTSTP4I2tol26yzmLi5cdrGWXHVJW9L078ZBUR1b3uoeMUIqJUdF9+hIxVS6
wp2tREJmtFO9nuEJsquTjIsN1hVK+QbrXpN99vT7x9eAXI5YxWo3ugurqcKS+bvYrfMPL5NbeSf9
vEtGcUbOxr1MRKMadNXGZXxVToUBxssuaY7AGF66Ci/hlKMTCE2G/2Y9g8EZYoqq9SKKeNygU6xa
8Sxyf4cWdelqgMFau5pIfuWJBKystbAZOqGaMmy4vAoNoykFpb3k6Rw/ZV2yOEXvkxLGsRG2ZGVr
IW+UnujIwrlf0y/MNivCd8ScW0QcQNBoxvbSKX59FFwTz0siA3aYer0t0yeEJnDsgKxobOjgqLvF
+7qFmfB6AbzRfcqB/1Z0GsSR2ytO5W8BdKSHsdxDp9vAWUp5Nbz/TDEuKDWmWU7hhfBfJoOd6sVu
FgHfJWg0Ul93eUWTlHhxFe/8Bo4ZM8d0cj9lhdqhYKOd/wwrOK63jZKaD1YlDvYDt3x0c0UM1ups
Q0SscRwwGA6Ohu6s2GDCuzCOjDqPuE/wc8n2mHl+QdpuHSUBpRt02e/hMs8pfeh/54gOojgz8qUD
bF2BCEvsKVZOeeasR4rMmBmfkDydha6MMxrXhCTwHxMuU83D2Rz7VKVKi7k1lOhhbDGWAl4LaeTI
CmQJKp3UQ+czIAu7HQI6atKaH727NcDwz1Mo8TZrD6DvBvB+vv3yAEbGHrEdZC0ZylDob4H6Akep
vNZjg4m6qr2xTvsu9u3AjkOr1VlS5XcRTYONrIu+uYKyWMnreaIWrUleSqS66F8Yp5gSjp4KqLKy
sjtH6yy0sr0hQ/ZC3ruskZjg9Kt1OicXx8oPF+HtoybAaOi8aIf4qfv22AZoRDQMN050iMdhzRk5
o9DHmxliUOYotixaAlAn8QO1x6bTeNyxat/kVfKEZUM111FpdPIXmExXQYghM0dSiHQ6vIB5RKns
SJpgI1+pTVJ9GqujNucZAIx9SWkUMeVFltyLgplpBkkXuPpDOpKvyOvMr/2uCqt+mu+Gu9tEy6fy
P2kARqiC5bcMIRSR9M+1zGMJmYUvg8hNgY6k4FX95PB8UsYVhsqW1okUFW7BSFdKBocYL2eSzFtP
B15fM2zo8r9tQ35y0jqkT6TP3rMqkb2vq7/SVx7K0X2PCZRm/mBtpUkpYmXMypi632JVMR6BJJW+
Ot/Izm2tWGqBaarlY8d03JFWdGH2A86AYO6l23UtpKwzMNJJsu2mciwefsSvZ7bBAFfhZt59XdHZ
qAHxQeU9OzZpQq081fek1RHerZnkdaWkaKTfusyLodydMSOwLOHfOkpNusOnLYFNRASf33TKZE8/
In4njxEFRJPV4CDsymUWY07FjRKFw3OOf2ct7BUdoVNZtY+gkCNgHsXusDgYtyCCWlA8Qj7cZM/4
XM82gP3jAhOp3unGPA1dHalcrrFhYY8bUHZutId2csn7fi2AMD1AphbAZf7JVw+kdc57EXOk3/TF
Q99UUV0Wu+xTM4UBPY5u7v/I6Czfrbgx06Qs84pU+8vluJCc7gErl7HZvWQEAM/3gC6vWI1dZU26
1iG53GdnT6IDbZxjMqLhEoWh006we24b/9xy3CKNQFgfLJ9dSxd1ZAuQ88nOCEVidfecGrBNEoEJ
Gw69dLZjVyslW7+NuhOOhby66N1dXEV7SL/M5Pf8WPPP+N7VnOfpbX2Cr/UlSuNLgaulJW/kw+0l
eJsthG9ld4lhNBmO0D5HfhOLKAD4q0wr8zuXUvnEFrMxj3x2f7JKj9tBCEHptjSuQ1HVQ7lEPFvL
yBl5x65BqF3TVY72/laHve0rMAakWjA3TS/7o8jsCDsMMFd+aRREBHfRKY/alEWh5XN0nxe6DMIp
bE5QyKe2WwFm4cbGE/Cpp3kP6Y3nFt8O4w/kAxVA58mFffDNyaxuwb8zkxwnAwhoCYBsnkLDDm2w
Lyv4S39TvOGALlNIejAxD6yHcgGJXxqYqKfT+Gs577P5XpnsMRf1FWCAxp9hVmFz9FLkrRMGutpv
o2x3VmqNnnJO8PxjcxKO54SkVTQEgRZXz9x7RUQLXB92x4okjjEB/tQaeb7kf6m3cqefxgeyxDIu
4nKmzklgDLKJZGrAWFK3WMGRDTlwmD9+hQc+TqBxLbvgU+Ols4Lofy4GvFW19512S9Z4VmvOJXl4
p8/bniLtbUwoJp/wkT6m2zBdZipaCAC7N7KHYNn21jvIgW1nAMnLVblvaMS79XmBa7joh0ilA1fL
zmIT8DEArPIsVIzuMJ/2Ov4/zvdzM3h0XICZmD0ar23vYmLlTemcQuqgLpEIFfVnUipn8wxXKc+V
4+iS+5DKCk3WrxRq6R8f+dQfXZeNrr5lOz3Y01M1dPbW84CxY+x7ABQNihDWXmigvXyq82vvQ6sK
TTWVYd2GK9p3qvhiKF8g4RiuU+eP4pnJX2rn+ly63++hmKT3LpK0u0k/8cQRGxAEvpxo4QVQmIGc
yeq7uNqjTKomJ2wm1tvf0VLIoPfr/5Hl03IbWlo4KdR1kUP9/oNh8ZSb1AhR+rLIMM7hecpqC2TK
YzDYt0kK32Fze1kyRla+Bkt3zN7C2IodMzPn5wHtWkJi0Afj3kRn0OhK/2miW/qnqVaITvaySZwH
oA19r5MgwqHwf+W2ikp6cKmz+fjXtIXT6hcc30Xir9P9yLQblkp3n/VCIQXQ6feRrKlykgmkkAIL
sLzgYkzJ9z/vAEKGT39iBgFSdSrMWqxn2XQ6kQN+93GdW/hGVxQP/ERjp7XExZALrWDVl8CBzAOh
AIVyq+J24l4zhbuc/gsfZAl29GralLhVCmXKEFzdSYVkTn8m/utu7XFl65HrBV+PurgouobhZSzp
JZVT/u3LCtflKP6+McPWZ2zdowli+zZTyKg8oFXodjAWnKqto4D4L5DLxoQHgOiR7w495AJTm8H1
/xLw/eGGPjhonqxZhFZc8Id8L43isfCmU516TvWYJhqJ22/s7afo3405xuxfl5vJm0TaXkcn/6TS
Xm9mJ/j/OTqlRDfqy4eyeWKyaDVSv08i+a5xb9H4gIDD1gWA6b52RswjFLYbA9u8tcwV8kdJztyA
z4I59yDwkzRD0nugrGIdza1WS4n2RrIcYeswt2Yj4d99Ei2ovN+FwiDFiUfKDdUfTXsYGXPyrQmb
y4gLQ7symFlbYi3xXSto5ZNes6o1YvGF1aZVAwU1ElQfAhTuSDMrKB7t+OR6Tscz00j4syd/WF3Y
hm3eB6fYD0PYm9POAsr71Xh2BB8q2o0sDvT0A5VVqC1ea2oNymSkySqAApyipBk0bt46uO85Tete
c+up15FBCUsaLWInjwKuDnngY+SA8yF/9Fq5rMbD//4iLuJqluKgbkZ71nhjEmAbbUkrO/w7kyhS
i1FxlnjrS7MBdvzV+2ElT6SW/qhkkaZOo+GOIBMarn6nOyJXGb1dOVQON4K1eIdcNPpwxTeY2+6A
HuLSlix9TjAjtZ5Rr5ayPdda0YRQUsGCh4EbZCjMYNmf/7mtdbrGSJW67Vakq/g/BZAxtNLqhxzr
tKpy3BIqpSunnsMxan7NIYM1yRp/4UNjor/QXkxtj8oqrA3bfWdRsue+yrbNdn33FU1lXn3NIdxy
j+amgucVBb+V2AM+Q4TKW4e4R5nT6Krmv6wFH6H5WuUxGn1q/DRvlDQUVVATCUMUe3aYJHr8RoN5
T97WR4Fg2AbELhHPud7+PSfnxQoS5n8Nt7hWRPz2SQi6ucJ3ajfFxrHUWZHhlC3dP8YwOTqgbQND
aF8BnZEA8uG4Ok0B1DGqLxQfBK8xkdLMNtgf4gxgUnOfnBnSq5TXagKqPjAArCd8c8SjDSKODhxc
YuwZd4WqAm2I7WtXichVyxVXNpJnKzmVI/3JYT0ix0yhbIMtqJ9FJ9Cq56brHOGa+e2nB/0XZK0G
arDPMADnLnGWYDdICBMzmwJl2WTFB3yvFutG7XNkxwOjPPAmLOBYVM/fyEqCQncYViRN7OKJyW5G
2NnS/OWW/4DFt1y1SxJ/lNBAdhkWAu7ZNDcA6P9RxvTBZNOIYpwMRRVhAT+R7bCqCDP3pY5upRjs
wDt9ZfhRDlxaln1Imj58vvGraAGYw3dBZy2yPI4b8MLQAX7pVv5LaKTD+47+t9GpGK41imGlwUBh
HgD+UC9mFeNkKkkMRKeTjfVy0Qq9N4uljqpB0jgF1zgIAYfOJdNI1sKsKrP62GGMYTx61b7k7joP
GgoPGEFEVsY1dPUzP5rXjYSb8TFxV1J067QCqTRADHCQKukbXlw63kvLYvBZeQU/dCl8Xh/+DKzU
9VxiOkoF5C3+ZOPj7NDpxNQ5AMgFf1wDIWGHI8/vK6W66ebbS9xHHbnFT9PPhKMAwR+GDaWIqx5P
r4poR6835QaxIBgxiF9sDInh+zfTie0BXqMPQ4qDiLw4MPN/mQQHwRGSVkQs59+t4uHjtZtYmdXi
MOlF0/RXsLeDUgR+pFVerpUfGkLYADtenbSVHIEu9mOeOeaymEDxEsukv7rWW6B3wrTxKpofoNne
kPIUjNAeU/Va+/ZpXqCU1Fvp4RyqUwJN88refuZTaGiDL4PBwK1mU4UGyeqsZwrxjeNcvvO25f1N
89YHH+S71rrKVIuhXNpxK55HPNCndxUOvnV9qgM4zWyWS1CifmTAPdFi7ypJ+j2A/O9WE52qNoDE
3azafFOMEmj1+Ul+LdJww2nTih1VoYZxT3OKikZoJ+f8ezgiq34F0V6LEQrJej/4LmS7fjhNJm7l
+1/b9ORiyi8nPup2jjTexPlgOLY383uPOd3TB/v4RgaPCiBZwbbhnrxtFEhjZ3lhx1SWFpfzsalT
rjvvHVpRROccIsXgZKTLWpRZd1tPkC6Y626Feffy3Bx9YXRxNCExV5qPwVFvImle98Ho7Buz9Zrx
996RpapKW8Paja+1TrA7IGsJbftnnUzpi3W9/Wn1qKLvw2/q3JbQrITJMv1kPqMiUIBU+faEDgzj
Xw3DJaq3iEEX+wKjXwrBgp3YKux/LRhni2enTWHyc9b4XbJGe0NU7+6vRaBhp61ouF+/kKm7+zp6
+Qb6QF3I00WSDyKdV4nwsiG0VF2GuTsUTVWn171cBx8lxx4SHb37PxYil/IgwWkxSncAMHo3FrzW
xA/+pwzoWvbJ67iay5bQu0U+XSfRzC29HiGeyR0X2RmTtolaFPnkU8qx7TfEQ8S6DchZKFLjqP/x
aO+foKqvu323tYpdgroDasM38rG4wj3mXcDBJ7lSmbvPWdJai8uOqEla5AsPH99hzp5+1ehwc+Af
Qh28YcG6cZZn1qdBZpT1c42bMNiAvOYEzojnblcecn4kk0EgBcnZotd/ZbgKoUXjHE1SeFZi6B+W
M8Z6VwGQvogXcEUz0HQOw6R+Kk6gcXjjXeCh0R21BelCoExo3FjpV7Fu0A0dXU/29pmW3r9M0ANj
FPgw6UEu2egjGjd5Qj0YVC/DMg7N0mrlGW9aUU8jdYEXIi+R4yYGpEF6a8x29iyy2ibkmfp7J9CK
1z4qIN2G7DH5/6aTD8nzsi2syvo2KnutPRzYiQD1sFjUhxBui2pbGx0hXWApfo2F/J+Ps0DeBios
4j5LmBSN/YAgsRMiN0pfdxB0z4Xn1mNJDdf8w2PrmcECUYmmG3STWa5Vq6efD9SkndgP0bExFOYB
plOvw+NvmArwJStKBhUEgqkHWHQngqikx/BITzB9lzq3idYHuC/3icwPX62j/AdVRZK7X3ep1Gpe
HQ6C7aK4+sKsqZrPznb/bnY3Z4i8WF07NhdWUI+GJONXo3Cv07UTBOSZiTeLBOmX1QKbCVjiuAIz
9f3Sl+PjDa6fhzh//rWRzDlxFnZj51x6q3tBAHTYMxSkOQGBz8nb9AxPNM+zGXTEtz/xahrnQZCZ
+7oiLpgOTuG6/1HfAeuR/owx2xeNbIx5VeVCiT0CgdTEQ6hnPNq9Uv/wFVWhjiexJj12bf44ZhCQ
KhGJscHZZLPu4nR2SbiwfWJfgM6+laotJpiUIm1SX4l7gVPAYVwiN9ruyhWuuFV8FTed7PWMV2KU
aA/Ay5a98ilEUUKS+zLPjWvfW7qCi3cq1jv2WQv+vYsTh8yvCGdwczlXx2aYKehvCpIaa6H+PXTP
oI9QkNsX+/14ncGPwDG74pGXayq+/sMSGeypdsQUsDVd7XOfitJ/1zj5J9Kb+JZ/Z/S5XBA2UDkH
Pyzo+LzKYB+2FWFZ2A9vSLhI2m8Gck7h1HeaLiFZ1Ox4CD9cTXVouETmxhMkYhxyPeYCSRPTZp8V
HiBiWFxfXTZxFEcd39APxz6/8fg5zmpnpb9BSkR0AE5Z7RB1gdTJ7QriiTb6FZ7/l+3z1N3fL29A
D5m+GkQYcFiTtF+torOb6MsyvRHPu2nox5CGQww4pQdGTnLcpRSdJppPrCmgOvve/zPhS2TK3Kf3
FVab4Q3C1HC89HakBsisb/djxrG1wIu218hM9ehiaineAk9S33/onsKvH0OCuJMivcrmuEkkstT8
h4oWKALkhqADgrjb2oKa1P0jIua2z5YAdvhsGvHautlgnSCeaWiLAurhhTW2PBZ5a99rzK6vtVTa
G6GYI2YY1dnvqEjV/Wg0o0y7j2KsYDz6oHNQnJE3c6Jwa55MCPuEbLb0dFeTwpYVRZ8SM5KD6IV9
ESpJ4lJABoFle21xtuMv6MhhV6HPBHoVAsQYjm6ZBRg5gAfCJDdhM0VFO3X3Oyh0bD/2IkTxnju7
eUW6NZv+Ow7858LNWINyolr5W/CBHg+TiZ2ohph6CMXGFf1gmdhvNSSf/pYxJSuPrAC2io4RcBYc
qH/4EQGprRUZurOFu16UZNcK8Mts9Nyk92kNQQL6MLXW4Vc9tm/gEoMH7bBPdK/Y28rfjji6z9yq
g+dKLkmnJ5h0+hZeiQdvKK/Ow/rHJH0fEX6tYpf60s6kRwQyIaZo0wEMZRBuWOBLk0DnUk0LPnaF
C5Hso28wrCniDwUfbfUfWji72KfhT9X4033BGN4WwoKGxEU8KiEmLZUHGw8tDqajK5IMOCx1CKH4
SoruZN+G+prVlQCKMH0GiildN42BEaeIaUrW2KydB0C1ky6qhOUf6UPLeQvUvJhRpOYXZsjkHv43
PgRVRPRXc1DE5lSQ5W3CTGEz3thdKtWTAor3XRtrC83Z2n1hDc9bLB0FvqGCOVStOi1+tYYWIoop
fl6VT5XrTvkOjIcCxW1zqPZiLV4PfIx+h5pJ2yplaasF4Kg4nEP1lJlxWCVTCMZg67pPsAmBgXUq
X9jLCy+NyFGq97NoH8Ltc4/Xh4819/Vb6LswmmELYxEgCXKm8jaBzi53c6QUZ7Yj4IB68lD2eXtC
GE+ziCaMkP5RFX/7F7dtkpne090NJi8v2F1c9VFKHF5n+bzS/ku3sp4fIBQ9gg9dfO6HrciKbDFU
B9S6IdyltX67HkynuMkNrzJV21mf1QfwSwk3t3q57RsgS8uvJxssF29wzC7vUrahy1iL9FdHfsBS
8kmVZwxzTgDhYDWtQVJx37X+JS273N7dcZ97eNhh9pfQSi6iWVRKBvxDd8Vr/BAowbB/MMIr9f7o
oe5CJHTYGYYDClXtfcv/fXbXBAGycXql/g+wEKnwah4EsfJcMlEtr7G5AEaSmkT+bMtDi8vi2o7C
tVlYoa+yzRXSZfRimOoiSMVlECY3V9OP9gj4ye1R/4D9KnSco5OIiaSkRNbul1AuIzukkuWUC78J
9rg4APwZQMobBzhWTP2sJ36jShJelw5kF6ZGsUnpJeDwLztXuP7wMqsR4a78Subp+Eee1dhI4vwf
Vgjp8TFRpfxRkKAj+zQGJI84uW0KuCyap6PWNiKuo2Si9EjeLHPrLM2ZEuI+8BWjqZsXow23tGfa
FXKkL6oFuNOXglzD3liiaJ9A5WBa/jSLkHmY62pdUUOH80Gk0Z/CWuACEnT5ZlOdF2R5EZjGeQH+
iXudCFvAn8kSojNFWwbJ1ybpKgrc9DVdCKRMGnbKRWpR+QVV8QO0wuBFboA/n5sSf9BtXck5L2QH
xWzSKDRipeRYmVT5VMZ2JSC2Y8+u/XhzR81LtzC1g9kIok9yMuQVgIOafVXS35pqO2VNJQf0qUBs
OcEUG3ZieL4If7uB6K6gT3JkerWnRMHwgaa3+h3Uf5xhVtRpkgKR1NuXZ12PZM2dLo8B13Dfm6h5
VvtxfEPDSXOwbl+l6HsfMLUBpzQZDJyUdPTJMnAUWEI69UfML3hpVbBEtJeN9Vymbm9nQ8I1vKHp
nwu73VYIqH1Hkbf+VZQs7yDh76A5HJyVzUqCBfgrChuqyPqqeZ4K4LBdtDRRwztxklpHaubLOMiT
UntkRF9KjqZKiLXd4qgU6TmRCp/X+za2Detfp0MTWmCjCv+rEkKaPvaNEvsb6uP8Tg1dyGQC762K
i7xDhCqLYa4QhYWpaE9N9kXN8RwaCScBiCwOn95JAh1ZF6qjDSXHR6yvZt0+8kFTOm6vCnlxeuB4
VzhfW391gy+mDqBL+kZjFEthNQ+kxdUbUr7/QXkyEAPD4QG9uSl3Q6djSyfIPzxvEQtX36MiBLSx
Hb3dGpcONb898fy2cKN5NnLgxgrXGTGb5YvGCUwBBw5tdiWl7TGKBIX1KK4QVvNWz9g+seDRYcYL
xUF924Zf21YTjM1itPSU+3tBu7w8b3DTTwOVpH83NRwj5eSQp51yR/C3wDXhrX9TdVP220FSSQ7q
sAeIe+p8Tf6lbK0GT56XaaxQw46faiBJd8g0q64rkTbWKlq7IY2OuZwSmnI3DPn/KJXEsTbl+aj8
RlO3mnqPK+E9RHKIA+WuFMua62oEvQDmEBhyUuSDqBCHkdD7jVKXaf4m8RFVrIaXQvyNSTaM+YlS
7LvWJcG83u9Q8Jodx3KB6oGc+ptHLO+sHow8nBwfGN6BbVr0G07anK8JMQUxPwazIBf7/h3z0h8J
geXcSKd9GWQRncVV79+Dcq6UhujQ7dQKTKOA4WKTzA4+aQlS+l48Skt+KenQP82+du6FxvLLjbHW
rkaXywA3MjWNw1sW23cKgJsOfT7luQRrAFKq4+mIYpqqcNViV8Av8MLsUuef1KQtPLsyUguB6nl6
bMOx5rK6r3miFLCDRiniaivzemtBpxleOI7lyCTgrwdjELDwwrzck0BioJ689N9aQAKDptMd+s8w
2fy/cZePgqwMDzAxZzNiu0VpgkQsQVUYEl5v2UYDlw9r+GHIXwHVV1ayYQ08/tibd9hRxAQFT9qn
CaRUVBqfqv/LrXN5So6D+ldTVmVmrylHk2OnYDI/NfrOii1KBpCJ34p+UtRCbJbVcPDuOU1ij7aV
eusAUh6cxjhIqbdQW32sWqqfRzjWhJWYHY0Raw66p/pltT/Qo2VAsbn6mmhBbOihBTHpV+fSGAKh
yC76be4jp6uIKP4X3hP0vSt1hdZPF1/yiaDBYDj/ruRA5sQVJS/jfudPkbpPTYNCywr/LlENgEV4
Q9tv8TrqetCj7errcAhBhrcl5wzUDReA13x8t+6N5+GuFXUjlRkF5n91LqEkEZPZtvEY6Ya2TYMB
chRWpdVe3pAEM0tWaJfFtl4LBfhsR0TfrRZ2EbOnvgMfQqQkiieCRkx+akaL8gjDgQ0zvK54Hgrw
rEe2xCWMtHqjIayQnCgnm+66neEL/g15uxcbWqhCjWuHhtoVYLikW4NTpdeAAWsluyjpgbm6aBTS
jKOIFX3Z4X+ly3Gz0Pq3nGSpTEQz0nBmqy07l92wLHiL6Mf+P5pj1687D5wEQtWkzy95iPDV68Jq
KkDiFvql7UMkfutwZzkLYhNSGY8oFAvH2TYrUAkJ5w80BY9uEOfZo3DgX6kOMTShElJUkhpLf3q6
1Gqc+gLgNsep94z37fmDWKTnveLzsrdUXlrrNBX8W/5QiVQbOnFGGKolJ/HbjZ5e71tta9pyPsOe
d/0u5yS7h4lIBeJOO46MZsbcA9m1h54ojIYCNSMGBjqlYftpPqFtAE91xLIDNuM7VXctQhbhUN4j
MW/mp9WEdAzTxAA+MJ5o3ooZWYN76kZx20VVBOGHUx4w1cy5QCOYsnRIsNEHybOVBGVclnXgSzqP
zDixr28Quv2LP2KKmVQwMtDKUxVxLlc+9G7bKFkMtemf/iPqQ8Xv6IInpR3gG+EviZVwyE/F6smv
lzYPLozfFOKtZtf42su3zdWPJExBOpwlU4GdvHM2xG63lajSoY8U3C0nkEZTSHuLSqBpm8wUDXz6
FwTLxNFFAOJA9meVTT27KXCkdNWokvoZ1lCO7UFrD9+UROPvxoCqGsLMMHZHgpktJZV0F2gwyzpe
CrbhWKoeD2rWZnqs3Uax8kZpRx15/zmZ7yna3l1b6Ybl437v5eQb5FpOv99aaQzyotkKeKzySnUk
0Pj0bZU6nZxoWZJJMkmfmY4trWdCRUebqAuIDHtT//f/ciJtfxksYaGKZ+zEDY48TWcLCuy98OwR
YmtYqYCQWDxjn1RMPG34ROSZn2B03lWLmpllo++M9+6J82pA46eOM6QUMPFp5lqrDKWW3qkOOOo7
4MG/emDALAAtQHJz4F7JTxhcMJf13hCPGUuy6bUzS1l7ppfsAEi8UzhWDFXaOhkU57jM4YRZ/03c
ON7CLGf5RHzedipDO4cToRgd5/k40psb2RYaHYyeiNh+HCrhL3dfBXjkIxtXWmhFnaoiHrcCSqIe
HaEqZNBgHzR/lFo2SQ+4VEsCDkr4bhUpvMONBSHCdS+4OLFG08/Icu8wKUS12gGxDr9dqiKDfGsD
eAPzi28awMiWQKGKEk+exGEiqLsnmAJgJtIYrhZB0kAKSHu7hwB46wmqKgKd/CGuYzkx8FkvLXy1
e4Yzd/azwHYXx5DMaBdaSl2H6lJKJf9948h8E6o6ZEaRp4S1rcbCjAXXL0nXJ6rIAV+7P0aEfRv8
VTRKs3SEidp50AKKf2nhRJBCyMnxEHzF2e/mPRY+mtEd3tGpkc9nvEgwh+eUs+GMWsrWiufWGqiX
wPa+qd1aDx7YoBDbmcB0h2VZm2KN4BGMCTQhvaM3DORzQvqPFAXBPopzW2N61DLTV15dc9VEprxY
fTmtjbvtouNoYASKWgAzrmXZrB1A2buum8qBHkjcWVNlCOq5pffDzg4j5Qs+4jwE8lU1oX5fek2x
0cWORkst5uffGdJsuD4yvnYoMr7xq/fa3zTKHJ8VdPPFrKmR2PpD//85BQ5CrGXJJZOGvK18/+Bt
1P95wA5XW55aeqGILgWfPT8P0IWBzzNB/LEJp6TtrSRPSRFtoEZMCTwecXAATt841ou/F/JDxrEG
Y2BGIouKWm8uUqi455wiVaeVeIrTO+DH47FB0DS4U3KUoWSjzvXIo09idJClyOSAJ8le1h1uWp40
y520AQZ87sfM3k7PJJrmd2rD0L7DXWrjp5RQ69td5O3UNHxIWzSFebG647HTqP8teYY6VFy6hovK
sxuByBApeZe3TPihbzpve5vfq1zxhvXPTaGtpzzTTK1k5tjrth5ui407oZhiQWbp+wEBr2ktg9sg
WRPjqxGNJDWNvOYBopxlyFtDgn/A363TxskdUdRLybWQKw9ihx9m91hIgLedQwcXAc4eubqmFLRJ
JukzQrC5klf0CFYZc9WuC0hWrC+sOESkRQbqj0+RKFE8BDnToonLWtqCs1dl99SwpVPjE74xE6L1
5M72w0t158paGI9J4bRYvvpbZ9LP5SslAA8laLd4mpSIG0R/bQ82GI2tSNl+SC0MJOjWMclMPnjo
UXeSu29GdrB3rqP7/1LQx+CygmamPlEBvXtd1qt4nNRwGOq7/Q9LSbAijWOMbB7dCK/jwBtNujH+
1Lv9FyP3TYx3S3UA0JDuYWyg2S3OR/7koltMrB12fdR7OZyxPObZ9pRU/vweQM5t1Hs0eXnPvXx8
755uhwOsl65NAGoWrwHGf4MxFyH+SpKQwRqTnWHwyH2AvNjXzdIZLi2SknLyg2lrzPsuTHsxbjBm
6hL+5EMMG8U5zttnep9JLi3S+gmtbYhIi25X83ZR3CN9As1eYgSeBVw9/LEbzXUtOktpJXN7XNQN
S4f9qAenexjRENRSN3FUw9ruNwhI6oNKpjWx8RzXJwCEdChBdNMypQdndHTdbdIJ+rX78l/RHkiy
wVbATjoS426NzZDZq0dUS2bWPAMHKDVyc5LQSN6F0lEq46AjL1Jl8ehlcpdIF4w3qNqI490T36KG
11pTE1qOPOx3ZmF8eCDb9CAutnE8YS3XxCTKmoZgS0SU9uu63PK4txlH8ZWjcAJXCvhtRSh0gl4Q
e8IFmj+HQSezeNvpF9RGIYiTfbJVz2ppWQkgq3wOashMrpQUVMqxG0lLKiFlUnjXTbR8cCeg4OwA
u1OKeoAdkngipd5YqP4TINMvw6VeCahE5sykcV/HL/02q2N0H5QrzYQfTIzD6LVV3u4BchQ+vOBb
GgvN+TL9X5hUt7o5rU7/YRAqcNXpyK2kXW0IKvYvLDgqzT7aoMThTuY1TNH+PL9qJVVoP9sAR1qj
SazZ5nCRNTEa4uecMkgnsDvEluzqJdZNZBjbxwV62j7ibj1sIzAYqBUD/hjdAv5AtzvtH3Cr/uGs
nXwRglwdno0BnR25OVn26q6WVwejRkxDcs5RUox6uAoufXNeAAxGtBCOTElXFsr7HSuyiO+qUPcn
Pifa3XwQszywHJCZMFsy3K8wILsMv8eui2oYD6NSWuqWNNxl3BkxJsdR17240EIKeIEaTIoChTPw
ozuc/hW/+pQsLKsgj0RytQMo0fTif4hLgJxltVx0HUXzyUSSmQbo3z3pyAe6Mlhclpp54wdpeKDM
8KYq4eG/JmSBB/QdGhes8/Phjg7Un6j1+eFM4SW6HVbbPAuPZrAeRE9s/AWqJqss1Sst9PuDA0KB
MAXJmSvQmx9Lgi9ESyZqsSFKl2bCQEAV4xFUMNgDDlQ9QOWCGdcw4RPlbB4Ns98fXtMwFrn1kch1
ogCsrmdfj+4v8xx8Q9Sqk8pSMDV7QoB2lxudGcEmSUWxTqyeOnWPU5aOHI66qiWGKWk3mFEwL8tA
AWfHFYomp8kJmgcP7OwjYVIPvTeGO1f5HV77FIhJPgf+fiyPP19KnPWqR5l/wWBw9C3ozAw3Hqg+
Q6zB8t1omlngjWbcLDYmeTwuFTidv7IvrLgbnDLlYBaaSDg3Pcc6urO7hsKhb8yKehPS+9OpOzmy
9OIZSvcyRUeUIFOeOGxQqUE5uzYq2+gnBSRCtMHbhrYrWNG7gpJRXRClNuKh2ZMwinEOAueXZ/4D
uLlHT6FzsI4YKjxxVLuhu/oC/iCpgIn5UAcGSQ2NZgnAksAKmgpeZHYHh0s6ohcfYLEmSK7p7e1Z
vn7i8pb6SwdGjamdly8tjlLjYFq6KLfJj9Y4iPoMyaaaTZFGvixsSM36e4jLbSjtd/LM3cF+aERe
197q2K5uD/VAMDoyKA1LpV2ejDk2H7OglEmmKQqX96wLU2IhIsOQXT8yel+AhrcuUNxUBjE6fqG8
Q3z/j6ktvUICFQNAwrBvqhlgYsmHKU9kgpo+DPFz2w7zseoWfj0kWFzVxuPrWaBW91eU5M3AYa+0
9df7f4rfXbW2+BQHrLZHtr1xc+0apLnycZZEaeCzPeyHN9YOQyjLGnSTgNQHTH8+ed37D+QM2SRv
akUW6Gr6c+ith+/i8yw43eXU9JfwRZ21DLxK3CIR4D+ozkM4+3chPV0J68Lrj4BVZY1GeNLRmjVV
UHpmKt8DtfnvidS+pQzL7dd0J4kLUHolPLjIQFD+lzHQ/orce2SGUcUzK7GtObpgswZWzujuhwuI
haQWid7iPP462OBYlJSiUUb2qOurjv2mPAxWKsSxL4+I2kXZp2HSlfxOzTgeDi5ljH/kQMlkTUOh
a1MHvE2yiTZBSbVQ1SD+hpVSsgUkpgiBvWcEM9Li813laDxHS9T6oHM8z6C3DjNW/Asb0dE6iM63
d1PESlkLQRDfrN5XrvQDb2Oy1wseixyjVy4YI9ba3yZLKp3qzzfVBn/Zy2dr5AK2EUNKuZ34ymaB
YWJTXBu2Op0Lir9cjfOaqedHmHkc/OoEByfcGySP4DijwNjVHPVu2YauxSI+epKsLpKLv2R0ta8D
JZyCEq5GnNRV+6HubHAri/3/89Ke6CAjqtkLX+qvxqzIwyslMGTSy1lfhMoj8DNg2/8MfF1Smaj1
uacyXN8IvlXyxcy47s0fs1/Ik3NuK/U7HI47OzWhfO+fRlfpRqeJttahmrbgWTg64Rd7bG+LXQ5w
yqk22EKlrJoBVjkF4hEJw1Jnyf20pryIl9mO6O30Me7E+8ZKO22x64E1GnkUvldXNbvK9IyaN5sn
VbJhhJrYyqv8Czs8mWPcVVutiIG2kaartMnhSCDAHV/Osje01MEDqykR251BvLJ9hgn3U7FGUwDS
taxoUHzx2KN6eiN/Te5bs1Rc0yAEDOrKFVVY7oG9QB0ciKCuuce8wz8ey2RBp4z+jEwixyIjAm/+
XOIhiP4LGQMBO6rvTmloIR5PefMnsXCLoVbDsTBoNICmMILcW8js26OuGNCsD63ZI6YbhYARew2f
pLzJFZAPNqFE/A852RClbGrTKezaBEGTIcn6hiQp09OzOUrI16er02A7PgX7xnfyJkJAgChlxBvj
u486Tp65neaGrWYzbEhud1+gmXQupRRclq32DboRcYzTzv2JM/mp9+UfebsPfugGk5w//J9q0JBQ
mrAgJqopRhun/rAjjiOn7SXro8JZcSQLRoVWE0vWAzhyjm/VteVhsndJNWWTv4GjrtFzj28KdebL
ig5YiuR7qtNFScRJu7HZ2T8jzbCwIoWGV5v58Dw4Nk6hgduNf7xhxX6pUnNYDTaRuW4O2EDO1aDe
5ZQ31wZF9upun0fBB/vYQQjpV/NWLOUmP4uY+5Gkh127p3XdZk8mndZUQfjGqvca9utbMki7m9e9
FZDt+U0vO9gFWe/OqxN6JmtVmYErxGM/RrsjT9o96oa7NxjRLO36S7K367yQc4iwddTImhzNLAZL
J9TciUL3NJBZ7LTg1deDpvARLXdRXxD7op2wBwsUKDVxok3opG2VgdaSwZD6afADKRenjuGLWvuq
8CVM5v747yN6p2j4/u7UT/miD09qODC3+jcVYTgrfDjIz3+zKQ/7dDDzFaCTH1pgOTgr7XlTKUvm
5LH/ezcPHlV/IgxiC1Uc6TvwWeEwgZDxealt9Tmv6CljTT3P0cVVru1+bJoBRl7gl7zO6UTVA7ZF
3+0OXjnRR3WLnZIe2kUaLAwzl5hL5bLTO2OZfhj3e46lXR5wOKCia0SkjazdCsQ8cgfURgy4309k
xE5e3PFCpHybQbU2WqlX63g9vK3dcOpEOZlLj3RYIySCOF5GN6rOFzQb0HucybTmZ9FaiYr5CtPv
nyzLRi9wO+HBN2CC/9Q9I52Xqw9o38OOnbzrUWHXgVunyjem+/F26oKV56UigMN5owFKBW6AfIwn
ESN71JHeXeDqeTykHB/9Ps42S4bVlYHI7sqUsuYdoffp77ELGLlMDGZRvSmln6dq0E+5HFVp0RPT
Ypc3+50GsRxwTNE0SBDsUW7EB28itVq4DbKYpeXuvah2ve6vUpxmJmUO/y35xr+S9LYkZk+My3z0
q1d5/OKRjGGNUPlXjAcrUjfUTcqmltOZVFN/o+r1V0+F7GQM9HUC0oC4u6JC90c21/WE0oneUJgp
FzDuDkBG5yTui/BW2EFI2umH0xLw9oYD4z0Q5mwhjpphRnggebORECVpJrXiVyR/Z7dzJAnU51XI
QcCfhfKNigF1FVZeR170/7kgBNtSFVHqKiqI8FDdsYJ0at1k2s+lSdvJ1qFRBgM41g6lbUmBxCzI
byC2pdrxPHiS/H5c2hJyJfChbe1SMTlgVd7jHO322i9TDX0/rF79S0O0kQOvK8fSyjfgGseC8ArC
zTuSr5zZnKbRZIsHclTi58+AW8J2A4e8o7IF3NNMWZKoMNRC8DR09t2oFSugZOKxImtquTlUYg69
4uhWzcO3v0Sq+GhgpSdXvgU07PFPEgX66xJmpm84CRDqKjgT0XkQxBnTPB4y2qbYcESbueWzSNES
LwUOyUELGN2FW6jZOrNIPWafgtWYimgc+gaMeKCNgCIQyI3kiiBf9LcAj5Kw7Ng5TBJVwi2Z8AMi
AgycMYZDUydVMA9uysMLuU9x+hqhKIEqgzcEGTiZGDUcoQvDOtyKKAlgJ8W3G37nsqYSk5HM82DG
oT3K3dxWOTQdzdt8nAI/WJTxhgUS350T7bh87B5SVEMkP7EyqGAZDOK575YJ5CJdJi00YoXBR3e6
MgmFsExmVWKatfzAdG5Ea+7XWZAk2DT6b1yPzolY5IExvYFQ34CkFGqZzbYurrOTi/rHhObVAD/H
OhQT21ybgTSrPH95TTnxdORP394AeJO9kJIGR4leqZb7IXfXzkwaDT33wI3gejcVVDuiXqXZkgaU
z2N2ldjMBsrWo6zRumiUlAHiXdda8S0QU1j1ABNYRYItZOndC88c1Ie50KO0+DH5aTPb9s5BqmPi
AtadBsCwRzl1X6aCPMmQdUkuOR4uExbpbSfLMZkBmGxNXOOoo7kBl9+gVci5l6B057MQXZj0zuOe
KdpDAP6VjvKg6+jxq7/dL5CU7nwDCk4wv9Wh2ot3hORUKNRZ/Vv8DtYntmVcW3M1n9g+V2q4GZ5v
ewikNKHPjVJGSrhKnn2oOKpbfVMFkPZgT1TFkbmQsseRcWxZQLh9bEDu/KbKRdMfJLfYr9HSxWG8
7QQXdKizCUibsrgtv0otEmj1w9apr5O4Iay7GZ0k0U7+CcdLgJkuaHS7ZX+hvtthcRXVgUc3BGZm
4fqgrcRCLJCTgp/Q6QpBcclUu1h356Nfqq7dp3Ihhg9bZxRD2uCYoHqpubpOcnlvrikhKlWMgpEl
E1ULytBozST+SDpXpL2GT2PD0JTPg/MFp7yHtHrxTT8zqoCWB0UHWo+qr2DQ5fn/dq/FGJwOKqeV
OHJG7bMz7/SMjA0k8ZE0GDHJmxn1TkKrWazwlOGNutp4l++mLcMgBeBHVKYGNAG7OXwDKxKxFUVf
drd+gqxZuLhJ1dSjv240musCDxUXsIKGYiccp97X22aoBgEfSFL+u+igWycIWbSyl24fJ+dsL/3B
w5/C/mftL1QXYiNQq4ATMtKc27KkXsczTkgE7O0SbKBt/BrSEJPqDzYlsRR96PklnDcthPE7zlIi
RoIsAgGthPC8mnK5IsFszPSQyZVFio+DwxKK9IvTxyEvz5a4w3vgYmMXEG78nf4Fv5+ItUMydCcE
8HOjcgLu9LM+V+G3Sy2q39fAF16t2fdgyyTU2lPN91/SAqp2EVxnVzrHE98kGdjWrBRRC7Ui/j7/
FFjCexpiF5N4jrmVYK9DcnIpLs7uG3GcvynHjv87i/PdG0TGLqVnKGEgYYNU0UxxfT4KUkJs+2jH
68qHP+Mz8J6yfwKQX5GaSW/GEte5qcBI//Bs6D52egKI2ytISIQv3ZWTI/AcHzY4k8aZv4PnhKhP
+HDUf3n8LGrTSrpqChFSHOBrVppgDSRo2IjbY6ZkQygBFOpChZoU0/WRKCQFJUko9bJhPzqWx1Gb
CHQx8hR5jN/JthRSJXfD9hScqDYzLbtDZoWYWBjMMMbv4IJMht6HCZQ7Vajozph5FIN8p121xC0T
6CK7ffxwN4KFICMxtdgXMZd1ko7kqjKvyGFekiJM7xMmaHuRBc6OO3aYiXsOooQEoEkHP8jsdMKR
qjiZQmRo9AA8AAHNen6N3KsRASbyYrS4BxFKc9e2S7Dz6WQx/rVWxQXyDLk7FHoH5epBeD/oGVMp
QNW6b+9C3QdHbtAXRqgi4TUGhUab6/1CUn0noKVDJvTD3OL+dzAPOV+wHAQKXw//BrY755XEQx9p
XTaYaEgcu84QRHU5WVZ93l9jpl2nd3nkpDSEZlQ6Jvm1Yo0PqR6izQ/zSpkSb9sglMVVzRjNbcnW
z9FPUJ+3ltxttxdtv5Fleb25nB1yGCuZHoW2L9v8uP2YCstGp3gcKiOX/H0AUI9i9/mLYusCBiAH
ML5EEgzOcL8Y7eWSeHty+oJH8MtDROKkKERG0w+hWWBDXUja5FDRzWeyz17wrglBVVR2QL4+hAJ5
BI8Fwfo1qdCOu7+lWrP2ijGkfFKJRRXr50ghaeQJuell4aXR4YKneiUisux5kV6cyqNTpW0RUpd8
303Oz8ULDhH2u2Nvwed+pwAh43vIa4GczDKRklhZolKO3DsKJm8iALEgXBfyQ10RIp+uAGwPxppU
/lBdZqc+lnyVV9edxxMEQKTKzygTO7IK8nch+u4OXzTDmBueFFzLCaBKFeFomuMla/QmEvWaOBLh
VYlkoo0Axq5SiVTM3Zxb7Z8x7rPj+T+t2FuLun4yv90tkw4sweTpa1qyCvBGb9MmtXFFS7C5TiQ/
tWV/Y/hFv8wQDMNrpjZJDDchOnVWaAwehQxg/qwaderqr3ZDP206LeXE1Bjo2nqLaZwUPM90xDp5
h1tC3faZ/CYyaU0hdUlzBAi+WloPBhVW6rPcRyMnGqG8SPBFvREV3wZ/ORnu/lfEd4sg9+NbZf+w
fh5d0tEvbF2+GkY94rLdlD9Rb4CRCljP/LpdnODJ8ubnrFZlC4fRdYWLctL5kpNbK92q4PZ706uC
6pt88T0thvyan7Vti+HKfoit8gzhdeDuqcN5EcGEwUGHHD5Yfd5GWPulwcGXI6QYWp187O2K6wsa
+MN0LHPibaVttwzVx+22USaRrvgFnNUrSdI43doHTc2EFnPTUJ0RZZunqcGYpnsuirhtmfijpM4u
nRvlepzSy1LhFdzq1dx/v6IPwNZ3SmRx6rNs8upgBMCIAEOGVwcXla9ppmLiBSvM2ICCamhZ4QwX
LW1lrbnUfQR4n6FNltZ9Z5xRVShPli5kqB87h6xBCOi1eS3yOCbs2N8oVDj+VxaGY93Az1HU/Yli
tvCxwsh8Sqp2IVfQp8b9VSSUHDIj6c0LQrdv/UUy9kM9qfCyN40kMicEpku8AvbDOqLj3MXE9gvO
v4RGfjs+qIexrGkEjmPCAk05NVK46CG8W2eLwpKEudtB4DQI3V/LyPLYo9D8W8OtAaYX3WieqdFK
zlducK4FJ+yqGPyKBBdpZgN35bRGYY5dL4JMe9ac/Iux+GOa4uzoPPzEHr03WmU7jBZcfn1IK/Bp
4QrEDLbexMwxPFmswGj6kLQmttPiP0uLdzzDfzY0Y5Rt1APkC+N0SurzNz12BewOmwmcb2GOmUaT
0fnOKk5elV8XMN/RYBRB8lCoVM+7TiV58ciSrMRN0iRR8VWig3uzeJtPnOzhDsgUnuWNanlhEmtK
dJ1QKcx4DPHsUMIVfdroaliU7IZ6PF/Kg4GQP8GqO4YUIJzP2b06c9G47bVxONYMryOISGY5+ocx
H86xPRkizfFveOKh1iJKzNCKUQPE12OY+xnxFdV1YjgFf5wiepe8djhLF2d/UGyNqFoEEfnGJFLA
mlpzCUPtMpQ8Riax3c7IlxVYeAzo182ULHU//OOpvM+s9HWc3WXOQAzrMV5V9HiO8Cab8J6CglAj
x+j5ONAMC10W3rnN0/txRhIB7dZNHI2Q/TLB5TK/kM/oNSJ7caVpSHTsMJm+khsDAGxoTUgxKxqb
1gE/SgLEg0LDn03ypRqr+me7lmDcCDmkd7E0YmBPxQb9HYnsVbJbKrZDCtobsi8l8pbk4qP8WVf1
5hnDZTdeNRXmpgKTNZW/8Kb1v1BZdQNZ7+DyWUnHGRfVe+/6pojBPzzbPCFxiPrRh7kvAbkXEE+V
DLMZ8bdFZRv3SZcHMlbSwLseg4IkreTN7tQDAUJCzIDySmjfjmRgjPrbTLk7hLSnbOuYeCxEzbeH
xwq0T6Z2FKncyCiy9v3DC3CH/if2ObOKgEk0+UAVfwP7iYFI8Lea1b4VMBzqusmZd4UEgoCGJZlu
f728MufMjcpAM/LCv/OckQaiOhvtOdqMHaXTw8iC3UTvyYD7eCdgUjyJJOpUbxKlUuCZcIlFse8B
Z3ck5YXsiarSMnqTSaPXePxeuGbNKIrluj0JA5UB5H2Uf5Vj8pUI43ncBqYi7ZpsW+JNwaSPkSHZ
k5Uc5wg0cIgzKboiztJXi0zJpUkCLcLR6MRh7H9ObwY9EXv1vfkh52iddf1Qa72WgjOYHjqGYltE
P3eJ1ND/P3cHWVymNg4JIFSppamrcOprvbMLrdIeGJRgnEs0oyMvmlZX8YfXGf32A+XLqIYQmGXR
LT6sU0sMkRyR3NyjFCocJs5Hmr76eZLczcE8tNo5BOlaX1yoDGKTE6H40D/pmBgBXjEJGRgMEuFq
LZ5bA9PX50yhJcpbdMR6SPOdzwqJBm66188A9oTvPudQCKFL1Gs+4IOTcrXvfV8vgH/PSgNTAE6/
fTQ4bR82jOzNs6a1OZgm/JlzEXBTY9/CK4q+cLKxLUGorEs9Yf0axjMnf02eOZwDGtMVPcq5lQCO
vRkgHSFlWVhRQbkBQk/DQDftXrZ40Lj/bfnTwss7FHiSMPA8ybZ7QtP/P+o+yxVJr5u3Bk7zs+I2
UD84VERcBgH6ZVwF/YbNbKV3lfuRuSbkWRp9y6nx8uYlmnx7S1TUu4M+jxyB9uQbIwuMvcrIffCo
b6OEI6DqlJs15Vp3KwvFcF6qfo3Nz1otQ/wPoMXYRQJnwzgmCLHuzjCXRm3jgRkaVFup1WpsN1RL
bX8sBppiyHWVlnLXM5jm0p6KQeQBx/mLCdq2c5HYt6gSBugyzXNLkJFPSQ8M3Dh+THThqHNbyIw7
LJKq1vhGBNMMeWNLluiUzH0wyoGzcQ9z1zhwT8Lkg1dJXkmU0rtz9gV78jsmWR6D9ziduV7OPRZh
49AgAKrpSFlLhm//KIJAuopQZksAL9cJImW3OQUHNLQQwmCPj9dTU9aS0ywLvS8HcZtO0BWtUFaW
l2x6tj9MjbMgKWEXD1zPNxrqJt3Kr95Agf8CLU8dXThCNdLW9hoQ+z8bFuSaeDgisi3+Cgi4at5V
CRW/NoYdSCJbTICnV6hC99nN3hQ/U+RsYGKxRU8/FL75QyEe/NzHjswc/T6fxVPWeJpucdSLelAL
jgXAzBB8L4UFQxcLdrpAzMlHNSGpL09FDNBanfCcUd7xQuoCPfLoLcZ368vdpNQvg/AbYM0lpmy9
XvjKbQdnlSMwrcrvFTVukehbyEyy6OJHOw4l3mAJZAQoHs77epnb1pXA4Fdrh+yAwk9V93zZEQuu
FRrig+LFvsl7AQlg03/0wSD86j7ILYChRCJJfnq/ZQ+osjiIBeVGGgLGoadYAqXzJuLNCIbuUTFG
0+ehwUoLFbOt4MHHKh2Hddd3maTN8LesVz+wr53Qyz48WzHoyl1x5DrLfJzTKWJ/4gcHXX+9P6/Y
g3Qa1aNE740Z0cDG+WUEVW6Mhs6UiNyqg1IPiyVUqsl5BMTc9InrWTi5OPAa/GMct7eYXu1xEwHx
uEIAP0xWnSzRwDqOXDMBwTBeDRhJG0YO6ohFUVlCNd7KDy3i2xQK2yWPdgaGMI9ofnM2sdaNd6Cm
nVYkEcgMx0UTmw9E5Nz6bfc+N4r0ygZjHmOGoQgtuqGqfCxfwA1ovlliiBQmIB9f+6Hz6MPgmhHJ
pwTzjgBIqQYmmN+luripYrFNS9N9BdzUUAgkUrW9bjAW0lJtJLoZUuTIpVtum1PyIQ79gz6wMs/X
AWfnRvXraNeXI3bDBwD5cRyvkLm09yJJHupVvdgxBDksZEyRz64n0ZiA1RgmA1D0b/5+Nyuq1VWP
AelK5lKe4jlOdR1B3M3ed2Cfs+/XqH2dFXHmpW/OUjfl4b8n/c/ptJrj0/DlGvqK2qD57EOPhdTu
UYMlQmRAFRAAccEEsc01xxZDh4jW7u7gBzeJJO5/b7iDOpbHyuUqatQ4lwL9kwqLobBTww0VYvTa
CFN0oCa+aiVCWmRbtjYXkALPyhVwoGSpZk70YiWvQ8Ds4KIEqH4QPqb0IYYg1TTZj5jvqpfEIqC/
Fg0Ja/gmxdGCtZD8jlChThK6Uv3k5eYV2Ji/vdyo1WpDjMKd59sFptd6f6Xg2gxTUfHoDTFmFH0T
HsgbZaZAUjQZv3hXKX7UKeWIQSxcTRHYGkzmNEkh+KKip+okd7wn2a8p/uMs6jriz8goET8Lk5RV
X8doatUUM1VM8wfsxsG0BetdaGhrgNP21HmXHGqnf1RxLqi5YVUeW30P443GMzEAHABE5+XIuXOq
CLDPxf3KuGISZ5DAagvF8WBIWfnaJPYCl4rt25wbd1VAYFKp0AEKSClfKX1m12dZB9O5kHR9/dzm
867LRW/RL5zjGcRQNsWkTKjVe73Zo11h5puSYAqV9nV7XoRGLI61CYmSFbJVYZO8+0WW+Sl9I1Tw
7bDO5pIKIq2+BDYO57/PRTskPj+N6idIkXVkdIsncNAhYKwerybNmNkkysNq1UrdjpzsRHtCORWj
rPQHQ731ZEl2uiEtZxIf3W6MDZrNf0eBotrahdnXtvDodtzZAlmaelvD8palNqaS1gta75cJWOQL
WlrT8O8vfDnRzRHBIVx16jdZqFuWe6QM7ai4Ti+BP1VK1CChkIubuh8bNjJD5rnsEsrkvltK1CIA
VZhRMF9FGMjU5kc5kKz1oBcbwiGEGn4rMSKtv9XT+Z0PS5Po5sirqfJuSTM9ncC+2766jXEDkPL4
e2kxQ0FTdxrzVjWx5NbwtI4CDxTbtgZOqMLttsJFNp4qomVEOBGo76WAnZDQtKWe645lzpl9Mt1L
lJH83CW9IOI1EHVR17AE5muR1JgIS3lVVy2N+8JWVm+2ZdyzgdrMynEe0r1foOuSxYzSLdAC6Seu
FnhdWDXibKsDXbpShuZ1Y++tqqu3NU8cQ4xu37Hn/GL0Kq8AVNbCY95MjVDAytgYfs31geXhwK6z
0nlV2gANeKolslJKKemWLPSCopCMQ4APNmkBiBt1x7IMvy6h8CTDkg7XOb/6y9hfu/hu24Brm0m0
jNTy7pKSFoB7eznw6ElWqe18qnwYXifFzDq552IxPPmW3yhEXT/r5vNjq22ZxiUGXT9sMuDdQe04
XJHZbSHhpXwaAQ1JbnlERlnpZQvdEzJSeSCUxLb1deTl5P+8siBDv3fKAmIB0qHj/prpIizA7SuT
RSE4ui+WwEQocoDEdKVSyGsuydU0bsbxIm2v6POaVdhsHB80KsiTiq3TiP+eTj9GynNnc1+XtQs4
KwPDlB4yM2GdaVy2Ty33nO9GbH/YzU+TrKYVBdCnWJlySlUdZRPg5UnOj2kbRhlb+Zta+cHRpTHQ
m8AKowFcAuWXt1q+mGPsHrIyVn+JLPX4SXvyYpGiwLYN36lZrbdwPxRWTVcTJon3h0nspxhDl2Tl
gir23tPRnmWwz5ICsxBqw0qx077Mmi338CEPvVDb5UNmtzSFSfDJiw5cOH0IQM2bzvjG6z8LbJmv
yDR2gNGAExbf05UEMLeE8a27FcnKorvqjzBKsCkPAX1tQAPbHvgFl5AvUB6uFp4tsm3rYST/Ll8F
jJQtK7oIfsi7SDFyYkHp/yAV3jb9fnYSFKboKRuo6/l8oaYSJyU22mywCdT32eWlirpM762R7IRi
6Eys1ZhFIACRZ5n1l55pRgV8IV1kIs4fXRwB4D+SIYW/rc79JWL6tg96o3iwHHA450uzFCooOW69
XwHh8mh+rdPpd04x/zX/YHjAp1Du6MMXBFGoDG3cQYVpqhnWHcKNFqamKS2L40em2zdwgaawFHE+
1i4+mmVAfTllCSvQAq6/cLaBjVBL52pZkLmB1izDPGErv625o+6cUCEFzKdYbuHovICIao+4QHoH
aDQ+dfG+OyWEdYJR6E46jgYAlElQIPPviB77Rt8u9ytF1pO3mxFs3l7SO2V+9KRPonbcSsJEZkyU
Uf/U3CeuvpexPpYbwgtapZctVekkaIA5lIhkQgS3//K8rIoyn/iGTgQdHr227zcqGJjxzypAme5c
pEfN/yzSptJRMCahbyEtupg1KxNzziXKnSN46dSHLwvNTBW+VqSZTKiOYvA5zhMbUrLCRLLJadoi
J0V3j59EOs4/UjAnRf/q29ulXegeRC9AdY78FxBAwk28WU3+/rErlhO0CTE9mIy+N2g6XQRFOHNB
THa+9qyvLC6VdMVDk4zInejMp84QLRBdj+Wq5yksQTWQnm5IuL+vi4PRibS6AADyDmYNaMIFfww6
0UEQusuceDtAya0wrQAJgiJP5aiyaODxWm9PL9wU4z294bXF+yXW00Z5CjEV56F4I8zDnjrjLqDX
WCfW8UhwAvXg2ZSrriGnWr/r9lUIus/5ZY1hlyte0AiFPgIWyBRNWK56NGn0VUkbWBZK6uQp6ZSE
9T3OXAt+B1NIimgx/8fAT7AH4mDeJ8pxOgK2gCBjyddrONk7tKLYopjzPtYIjukbE9/LwYu1Oqek
iq/kDF2zt4dC0I6txf3XXgzkgkNpbqoHlfMqR6Jc01L8bbJav6WDZqsfmm59Xm5sYvwe00H9Wbc8
tBmKP/1IZ/atlaNQnT/NY0GxhyqNHrOAmzKfVf6NvIeEOh7cGcrVAXaPdr4ZjCQempwSnwQTlfSf
nuU69ov3Qzlq/Pqjf1+H+mZaXNiLqODZSZ0JDgLhbjxHP+WLYBGp3YumfrRvdAfIpSMaBph6nCph
DwkIcNkBY9Cm0uiOYXV5PbBW7ITy4H69AgRmn2ObiAdL+xlouzmpYk4fnlpZdGhf3F504nvaPwFJ
9NswrtLUvTohw9U5P9GuopU8hrq3LfEwtZUMmsNcFoVqv1m7+T0VWFSD/N2K7fw+2vuHJAPQGOgZ
Nw4ja6TkDiX/8ldrGqDifFldIsFuXkoXxX2wUfQfbSDeoyV2dYeKiLN4MrYlfG2L39zjVJ95hZF2
zJHsEXvbRgGG3fB6sUJx2h0tPgAaSEBptMVgS6r0uZAc1HOJOwhokLpBm5TBkizkbsmOTBxxXjHn
oXkVz46Dwdr48NtbIbfYjvaPk23gMpNP6KuHox3C/pJdYx943RfsAIJXycMAuTdqZsxaI6GTeQDi
KpMZqRKvZl2bbmhBoEsWWrIhBc6r33LhAxcOi9uAJp5OPO0X7jHF+08ITDy/8vcCtcV+zzvXNarx
nfBJB3qbBeiNZNPGzhpHUy0hNM6BwIMfdLdGXX5ITry31gxBA8P6id7moTjkXCIKCul8LdyRZpt9
foOG/rFJWy00fL6c9wDa4Kp9i98WYjGOYlQ+/GvAYWzFfxu+Ezv4ATQE4UkPZmbGRmN5sRQRftfo
GYVX+w7mNpaw6pbPpp188vD0rwoTgazsm2t0l+0l7SNn5mhOTGOcQWOfQUo1WmqxK44BeeFVKYHh
PaJJ+ybJS5Qrd80w8gQgQS14I228Z2+CecTTpoh5G1UdmOULHB9I0NIQHqlQ9VKQX2PCThlpPKDy
TiQuqCwU8RoPcyegBUwgnn4d9EzS+NfM1i+XHpONlxvQnNAud0JvD0OF12Mr359cnGDKyMepnrpO
mEF3HjPMWReSY9mntN4ZvxFldZO4MPE9DLZ2uxBdlL6/RTohjYP+H6I9zLUX6vTcp/uAu8q+jKLQ
lEjezfnsTu7oKYSRUZUrMBUqnvT506YVjHx5nnrKKC/b7cpM2NXKG1djQS4v7MMHTzBj+ZbV7C63
txWypjwmakgi7K8vagcejnCHOoTp9iSc39lTetLJE0uZ4FHbz3OnOmRk6ArXPlNgLv48I8MDCUR6
DIAsy8a191uYHhM28rhgMDIpqtTuRRhF/NOgkNJrTvNtXTz4EXL6wOJwoA2FNSWTvSv9+JLfwh/6
wnypks3cwhNJIahkc//ZMhdf3ejvC1Tv6q56pHji+2s9Ql21et5w7QAa1geoIQej23US2FZ9csOt
2dgvwODZcFmAi/uwAk5qEdgEjHRrVCLJ156M2ENg8uCYT9jAiHdFU9B9W1iYgZoZEEncbKjSJXEX
iUkewHejqWHIf1l7ADiXnhcJ5oj/viDHLgPW0Y1rzra5TNEHgrMxUyz9YQKI1mpgGlgZ8t23/taJ
rLu+i+NXmPzEqlnKRkTiq87lyjAafwxZwCaEffMnXSlyGdwFcsa9cj56gBsw1QpAARDppq4CQS1s
v2ehfolclE3cjfxoy1UjL7EmQxT4AVCqew3Gr+gsOCRb5jOTd0F5dezRAmzHYL0RjUw40Eb5RO0d
ksSFzJrUybLQ92rY4hwPgQUSgh8fRA6hDIooLvc6go0VJx0AtmireyhRpJunkaEYC4k2R4I6gNmu
j5UNOgFYf5uixZ1SVDSBGzYzO1BfBNs/TkcgZr5lkAtiHwQEDekz7Ng3jfYw9bbtJvUKhFccgdPj
3yozl0Q3hQnr2pRsA31WwVxMCcclInCDTlZEQB5uuP//lpK7dpExpjr8mopjEKgdwO3qU9mJ+2z7
PdiUQ3F2CzQwfr1AWYUVTkEkQal436SOXDSfR4RWurbVCSvRVGWI9MPrPoHirNrhJcAFuLUSTx4V
Lgm//oixEaHF4fchbJHzgH7SFBbIKGbgVUAzNCVWU+q/ZKPDVRNpAMqQUkVNIgP1h2MACK2+gmZH
cAHZTrsXeGGPFlOsjAb3+wfMirpd+u3oCJ8Eo3NSzfr/9QEQrcF+5ERYGJYbKS4fqhVg24ulRQxn
2yjrW7s7sMxtgog9N3gS1xfaeWfaXDEaKf77J/No+dgA6NHbU5g2vUMnHqyauCFLS95moWQRWjzU
xFEiEEyKjiXOnSQUVH70SF0Jx4kA65xc76fmDqYjD1et5KW9o5CWd0x3Q0nXZvvk0JxsQ9sAesP1
K1+3GVR79M4cJxOjkpUP+hw7zT31RjRXTwG6DAPgbgCDJjuU2avETbeE/A7k7dOBeK1zcAIiQKuW
2UC37MLfR/XXzQaZ2wK8y/+RnDKXefhlL9pOZR3KE3gRH57jOXdv7tOeREwLRkWgIrlkwRooxRKi
66PWkrjsmx75Zxl8ZKwpDS2PoBMTLjKCMxPZT4lPEfUUJONyK66nnxvWEZNODt2QGt4CngD6jVe0
klCo4Vb35wAIHIe2ecqlq/QmokA2+IwToHQ6LuEu8AHUpTENxgWjhf24DJdO3jQCUq2vi5r9YKnI
OgyHC+ObcaBle0XVyeC2q67uS4ftILeuiZIAe/p5UTbQ1OS4y3gwoKRu+lsgTKSQsaFNk5WJcMV5
EzDeCjVVIRPfDNrAwdt2YZfQ09M0dN7e2PkWvNrF1Evp5ZVQIJ3bZRumx9bMRzz12NxmCvkPUb7z
IbtHOvuBgn20zuXXm2f70Bq7PQEPcsBjvwsT7ULDIGsZCVElC3QKJp7qaw9fHYIrVGmWvZjhm82e
ugMNeiUn2TBvhJ/GD9jUpierUB98Obotdoso1hGG4JHYDuzNhjrWEvwAMprbdJWGrv7V0C5MlZ7Y
JnWM/Pk1A5QUXZ3oDZchMkC+L1HU/3GtIChS6GrlqP545HM4jJ/0gj9Z7EXw1aSx8xCaGpAkG0xy
PH9o3DmGO5WxRWKHVWKXQSueKi9+rko8NWtet/i3KEAgbJYMwKkKy9E/cZA+vmUHCaM0Fz8XV42V
HqYha8Cp6dNWugp508lsbgkG/tWDSu9F+X8eAO2qtSTDtLfPwcUdJdGoKquKnAuRej7gIYbQTEyM
eHRrlhxcIywNnFVB7sGv8GilD1TZCrtxgQnf3D+OBI7uVFw0pDMEmEcCi2KQ/MCGGYBWRVHYGkbf
h54as7Gop7MEJF2vDXcGORx4q3a38Lu73U1OVFzkec6KPUsmrgin2pd7N4GY7pgOY8KlDOc49fwB
vbKZ+Cbx4PBnT/wOYDgpkDm/u7X8sJiF/jMIXHNDa94KkEWJpg8vP+cL0GI5lG1UwJHUndCoI9hV
WwMXjh/Nut5kLPbq7PfIIpx17Tmxe9W0Ib8GNexlPmk+sDC47HsKseFS/7FBcnB/iJ8tq8gHLOVg
c9K3tCzBVa6zAAiwqZlGltBE/TnFCR+UwcoqPrTHwhzETtsOnw5VdPsjvkk6X819ZbyvGzqSzM9i
oTiFiphdJstiOqdAkLpitCQWx3bym71W+YaRIm6KdaHGGB94L7V0mwSYSnPCIMJ3TOSA2TiBw8mG
zfq6pOGouXwf0aTc9YswodlXvh1Ehmu8gYaEuKYrTaoJNF7CplW3wkZOPLNjANgWs/aKE5rex7ZM
zuPFqPTKumcN7hGjh9osLVn7OBYq9ZqaROjGdTGPyys9EHjA4GYaayQVJVPs2+NKEPIpt/Daf1ZU
9pMELDU9tSW+0wo9Thp0s4HSYS52NS16pQAEsZr3Mm/CH2tWIO8cJLe6uP2WCDFlW2MqrA0Sn1N+
mYrgo2z3CbraErFCp/YExFa/JCXCZRaYs1YRntBJSTVEpqtKKLMgShjg6dbpBdSJZH9dMVBCdPgy
kPjM+ne321sAtNONlrg6GUxc4782IMEXVLjraIjWVqwCq6/zrfyqChrB8Lz4s1TuI6Bw5LnEDpA1
J4fL8xjrlXFBqOm3+XM4mzNchgSwpZZIwkw/+nOvRztRlx6JYGK9JVi56OY6U0uzYPjp0LtxwpXb
Y0g0vbfKAflIFQd/AMBcDxDH3/u2D/xV8jQ6ofx0kLcm7QCH6PkODwn3HHoJylbRB6cLWUDXqlZS
d4vU0mmussGpxzFhLu33In90UFgSbS8rFN7hh3RG3S25T0vHbolDDI55ygu8HkB7cR+UFs8A10o2
4dtVeFgRT2qNIr5MIDUcs3GXo5SGV6jv3jkHymnS19y91Gqgm6IwJ4j9FU6Sbsp0+prn2Am56JU3
Ma3b3pKutd31ryS5fbQW5krgh3sP6IRdtwnfXhZcCW4ZcqHpoUnUcw8Td9rA5/CZyPc3CB+OntwD
Vx0MTEvENj5vfTsHsOqZnmgNkfK8TinWg/2vxseffPo7n/sLzFvXt8Y3dhi1uK45WMC03GZXYT7d
xYpvXIHsFEX55Xwq5ClYXvP0E37b7HMfqtLMXMqG78mYpZVVn0pyMEmwaXm49hdzpfUNM/Nu93Bz
K7uUX21o509hKvp4MkD+C/6WuR7LGvC5tSgLjjE7FnCUxghkSm3o/4PqNhQ3YDeBrTrxaemZZno1
+tuqNKVxvvQT/BQAkEVb5ba+hiatvVFPN5QVq1+tQ02Vr+kcqsxlHnsfqrrm1JH3Ja9uja/FOAjd
dKKL02/3FbBjj3ReC0GSKkCv1+mEPbyYwH0/30TC/OSgqzqK+ZNn5v+tFJ3zWWIkvnPn3uxTJPpg
G7ho38aEAaVxU0MHakr9XwXGF+CJEWZCsrNTdklF98MfPc2zdcU9lQ9aEFZURtQRzI7GFibD5yvC
nF9XSjLdBRfoSJbJoeEZR4l6t7wVrQgo2WXjdOUfnsy5A58XaEc0NwtQ2VrKDG0recAj11Dmaae4
kkJiUUyQEzk26hg9KqmTaGy9rGUP5CN56n3w7ymUe8jR0zu8g3UvoOKq22td4vQqrJgjWtvwtiY8
TXzhpw6RykgHErMXB1xYt0/6eisQBqHqnfrFfKPsmjYbkxfY1Y3BTVMarMiqEOuh3w9NisqkcSYA
2Nz8dqebksHcVVGQ3vdyhs83JnKFZDzHYMt3l8g4yeYIpEloLi6kGIR5MBeDnnOhJiCIJpLssagZ
RFN7yFTs8x83WMQFZpMeEMIFFoAX0pNrvCZbWJyyVf0HQ89iyVNl2PGD8YmXRQZHikzKbKAuIvil
Y9Mf5OQO9YdIOgb9U2OfNwiA5QDAhHrRhTbDQO/Vtriy5W91Z+7bV2BibEGtn/xkXSrCM7QZ0v9i
KPVaeTKWK7SkAd3+rkNs5Rsy4Nl2IzSVc2APB6CMSfn037k/K2pMiwxrYQx+YSVn+Ytn5y8RHGdl
JShnKD7PQzTXDLY0k/OddU5568+lh8ADgZUbbkabwAPdFw0e5QR+r6uNnAeLoC2+wUjtVcN7QIEO
OIea6Rc4OWwJU79mb883v8a0fIH0e4lo8x2kevqfey0N7eogs8Emmq7exTUUktrjbOl2E2I5B9J/
NzBCsqdzbS124yC53Evnr36IXeGEldvbImiPKfuyS2syYO8o0pQ1MU7Jhkn4T+evOibCcr5cHgOZ
hWVauYdo45jUGzRBQIA23+hs0bn+OF7dGTbs1ng/SHw3v/5UK+QLh6wggYrPWNRIrMGT6txsFgqn
qF9jK8reD4nJRgeRYHTMSZwI82MDFZ7R3blI0r9GAIFJiixC5fLnUwnsHWVDSgS73Ys/BDnWtLJK
4wQ6PEKTn2a4DON179WpewUPhHP4YzxHod+8Yvw8UoUWwUbYrUA2rloAKOjab9jopUizF6ImJDN/
lY8Glw0Ayvh1n67+bHKIQtLDuB2HhdsOIATLpfP0R2Rt7SxXhXpRjRsiKCJnwRndTBGhPjYKGxYr
YvRUwwVea6vh/wd+M8KLccFmgZa4+WRTIoJMdQLbUWZzR30CghFXLb4ezYk3/CzVf2lWCTibLB+A
ezuy0nCKfSmpElBIhjZahwBGL9a1mMQY+rEknbdeSCKCv1fQV6T3ISF45YNzNs74MDWghW4J4F7G
byiZYH0xawZfFUpMljGDAJlEVb8h+ZZw00ccii4QdfI/FzcUYoMEM2a5R9u4FWjBn361EqMyEDXy
fWR6mw3Vlm7G6J/0zJKS4CrKlE9U6gDw7L8s+n4BrktQflzb2vy1H6OpshaDmEDSH8LY2E6+HMue
lgcPocKoYd1a7ATKk6/xjWMPgf4sNILeXIA9QCq1aG1Asehv1JN5yYJO6zCk3nffsR1AnMpzDh0j
s+NgmEu6+LNz9KcTrLxA/kzPT4I032AzWa+0mybeeTXCwLRa5T/haQDeWPczLU1KA7WO/CwWgIyR
HswIBvqiObF+xMT8D9eBQ2rpXUeSS50Lfbg0UozPSYGdb99WEiUU7Qzt//1i5gnU1bGyEwpdO6Lk
vohvxoUlttF9UG/+oWLaKZjdzKV8vHL9yOHVONwyvU6zZ9q+KtXs1Clof89ZOlSFnu2L6Gyb6M2r
t4rdoZxBv8TUnCivUbGYdIArcdxECHrUpZFRjl6uzkJExadnoW8iXsLaY4NUbuXTj6xHBbO18VA0
SplIonhSMZTN7ypvddjDk5xvbNCDyjuMI0FrgvsdpTX+zcaItL9YHqD9W6QYG7G/Bj5k4j8aQr3F
aYnvV3whi4Y84N5cynFbGxjP5frJtxIif4KIh4VZGWL1jrX6rAOifdt2plwuP3Jj5gD/SEv67TU/
S+Ttq9Ssj4ZZ8kwoROczvG9C2KlobxCNIwKzbcDhrX1YGhqYIZxc3hrroA4RuoYwDgWFS7TEpCo6
mhHxbpIfn0MWfBZ5Tc6LmCewGT3B2iXONEPOG+AmYNNRIHDz4q1nq8/C66pxePEVq+UasL+5hUrN
eyv2Q+5L+OSbNJnSok1n1pCQVgxm7ncu/skCOjTjBN9JEEsG5W3c9T4P18EJKwD/mSXPR4FOFT++
/hTfQOyT44qZ19wwOjQTDSS+xT8XzW2JE9MkdMslqJ0fyLrQBVbPk3W5QVak0EThxoSh6wyEK7Xb
hWnyz9JTaaRJFSTJNWMqkjrhabVlzh7JEN2WG/sk7QwZUwpBPgeCQod2PwKUe8deVLwe30TRq5Vb
NaOofL5/XTYPuemGY2KJkVlnVFBGqysJ5V+8i6B8nnwlCeUpQ3TBrxwir6j/7Ok7hqXgG68fLzKP
mQPZb8lZYC8Iov6StYTcDhTyG1so93taBCDfm92sC0gK737zvsYgOxMqh+DewgJfkxGn2bIjSZ+7
axJwkACB5ZHNQY8qqMUueAoOr6Njlx1CYe05bwAnNh+kvu19iatXMs2ME+rtWgzjnkP4n1/OnSMV
fxRwtHzKJ1YTma/IsIUxIkAh6whrR/F8Bg/hin/1M4WEmdwMcyovR5GzMPDKqVxlUF8V+26714Ip
+dryRAY72Nn9KTh4KiHyahle27086Qjqv9C6MEIA2ZXc1ftnnhVuQt4pZuvXZYrLJ4pTZ3ySJWMW
Z0Q0+51gIfVeN10wEAS0ILjMJIT4zUVqIVEKq9ALdogI/LwYeP4uIB38l4FdFi6CXPseLiMoP59O
lE+RcZHIDrCubtLhy0+CXYUvpQh7fpqujqbv198fCfIRodPuhZb7l2P3mHJHVF3uXW78ziVRQz+f
FEChs+ZP6X3HnxT962jdKyoZprQv9gyfB9xVxxx9I5XcCL8SsbWcrIOMj0wCJjAYpaz/lVMpYB+p
gXsDNy0u5v4hKasMKlBfPed8t4IjTDXMME+N0D93VUYO7Hd+bDa3BrUdhVjrCOnsL1dJz9E0oTxX
Q2Rth/2yZyr+3KQ20Cf5tliQ3v62NkeZAkq7hpNg47Q1O8dP3pGu9MjMUlDu6Uc1L3BHxN5wLSdu
BYuh2BIJHdeDbFNr+SOoMR+u8SrFqemkjjEWB7b9E4IY48wDU4dLlff/hv74Tr+0frF08dPu4U0V
8Uk1NfDmj257FagXS/vHi9NLAUvfKw3kL4lWrcJpx9zX9ftX/OlU7SBYUipr5LjzMVXCP0LwIkQj
KOCs1jmlGmlbJtuwXNHD0LPfXFiXi11t8GYZRkrQb4UG7j1Xv9EnX0oyeemJXC2LYTc4LDRAPxLD
OG9SkMbfGJxxoEWepoJ/R/ShNQMAJoLNOw0od+3s0SXAid2ChdRRSMz8ZsEoK/57DoBav8f47oZp
BzS+kxHnZNrb3Hlul/68dVsbRQVTiUQc0UjSle+R+vn/aA8O/iWmouc0LaUex/DqBn6ZVVZ5iOtv
ZMwRTy89X6D21/gEppWOoG3t0wg4lZXYvFUUgn0AYOr5dgMc0UOj03tD3zQjLqfbCrGe0ft/QxHO
evq3sBYjDaqHsJEsBxL6j0Mf5pPVTzb0DC4M9Jg2ISu0mQIHqczLb/QwXZ9p9to8s2OBpmirFxcH
1b4RGHK20wGEQ9EocOOf0uQRXANwkrKnrrnkl+VPGqlEG/EiGQv0MTQBZBaQID6j7c6ukFxf/bNZ
nHdcG5GoSLK0MmrRRmDuQy1pXRtK+yEufxzXv50Ld6Kj8Y+kuPvHDiWE7M9bAknlPzgPfP4a2jB9
gnjSs2YeQNdyg1YmuoeFUx7DTJeyG0igSUgPNGZGWEH3rwRmMNJ3lJ9gEihWsjXHW44qaAegGNT2
U5TOt08S2k1J18EU07CGyLgAdlpDGNZQC/3S1HNSca3mIzSC8+m/55Xq9oIVK+h0CVINK2WaqRgq
u12AZ+It4EQsb2vvWthE7vWg7Ue3+3BrOszBCEwoK2UqlIMFKH0ZQ/KoytQ2GrnRqg85gvHSObnX
D045mpOH3f6o3lK8WZ7XijXej4EtWG1GemV4GSCADQoHrbBB3iEo+TS/Fi6pw3aOIDwonLteXt8v
XejJRTnar5KJYWe+ZNJ2PmcJnxD2M0GVxtw2gc6qKtmkeR9XvQXdcevRsin+tiuW1FrM/Trm1ZB8
LIYkSy6CM1jXVIJLV89PZKseRrj+16el7IfEifeuPmvGlFhTV+IAjg4njHv30iq9RqlQQte5SzIl
kERZl8OnE3M1773SkDzESMm+gZUj1VpgG4/LTC5oucIUL+vTexqpzdq2LwHcP1GzKKzCFJpcl9vh
RBe0MXOiDNbMgih0w2vlTL4MoAvNZk5kGqm0fhU4kZiGG2jqKr1ZlZa8nGpiQkXnf7LzqNT6BQUt
Obm7k8qQRhselSaMkIqKq1h7GiXhDlkryCtOJ2M8uOS4a2eyOeBgjU6ZItCyoaaRX0zVotnHTzHt
yteDtN20cD6lsCyu3nZTclCAFVzQ3l/8kwdLlDN/8nsWljSLnKsaylLGibdH0JnuFDfZpqmKfSwW
SuleCkXWydLGgjeJ1x/LrSUAMKi30flf1NTce+9G+DVhLaIyjUUakQSC6PapJoMk0aRHxPcFRHMz
WBfGY9ztwz62jE2qLkZfganOxuU7iVyCKy2qNQos4G5ekZPc+Dg/Tl+p3+xs/lTih20uD7/iWD57
20DMEsRhtC2z+AlyUqFgeQeu1Mx9RxsoKPAAsGEIm6vyaszgbuFtE+bbSJREbQS+LtrcAW6H8nbt
00Y2e+L2W+3jc9Ak0Ji8ePBW6BOt3DM9T/EZY8jFuUKN1vgbW7JupdpzKYv/HjftaAYCnHE7pBRf
B4XmSjQraIIoxLxiCZmVo1LvCFhrc8IVJCbwyzsKL2cDzIqfIvUB9uVEYa12uPbgHf8qSDv+iduj
HlLgA2lJhsFrpuOhyg4bQm6gkwhAMyxy8o499XbGBNvM99Hr0rBWPPO7DYBBHfvXHyEPQjv3MRGo
FerrP2YvXs1Z3wZGXzCkUfAOga459tG6p3nU2t29pY0zEsgB+wgid2U+AbnNwmLY6SVlWznuv0r1
nvMwI19Upc7XEgXQ8bj2xiQRmnbc7SpiJ3IuKHSt9So+6oSzsoVwFBRgzBb5qxqEC6IPncmpxs6o
8dMONHN/7ja5azwar4vEUEa9iKFsQ9KVLyHpbtJ8o1EbRNlid+ROxHbXEFV0rGDpUFGqpUmr8iZ5
mYgv0to6um0pidX2QKCxs0PEsD8oJipgIQBHDASjNQK22h+32J5iwNxfermMpwsaIWhbrQKFRN4X
7E2U8Qksr6VR1O0N4CUKH0IO7ZGvKZydIMxbHII4FM7R3ncTbJjXuRlN9evBVE0qr2dkjjIVF5jW
tuOgefWlDety0++20BOaKUPJDoLQnGIV2UBQyqAa8HrZtUr8BXwNG+Vc0IAW6DpD4bUywkhK5Jbb
hmxoVBH5z9juSbjZp58elcTlhoAngWfU70LO6WLxg28MfpA3WiaoGpAN1WGJ6LuReE7WDu0H8Cx2
8ExZZ7Us0y0aSucVtyHlElzOq5mClTiTlwRA6VdvYjnDeliBQjXa/PsLrtEp0kJJVUM+2c46nMPp
jSg2z/+AhW2eIuF4rOdF2qjbG9OejOZLrKkAaGcZDm719DhLia5959iABwTjf5ivO9LzlO71C0uV
D2P44r7hIBv6Wk6xlcZrir/18pvvJG5tKruy4hnhJNlkSCYXXO8kGb7Yy1wIm6Yjv0bBWFVT27ud
9d/EccaSoJjSGBRBrPl/W0hqUq88OYGrlMXqzWXyqrYf7CNRe+dRPkAFNInmv41oQUqQ6hhza7e0
TiOMh0nCd/6ps5N33Jnxcll9YpanUZlh+tiBuCiUmBTuJnBTgj1L4J/YCqn8NWozwPzeWnxwtpQq
UMudOo2dcySTErn0+6cFeSxr0sw9CIgAuiueGTmOtOOtwJEmLgIG9LWunf05+8Nezny1/mwxADNz
L05xwECB/gDGx7n3DxI4I73+BRNyOo0HpePx9ykygofM+FurcM84APaWblaeh1wqNPfMdeWGVZsu
d4eupcGiThmN/TH3CM29MYNaO0jZ97VSJJlIEdNPlMOKSTsgG+C/3YM6KaMF9Q1kbkwglHcjbxZq
XJrxlSRkURvnvvp0nTDiBoH6MZNk0cnG/kVe3/h1MdOyH+K9Jgug5+/Gzh2n9vn3ZYcFkBR8NGs4
Ry3CO4uQIQptfPsrYe53dK2VTsbxthVsbngCedCbILI/YNIyevMN9LHf0zwF+8MD1/Jo4Rf23qJf
ffASamtfrpRih9/XYiWP18bb1ENprb+F6PCXTauEU2rTSLgSghjAecZof3vnl4dA7fEk58iG4dLm
nVqq2U04VHgZVOe6oB8ID1q5wj9D3jo5BUQhrwqBxlow4qU2O8kBhJ47OQwtOYYU0xDi4qxTt37w
gG3d+bDk3VA3exet4Gyo5YWFvXFN1dlkTV4w7jcJqaPdmYkrf9VogR+RJsZtvYFgSEbDEzyMx/PG
b3YmrHgrdmpDIoIC0KRDK2kFKgoAqMvVdM+bZKggJLmztjr1isdEkvqAJly44ypZ1Tkr43s5Liml
2aeHePWy/tXzJWk4l6TwLLieiiS8uCGseVJF2HJF5PJURrfqbBZAnalR+xqaVn/LgVBfCUty7o93
JSrhq9juIzvGgU9Q7tclQ66K0/VACvWS0jBsBzZfLqW8XS1+iFVerFBFEJIW9Z/R5od/r04LxWaP
gGnEfyYBtlyLcEJXCwJFazzfPM1A2f8T5p9aVaa0zMIr1pcrOUaYqjYRUQB4McgoHRZFs/TzvEP5
FMMotskCC5MGAzYt2wRirmoVJyHYFWIQBk05S4vSyssdrnLlGGfCeaShIjuke3pDJk9vVGE28WHi
f4is2hKivm8qJ6kO97VIgjsOuwPHw+H0x7ew/sbMz0ZtZor877ZnjPEQlb4DF8/DXTTM/fj3/vDq
4OWiJQrvVT2CmtKMSb4vsv2FUaaFIKZfBjerX4Pa3HaG4LyRMZdkrD1ASoKDX2B04fhhtnyk3WWs
S/6DnoTMFSsOKVtJgifSkhGBuMWIept/6tXPy/aC3+JSp+AlZHp8T5wfKWoWALzSoODdyRns8Mmo
rQgY+tANTiSkBfKUqzleHsxdzB2W2nztPFUdCD/NpCHGPEsmg7s9l86nslkiPVjdltqM71ygPrX+
e9qCDCfZydXyg/jjv0hp7gZrMcAh+OWAudB6vZgejVOcCOTFl9ELI+fduAL7xZ7p9ZcB8mzldxOo
0tgBKRTiItDCVe/JME5wF1s9r0olha7dPQaHaPJiGHzvJBllMywkLKnkdA71wVaRv1sc+pO86fMz
JF1NzSEHFAgZyOQzCM/2+f51BJSHcRFfqlDgMh31bCW95MfGxpEav24NpllDTfhT7uio/GRs7h6v
nIBE4FBFpRBebVOLrMXLX7KOqoybfeWZNnbS75l7tt/elSXeuZQXrcNwlEE0PCVr461hCQUfQpf7
4jXlSpeZDslBlfSsp7JeO7WLYHvPVUoW7SkGcIVvvBcNVpT4qTyXlKQpnwKhF4tS9+uLLqDl/7C7
3nw1Gt7kUFvuUGvPxCYhZvnUd/D8/crRGDkuwzH9rIG1lEyfwJVCC15VHvXrMJb4rO05qLh55JPp
SBACw+j4Emmc4DPyToxmbs8/GXU5LrppATcxuoHBONDRSzKiK9aO/u55qHD0L6oScPNcxLRuIFln
r531bFXq4otViOP5NWeSy3Jh/ZF5MLMHSQj0iTh4r9QNdzAjDdBtBQUNxMktt+sgq3Yp8QXpHcRk
c7fU1W9Y79vu7us/Aa8QcZBHyht7WTJj25CLc1wlf7jOiNl2O9RILPoJdbTqgEkb/gnFnpoecBqX
xwD07FwVIdpEdvVIPOC/U5XyOEtYoLFUqo4MueM/fFJ4VVDwuPklyRwePZrXd8Rv0AdjYJf3ivxn
oZmjboWVbWw5tfLJXInwIHvUaejtBjUsMPXPbTAefW0lOXtYRQelPymLCQOM0gwLiI45SYBtX7ut
Jpb9Q8yIIf56HyFUsAo4v5dsxkyFVXDy1fbuU0pidMDbTePdB8Km4b9ibukOAjdlnC5eqzqYOFIw
lyh8LQogMDDs2HRyu1PXMdqCV3B0JltRWXiLurqR4YTUUu7ukBW7HjdR75V823w+E6qC6y83esTK
yQzLjlOy/b/u+BuDygJqvU3giw7fECdUNkGEra0kdKNRnJl6eZTqdL5g5OH387YzthfvaXYSswzQ
NRKA/QDtBaUvf5QtC9+0HPayr4KrO6VR2dmORLgvh20WFyeavH6qeS+CJHrkhd4mC0cJu2fhNsda
vmImgIq7xu1FL9dZ+bTD16pXOwOMbFOvhLYkXjqGQ9VQIpfqd316dUCLPgMpO3wxx8Y/5QsRKmqO
CIhxm24LiK0lp68zzHRRiTITn1jXmXHh6c32BeB0nGepvoqwMn2YIpnDGGXV7s6RQS0kf3uat7ca
/50XT4bRo4uzYrMfLn+DREvxS8P62A1RCTA4bCYFiYavRMAWF+ELv6QVDNu/EJ6aagm7G54bYpCC
wjs+LFdx74Lw5QBAbqODsZiloItLxUvurpui4cJfmHgXrfH03p5lAjJxXzxuv57kbOPHTimOKCss
0TwJUjw7wU2vyzCtf6m48rvswTQ3bdvjN3VuOMDJcKFgw3ikQLyBtdTzdcpK6NQtcgjcDbZeYVAD
UXA9/aJ8eCxDT1FIZ+GCLuP7dbhjDeDj/eeQA1cgIE1eK5bno44G9B54Iz4RFUgiM16oCpZAJGkZ
vZIqFz6iKq8g3LOvvFtHwpA62j9rONRoQWaVook4/MzdmMO4paDr1+n+f5axsxBza5Vf6fkJw9oY
C5Au1iZI0ToTHUUI2nbWqUMGVABXKVjU+9hKJMsJGy5oI9wHdU+aOfpNJS6qJejXHqPxjG1cRUDx
nQkY7DB+/onJx/414ZP6kksRWCSMfX7uYispVUPy/d5ONnlbikEOsp07obQ+/IFW01VzXcfIfCEh
jAz/MdeW+TfY4jy5XMRdNXsYBHEZtGRcBwzwGHAzwAN8cDb90A6Er7iA0hxOxc0SYnD+00tlMLTe
+N5y55rjuvoA5c/3I387mNpVaJdy4BC8v7yPxr35X+2EnSDDYuDeLlsZvfHO+Cb475JKrkOyjMss
APAZZKpVYitIwX4mS8424Qe4mk0VW1ASu4MP0lpvC837EwvqTQ3QfPZpTuaXyYaDdWFOliobZgpR
MoAuMBd0BCnJloD0u30RpEwuWjd1fHcByU4cDDMRhMF2FedGjU6hgmUQa7kH6H/xdCde44C+NauG
idjW6uhqTh9K7aYl/GYc5XkQMTAcnASzk4xf0le6gcsxd0UiuA2HMHByunqMnaX6Ey2D5v+YnJoO
IAg5EvfZ7CS8ALIc/X5wx1iv5RnIpQheab0SBbM2kF8bLw7jBICz1WoAuTHB5OuemDfoWLTMEJZ3
6TkrrLrHehPrnG3gS0o2M7/q0pIEEawGU9GehD59Veo6an02R8c6bb5Qm43bIee1S+Y/anM2YCaf
G3Fu0WTcoAAT5Z8kXOWhvPtUtx0FY7i/8l/1k4K8M1SQnmdLrJZlCXJMIEz4HwYAzgzsq++TWxB5
vQ6TsaQ9rsSEi07C5n4bKEGNbkQnW+GdM6y/aOseT0u/sEk7k58ENrJ2fAwfbtd4Aiql4OiDm2qw
ZHs2TL26HIicgO7nJhsBo7gaH7FVsun3E8wDAmaO/C/GxY5u8kD3X2OgvTc/N/tmd7zO36foFQpL
WBVKu2eYHnSqidsJJ8oPXMuwFcY92EAGfUj895kudkH8cw+TixZNFGOOJulOj3ya5V8qLOxGOdvQ
TY2e/2vCg+l6ulP3qsgqTIa+5AgC4DJww9g2w1tl9uXy8fb6ix98P4VpttjACoWvNGbsNOp5yU3N
hNwB7b4wz16thugfNa6PGkAVzQyAYN6uBLWeKFPG7rFB2q1rbL4/AmDEJl/f29/HIuNSXN1XeQJQ
exMX+XSstzWPTKiv9HTcad4aLBo4pXTpoNyRV1SrYfbV2nkJ8bW1TrJWFm9/WQkYyEQvBPsjAiZY
UfOANeG0BI5YrmD6rAXeTBLEkFgIp89KVvrroSxW1zDosmGeiR8h5MyNlCKduzqMRnUTuoa9anlR
yzNEY5DTup/q2d0+VP8pWBx+zkgYtfqwcEctTeC7anaUBxf5a05I4LimXBcqGw0+fsD+UkqzAna4
qQxt37Xs1/9Za2HHuIvSrPzjegNzzjFkVSekAna3v4LdcEa50eQMQbHah3KE+mNhZhVausnuNlk8
xj+6j08MjoJnsyabzUpIPSxssAStfvTLx7ksSKi4NFJrRyUd3IebvC5gHiET2tvihWR6oVblLsGZ
5c7a6rVFZy7j2JaQ/4dNABGcaXF/BTkKRppEGLmNDJXtAlDhrM536Wx1X+/OXPMl/Gi1Q7+0I3hA
T/tlO/CGDOGmshpvkZNH0xQVn9gm2fuEauQ/+5R90yGjZtoL+YiihskVsgKHYAbo5lUxkjx4ysZw
Db0x0tVnWOpfAWkR+iwNxOyl3ZYdlKfJsoLwaydkAHcYFVU20j7rrq/EGKQvPjEOT0Id4C01cc1i
MUFQNv2z1m+7fVklpQtefrkuvCZ5bJLjD9Z62DYiF7V2Msb3BMr3mLMobZZ4BsvPJjMqFp25amD/
llrk6fWwRSkaaiVIlA2N9ivRt41WZ4AOqPOuMjHxNpJvWL52SmmQac46PewWAE+ncVDSmL0RdP0T
TmiOBIvXJH+XaY/9tddNbTdj3yaxQtrUvcJZPFGvFZSFBj/mDtHQQHQrSQU1PU6RNLAQzzny2kWd
q1FJeXdIwOWt49RmiY4+o98xqlUT1QE8recLv1zQMyMwipR1zCaMylaVd5GaQ/G+dRhci3IKlAff
cwEwJZUrtBvHe9hw4GNEyHAG1ixN3Bsni5QTN/DKGVWKnLKdugJgpoxuDbtKR3GfIUBPTPxDNpT8
2NsObkOcj1DNG5okTij27d8aogIS2DpHJJY/yosVKr2nx5BYmtu7jBofa5UMdYPiwY5F/90nPTHl
QyUs5Zbf7dqRcqafvkGquBM6ZwOLjZqmrllq6lIXWvQvfXiyp3JeCPPF3a6Rahk20OzhbvULByPC
j0lAivMYF6Uu9D25MfatJ6DIAKzxNOxDl7NvEySe5rQYiyB9oPi0cluUAC7x/PQoRzfxQSyLG6DZ
epJwWQX6PJY1qPFXSf1bWxiCkMr3hcV7B24y3dQPtBX43gtrzclWbEJd0VVgtYYrBeilAabbUIC9
7jjPY/6hzX3048PrlhcGpRLU8Ho+akebjWpPDcUR7R5ZMC5GdyGN2I33+BLeo8mBWSfMZXja2Z0U
/hylrUI8059IRoiWAZyb7rFelBfa+tX4jAlRAJMFsm+PXPuE35yPIwCYmDqfCZtcD+yZGG7YOvXI
tFS56iqXNSDJMSD7LYkaaj2TBc0Gg9Nlb0EoJkX3EPEZvFvOGa9iIY2jKDfTHUcvYMvS18kUW8mg
VC+VW4zbm4VkE8jFwZ3LyNvS1uvixR7ZaoXh+J54nh6/VfJG9m1sFp9plmxhgGrGwbpvU7i1CZVZ
2n6+LOxIEOaRZYZk8uOigwT90MfKWCZZSBRSm6UI78HQ/0j05CyRJbKntpbwY8IWYyKzsfAq8F2r
h3Pg8aQj3B+K1Csttg1U+jDxCaVRKpdA9wTyFU+n+xqnhmMReh/mizhvOUgevkMUCxloFY8ZQU4d
7L03QPTk1Ym1ZQ5yS7c1F3KC63Exc79NnB1XK+A4fP9KXLN3BsIl0f5p3kl399AsP0G/LfC2pKUu
WR+2U5FoB2I3KNcQ+q7QPmEbdS5aE5b+/Okba9SZeBcSDdYem9pXpM5yKTU+9juqAK1rGT8gKgkZ
wZwnp7agnUNdLR6E1CvGYGDNtC7/0I8ra43lJqXhvujTQb5jdcGpb/Kv4sBdMi2PyK1bbSpNaAsl
zHr3Kf4xy0EyuyKplGQ5AaAqmraMzhhIGhC9U1dGBdWIlL1BX11cwyKs3gYWwgm3QeVSXSqYSBBL
X3Xv0TxqA4eLBBQrpOIRE9X0U92MgQ+AaBPn5znhhqM5kktgNUfQFRCuYYpfXOj5s97ULd6+V/q9
5UTxaZvqz3/rRJdvyFo3eZOlSegp0bB/yrJJdySENfZ9bHvTza0513ezYsVG42V6KvTE78++KC2/
lGExG+7XuRZwza1vkcV3nxFRrhGrse16VBxfkF5XVuOTiZckncM/FwJMU6VhQnL8EtByd6S3121v
qto+E97tIoMoPq0YoSrEKIL8WzwEfHHfDb9u3uKt9skxH+8hkQS/JjPgOkmYZdwSTP41APQx95Xf
7blEa1blqs72bhqHEtK7At+LG5/LqT+VDAMcyJIgnXSVRjbWmW8rGem0jemp+F1cNKYdgXWmCclE
ws2HRafQD60yrzHvKETBvm4Fn8jjC1FYOK2F4xu+Z04mZ44GBzliT55TevQnfl6vr8yOxdWzWG/l
OEhEUWflwcraLUr88AqjOLMdPHzCf2HTQtvFRWtSpBK+0TpvoDIF0Arv2bifhQqMKoxV4u9jaJnI
oUCCm5zUkCHx4GIFBXnL89SihxSqMchib6/uF9qbomwlLl3RTQlAUsppaLJz89v6va0EOpDHe+W2
7otT/Fi/ziHgaz3NTJeKUV5Ty5s5aMvHAKCeGdSoFwQLN4XN57sTj6cQFG4JJ+Ynx9fRFvPr9ucs
Mfd8wodA6/0bdDRYW4nLQWUWcl9m3IUJyYY/SMiGwwtZGnG12GYfZ+g/bj4CqBhwEWdftS7lA6rV
XFTrhmFje+BQMQo2bH4TfpHkoV9mLww9A5B2LtZM0pM4gO56n99JDomiucOThm7Vo4l39CAPzDIt
NW07qBf0HKRrhKCtupFILmKaOa0P9Dpxhq+uC0MxB18NcLh8PLuTKRNnWPO5DKU3MuXMWziJDA7P
k7rM6SbFDmwVpAUpVg0N1Qykw7owyhwD6QMsZdlCTviG6JP8sfmaGUBci0SPHWuxdjeSrRHiYpel
ff1vEkDZhmYQVV3At21we9TSmFZhRjq9XKPKVgfBXwL4UydVTAqxlDHt2aedDFe7Bndj1QbPm0FD
BGLeOzpt4jfrP/W1zSlN4Sg256QljecCzwDvGwh3YAng4gDahQLYiiTCAlf7hYjQk4CO81SI1+Wj
J+PRRJXe8FKO5Nqcr4A3lOM+R00487jvDVF6mVgBNN1I6ekVdmji/+rR7dYRPzZBNDKjoIrv+ytS
Weefky1AsZQDyUV8GE+6NJwp9zAyY+jkqgLf0IyJgVzcZqs1Cwj2AwwL8Ict+pd58+BLAhOgTEGX
fFrfKGEQDY+xh1iJWu2jXtzbZ+GSqQV+BUu+mrOE2XqKeoV8CVxLDvIo01OSSnJneqnVF7YoMEW0
qWMKkq0Od66w9OeZttGyCwxV7h1SGeIHBApdsl3xGmiyumedPUlD8F7BJdmFBtbGqj3ogIs3NovQ
BRtl39VdpSSIb4bvjvL5szcLtjLvoYyzndqlVsOp5+y8sf5waw/Mt0sy+JKTccSTv0Bo/yysAhd0
qYCkLaZAuYT28hEwnTzz46COnyOz9R5NlMigUiO7uqfXdNIX9Ezhf26q/e7w/27oNMh9/dyv7OPi
plpnAoPntHHFzM8wQGjDaFnhiyMmZDYGpAv9IwyzIxtjZF0WCY8+r2s4MgdY8cMe8x/LU6UBXaZR
82BvH0jvTgGoLcwFaTNlU0Sr9XFuSxXYyTD6tonJxU8D6ch2o754bv9vZKCaOieTGALFilE/mXa1
qQw6wHMhmAxSPocFBGb9+8psmi+Rmqodb7J79l9f1o+Y15wppRCNJwfjMDf4G7uus72m37z++FPd
b+9Bm9SqCzEoxlmUYfZxnUnQXug/2jmKd6txXDd6hEjmr3LlYWpPepAwCH5a256lLryURCNpXZZE
HNJmO/v7HQHyZ2pL6nBSpc+Yijc25r7P78RdYmlnYVYoOi/CCLsnEu/9/D7AKRoPHKeH4p33+oWl
9/UpFBavaxIrKWIjiWkMkOirSYPlrm9nnsUaOA6ra2ARLxo0PRrXugFz65TyzYOgR4W5yUwx9jFL
h9/d847QECQ560y2Wrk9yIzbPFdUgUq8GFGaqgXfGedSY4swx2fztKtdltQIHYNUMYMopi2rAkOF
SRIeTYLPDyCsxf2U7US0iHBogk8squP/v6oXV7VPENB+nEoU8bnauNC8F495WOeDVqNXSwAT6WCm
QbtgfSYHJY+AKCQSGqxAW/w3FXbFBAqum1rxapJYombYYFo6Ve6/6KaKIZsKm0nRURdffk17WgjE
PkxeYGM8447PwyEi4kSnh44c7sE8OM+GxySGBaBTNg1r8fkFW45XA2SeDkjWGLaIdKZo9d+9Ucy5
z6zIACrIu5dVMOwpFPUx6NyfHPelQ4hcr5DgvyG8XqE+EerDGP3sNJ8icbP9nayKPPaBxOuybiSM
Tf5r/7lmsxYNrCh3mGRGrv+KD+c8NC3FBRn+DLaAOeMpQm66Y+xs/peG2BKb2TShz+3lKndO6aNI
FHZrMcd/Fqk6UCLUVOGxQypXK3jWOUi1eUNGBNlcLCrVXbfu18YYngyOLC+6dwSOEFd0agQp4AXN
uYPMcgyV0gORERqIzj/b7thEzx/+qa9PzdLZNzga8wc2BCXkbD5MEJiyT0Zza9OyRsPE9fTONgTf
6V2bDZdMF+ayR3i1iJOFy8Qys+YrmPSxNH6GIIzRxmrx3hG6fB1ds7D6htLE19caxExhc3wyn8Hn
gsG91G6trk7DBv4ePTtsYLxLB1CHlOQu88LtxwfKW2H96d23kpcwQd7ZAhhj+zjr9VRECoJNzL3l
Q6Vyh9phyOO88WphUOJSbpURzTv+2Clkksffix80spWK13mccprwFU2EX7QDI+wQJ2c7nfx4O97a
Q/e6ovR18qijvqXaD7Tk1yGaXrHp40699OgVUxuQFcQfZ//G0anpwDbRI4UU49Uka/hD2PjV6NS2
QFcL7lUYg/TvMMPhMQinK/9yZTl5GIOjHVuMrFzwY+PRsV9Q5WegRmdSxGCfAOWiCZWVXx2GMH9d
SIOQF7MT3z9yjQS3zx5QpOffwq9VtaeYOzsYJ16w7UbYMnkUHWxjo0JX6pzMkmcehT4a0XbcRahM
hFA2uXd52fwDhaT/ucouJou+Ydh0fL4jK9lUYY5ehBAdE1+bBHhCopa14Ytw/OsE6fhW07pV/6Db
jemMMSWuD8vnTmtDY24bUbzCqaXDVFnhYgoyt5NiYxjo95TCdFXO996mMJjwYRZRsbKbm3YWS1/R
Y/n25s4nxnEY98gV1WwDc3lBDIr1GazigL0upPUEkh7UkV7jEJpfxmPylISyjIQQiDZE/345OuAc
PvbNCD8vFSlcegk4oDnWvkukHKY3DjmM/vnrxUlrK2ZNKVlMzHoWMSnkyITea8xb9MIaSLZCcM3U
s1TFlGutAAHKMCawFQWZt23kYDbqleRi/kRX69XJQi6ErEZxvZE7tfEPQluikXsl+9W2BKCZIJ7Z
obAd5gubSZDtKAXUe8AFZJHUuob2coyBErR8UerJlfqUhZcSkhchtpXXhjOcEDdMu++Qlvtin7si
932tFuCEpQxZ76myypqIL5pBkTtSnhtO7GxDXg1IhNLrf7yHNa/jwuA2Z0xJBFocECWt89JlwKfL
dZYi8ttfpPCAwj47mr+/Boxs7oHt6z5AwkMaWVtfo8yBqG9gkX/UD0c0EZVUKmUKzP3pG6pWTewa
X8q2Ev5nWRGt8F/CH/8ucFhh5ClwiN3C7P1X+dpEiCXycfXkhSDwH4QMYHzNx1kSPoJswiyIosMd
0vwSZBf5UdRn19wUZO4HqE8RrpEeqHMr425arCTuOAER/b8hvZiY8y0OB+lIcyXfxDiMPzWMqvBs
PuSNYmsqME2AYVLNf0EqmHLDH8dmoMHVpYnrIjVGbrrCGyuVL9x9h4zPVPJ+u1GdOE8mLxex3IPs
IPUUy51vCA7VWcp2eBII1NGMq9gWMKBQozTBXv9pBqZ254xRfw9z9AXDvxA3bJTSVJWTbpPMnyEM
Z4GqqdQnoZbW97kvqRIazIZ9U15ypfuEiroxw2hg0K6f3ML+4/Z7g5lZ0LcZ3D8QaQZ4MyN0z7hy
Ey04Q3MEdJS4S8f7FVn2IYfK6mTgPCH3mRd1ACPfZtSyA7kE73FQVIoT/fKAdlRQP9igqOW+OuUv
9F0PeuV1RhrRVV0QaBwzhEgTvHhv7wE+EY07y0Uu+jmcC/L/ua1sbmPvUUtNmcFN03Nd2c2+rpUu
P+tJk6JqlfYqXySSOuqi120OVXiG0Y+YJFQdM4CjMSIKoIrm6dWyJeBXskKiNnw0d7bvsiXTqE5U
bHV9zNTmFVSw1xX5PaBpZ+WyUGdgVSDcnXaZcpKCX9sOM0myjTmnwfRb29gMmY8MID/qPOVoMowO
QDVM8rLHfyuefkvEBE/aPx5dRvgjF0XQeDnSRZ7tuMwj/4Kca36bca9g+pMCU20P5/ZavPS3nSRt
lc2XAXPYWzp9wgLb6kAwSQJiWWSjdZjEYmoFsJhhAtlBjZUa3EbZDzU+sGKf3DiNUDVp2EEyFgjt
w816gibyuO8WQBxSV9iNdUCk8r/k/MpqHSRj5Yl10SnxnhuxQsRviKk7v2MRzlB9Qk6vHczIQttk
4Th/f0WRoE0zgCxLCqO6CmVogVrCd+lSVQdk194lzLts2YzFnX+Ut0UvpgI01fF0q7hu0bbC8LgD
CRlmQRbRSqRQMQnUnvTLENPTwlkqXLcOJqeMdUU4n2HjianqDU08dPc+yZbiqinhcsU1GDI3IOW9
87LP8pGQGyjc94rpTMcBzJUqzb7TgTVt7q3LOzsf+vIXoCgfBDfk1FpKqkcdo9jn3IbpHgs/uVcN
Sh28OBksB1CuOtm6q+n0vN6t9no3Mq2pD3ERQkxWlrHO8e7rXQyioXtC8rhGhtp1JKANaCJFLBdM
R+C/T7CExW3YfNN8w/xRsyZ0kFTObUSZ52LD9yCPofTaHN3XT2k8ggAlihn0UotGkNs6W/crH35b
7Pw6+OQ5CHCdrINq5H5EM/AhidVkHZxkrHM5tY+N58YP2kTqGyBWi3uN05zYgVsxOTWGMVhYFt5l
cqeBnpQ36qMVhYaaBTFcxnOJT4wE5Lp3NABOHGGAg14cbQMRH1np0BuCaMwWUnuUv+MiZad1j1bx
XqJOJU7eSNSyEejYixd4VM0LcTC3ZsuYKJ1hvMrFdz9cumXTdij401o/WVf/8ORX8E298LoBzd8o
XW+ILCZHbQbFcHLPcwSmNEYA600XPDMAVhk4q4GtsVDCm7+0JfdQDR9aVXgSolGoOjKKpT6hNlbG
4GzqfZbx30L22Nacts2kLbdvKrbcdDaBKtevPBqt+mYqmL6ikdBQUqMDF1CTrB9aghxTPrbYsFmp
h0FlAEFoqEkwn4IImJ2NlcdjBTOJPWMb1kCb3Zyxyzps1IXGgdxBBP3wQtIk3mMwYOHxRDTUoIgH
jB9m6mq7q6ZJBkh1Y7Y+h4OImJNjgBgIqNdGinU0h0OCqTPp/sB1yJApeNpp5CoZQVSwXTmVkNu2
wNRqrmJOKTI4y2nkAFLG7btLrbp3BIXVl9wRBUmSTzsB+VQFngv2b6SU0HCptWqsxkxfy+PMdkRB
rX0r/6CZjpdyAWU5yXfPS5Hdn1/h1XG/OZrF68E/a9H6gyBX6U4f1XUpJLDVz9ZAEXFgp7H4s3Dc
Tu9G4EasiOtWK0tXKZPUA4BhUCzyVTaBesQVTVVykWTpfSlnD3KoLQ6Ltbhze97V7lKyuPaoNgpS
QiKUuNCDiIeTLAnHYie9EgVSC6iU4a3JWFokumZ53DEB0XSP+eHz+iE9YlR6fNXt2b4xTowlgTZK
uKP46jRTbWfzSoOlHfiKspql5/cTrBLvdcTlNDPaZ7QjOhkN2KIanl2t9u0ElL6sMq2ka6mRJGCa
hqOAPFPczs1GKC4l0KSYoUW8q1uN0pqLMNhHg0Z8AjiqRoRV7q0I7ioY54GLNvCMOtoYrYK/UgB5
GyFfcWoYxO+ucZqjWT8mhoKNarDQ1mYqNaSOrDt/pKQSoXbt5nqk1G2lpsx+bZ1YLd1iS9Ln1Ie8
K2gNAu8wZs1/Dm/OkTdCtmURq5M69e47bs0XluAiH3Ex4m4HFSc0x7dZ6fdK6bRXGTnI5T1SUOlK
6ZzS89pwLxTWmUb5TSDNYEcmSMNDgTep00sVGdzlGOaHrKZTv44zGHxf+AC4sNyzc+5WjXhUSMLy
DqXiH8lbdJNeUTC54YERt2G6XkKZe4pzYjHK886RA9r/rrKSNS0+wY7hN7DzeITygz05llCKTqrJ
3BNMhvLAxm4pDHjx6tmoc9qu6Rpc0Re9IKh2JhAyjvqOBtJehdPmpHGab3+qwTtCU/ry9hh835qB
HhKsyAHVyt9UmUWlSNl51nHDEnLfmLaqseaa0UqVMl/JXvswau1noH+fCBN3t4jdmDJSxB4+JpmX
mGldUR4r6YqOXpnz/4YGGl4hfghU2LoJw9Na+Xm0Er/eJZihIoncUrqtiwtxCpkSnGjF4fHqHbCb
UGfDg+CMBNJkegdU9EIvaGPZ5Np5ATue3vWUZzbbSzyO74XIMsv5ZQOPMDxrIx/ZgmWODUBD1VYV
oGrLxkywxxC0ZtUh0ZDuIXhCzygl49By0pGbYR58hP2zmYyB0iFU6jW0Gm3pgRhYTIQFsM5w0tph
QeH6p3blANFO9JgHEYWDpNDoNhQc/FxtEAAMdteIpL8U4hGeVM+I3pJ/xVN6srTBGg35mrANejS6
DLnRjwLqfi9OR8B93qleQHg9U8w4Ck2LPY+GZuRS6As/f/kqfBCXwdP6zhbuD2U+r8w2Ny92nry7
H1p86Aze3MvSmLJu2wf31bdqGOjfO1aVPPyXJf+vMzcYucvYA32GGghnW2kP/Vq26UBNHr3ngXH9
/xP8vgHPKNedBjnvtyd+o9s9d4KP4jYcvNTmgx9bwNIhmwJFMh2JCNh60ocXIHsh/OFr5lqybRhX
BFmcoiBq91xq4K857MIKTceuD+jfzIltfpe4QCb1OKWAwiXDBdMwJroCVRkQMnrdeTlqIyizwh8H
RBkfoliF+U9MZvUtvEaUJgFtlnwCkxrVToDLiUy73hsQfu1BJvMi8FTR2fgFRKf9YamY4amK4Yez
Yex2APuTX9Ni95BlawRvMDrYJEfS/q+7NX1enwvUVDboRVO1p1eMeeuJjXvv1cZEX6wsozGgpQOK
LoxufixeRiEK7scxlbGpL4tMzugAi6XPnRHqRUVXhd7Ya0tvGHNxx3XjueitAfQlO3LHz4MRjPxB
XsFPSEGfWkbqXv0fUKFumxZP28cnk8jB09W+cb1OvxtyFDSA2aMw9l1fLmPvBtZ0Ge9FaxYx5ij2
XDR0JQPR4iV/MjK8ZYWHleivNRHcm4RaH0GvrEbeN7GW4VdQuRIpJhJc7VGErsRkbbtDKblWs8kC
5NWSVSMHri0Aw8GnvIVgIhyFJPP4al0rcu2+GNwS4EvX75t+trNHaNj8NPQ68syYLpScu7UxTA98
4vWlmrbgqF+vpjhjxnmnWDw7lAOjuvpTHF6msk9HN8pMqA0KD660Q5bs5+zWtEn8tFr313TGOyln
NdAnkURRi2jsb/IrR2RU7Hoxpvlp/gwICOiI86ysG+dUQFkU2abxdfhZzH0yiZl/RGMg2m0qJotK
LwGyY3Pfxb+epBsoCa2Mh5ZSeVuReKrHNthSsBzSLbzQ4Q9TS+DwrMRso4c56xTZS0e+kdbmpPr0
+s/a5gtvcHBfgIDd1smsU3UPhY+VBJ8CiPePlUtu6bwDlAi9IptYpVoOAw6rpx1+NHgbO2jXJMv4
6jo2CsM2073Fl+QxJ9/3JB0erbug+tGVibLVr2FbFbMwYmGfkT+9Sw/pGRhLgXCtmQW3ChTDexr9
4Jj2j7gTlBRWsAzBPbeSko7E2FjllGpf/jqYh0UCPre1+zXk4YWo31PmFv0CL67FFI5REQnKc96T
Frmuh5zHPIj3U0336ShlwVIW7Yz54W5nmheYOtNdQPzKdVQO5qplCW0UGhWcQKJfs7jWnG5LbyiC
3oZRoXw9WrlggJyQMaYFNvXrjYT4yP9/HZAX7qF1atwufycbFbtKgTiSVUyhNACYhBnbCeKwxkFB
DLN6WioOqX5Goa6dumq4o/+0k/TafrWuONytWjBt5CcSba/UMGfqSb4bQI6gJAZHDsxO70hk8elC
6xcGP9FCEKdkbiIbR4HspE9UT7I1w9Fd6fwQWGLr4xnLekWfGm2+AqkcgygZe/F96USBx+GcjJpm
yiI/EJk03DwhSSEVeNIeRJnK6y53E7WV3zT8PtAB0aQY+jZce45isxIpgGvgFnyBobIDJq4hwrVX
3TEbrqsr1i2kHAE/xvgHCCF2SQ2e5mFGndVzDNM1h26cyuEJJnT59Mz/NSx1HpytdcmBxn4Sw41H
ax+hwBW4aGWc/JFj4MBfYnxCMJrqI84iwXgkBOG49Lwt+6HXqIbs3+T6JbBqnFSRNcxviLS+qN3+
pHCf8o7LO7Hr4hNXhka6mm+x5qLJPVIaZlaWVvDe5pGUzHIfDK385Xap7PxOcEAl5G3J8EoKdg9X
AwK2k+2NZ0vs0/7ZCa+pc7i9cI/vKi5AWIm+wC2JH5NA0DeuJV9Sdc8HXcYX9SadAEIbDh2Wgbzc
qZ4hOwRJnDN75zZ9WSSK5kpc8PY6QbKOdUIalxM/Hu0NYZx5qi88KdZ1+n+QcTNGaqM0+GzAgYE+
qMbmmaWHVd2gbP3DBCcQGHd+o+ThFcV3xF/yYt19l5sWWH2faM5lrcUFg9wQJVAW3A5rPs7xPRWh
8UoA5X2LyHwbFSp0RL9u9w5FVdLnejonz/X6B5hXTHXqrHq/OLBmi45J9YRblBaHIz1rEclMNtX0
GPOtxz2df7qMXobdgvYJx9NzRGlPUQ2+EdOXuWgMvdE98faLJyNYDYqGm+VXjf8/UWZDk35u82sd
hIwKVt1UvdShtHUONWi8g7l1qnbqpRg2j87ixamswpNIl5ziapBZRgA539E8hOT04ZCF77V2ODza
anDJb9ERJ6tizIkSd/NvSdR1afN/5CF0zc3+1n67KN0S9hih+2ah2dcGYx83kq+4FDCB0bIxsxoY
fxau7pCcRWQVi4zdJGVKU2R5N0qGiBu3YZ0VTXSHS6g3oRnxEVa1haoNfEzoIsiVBmXEhTAgK6/V
UMRfJ1FDFLqCNLpgVktaocNIxsEEB94i+lH4GZiK95hInYQldJEr2mGlCtIPH7QSOQd6f0EOJXZ0
aH9On2XtYS/tUoXx8eA+wmYsoEfLmmPKs0mhvNwUOre+PcAag75mWuFL7ctLao15REwksoZT9A0w
YNxruMFU1vr2PujrgBvVAYi84LGZLYXm9jOKod+ziX2CR+mhZt2Drrxdd6SHsE6Ad6pciJkgj8i0
vICO7zVLSZBpfqM6vqOAp/VX7/Lj6vrFYsf+hQgvXEJ1+fPmCeA0Qe4K5W8iyBgbPjtHSUh5Nt1m
gZbJ1qyQgA85WGf5xiVyRMvwZmebc34/s4tqMv9WxrUWg+ZrMxn/VDv6whR5gGLaFdFhojpVMI04
dNh3NloEV370JuCGUEIDcwEB7RJO4POfaUubnfkKEjfyTP1kMgccDJQF3eGwHoHy5Y15YxAZgnDd
olVbmJHFIV2BCw/E22NFTqnUHX70cKVMqYLsX5r2ehQJn4LHQLMb1BBod9fNoXENx+djQZrZpi+O
KOKvkonX5RNZp8Iw5xjCKzBgm7KuxiLU1ipGHiwTDk/NjcLe/sLYfhIaWailpDPR/Y/ICxolDkva
16SdHYjU+Voq8FZNQXR20n2t6MSDOVR72ApbZbDGMZmwXulqJbMEHa8d4uwCsx4W+y1bR/IaF69c
xObD8Uuc2OvFT7I62uwGwQ/WwrRR4fS9DBQEJYbxghEwJHsCJF99Wp6LEQxaAFVnTFxmvggqPuZj
tLZ+FYsvJ9d2l3BP69DJoIOhtjNVQaFItgAg5xjKMNrA0JAg1ibugkdOnWyDvJu8sN7ftxu00qEs
/bLlg+iNp7Qmbd7TcRZtv5n2RxgyG4T2peOA90SWQrJBNe4oyZraIpOn92FW1WvNhHxaIK0sezUo
SPgWkJzpH2O41abpiKVa8Bu+kpfnpf6Rb4qeffK/0lWFRq3E8xS1rKq4AZSM3kM9rT14QcZd0qMq
dSepQ8J9dgrMxoXmCLbMnw8V34nZdn1T6zOYfDen7ZQZqX0NMZk6h6oMUO3P7nZK9jp04IlZNO+E
H1NvkVzc3A9kO9W6F7Ahj/UfkM12lZxGDPQbXDgo4Z4u40NtFmtICeNqrs9B0dleWMyhEROOCCVO
nfA8WDiPfx6IFt4z0MlLHPb8IRaxWTUQzM5Zi1B2syCk7OrAzHLXMwbh5L0wkaAGSZWVMDH3AkAp
P2qpQhEU7FvORwS6eq+bw0l5OVucBPMnhl13thEpr1DfugrZp0bn33FB6S8Shga+UOOGYFcMvPJM
bzQug7pF6+wuJVdEBDgpjiycAex9NcX8d6Mx4QdDIPJexUkbAotOjbGA+sgaz1beHbQkafMlTNdb
lTwTWM2w1e43EICy9Jkz0xKgnKmiCSF10sos6xAH7v1iwsoiFUDCKPNWShu6RzUawA3sYlnElPJV
cv+jxmz4rorW8c0oytABKUL06+Ig8LoMKUYLrelaviw7Vb2QvuhcxMONNuZl3PN7VNTh7G3U34CK
ANvxDeVu+zNwKCXNVNduE4zlwoml7NzpjPsVgB3lysy8ylft+u4Iin1Tl3QGYE1ooKa4chDnyN4C
OF41H22lEs8MTBGlmTNUvyuvKhq3qFpN8bGs+nmHq6VRatztoCa0dGGDWdxpxEUizfVvb5mY72Hr
nWw4sHkDH6olpVwsDt8h9PvU9vWknUd1OmonYXVSJHwHV7HJBvnYMBq1hylH/ECKlWBJfj1qMGks
RAYe0IW7qYHoGklLXYKed/0jT6uDnnL9tQpa8muZGxSmmFVHnBgqbWKKDXKVsJcvzvpYeU2JPBh5
ZmDc/1JPfdfs1vIfp0bc/ReB40cF/aCc+LEX2J7IIgR3kjwjze1Vzd/6A/2vL8flZ1Xk36kmNvtO
EPzUexZmts5H4JiBgQGhyPHNYP22HJ9NYa3ghHrJolYOD0X1tEtqsW4lyvncmFcyD2UAjItQSGcu
dOuAgWraWrYgmcBQrk45lXcKb5U9AjMFZdRN6MkpZOXaKV15KfR1WN1SoQmLqKSRTvzMOdBo3Lyb
PVH4aMwPV4JsyQQTBU23MYL631mwmAZAEOEwDuvUjUaa6qhkBOZeSbDGtrdUMwL0dzYicOdbKEef
IdK3Ij+MdTukiGkVs1WDse4zujjUxHRiVw9dsbW+/7weYJH0VuRk8HoSfDrAUdDoz+6NDgXlDS+S
F+CNbdW78moISKJIi0a01fXS1pHDAaSNO3GhV/Dk8+EGD0sCOakRlMpguM/9BEJZqnktatToMD9Z
Qefe7manuwQgqtoFnFKyjGkuz2LMJzVRGG0b5plMUZ49AppRSIA3XUmzSyoaICGIFu1HoWvKIq9o
Ns8czYyRNlLonZdkRnIFBka5RetYuSF8LNr9f0bB0Rw0+FBOqxFyiQEWontNpLqtW15SrEk0uMIe
e1jqH0wbHy+CNYRbB4fq6KcS2cbWubLqGwh3sSRizJUWfICDTQ4lRaECEpr/eV5VKDe1RLJlx7jZ
qF+Ymfen2SkG/R1jQv7nArYn5MczTbzgKXXAvPbhaCXm8uv+wkbAuHDc6bzS509avYDSKTYe38Ly
p97TAMyziuyMFcvQnKxcXoOS8UDqYiUHyj5vW1Ii/qu5lFfzIHqSDAkJ3opeaJSzzGBoExyr6tJm
jTMIYuLyDM92faSdzBFifZiuDH8m834dE/mntkRBwLMQMiFd8/GbB/SWucXkVJ9NVL69nyfIcIH+
XdOwypjn4HRypt2Npfy14YyiGqCDhj83V1G58JLpiLT2tvGGzH23RS9QUFSUzaJCpbTNW47zCfaO
IMSlBtDicmN5QagOH8naFd5++SzqdkuQxUS6uyPmO6NYf7SfGguXFyNGH3lHqRbrmvSFAxvn/HAG
mFJjYIBPH/SrcfY3X5JO8vpSiPFbjnPiMHeQaHAFVFHjAYktkAugqqoPkSfutaLVlNwwHVVn92ug
ewmDdFPheyxBlI+oOrAyNzeyEDKPaJk4MEZcbMxjUmE7EFywAqYuVmNruFH5gUIKtwtkvMFsN4kh
eaOqHE4qjghgAxntrRIxW+OJgk9R3OycoYt2Qy6+EmUkxbDpTkNLjWqLLw11ytvG4gboGOiSGLaD
2i5gtjD8yBguqoWPfo4myw26yGYjypG8KJbNgMULVf0qGbuC1zIQIpwqxpPgI4ANfGjN2vBUb2cq
OE2RaQ0FH3ddk1mg3vem6L3NQtHwfi8R0+x7MeqO2snGXbjMp8SMw/+6fnRoPm7itAPRvD1yh05F
1GeGe8ozyf9+UhIKBjZ0h99NfvQlbIrNotDoeMlpRDyftBEB103ivbKdCIpIQ80F035uk2MdPbXw
PUsKQpyAXyWrirzUJXiwn1a8kOa3sWIV3HR/jkShxHCJ9c70Az4UXdN+TAcpf2KYYgwq0SGUXtbX
e58zPg07nXqiFvjKcadWNWQvPeozkeoojKNx18rOum9r6ifItNjLl/ufjyA8JiI4ZRqrSWy7M6aB
9BPyC1C5eaI+ncB3exTQE2+cp9WFq4Rd6SigZb7EdCPkuUyWA7I4UPYHRArIQWZND8ZNpmW8CUeh
RVG2zMOSNJ+LAHE4fbPx75b9Zqo6N6lrdx4akcF7wm/zWF1p7jyPJHNIXP4YMuowGgBAQtoH4O3z
TCb5kxwIpVtA04nAuElcNTdIKR1Cc8yzy7tRAghONVBJONLt9bYrHYMNo+r1CRE+t1Ct1bZabZwU
+THmQj04f+A0ElM7ZPOr/bFAtL9f6Dmg9R6DIGdKzjuTX1OdhcapqOdaP4wYevLcRStELM12v92M
QtSsEnpKM1gvD4jREvpdAsublYuOHB0rGt62vDXcVFagAVbq9r/8myDtc7iUF3kG9Ov1dv2e5SeS
mxGRXRNTlxDXXhmXL21t0psqZdGg4jwBJVbOmWlcMlrrGQ4FejpwXTw1dQOy/1uNq4KrGMKPbQAo
ozxuKTUeevnj2J6c6Yli23YW/F5mlji8ZvnBJmAP1oH8KJqn+ubuKp/y+ee/Pz3uZGQXGG0dkTMd
D4klnYriHOaS5K+BwV25gEr2aIcYaT7WzdlAadyoXAy+PZr96yxG6ELmvNtJyP/dsb3jbH7SNZA/
hxX3ucHTV5jNjxUBl0CIzRypArfNt9lmrQYSpA2ugsIYzCdrToSX/Q2URvNCIaSx+1yBYVcjaUVk
+HVpDS9O83D2ijpd1uKfdUwCTltlY13BMUI9nEFoqf8Z4jL2rgHgfOD7oNXlKdi6sMgOG/7H5ku5
+/0QPmeLyNzEDcNE/xZ0OKOARHv+R1aOyecAh7wsxC0ZQS/R3UwfQdWDyKdytEW1aGZLKJafgFlX
HwYKDaOnfIFdyZkcRLxUAybhD1Sc5tMnTnTRvuKqRVqcIg6WYN9sHMDASzYNJSKkg84wh5DVOD5y
oHO4KewHPdg/lUjDTf2YnqYp/6xBieN5KNjbgMJeJu8g5u69uDZQuMlj3SnOkdLWxB3L3Ug1K8Vr
bb3BVREfC2ydtS8NJl9EgZnVJiMGW1yW2uZ/lPsW9gHxj0TCLo7UWijIvmWKk3Fn0R3Eel487wnG
wAHJgKHchkc7El9B5CfNxJwJNA2lYgHM1xllSO4uw2GHA6m7Aub/NW8MgLobW1YFSbXo7biiuZYu
cixeIQIz7lVImT20nEsSFJ/j+rr8AbqwB2o3uOXvoAL7jaVfN9wYfbIwbTkgF91UVx+H456gEZW5
qbiNUMbFRzT8NszMFfd0631R744ghfvXHO/Fxe8tPTXyKKTKxPL0Z8DwGcK9EYLlRCP+nhL2Dnbp
EVLTpwDItInhH3yKrRtvwvV+n+FIrn/r4q9BPWI5IFbXXoermIv/r7RzhmiaODh0Ihte+Od9PZti
kf9/URuzd8PUsxD2+1lDTf8OYLQa/yrE222WM+fMlL6RBZ0aAH5c8KYSfevXudyNVIBtKIOh0ltZ
a+qSJ4Laor81zXdRSYppZ78da9CipP5S0aabaZgxIDh010qrpl83t51cpL+re8Z1Gl6yiA7wOj+j
SyVSxRji1G7U8nZB1BmJewogVQfkpAncdg4EYK2bwuholYKxOqpgwifsACgR3RQIlbPOvHTD812x
myLH+PlOPVxb//Bjc3ciNY4F3MZ6lRSnZHk9Pej0xlcdsYjYAuRsTjXEcqEsLw3DHwffkAFVoTpS
UWdLF+X9yL14sFM9PPSZwCFwRikyJk9TM1FBzAf0fuIhlqgn3wmLXbgV5EUmlxzoAIwAaCjqAEoc
vJtc8UCEBGE9sWWZ+0D+L+riGVv3oqlQlk2rZc3kD7vPXzNdfKGBbveS4uAHqvzrZW5jyUtR5IuL
FNFqdQtzDCFow+kSj4mEg3n7s7K+Z9cs2i0egY9w6ccLI0Gpf2N1jhg7LUInG1kADuQx1ftZ/8Ic
UQw9ZX6dTgyv5oDxjCYuRh4LoKcw8IyLJFzok8pANXys7oNXIKMhBf+lzpDxL5mS5pDK+adFxDmM
cIsfq7eJNwtlJfZDaVceqtfChtE+Buzmh1n7K5ldPyHFTjRz387LOv+De1acodcUlzdONxc3mIOX
Y7NkdTTt7gHtFTO6tHyJaxFOdHjDXxzeJVVTuAJi3RyO6f+LJw7VQmr6HOZMu1WJNHoRkrPBgMUr
ZM6KjTLkooVCnM5nCzB9Jox5NbCelk+IFIzbJp5foHT1008ZAPBsjpczy5A0KMM4plagnalCGToj
1VUCLuBU3B5DY1kngvZeM5AOfQpqbPC/yHqxjFi7Tx/U2yqNb4LDUqP4e33VWafFfyGBapvu1/9R
y0oXuCocTh0G29KBYAiJhdF3gaNybAvleyG7I+ffiJNrhhsAQamHB4v8A7xChseFYnkfrKvC8J2W
hSTqXqOmZhJLOt3Bn54MSUMli2vHQuRh/W0q27VegoCBeO59G0CgSPNcEIj4LD29mZc6RyWIjUTQ
jxvLv/gB6v40mdqIV1MMcpNRktjJ2qadkoEgseSyG66/uUaPtECSj15H8BkfQ/eXpADRsNER1wmg
0bVMrCo7dL2DlLjHfSTtwXTftAaMyMIe0Y2WPjalZqTehBxFRH7IiZv+HHECd0+aLl1v3N1MSXdn
0hlh1vYkEHHMiR2HLwXD1zK2YgVfg2nrelD7fjZ9Z30ZjihRskBM/IECZNgTdhTzkCd87EKm14ON
yLGgJ+7bqsDaDUw51+THOLOw8Ft3CM8Jnhy63tTyaKZ8pniDDZNLiUdBYeZ8O1NVHVtVB+5OQcgM
FcGPCcEInoNahAOL40gFdwDpj+lA/eQBGmK53jRNSguU8uj31nbQTz7temi5GfFWt1jaHDnVzzwN
Ztju5L7JKs0gs95qAPPs2vgOqNooBKbBvcjjfxlTDcOegZglZMy+f2W+/JkYTYMXN5l2spKQjzq7
aJkPZKR00mTeMpxjTX2UmVWulgDokAeX7dvBSfPmjZuDRnXN26vyxdpgRgo1S2zvT8p7ktjLXD04
bXWwBCjwhXOD1OhAGMB/HID9dpucMOSU2aOmiJAk89rAjAFh3ruFWelzzcIkdjqcc8AOeGH+v6fq
bwP8dNEitrLVrZ06h2ch51N6PWCUI6eZu0cVXIP43HCedSiPiO7A01/j0UoFz4MJa4wUj7R9VzVt
zF/UswR+o6mTP5ptGozQfwOHxkSqsy4wMpn6/Xz6W8oFpMf/9E/tpr1M5yAMhUc3UPltNUgKdl1H
3Vun2JRuYERScuFvrHbl+P12mvu1zdIRrSEyT1Qrm4YuOaOuNLc4zegnIHHdeKHC1wUbPAVgYrLe
aDhlchAKIlYz0f+yocbVh3Fl9DURiVGLSI1G+gIS6nYbDFyE8DsY9PZDfzasnMKdatjUiCQvSEQ3
wOz1SFHMeGVxP56LMsgawbKZ4LSMlkHy9RuVGrWef2T625RYi0dX5gmKbEAv0BdLp53ZmsQ9Ne06
Sye7686WOSiDyb6za3ZDs8nMrHgzLZY0xplt9yrX12wnFqMU9yTg8K2wwjMnVWfIX9bW6OyL57I4
VShL76CzzM0gohwm7OjjCXf167bnu5l+HTTxMOjceoIIEweN1I7t9Ag9Wbg1WCr0+LMzeFsp2UNs
40e5xLVNVFbbRoBQ2ePTOfONUY8RLNagtdErVtKrhRduD/iTYCQUn/pxWB0IlHjgQ7kx6lHbT9DY
CbyYsyrMNhPK100wChzat8BFq/4SFYy+UoNvowcTzJLjHeTpRl7A+/vwRYsqM6naYv4MLPQscD0q
TV2RJg2jx8izdSBy35FgPFrBVg1GkKXRzJTB5M1rv49v3spFfBeXzYCRfHRzJdkbGYrcC76OdWIS
fgMDOn8Fu07UZ7c0Q5mXf9l3xHTdopBWDGV4gXPc4mCSQJDKiiyDTR0iyfErzmn5OvKISpmsZZP6
NXMimSFQgN2TMDpHSlseYjgZrW+K1W+BgrXWJsbVFsksOYQtMU5jrjjmMitHlh7T3dCYLyFQ87QM
B7QgvY21vIaww5QDIhKv0DfpY95mbXXGR1nD9CN52TlJ0bO2zZvtWeoPBigN2ENh6gpFzIStXbum
H/p1ndsp+ySeMTWK0yzbSktVAjL+qupe8GAlVy3JmwZ9os97Pm5cy/OXcXiroKspLhYM0+I009Mm
zEaREa23VDTax/jk5SAy6KVNr6kNoqZ3hc8dXoHroZT1snpC+wz+lu/Wo7TG2CjrBkmOv3it5Zxi
9TBFqfrwjZu2IjRsSB78QD6z43ogWOOC+m6PD+B76RDL0CbtFoxOhzRAxGQ26hNxs5G46cmqWbrp
kRppAmP7A2tRjiHyijSVbj4uV2/xlgZVA59yZM8fKeNWbVWsCVQcjWwqsdnYbhWqMASlfsh6+NMM
xwi+9okUxNiNw5PLutGxqz6MELKVW834VKD/Bq+PupsuQY0qBT5rA5sabm2H4xF4hf41h50SUeSD
tB/K77vk5XRFaU3WlxWW1lBKajEGu5AAyDOLw0+3+YloYiLGpD4DLn117GtaEjJqEtjX1yig+D3F
DxWsS54AEQFYAWUZnImSzniInSTWAw65HJBeQ8hvc94iayDc4MGZ1WgAjo1e7QLd5IvpTyRlQ0JE
0zeb/D/Ghb1Ub2jg8vKW01kFYmQs0Ty4gszlAHf5Mh+JwGV8brC6m8z0beuezkaUYvoQ2lbSu8M0
Id8C2CELJujkjCM/i4vWKOYNb8T8VtY7tyfe37wRXyRr1uBRGL1V9cHLRQWBif64Ijx3/7VlT5rz
czmXIANtJFGVbInfGtQNk4HZAvxQJ+ISZeTE9yPcEMq2DDH5cNSvzY2jc8Fs5Hx6AC/TJUrbNDJ1
aaS44lot3pYxLEtwGGYG8Im/Nz9hmnQJ+Mo66KMS3yXxnLHAv80/Bjwo2Esh6oOXgJGXFW/dxfjC
bX+aosUukTPSEIA8WvaL7e1iP9MfS/9Yh4mAC8BNrOKvW4nB3af+ZoKV0+pZGgEfThhiwSwu7yN2
H6wbXWqD+kA8eHQgVPAd/5oXuDTXX6aYYuW7ikCsV8cxRQaktMpHWpQNvv6ckjnnm3JCMZ6LbiPi
724wYktpF9cRhuJPnUprMtRfmNZlgI8ajZFjdScCSgQFykk+pfES11fifYag0id1HNW53zU7pnY2
xatA1UPP7bRah9/Pk9Y2oe9iHXpvYMhrXBw+9qwrpDWRRKdHlgSjgxS2Oee6W5wxH/MSNShqEH3s
bYiLRRR76xunPcycUTc0v7pmJuvB0cymlTkzoUGZ0QOpne57Kfqv4aaklznKtyfG8se4KXuW9As7
TNdNCnsNcH8glWkMwoNDqXm6XcOyPRbRSB/Q32okhSJWq2ag2bGnRGrGeiAVu8SD5VzeCDgadKlS
V79sb+cvJ/r86rt6jeITqtLmvCtqDK1i5OQWMvQLNWZlnTUxGDMCt5vfFVL+Z28TpYsKUl1ucOZ5
jjrtsSCserZUDdfos/9Y1mh4eqDUyH17diMHeP6wou5F06L7GTYRBjaYAZgVeG3WpvrK8ceui0Tj
d0vCfcLUrpTJZ/y98C6zvt0LPJf9f2AtxOrafc7qGy4jiK5nAWDLi8cbJh/bB3U8iIQnEehM++p/
pafWBjkLPFV1CKvhUoky+hiuCmor5v8S+9AvwUg3q2ufuzTx4OpwimWN1/qa5guhIrBQ+JiaByIW
4uHUZnU/zLMUkx+1cwqcCmoHwQ+bePo6bk7zjUhBDnqGDQFSCVzkc4QFC9B01r11NU6/pTyMp+WT
6kBsU9o853oG6TFqGT97grfEBahFPDvg1y1wpKQkJs8uTkGs0R+AA1+BVyWyj5YIa9a8mzLMvDZI
HRgcPkXONtplCHF7K+TYW0xhyV0A1qdR8Hr8/om6LlAWCRISBEjwcC4KpPU0wYz4mqfUzM3Hzuxx
Z0ssYkkKxbiOjH1fECbvlpvTc+VyQYTH+r79JKfTy/tteM8jTOUGvsms/MfsOVwL+SsS7EwujXAL
jGpbJuU+0f42WSBsL26PByp76seZEcZQE/d3Om69cWwOQIuW7Yzp7bkmqBSYAciav3Kn3kyrRREn
9TMPZ0w2d8YIN/S3j4cSjNDK9ISimKYZPsNJzEK0HVVvwUAJX2wiO1RzcYXxEkuMpKy80+rzYgYM
3weS7TZQTYSZuo67mlrVf7JnhCFj7mFGzW9l8H/A00nNRPd/9rSIyzxhK7O/Dazq2SVuLrq0Ilek
xyD4vkrgop4PKtklD4nS67j2sOTx0Szh/Cq0kxUWXDwaiYntGUXphIUoYaXfOVPZbfrt5yb0bx7F
l+c4iJxzvCfFzD01VHYCRNt6lSCJTaLrEUxr4PQqD8EOLWjOA0ZVgLphFTGmkbd/BxzIW8SD0pZx
8NUIr6SBQDZvvmJBdEQt91SM+ar1/fdjbLCMCskGsB/TE6egUmiYQGMK9BdP09xP/VIFJmZWq58c
0e3y9Ic3/XoppV59YbVHfVR/OwcssicLnGrFIxYtnQCVdssQx5OVJP+XWKooE8HVZvPFRGYm7Ge1
vQP2dZoNIbE68Jvs00VRSbtJxVezYmmS3iS/zEIk9wmKEn4kCA2m9nA9xuRI3rWmRz5hHNfu6fIe
SS4Y2UTU5q06lzrqfciLfMZXk/1C15Y/v7xhUCjhA5dGq/sCyXWDM1/DUj6iBeoWcpsx6pBiNIJZ
XYK+ARtO+7A5GscVLdk00JpUVTuwAolaeKlsQR/xiCYfFr0RYzydOJ9vfwEBPhJTO0T1B8jKRPyW
r9HX2NvFVYV7VIxMs4UVv26kI3B4U/kIMUW3cv6eRICqFJ12la6sP88dCWQXqOaYq7SvXGPIVI2z
YcdIbctRukLjCQrnmsIP8wd7kEqR48MgJ5u8xb/dFzi7/o9R10gWMHDY6PThURj3ppAbwJAWESxP
mckKbJvQYHpiU7cXnKc8bXueHvb6iRqcKr4BUTPjsUicUjsmnv/+T7A0lCSvz6Jhd9L0cj8sm5Ks
FZfYhj9beK5iu2/DHYiIpS9qtacSF74aAclnOPoDTneMsjT8ZiiXME8iZc8pX6peKjIdQI23layW
eqDFAd/vUsX1V5koEUKEOIdNUI5bBR48kv2aTgyJiOdZtTCV3k+8x6AvaoQ/PHGEC5DI18920iT5
6yq8BXx9gS6GgiFu5i5/FVopEzm/ZCmpZYLjQsQSH603eI4MISwElnv2mjb3mTcwlLxTcCoSdw/d
qe9RtlGKrnT/idNFovS12vKgtUauB7znb8/qfGEMfxwc4ySYbQ5f1q4Xd2kBNx+1znP2T9wFCGF6
8kBpQi66V+2WVpma+gnywgKGyjDLy/F69AYIdBw3m5WRNGcL/hAyub1Ogo54NxX72OVsH4hBjrv+
vL9OO/ZZJLxIf5F4JFXPds7WenBFyWZmcVPoWGxfWLX/2J9UjBesXhXmzeRECyJvvX2u1PuvmUyR
p1+jUn2Mqu52lI9Rf9BVAhTPaQcm1yCToNDHHn8E6vKExSMSrzVs5f8xNnGPiZm93Yb3YoewnFqN
pOTeV+75lYnDD08fuavk6FoxXh88i3LVGW5ZaRv75kqSKzUm/JwcIkYo224kN/LcNnk4lWU9Q9Sz
3cG1ZG631tw3LJV8RLBVBuwHFqGLjXrJ8NrLU4cnheuB5GHEVIL4PiDs55duwEsGO2v03BKP1u47
SME7Rc+9aXDME2/jE5JlBBVp+p4Ua2Lw6ocMu1bqglOyerxCf7o93qfS7O8/e2huFIts2hlRnB9I
ZljrrHP7EDmv0oy1cBTQRT38qzCvOiuglNPYDi8tGHDNwWi0LnG+vWFAdwLET705+4fhV2FrWsTX
IlE87/PkMmMvv4qNAO9G6q1vrgsmsnsgdt7fxeoVq3ckzeqam5HDgGNiEj8YI4twahfrMuHFalzd
UMaYicu1Soz41nxGFzTX1y4zQ3RDCaEQtiJKNDoCoGRz/WQSW5FMeuIAUFEF+SfEdlS6XGb3m1eo
BKUaktbPKp05QQpaH0aeU5pa6WncY4ZjL5rmAWgRoagpx0d0XyCPH5N0oNwXvlb/7XJQd4jcimOQ
xjcEbPUc3mia0rfRItNsMvQu1FyDACyPacZ4avAPC3aL3c8CR+tNl00V4gpv9dNbJPRWxivnih6s
abIZq87mgds6IjzJ2C1ZsTzmAXUnnhoQQjkIssLwMmUpbMIVTgsjxTtCjBR8A3Q/PAPD3taBeZNw
V6NlvoUU0xP+MCZchC4aadvrP+uGMj5aMoEsWUNqP1/k+Guah6Zwlhn75zZoe6iceqtggS8TYFU4
hiaRL03QJxt8rNfbbxU56XtgLGcAMIZrBIZWReMhECz7iVEnqtkedY9ABPzBwsmIFqqYFURBVUiE
mf8QPgqxskInJg6lgxCSTc12w34lVcUdX+OJDgysEDP6apP3WT33qUPq79b6hV+itzUgesbItWf5
2knkxjCxy2dL8GIrkx0UeD9o1qYCS1wURpdGphI8/6ZR7MPgva88YHSEKVDnH5wdj3LQPCCP1Pwg
T6aqKQIRZ4PyEqREWHoJOr73Y+lGEn9edIvIhq2WNPX7DGNf8Qhzk/3PrR6YwrMXT4sv8L5PJL5c
9lemQdNCZt8VwdQiuoDTR1RFuDj0lvDg6GuebT8ds9xH+HgmflG9xGm6o+1B4TzJbI2SUHXMnzsy
weuHsRo2hWOwZI3k6G8rlSpAUHkrMWmIVxpWAY8UDFX4+h9h2caY8zIqF6Ygjk+Unu4eykg6pz0M
qQIPYi1kvShmYl8cnBfCULKMDheRJqQibL3O4JG6KXfbc68BJBvCiM4muhP1ypdEALUtAUzjE8H/
KjU4Yk3X+qH5M9GY5Ppg0C8569KsUxMRR58TNssI/DdPMpp/3d6TEQM9ZvurHDfsEjugMd095e/8
jmFJAzKXd9dcMeFsl47/EfQQ4pMh7Y5sruWEYSev83tWK2B3wooiOa+JDRYth2Es0T6SPZIJ+7MY
JS9CTf/EXjKfsEKV9hxP82QgCtbZCwi1aJAJosGWQsgel9yzBsCnHBfMK46INAwLHJ8KwDNBy352
Ib7uG5NnO2GIKMUBcWt99aHYtpa4SCqCC43aarh1hD/4JoJ6zwckjcBUq0GReDWdKw4GE205Ci8g
2X0AqWEK6bIGHZ05uN9ELiSSbV1bYTaHL4itMxIn4kHW1xhxVmwiqwFaKuTKBe/xkFRY8xRqZKLL
dWl71x+OVsZnZbQ1EROqK6b2Nh9Y+bQGTciIajQ63SxSNwwgKDKNraozQgeTK4BdmeYJae1VV8bg
fbZmSMIIMQbjS/9Pyx+0WGnjUN8uygimQJOEvQR/rctD0VRolqWBqzlc7LMpv0eqb7/SzM36E530
G/cL1p1JpUgL5pqH/YcGFPDpIVNwGLXG8cgnmb3pbRFa2zJb4X7Ln3Qgyolw8H1G/TvGlhEkspfs
Ro5P2WQL5DKpQ414Bon2dflD3TRAZjKRXwNdSlA7VgCLYGF1/K0edbgBvVSglYWmQxAYOHG8glRD
l4PsQTIp+ahwBF+dLuivgGaFe+EhP1ki3/jVV9Uw0DanzLVOgWBhcgv+0aKGSOQmq6UjARmC8t5+
mccCRFc1MYTIdjIZSpqyAIS+ocaYJWgy0gnSrNQtLD/n4fJGNKx93WjZSwxlDgep1htByd+yfM7p
NRAoDUEVv1GfK0k72m3DJEspoDlqlyZxyEW2J1QdDpG8/38Ek7DyW1M8LdltdaLnLs9RHcKbuqJ8
2K/fvXWA822zmrwEjewemxbbgtvSkrP8Z2o08gGEBjS5e75x4TkU+LnSGg6DUK5/ZorIO5jPgkNL
JOSfnwtxxuwMrq6rO52Q+3wsxxYqq5OU/fNyrx1dzzyFFHZw7HQbcNMURJ0W/CmVv1K81ezgQtC6
bEvYfmfuw97l3250WXY7//4MPXRgrM1/jU2W1JHdbhn536WkILwdL+X9rm8Czfi70DWGPe+wVmCn
GXC0Ek/VGp6imyvnuZ6tcqM+Iwm9H0z4vATF/g/MMjfn0Yzc6+xpqgy7ZrPlqsnE9Ppf3pLXDMKz
V8U2bGiO+zvVd6j6aDxvKtBqHkyotCfh1j3m/UF66+EjxQxo/pY7DBLYQOUlzurV9GpQwNYT15e7
5tiJAEy5WnP0lRjODcpUiP5J1OT29WceOXeRto+eb6NXvAJQZeZImQGyy4nJoR22K7DCzM6R6Co6
ndE3zUXt33k/qOQ7KEQTjJtqIDpzvec7nfbbeYp2/7bXtyAa0t8dilr7uwQHdnpO//TE8NFDiuZw
zWY+YjwkqqJqV3D9Db07euu45L1MqNTPozc37UUK/BUC6w85bfUpAi6qnsd6I4ccDO3YGabocWuE
U8tv+WGiH3DSfkMKsBfxz8vulMv4ExomG9Dn9q3VyVVC09hGYzLPHU01uHmxD1REHFk0vKqLWeEH
aIaUiNKs9ZwZYjP9tZos2vnrUhfgc6Y1Lz9HERoLSCYEM+lAohrwftAFIk83Bnm7Ya5gsGfmckNi
Mbfl+zJPIZkpjMVkeVoKb2vo1SRbaXC7Qr6A7zuiaOURgr/d7ikhg3HCtEpyG5NXfblpxs36nCSl
6SlxMdXaJ/zCq57nQBtkFAbyULWFLQJO9R/shaaXKQYehLRMqTshJnilK/j4hggO8C+YMSUpkZru
3O7hssVa8FZ7HLYiJQyXabRX8yzrOSqauhp4EIphhTuXpTVGHLEg50+W64Gvold7v+5NEPk3QERi
u3UbMADdT80MobVtVI+lcThbp5qLrDP4UOEFu40ac2nAmCpLGfRQh2EZmCncDHB8lLdcrh1kN0+U
g3rTgSz2os6lNvzKgv8fIW/kTWoPe1mFCi9al36SXR+CAuLwK+ks/PJ4nAErVo6ScVPBHT6pW/Ng
9CQicRBMypycE5OhqGCixunL59XJwAOt1tmMDziAqxDrhnanptZGX9U/zH4nziNBCEVhWnfBs3+i
zustzAvMz++UZrahv1q6KP+lSs0jyq2/bhd0tL8O0uZRZns+9aTiNFL59pQvnK5C9S/NIS83EpFo
XGtcLnnq+WLbFz7SKiKDYR4r+tbJFRmhzyjnmkfi9ASOFDwjjq2U8LaKWX/DbXPaFqpUaqFOWObk
LDAcmhuQJNMODGb1vuFZZ1FkQx8uk8YuUSb2XjQbKBdUsxS5BadPAqZqzgli5YZGwvuOZn2kIxpl
7tj7nHmWHoSxmfSo17lcX4lYxdP9srLbeZhDnXObcMa9hb5OsETS5Bjqv5v5WRAwHPqIBzWM58Lc
7IlGLv/WWvfe4WkcDIPcRkAJzTwR5fdqnaecBfkJ7YqNx6SfA3U0Z1np34bZbpa0pG4LeSAWxd9t
c/fHVb3w9bgB+9dVCvYUBZ/Ee4O2+uIX6ydYKsGAWk/lO9YjBs90w2b78FceFJhC+/M8aJOXjWMW
h/8mjh0a0Kep2TLxi/FS377x0hGGjjdwaNim+ye8ePYEcVihXHIc66b382z29X4m6fLuDsehhCkH
AA7CkzZX+Ma0oaxPotbfHUEiLxUzTXrqqJyb5xkCNYcZ430RFz0xn3g1Z2e+tFGJZdlF/NqKpHHK
s9tnY4zmNtNZ5WtwHMAaAHhHvp+Z8utVZC/c23IndULqR/h46YOXoj3w7wfvS4sh0lXU6dY/EqqS
OoT9kJEHMWooxKc0geYlbWAX3FawGWCN8n76mnBtxdsVLymezCn3d98D9T9SiX4I5jWQMjoSnbNq
35nPjefThotmUB1/4mt70y8OC3j4Ugr2l45qAmYoLC1hFduzD9tyfslmh7LEPl+LQWbRsygECvGa
oys0eHUiWmBz4nd+lK4UvtEITf7QwhYESLosvHXQKgdlZ4Nl4k4iQgjPEVMpZ01EEASy1baObfEc
1gWn3oUejmsVznamRWOE6YUrJvdyeFuyhb8vCnEKCJSrTd8SgimnDf+BA9+OX9wRyJj1kwR4iK9g
6PWLIZfs5NKP5CS0/3A7AESfea2CCbw8lujGIikoQaOW3rxQaVHJySyefgaLxsm9BlAFmFzV15j8
fGCduSsAoX8HStyVbZx1yzK7SryCNR0IyqRQ+5m4rEr046BCK9pUEUKXuGobTen/MaWK+6Tc6rZ2
jgb6K4GCFS275uYSh8QMziw2GWqUmNuOLeCkZEDDeCIs0Roo0gHinuRC3/sNct5Mnptw9yI9Rp/8
ceK7ODYtObDKnyjrWcmqdLBsfR61U6491eoEOEFETHN5CdAhxr+fkcYkk3QGW2ybAMr/uYJcMMPQ
LX4VKevGJnwTXlU5bzma7DPtyu46doSoa9sJBCmYVo+jr/uqeObfb35QGrBI3XWAe7QgMA5DzyHW
Wkgt2+QFN9Nck5dnXt7OHJC6RSHf1CSru+zfX8aVwSD7hGUD03Rd39mco8XTu86VsAp9hslTT/92
sUYEhYAZM4uJSxb4+2TqWrrplvUYWVe8qIydHZhx9Uw0V4zE+8CcRUNIn7aE7DxvJmjlSjZpf1TV
ow2TXnybEpKTZjLY1P/TXbGZzhdrUpjCB5rS9BoDv7MbnNdJa4Q7I37pGk+rAkhU9TY0r9UXvYG6
C//2umTpL3bhlCchrxvYd7yoNRebqt2GyHgAh/1CxgEuIxFRVtEM8528B0rbe/FDZi0fiKvaNch2
xikhvtwuYh3AxSMPgmtFRTThix+X4BhlHRGO8OKZdnbP1sKYKwl9KvHXggaz3aBaDQRaNtb1MY9s
SndmTkbkxljaTvbY2Lv4lyq39Dim0zqALXUdoYd4qly1BjdI3ENfQFf5/cM2thki5eWGJAe75Gwt
09tFmjnqeMO5XamL64ODsZCaAj0/4hWYOBpLCICLe4TWZtuaJ1CUgPuVH/kA6gMEw80XixgEWvc/
d8K98LiT6QSasCU0EAOYhsXAPh+xLNpMknC3NVfccROwNm/YnYan73VHbEXmfDdoSrBT90a3h8zv
j6qYhZt6hjBYGYgonAVHa57M/tyQ0Szg4x6sa7+ZoIPgibKlnovsqRoGw6ZpfvWG6hdjHjvDKt83
r4kZxykp5Q/EfEfTa8MqkAXzaUo6WcQ4SAmZ3Mc23LCSaE7PGhBJFnCyFN3klDLMaj/W3B+blVNp
vjKh8nd7GyERvzLoUBnb8AQObdrJea7Dwug+Ehw9oVw+5ADbW6FVmVuKshbL7N4cvKcYHBkOOKDP
u06ADnHTne3OZzPBycmVEQo9icEam0AOKoYuaVUB9wmCfV1HIHoUoi6kjn6d+ESSGeLSwqHVLQ2p
GK07VhmooMnVk5KWCx85c8bY34NW0VeCbzFCME6oNQyFYIM8mTEowkXvTkGNxlNlBtq4gNngI8Ys
00jBYOnw4UvKpL3xPKB1esUxRCb+BU9YhCZ/kMM74U15YwUXnSX5aWvX3CAJRA/LrG9I+2HB6Jr+
sG9svNGEBNYcltbKh8FESosLw16GHFobYEGNxIL4dZKXRM55vVZGILDjoT6QIFuFAvYmpxMk4kKf
duKdQ+StiMMErJ5cS8qZDX165//5CyXU5zurHtZuriOYjcv/oNQZTXjMHPFwW30qJ+VO8Qn+LhlF
LomDbPHVVpmXTvJLO/XpbwUteYwvBj7bMVNPdIChP2VArXodKzJ0AxB1gvcbCooiUjl3NUaYCsvg
u1FzDAPN4qlljKaDjTBeuRqb+ZB+ZwxnU70TulOlp05syARG7HI3jeX+7tcj7dzrMXS6hiP7zy+s
pg94G6NZPQNNT6Xiq8svTqrWDxhA7Ggnd+U+bzmWAPCzzYKwl78uVW6s2QZklugTeECV245SCT4H
ZHyRb3ot+BTWjxbz2Y5Itx3hulDs9gtWuhFR1LmvlX/O6Xqijvg/tRRJlGJWx5BlC4sCjuo0ncxr
Zs04c0EShYxiKXEM7XrgU+LJ7gK9oIPycLTznIXjjYhcRFhze9vwXHW6mPu5V2Adw/8tfXJmELKK
pKb4xb2H3FttvUk9O7nNFyxkgpQGz8BeN92nC643FN6ghcV5bPaxrA3I1zojvLMRfelc7gMNXU09
8LecIUKVSPqnCljCj66BZiGS352u41Dbb7VtwjOxcU5SwtLR1NpigWHY/qu8sqiEYFlaEaijcabt
syZRLzOv33ULMGkI90HDDRIuc7cqwbLxQhzuUUGIci+8tjhaz0ZG+ZFDz9ub7tegSGAg6zo+RiD4
onv5HNScqRrIDQmnL0pE76TZ5fhIQc4JTTbIQ/AyteLVE1I8Jh0sfd62hMVZTWavXzX6wwJwLp5N
iI7HXlMPTsBd0TvRVzn74GAh0khKm9r/Q7lzzGcYZCqemLXAy3CBJT7DslN/eBv2kYlosOLtOomj
e5gHZOgV9aqa80OpSJg/qMUtCaUt5r51kmEpRIR+tPekp5S7tqoYS6hBNA0q2Wp5skyn87bGgTy/
wLUqWbruUqZX1JfBDeGH/3hExKISHMzTzcfLjRO4a0o5FvqMtl1b8bUO0bIOUAto9lJJOQNfRz2r
KON4c6ao8jZpElXYVDuM+8WrVBox3097w/SuAEKTAC6nwwP+cN2wHFFJ0Ky+VaGeNlVodk8CBHHk
cB78VZLsb0yW0WOJ4j4gBJqAwiQJHlN+eBY/UBayba3CZxbH43cnO8yK2Lb9IsVQwWSPtV8axxan
DPsovZ10NtvVMMN9N3JAbl/jgWznyGLkBrWEzO07/5lBIzswHQ+cEyPzaQJome9GNj8e126Lo2Q6
dyKT7Tr8CbtTDzGb+uzEtyJ++aYe20PJpp0XyuWLPWCriWxHNe1LZ0lxefe8TrdUpUqrY/6JvUKK
GCTmNK3KQAS0klJzm9wQM/NxwSZuT8yC4Gzc3vDq+iB/KzCsnUkOKMB+gxkKS5WD35QOl8lhkorw
cFJ9gzy+Hh3VOCSljd95jTI3LzJQX7kMgLX17pn2MCu2Iw/7IDoHc0zaHlBrv4z9pvbYx5lEQvVQ
FAwwwVGZqG/U9jMLiMlwh2r0X/y7pxHyzyXmcidpksn76lxvOJut/r3cWtXaxU9R38ZGs94n79V8
Q08gOr6sR1uEA1W4QTRs1AYnkExAfTVVn7u/vZ9JOr7DeJ/Mxk2BICmGUr1t4AZziuGBBiMYT0zj
oufV01uzYB7nFBiwZLrRpBujRgJjA01gxYeT24LV1nkDX5HC2HqzjPoTHahzLox1wpG7umM0zj4u
9jhoKa5GnCom1pCNTczYZqoWbB9/VQCM1a+9RDzwRNX2M1m9fQKR3N79r+S6XLojc9D5r9pALCRP
pGk1LNuMoELlw1okjOxlDX/pJ5ulA3dOTeqnLjW+g0B1Z/Lp26uhsnWLpz3LMjhWrEuR/D2nq4T1
3E5HxYZK77dhQPiD01LQHl1lUanVSYCLflv6BLLjOT2Y8IorwCrkLy4iIDUBOWVuZqjRUFRwhceb
L5pBTMkuVyvpNaxCxJ5SW/YiF5qKMnGhvRFZtatGW549hGgmf/O3Io05MOcT3FTobd0nAYvIBesE
Qwz1mjigbmrvO2BpdcTVVzjCyJcnBFSof3GC2e0b0+nMk+oDM4qIWk+U6oqyRNnlOoebIkFKGiY/
w9IZCrXDl8ByaWScmoRKem8v/D/Wk/tA+bLt3AI3XP4J81aGtLfJVOvx//97CSD3pi8gHkmgrk+5
a8mGewupm0+XgD3UNum2JNtOXaT8mmKzQMcpD81rjpI1iMU9xVlUNbVDlq1+ynN6HIWSk1WoP1Az
i95seXQ0hk3spR23MG4xVLQCIOquR8Gop9MottwTw3lVHpdwUCLxJXnMS++wcMd/KIIjGTS/eY++
nPnQZMBZ4a80FE6tpBb3wA9MYIcvYpRAR/Qe5QBCBZyB6cSzaf83eZMUjzPPSf/CD/rOri3padTo
m6QmxnaOX3uixh7FAUyRWJYnXXLZK8cIcYwb63yfJw+op7aiamxyyB6fmvk6Qd18PHyjp4aW/NI4
/7XESA3L0sG50h5K4X3RbWUAGfUuULSHdiAO1kTBtpwS5rvwbAKZZtC/h81mSvZSC6pHHQq1kK3K
HVcxoU+0xOXrcOXmboCsmIjx612+S892gC7YGjsfJs/SOKpg67C6YQCg3NyWNDYKewIOJFg8Nkuy
wJX2KjIFDhkDp7ZgVvXJe96/190FPgVWPighRu7TfI2FJhvVbg81QgfdR3jhpZI4tvVDIlNcdpPJ
op8B8fjVBbXwfqCmPX3AjSlw7y3vzJdGwHAmK/BgwO7g2YeopE++5PbMY5zvDQ2RcCR8QMEcRowe
yUJjIVgD53BYkfpv/FlnF/DNE4soVnwcXSPVm754pWGy9Q+W2esKSHlsiDWPeNyTkckrj/jkXjxg
FN7ZhStf6wK1iLmqX1QUtYP8VcYW5/JxoMYXX5C0SaR5NE4XAhISHEuBpRJN5tPWxpwrxLeGbS2a
edGE9YhYgwFIWlPgBFXQ5Nkd5Gc63eBv+fRQcOF7p3PoJlbX9GLLzNSGulpdRntQVCm2yfF6nyIz
Uz5iVXHLN4eMLyEJYtCUeB42iR22geWnviYzogzxnHj+YbqIGQZtZ2RwlTQ2rtA+kdVKDaCkJC9i
A5t4aujtHifdloZo2H1eUfp5VbrooOYEMno2DAlRhrfegoqWeCZdn0XgGneqS9+TnOpjxyYy0Fpy
8iFFBOiEzrVr+iFgr3hnHFrGcGjnsPp/+Nrz23Vl17tU8AkOxyoe65XneZxfl9D24zOlGJuRdRn5
t2uLr9a6BV0Ukc6UxsTIVETFU/AA3WIDg1Q1NyisirboX/c7ZohHXQDB9BEvuu2us8kho/WjJ0XU
OPxPMY0Vldi3FKjw/aae2UrxkMwi2/0JnnqrlD2dl1HYByYyKgKZMnK65TaOkpXx+E5rpSGrd+Fe
5RiiB0prvHi600tVMZuzKyd0/Mx0ZXZeVwXeVZM8T/pC0y1ruPwY+ya54mVWQqXrAJ21riPH+dHy
bSVxkVpjfCVnRoPQTnU9OZY/pmAWN/FXziyUmX63uSDD/imTfL4yLx+pxHFv4eKgQGc7d+rTZgG4
pWcwBtJ67fpI3ucHpgwQAc70BIaeVHDg1zVIH/Fvwoqt3pZ7x2WEYnqlJTkXJCdB+RBD9jdCx59k
BwecEeTUKuiqcJhzdgey633pFOybLvc1DmDOWwC7NytKiadjtoa5J1SCHZtFGwArda+bMBwbDPWZ
h0aFcRz966lsKfvzBzSnAB3xgdwWMlxfzXkzjUpPAGOcMYA47LFt+yFCDHsMOlUC6Lug4gu9Lh6C
Eky9ZFJ9CYvT0F7vQNbmn4NYIAaZPCDSvXMFGexLqr6u0f5E/oxqUw1N44cYr4w3mSXo1mXoOc/p
WceUeyoQNcbkS8VWeGUZgrhE5+4K7bcAhetjOOLMrBz12O/Kcu+j9Y7OLe0K0QRimhjMEG4WeE8a
pqXgRaJZ6mY6xmdfzntQfMdFrxY+PnzP1mTnlfxptpgdqxWa814ICUyUT+xi5YIhCcL95iyNCXLW
1J4mqAe6K+7ckMKWbuPV9CsKqtwwrCGQ10Wlw0X/PjLL6/DEJhrpsDCtqm8mS/DF/wPgIS1kxTF4
kMjrPMzHKxxPyhYPZD9ofH1Ki0FsUzjwxgaozQkPQnCw/rwhPnl74+/GSV7SS/FSGzPtaYX9UIPc
Y9zPWfbDMjG2kewd3t3N/NX/LYG/agslvfGtgXvqaYDb+5RZdPxOHxwJdvrI4ytYDnjicz6x+rV3
db/BSlqM6iS3lJ5BAYptuZRRVu/gGVMRmMiy1R8vj8zPFCTIw7m0fbjWUD6aZXpeBm5HF3d3S/Jx
SBuGbt1iefi16KcB91HOazE9/v4M+9Qraf0X4b3GLm4Jep8/UpT1sDeoB9EZM4+L7bqqxuKyNgL9
8njTF891bC0usiARaOh9mecEudPJLiSVMUW2qzwyonuC82rgo+P++Z1T2quCLjvkiMgDDH5EgnRk
2BcoKvy/JnvXMF3zHfiwOi+WJTbDYRpySAqqQ2EGj+8GYj/azco2Nyc+Zkap+YIzROR3Yc1Z9DBi
iBOJClTK8L478q2tThw1i1CUU+Ep/oHbvX6hWGPFfUO44kL30vjzEYXit/s4QHvAzS5VH8IeUf5R
mC1yFg1BgAsET9z95qpGwEu21tTaU6x3zxWwO7O1iPbKwlBnscaApUU0nW4CVQmOXrOU4/tQGDgQ
NFXGpS3ron/z/pwhTuVs03XmFxs+h+UtgSly7yAi4TNi5z5Y0idFQLl3Kis+6w5YFNnBZkQodR1e
d/zuw+kHOXoQSxUbV38rXG3KDCsH0zCwMnhXug8d8QIAHTFK+1i+IP06a1J0zMqJrdJeeVnMJTHu
inbvWEDsHzp78fG1SgiNoew/mVvsfysCulcLHpCHnzPESnYySWeHRU3jJSDcu0g8p5WfHVsztk5T
PeJ5j7ltGPymksvNrmY4TKaZiat8cqOS8Q5SYNV7V8H12dnb3wW84O3EvM+xq491ydvLE+yIfgGl
1p9/5BLznNtmhXEIrHiNbDGrXktYolCGWHwzjsv8ENWWXBwQtnuwSc4FDqAwJLZWgzJd21QNaWML
U+bPeU0mmvClldcVle1F3yyJbwhKtS7OyGmpSEGcw9zNF1UlYh8DSAqwACiDuy27FzxKlvFaA2U1
Qj6XimqIZQ4OQuNrLpYuCuP6JER2GglAjXnwaAeZ2/1qWlDFGa4b1s3JSDjJc6FrQB0RtQ10M1OA
LxTR/gStVDiYFcRyNwBM1QT4o1G/CubYldR/L8P9G0n1A7oi9G7iz5CSEq1ypxfowrilqhY9zOLi
pIzzTdTv4Y1GEkyFyiIgpr36xVk8db36aFEHigLS8KTO1Iis6CqZICNj3zbnDOTGNQdzYjPRpksJ
hpF+6UUAN36NJzUiSfazmD/DTOoeO4/kyeRroJq9YZ3o/LDDQ/xr6fkA523HGuFDFHWgB4BPqImQ
z1UWYcEN8gwddEqJZqXnnxj2h4K6plOScVqgzEBeyFkSXDU4/eeXbG8grHdkQBFctRfoNw7iiGF1
NST3RuveUoj6y/ymATTATn2r/WEMj5gpMxPR/6beVtzV/lZhiMfuys8tkjmBAuF6eQMROteThj7I
dHhpWy+5YerS2FgnPBWpE5Vhd4s5iDg5axstlHNpj8M5wA9iP4cdMu98409xCXbgkXGQYNjs88/M
vo92Ff6AXZiET+t5TrKNoIcLcOutqep6K923EmxzuebfWn10KRqvdm+KwluhVFL+/Ae0/ONSg5Vm
tn/cnu+QHScT1jBD1Fsc4Ujr060NKJCoJFZOmdUBpxTkCdEC1ouLiqcx1QEFxUjMbokNdk3O9ook
Vh7BJ2RMLw0/XL8+XwCQ7jbNn/tqjx5bX+SelLZoUCXhY7h9RtIIWZBPnTvTVNMKWhVxpbzIopSV
EgQg4GesG2GSYCgtHXDYGhbHCJ3RAQY+DMb0DtT6aFZYiyAFZndCSF5dBRsq+8tVa7JmbsYLvBo+
7uhBA3JEfS+gqoZR1I8UpsSXmm6dgDGRQ0HBXwVxK8R+sxouZVctRJaafNYwgxdJJsattBrGrO8D
PJFuYbev4ErANIAecytFWQuE4WaVj+IjnQw/9HYNcbttyKXAWidtePbS0BCCoWzGmUlxwktxaIEt
1TpWIm39flkjWCobW8BLIieIk1/aaGB+rZ3fCfb9ELTztioPS3yuV6Uj2duxECDDILE3L0kmNIrz
wpJ59yuyX+9wbY4Ds+g/0wNp33lfKPPCKFZThZNedEJBE7dCggsZBzHNxNO3b1d7s094ilXGIz78
Qcksv1mZxJDHASJgkV8EH5CLd2+EsWD6DDGccr3/ow/4SCbOwxeoMvRm0xVPtwcqF1GaVsXEkIYv
8qACW6RhIcq1t6oyf69rpnVIYtmXr50NWsm+LYREUj31tunVfXx8FXH+LqWe6YCNQTj07d+LOf+z
AP2PWesHNJ5cAlsJKaod2yswK/vA6gLL/3btt5ZL0239xYjlmnn+GWEBlf/qLP9YuYtEQovjVr47
ocad8XtgrOIJ0xb6A2FT6fEfVUF7ekK2TJBWD41nK/OVQwqD+VVmERsPAQnnRZgtvlrHbY8pFqD+
Yprh5yLp18yN8iGUjsX9KbAJ935Ylsdqilla1xDpaCnoFw7WEaGAJz+F4HPBWRLo6/CARXYz11EM
n3Kou0rzU8rHsvuDJpjlSDUDFiPKtJWzCynJu2F0bGj4TChno5Ym5vjhP+9vDpPeWaq0qO7P7Kzy
L1QS83InthqhrfKIG5cIezQDCg1nC2cmxdlfOGQgJ8UcGhhsj58XZaEM20/ALrld7IFU2Id9/Kzu
CDw39ylWRqfvprkn774VsZyGjwDSyZ+qKVazgCiedwC09AdqASF/UZHvrU4jHMEStdXzvy1HBL4L
6uj2TthIC2JLxEleI/azk1xFyEZCdQcoXDmmpVJFbqLkaXvl5EZGKEiHSD0yyduil8+jXf6er8a3
sAKX25/Xdzs6by1of/nGYO2YEUeO6N5Qg+X58F9NIrrUGo/NVbEVPKt4dSPw30/HngP7SX6NTZrq
4qeLDWGdvyWlecdYbkG7BMz69UiPWh45fDnCBv6LmG1qtKbKsJrSsMP6iDINM7SveH7xCiZ8QOzh
+2Npn23mcr8Kk/BNSZYNsHDWaPYQSgD3D24qOf0P8B1QhVn5YdVCSLJdMURNqWF9WOXkBIe8ytFQ
rktS3hZxOfiKGhYdRxnZKhBnIrnvROglRjgBnMYeaM/31luvmLL31p6kjbnfv3DIh2rpI6jaxmrL
zUuY8upCwH9DwvVdMXqZr0RbP3V1sfuSuN1cM6r/ZKxrt2a6KQ9bDzkSuMMZLi0tPQKfLvX3uaR7
q8jKf8c37UxihKgK7XrsAR+uKhkmEuov9OYdpehXVaU7I129lhd1AN1CfYxcB2/7Bl2M8GzOuFVW
nr2grZfkSwzz4qhDuIIegUk/5z2EybFTMwY3WgHGD6w7a1s/anGKSL9IMc8CTVg61FtiKYsypn5D
5VxuWwijGpz37xfjgiBgyjYhp2desmjsS/6y94qwZQDL2d0Ao1hNi9IuJT0zbauPVSVWALQkg4ZR
Y0atoZo9OTN+ozx/c2UnCKRkkIdtoBF168pMdZbF2nDRZln/ZqVaEiNDvdUCuHm36/BcXGiRT/VM
ZoXJu7GNxogPzMNExBSn8uhcxWBV0cqe1ygZKCuuKWkJrllZbpLU1H+y8W4zqJp7/rarBdBbPkSd
NQuaDzcmC40ouC+T3/zimX3jRUeE7SndKfVxLvVCrBFTqPD2a3mYWg/Tiwh5oGlftJ/iSAQOgw7F
mWheFvXLFRjHmW+DihVHL+Ef4qJaGLSmZMb/wDFu/WOihUvAdthlX6EO7zysqV/cCV9mMvoeg/AQ
VEHPzFurXkcE5oYhyN/sGAY/TBvVffH3AkpCSvRFjUuP8tx/xWBX3RLRUxyHYdz+1XL97SIziRdV
89ed3/NXsrTPhiXiFwdC24JyUlp47L0Uqg3QjCW2xc7oN1XqfwCTXhR6GozVGyUuynrCoNvGJw4P
YSc97tDwSxW4+djHpg/2+WdS9hHQI6VdhsGh7STz574OKOvPWOcfPeQsCAthjbNkTsG1nTyL8aoy
VhQJswIuYGAsxV6rvsV8gNKzXvZxQTjBDO6JrBVkl30dUv0+GTXPCAsUGGUSJeBcl1CeXoPOcM1M
ZgbAFqTWVjCC+b8yrfU/RCuQBPd31s9JqBf+8GeQqdyn5J9xMc6l54aG2bE/jTlzg2oCZSYL4o9P
WvmnaINqVRhpgH3/ZCsvR7g1f/P1dQM3ATL/NRTKeE5ibv2BfkA0CsxlIH7tk2GErHrlbS8Z8Umo
KP5wJxfyzO5kKNeCACcx7uRmitloy6k7dnJ+sJ88dGrwW3VjiH59nfzSpbkLF77fDkRvp942NU+W
LVKfQfTc7cpfoff09D2YPGUJJNsnx3uf19X1RHOquMb1X5f4OvpgOCpMlhM2Izhc/fqBDJLFsZ8P
YUW3kNXHORn5tQCXQYi+FBdOYge7tHHHI3XvkcRd51lRNGUqLs78C28a2gL+TXn7xWeRlGhhg1sU
xKAxqEmqhqouUqimNq0lEl0C6bQWd5kmAEwVD1bLmdR5NirerVDsU9VJIl6jTG7AkIVhADvVcm6p
lH08tbPWm1HrWzm4aJt61mT4389ov5Qs4DR/vHHTJYOVmUOw/+Kx53vSAgL9hDTqVJIXpkSZMG+0
1pEHpVutLcfIzFdCuXXRt/lJETnQk+OZlDhxxH7gzZlq0gsvjAsw4uhsTbycEmHeOmL248B8/Tdx
IHMfqdx2lnGGuxLJGRcabaqStt56//73/+Tau9jJS9/G8MPLjEh7zwz57lqAc2yLcvxFZ+aiHh6P
nScHtNBBSqBIxtkixOdGI2Iykg7iIH7o2cBfMbwstC64d+xQJ8HIdL3uJw1aHpTAOWRIdYJ3m55B
ki8NQt1VGKA0LvjRoRsP/qUm0vNnTAasaAmiJ80+G+edqZCn8YuH35mHevr/xZhWV8xPSfRLjbio
QDs2X9weTBCOCdZzDsBrn1SJRPqA+GSFUgjuhI9/RXMJER+b0Jix+kQu7u5E2tWhd8sZ01fwcyMg
IUvnSEIiJ+4w7bzcJnbAH3K8sSDIewJ1F/3H6e0zaacqqazubCQ4lxUXiAh1MQJsCgJphQDYhAjK
EadWVX9cARz63fR1L1WypVPfMvkz9GyNwJ9FoDw+WZnsvnCCzus2p6v7qAYIxljavJlDhrF8+mCv
ENsDVH6Bv9Y3lnBOsNQs+9J/c+4VW6ybap5zkN5CNo33ZLl0UZ6MULO+kJYv0h2MKwHgobB+Aeix
sFhAi/XJm+eu3otTX2KeUIWebOvli2XY/XHzykHQGW69fIsueOvRi5j6m4DR5Stsj06lhiZC6A7i
7lv7fDqVGik3/ofidsWUrEyJrg946/sPFbgObRK0aUUaVxL5AT0qblT7/9b6Ab7A2gaqRfid17H5
m9S6FXo94FyCG2GRsse0aF/mLXw7FXjgkxLuqAaTdfxYlRLt908I+wOu7+dpbN+BWeQJ0i4eemdj
s/zfmH7j6TQEuSLbmjt8uGYqQ8wAKQfCfYRrX3m7i9gnBwq1Mvg21dpHsZW7ff0ZYajelODKBFPh
erIQC8YjIa5dnE4M/2NBiaoP1Lf6pHgZpO+UDHYy5IZLUMxJa1I+493OFzx014q6eJXLltCE5NA0
xdKcF60Z6pYZrt/IWokFI5Rz8O+CDTCGJ7d2cotIvZZ5ftODrlYTC6fFhyL4N9ueUmQaVGCTD02l
6HW44/zgO5++HP8/Q53mvmZsf6A7M2s8PaK5oXVkFrrK9ZK6ZxAgXsY7vgXy1KneH6W4X3lO+gXm
pjAk+z98GssYG1V/A9BwYOM3BOaIH7TClSsbAaNqxbWplgx1u3PoWD1F/Qg94gyItZdmMuY6NJGr
IhFnVKyNFG4j4r6KeryFo0QWeFIVP8YMWG4L7Es2yct4UMRR3NUbW7WMPnC3m725cmxTdfsIOOKA
QbFU8hHYqS+rsQ/nuiPbbUNnhqxbgpfAuL+gd8qvGPSLkBFX9yUMi2iFW9tmbg/6Mn8M8TvU/JYQ
7D6voGAvNeftF6fLdSMaQrEpg9gv6mWi7SE/1gtCBD61wK0UFhBc7CMQSXWZU7KH4hriVCaRZuD+
BxUeaYibYN6S/eEBej/d2L5N9B+5hWclxwT3yjlhLHfXimw24dGS05d16MXVbGd0NwLqY/FEpW9e
hF/gFnttRoCRC0/iI/mYJs9YTllMwCa5DiEpr/z9AeEkiE0RZkkTSrKoLVIvIG2OxAO8kGJIlybm
FeLHJE4bMGiF1jpiAsc//GOAQnl6w59pssGCKmawgc82o0F7mAcqwqOWbYKpprf3h9asdR/JGkG3
hOBwUXf4AZ8pHdM0+nIb1YskR+TBh8DkPsmX4HbQR9kvspZ65S6erQm3ljIJNIHk3nT0QkWY1A1O
FfAh4hlkxzL/xKzE8qtzlul0YmkSNfRFcgxO0Bcu57fq2HICVP5upYMVtk8RE1RP68uL8Omj+PBP
rglKEpvyM9FgzarQa29mIVlcY1zdcbbpmwAYKw87pzUUAlKeIVtX5D6ZVQbXm1qzyGOQB+waDtdK
EexEHrRTmfBV3j3a2D2TGJUGwmGaGDgGxj0QXV8SbTFe4BAFiIuJ7HlnlWbO8kQpmRgmAACAr9nT
HV5BFVBbV9KnbqQj3weOYaLrjNbxIl6LeeT3V/c1DUlraxEwKm4JUowPlVVZI5viIEcg3jPBwtkk
N2SSgJyW7u2k4o8blfT6AmJ8IjWhyMkYqbl4nck1SMpZBLMzC7JoNKDbNCqcTbEZweaWrxCMEw2g
7CqbMC4IISQAliO/byf89KZ+P5L6XhBjsgAqs1HRBprFUJJtx6tBkSEyqstYRM6Z4JIHucdejwAp
lnpECNkhqHzPFQwisHr7aQwsL4X0qatkgj0hltwkSO7N4xTollcs2p9IudmGVsomi4FN/nKnDj8p
0sj74+Hrqk5R4Ik2xQ93DCjLCdVEXeRu9M4nJwufyCpATCVoyx40l8+v9Hk2omKJDrlC7A6nCRGq
KRAqeBA1JlHvVFJVHyDHQ7vIwz+0kyOdHrS4pMTBCkUF+LXa8gW/nIgW4WU6mq39HjBYTZwTBOBK
pmdAvmPSNP2jy7hUAzKqI4RxdN8TIfdFd4/dAa9ehKTuDCoY1xu1CC84KgVrJGEuXgqpaXWXMDdF
vVRkfw7EoVmVgoU9Wa+bdKXo2jgrXCBMRkJKZaMwe8IB0hHR9dNFoFWkynlrxGq3DFuo5Uyv3I+b
FkFf5yjLCtob+KudggEyMGeX/VgEQHAtFnQD0mPyw99xUe52pUtCoD9XwaoaIjdc0ESUt/PknOZa
XNMzE1jCAV7o8uSfe4YZvxm7z0NOHXFxTqrcAyRicrXf0asM6ae9SQ24F0r4dYBWjdK2PLHgXRI1
f77lDfvRV+kk6C1rlM/famJmTxbCi/YMX1usbnu2JDxBC0c7+reC/QxvMseOTX1fDvALyNxqvjpt
6x+xHdZqPYesYsavkaERhnUiBCxIrwn4rFUZHPfbVoVXWaZSesgMOkY1TQwPwHktp0XgZ0RLYFZU
u2A1ERnP3rfVYKcj2iqL8Y5byuAv7EjxRZLjMVSCC85xbI/+6OgezhpZDxi3f1/ruhLPL2vWx4vr
W5ZQt1SG8JfJDLrmt58FINq3NaTANP2YGYJJlMBxEVt+kW86KuYP55Fzc5OzIQjmuaEedHK8HyVb
kTt7Byc5S4tdiB7Grx+Vhr1wToRlCfy4ThAjbdxzI+C572Xojdwp7ic3nh9wHAeCr+dD69GdYtEO
hlI8NAfYaxi8QTGTnYTMGyqkWIC2kw8F6VCBAentNEtiUvsoVOO03TJybMrlrSxuVikBxrH7ZZh8
OkNleAjQeQJx1c9Chq2v5g74uYIFy7SKb8DCdgCD3wODPz8f2PErHTD/NZREPZMofJcCRkt5vZVU
qwOH2REkgvx7ZGxHdlQib+A3ep8VCi9EkcVmK0EQTQnSfX0tNmFWdIbysUy2mT7casyxTYGgoBxO
frUF1z5o3RewnZfoKFShFagIC6IpmIbo4z4t74lT7bjNRBbvLgAu/MV8iQCnPX8XxFq0Vy1YitP5
QLJFYzzriu5mA85EMcXrjrmAKU2OobftwqlnDGkwicDybT4tYQ1Gpyw0eGVRQUj55X3EMYyB9t5i
XXJyFEPCfd+k2jTdN+sjtngJZ5AEz44eNFou+6eCtnEe5RGmQRd7cKws4J1/1RgjqK9/8yOYLTSX
jp0xsn42oB3Dva4e+Oqvl5CRlN4D8HEtc0ALJRCPM6uHeCo+HZT5AN12khqHqaI/VPeDzy9TTqoI
DrxZsag5AbxFXmnVaU+++D7M+UW7CFGrkppFr7j7eMbHqlMcwprBPsqlUwyTW/Sgg8p2b/p3J4kp
YQmXOjSe2Bg95vgIfu/H2hKrNLY8AnzjetmxhNmQBZY13IHqyPTux21r1tCRsB42La5eLBw7XKRQ
EVtfws0dod//WznzHJoPJ2px//uIjb8FpX1P5KaUCD+uAkucqbzCV84m4mAPGctLsF1VyN/u4GaZ
NVpMV62RXOebJnH992Vw7RoCrwXHlvmibfcDCWO7WN+3F9/vgfheoHvbKBl/5yaXyW5ZvIFMoNNz
ANkeXDOOtXNRF9Uf7vVAOvszjP0KiYc69dcPm5GcEcXzKg1IBdBwMqpxlhKW/nZZ4X2cvm7TkIg+
kIc65+LrnUgDcLBJDOZlem589mv+AVP06D5Mekk/XBy3q0xYxswz0PctfAHQuii1CyJuRN6O7txa
DDklptGWxjO3QsYDOAHdUrQK0r9mqcrSm5y8G0YpVavC/IpM2LN/6dnzXeOmWNYkFqHxmL5ozSr7
oEaFmHSjawT9COmOlGPSernn+wTSdGYLcvM7h+h4r4Rbzj7LAZg2l7TYgXEvvhASf1WHfqbKxpDE
3b23x79acfflaN9rZ+IeNfiTKaVxMR7BX3mt5+Z5Vxu28ZwVfwgN15ql65BYuG9VMIa67yacNWYh
phXlmfwfh0RHqkGsRGxEd926qGDlEFvTGKdCS6uBN06KHNc2iNAHcdeQT6HNypfjGkkStl9MnddE
DzHtfm4zmjlyp+lGBMwPGP1Lo+CicMVdXLKp10CaZKYKlMPk/tmGDXp7dGl/tcwjK+20E/AVcjfN
WOqSdeqPdQea05uQ8NMu+ol2BFeEnevWAAaqs0A0A9d1SAPIC2kltSaUcUSCU5+rJzfIRhtD6RCJ
kCkatNUSvViAgI+/Phr2ETo7uZj4Vw/RtsSz7VZ+e0OJQ7pynR943YxFH+9DEBx5j+DVjEfgBKYC
4NJ8iGuQeFdwxJWyhDlyc7Un1kdY1IPNqxTmNyEv280GzuP/11G6IixPzIQBuP0bMmodAdPH7upG
iFRfnHRKUCCnW+FSI2pc0kKg+Fs6eyUxmGIKIzTuJK3u/4LX/DcdAl/bQFpH10yxQ7zLDJowPSFQ
1ph06gpn2HBmbFyQG0nT1q0J7LfCKLyRw2R/eXT2KSWgQtqAMV4aTtXZDiHy/8XXvfWjuKxEj9V/
RbJCva6Jezo3jECnxKegqyD7aU8TqYJEpJEsLtUrf3I0goHK48IYHEE/wrHgoPHAGfJO5Fj+bxka
CPaQ3c4mFlGP147YXA2/iWRu4316p+rsR12/7pmbuoAEWBe1mIKH2L62DwpopoTyPZSWZVqL4q7t
8jS8mORddVN0oD0weRCdcN1wK03p+JQui+JXgU+SZ38F66Zo54qAfPeY5B3hQocbG5/A/cVOQqxR
gDMVWBF3y/r4bPwsVPIbjYk3RWmIeRMUXrCEpoQDMW4bSiju6SEbMdrfXvc3BAFmsKIOoMBVHP8g
K7djRsH3U0qoNaEiI0VWOE0FxuokNIjQfb5k+W9NPoNHO4JecdSr+EkVG1YTp4hjkO2W4aMxiFD8
CRDpnaxC3Bgev4A4dK7fWKiYMF0mKC/uuxah+AEsCh1tDrIP6wuAcORdUjQ3v+216gD0qfeb0Eu5
7Su4NuwbJBLKX5HhGtnbAmU/FSBAuh6OyqQRUYMw9oVlZdVBozub/88ZhTHcCGA9rhBukJB8ufBX
oEUMp6rPn69Y0dy//lOtmG+sgfM6F1rD3hm66GH6Ny8d0Z0iqZMnKWFoc//uXI/v3uyM3ZyUvRCf
orqTG31/kukChRzddoL7gM/azJ3RjiV5LsUmOmWvZ2H/PjWVGJ3ts2oryL+LrHapl10rsLfYYIuc
Uxp6r1VvkU7ZlwZ8qaoJARSsZd4TXwPwKQ36fs1C5fnPNvl275/1pE0V3WqDvyXRguGiCiflJAi2
7N6h1ln/FuFjH2a/u6wLt06lWe/fE/gcGxkZ+XKJwwWyBrT4A0CQ19mLdZwvmOhZj24uPISL81x5
k0yKKfAxC2zNJkmLThKRe7GRtrQymF5aCPvJ/BCrB/N4nQ9XHwr4reE2jWHjhAQyzoMwqh0QMQjH
+ZAOGWbrTryg1C21BQWwkuMm1b8cv8/CBmQByvsGz2FIFbxpFEbmGndykXVu27c1NASqZdN5zTN8
TNpiZTuqMTyc/dSolvOz3riLj0gtmlY39eY7gJu+NF/tgdlO3t9tJxE5B3Gwpk4wTUtWCFbJ+14A
QVyePT17bXR4F++w7HgJ4wV/T3ismCjDtrADK8ApPbgKqyD5uqnctyi5Un+fQ2elvJxm3vj/wmns
gBQhPljruU+3ONqm30sQb8l8+t05MhZtOaQyY2gfmyxpP7XjSpf9Z/E/EmLfty9HWv5lJeiV1urB
o4zp5lQeBZRlrwIhtLAeGsX2EF95gkzu3TWObRYp5uDW61q9I34BHmzCWzfV8YGN9CnU3Ab44Ouz
4iJ0R6mp7+xKH0qzgtoVQrKcZaGRLBZ9/dp4yhS07iiKGd4Ode8syO8/ErtwqbBkVn0qS3qlrsGv
pk/FrWNAGU7iQhgoFXdXK7+jFqriWxWvq4fKRXRqI+Dw6/GDne+5Q6TKbYGFpUCwNG3SqWt0F982
96XgnjrDDRrLeES/BZzrmovCtLuZkrY+XoDKXi1h/d2FBscZQ9BoD5gpz4eivv9iC2Da4/hrtwvL
T9oMWPrtSGadcWYiULbHVnEV2sekoO+hshyfnqJUAlF0bF49VBU/JoOZr6YSkpN/TT+zkm1aVcvr
FOMuxKaT7m9YYBPJ7s1FDDfTuAR+XIiyU42kSsCFiJ8KVtqZUg1TGMdg/RlobTpvKY+AlBAz+Ouw
FQ+Gc65yhqgqA2K5JBLz1neonjU8QlPx2L9EP+XTK4hQsLJJdEFmOQPDuRTcSSAe55zzEmkdNSBH
A//YpJceHr5/g5EUw7xj3861SCIv9+xMcquN38BHSpuBtoeF0PR5f23JSZ2kIlPudB8XdBC0ZndH
CM90b9mLz1srSEBOrb9rxG/XDC/bAZyA+ibxzL+Q5fNY/+5OBBK1i5fbDqZQ9ZpVJQb3bx2+7Tes
Dxx3Z+xLzDvGaNvkJI64+x3Kq+6d5J/rgeLyzLHJ+s1d9rnnsZ5ijhmj3pf1B3bXHeLrgeacrtzi
3iE8DCT7r+asbdIofQwRvMWOQ1MnvWhhy3Dg3GEfkCYRLLkG6Wky7YE5OevYZ675EO/JqZt9t0CP
/PXixv4lkritG87Fq7U5qC6Vrd9Vx+2axnTepGO58wt6QjMc7TD+9b9hBv5f2DVL3OygaAk93bgo
QA2IcTLpWmiU2BN7P8/9FgqYNg8MWq8gMrZwkqUG4QsvDrHY7yrjrtqXRmjZYWxVcACtoUWMzM3x
tHejrLfyxr+i6nugtj1W7yu0hIsNxKJAb5aoPiibA2c9FzdfjwtOhFtGQElivrMQQTEtiu8YE+NG
rhIy99jYaarc/z2cJ++/x4nFb0i/9f1+ixMNNQYRKRJ/sh0db/I2/asjbyJ/32KDHpc/W/93OIha
+RvYtdN/1Z3oY7xn/fh+tobL2nGjuldSIZKFQH4CkvXMyTk0Nzx2SlrKjGlArxnFtXoEqOc+h8DG
ihE0vlO+ixLLsFEAsZ205fkWl461apX6xSuuUBNEgNxLcOsReXpwxmyCxjtjMKtO6dpBJEPvMP9o
Kgw/Tf4dDBqTJ7hJrN+xMmv3tVUH5RWohDbuHVFByX1VArP3/yyJaUrDo5cH2lQk7gNF6UEVs6d+
U8NJQr6WIKnnO9LRKqPDTLsri6r5kbpDvqk4fMcBxaVk1Wqn7ihAO0223cyGwOecrqdo4IjGUIqs
B4FL2Y0CIX1xmjThYFPGXebvuMYTk67KY7xmr0vqIi9rpL34rV0vV9mi4/2PvRSwppgdO+nReoXI
ZDGZauxuZE5MtG9YJaYSj/pQXiLzOEPb8gSszoIHxlfrARGP7dW9uuwPHQrivI49AtSMXsRBSTnX
9bifInRyxb5RBf9+8y9eqnTF9oEJWUTRf/8LwOq5j/yPpNttHqa3xcdUeKwev4/lTVJXGzhBttyr
hksP4ECkRGmH8X6Bo2mmMzgtzcqUo56l7OtSaunvJkLTMARYKrRmjknvgZGqKvO8CeyOOexW4xPX
RSzpfbiEkTjhhsCbLHdIS63dYeoe7vj8S3s1Xjnhoq//Oujwj/y40NaVknPv5RO2FS1KXSqglvUo
55Lg51q537vG5bjyEcmiOUs26y2GxwX3LQg4iIcuLhqM4I6G2h5Vqjh0IQbyE4Guxo5OZqah57dA
npKZCrc/6RbBHoQGQ/X+FR/Aqdoj0+hNmrKcue46AJQ7fujgpOodPo6Duli2HYaQXgrST7c1P36j
vkD5zsN2BxRm/pl5GAo5YifLd1rr8QSb0vguPPA2hs4FGmngVC3oYpMkrrMFY3zpHLlfwn5jfmpm
f2BSMr0vqYccgMRdoRCmABUfvIeD0qLfqzVegeV+un+AAxCggp/rBDcvCbjYuHkAE0II7pFakYt6
jqUOshdu4v5w4N2+UmehxvhAcI5kXzDnxQ6MiddnYvHi9qfnqJHyczrAJi82oTryJD/vYW41X79l
wc29FJHyuwZJXwn846AtRQOA9s6XAtn/SwoAb5jQeMpSx0MP6SRzLqXQ0BlhWZxlKCkKxsud2sRE
R1fRY0WCArT63Y2oYS39zEJb2Mc0pz21Xz5TXWw92pJLak2cX6VMkzVQqxTJagXTMohSq87qUxSi
WfNODXB3UXSxMXigo0k1O9FRmuXAdANRX4FOFkuQmmQiaEunVOHZ9dkjzdPXBdaaDUiWCzNNBxBm
XgeRowh6X3QtDRP1otvMlQ3yt+uYzV8deWofRow9844cu2mB4L84o54n2Huk+xZ8TOW4rlYZgQD+
utqGPCpR1Xoap5KSUXozqQnIstaSa8v3WVFYJ+za3MV6VxDEEWOP6HeCEpNUbN+ZzrjvI+2p8POZ
VfuOeDrsYm7fRdEwYyaWajg2U0u0CBLoTpCNfHL31o2d+L2Gk2Pjbcf4JVVr2tsD45cd5Ij6HsaJ
eSiEXCSy1CPlm/Yz1v8FeCN6vzDlHfzhwIMKz1st8fAlxlyGzYPEZCSJ2V36PoISDoV34LP1nxVm
u/+fcKqi9FqudODD/wzwqka4qPO5VMC0sMVVxyarkS/3ZbFgCQh1RkbdL31U/j3HaLt+p3mxFx+t
I+oF+sUCFr76zoLZfPYk4XMQyfVHmjeMUOnoUjDqIdRaeeZdJi6dpj4Q6D4jQu9DC5MVjS07WoEw
qRsGHdPNQeQNnxwhELmnq/jFtjcuWmNcfXXTHTrnrX2UY/sxhbun27KdCkoXV1iNksKAdvoEmuIW
ZAnL/Pe/7ov+4tOODgkNQIKN5/hw7kz+JKp0cAIuXPjW06O1fqvk+56bWf3wJjcsvQlRpGFU1I7r
HRNa0MdzKqEME4fNtpoXrJl0CWOI/CeY4uYSco1NmvY7c4+ppahdvY0MqVNENMXMotSr+luBb4VP
3UPcoThCyO2i57INjXq+A2BxYkbFgwLiDQgaPrl8/gkvwe0GNtWJwE3VsT4vVEJWzz+Ux9lj1tmz
nl8yUhJXkRktxaApZG/CXoBJZgjXLkz9mgUBsLI6LpqsTXmhn3HSUTCL7XM2IsooHXpmiFz7h/zO
aPtOW+/IgnDG89leYrl4IUWrLGOXDd2+67hAiRqho4iwccacHuwMQNIbULJEp5OUg8QG/2irlh3z
z7yfhNmskgP2TfqGVkxbkjwNXvVriD1qb+axceDv+dm3R+CnJ7tCNyKXjew2YTxVyueHHlfHzg0k
0SPpMgvwhLfljgVVHiSRGGQWH1+mVTVxR7+p0jl6qZ1boD3GXPC6zd7DfB1nWXzn+WbL0mxjEpVs
NLSr+oX25prragH8deV8GMUwjJIKgRIXXDtMDG83z9E8m2Mss3y3setOqVXWjfntQ7gfOtoUMrw1
eukWpsYhZ0YcrJ59Aysuc3inY5pUiRdoJG7e5Hu1OncP37C2vkqRqjGbukgEIEsPqMe8Kya9TcpI
KMkoHAwbFoYXp4n7kJK9q8tThSPGQN9OhxosDD6A2dSDoB5zkqP1a+F/axZEn8+gEmhIgU9/WU15
5lwFemAyErcD0xtuMfUj1Z5CmHAOSBwwT2Atn5v2LIGgwioYbJRfASfyRNy66MdOLpSl5K7pWb8w
lamDbter3A6ReYPTK3zJSMzmf3DZxspCYIz2zOKJwh0FEhet4NBiB3m3xerujHNZPqvNzASugrHG
8l7ueh1OracZibkYkd80YlktzrGMzNIj8Ron8po1IAMS/Xss2VOw5uu94FxGq3QLGRrGW6efWiKO
tlICAaCCMoafjeTe6ca4tdNruNxpV+qXpXcbWqlSJWUWWskP5i57Pyi9yCK8uHOQ0v1pkweFNq4h
OpezspSneCzCoISGvKH0KEgIEqLTpmT7/8+D2eFyPlV/WaQC/m/NrDbh1X05re5ZWkprOCCnYnN6
J7TMO0diq9qEDOT5bCp9TMEfDpB9RjInAqZDSZcuzpivRalmF+t7zQjqNaIgbS2oy88Nvu5F8LKH
ytuezJbkUkuN4FRAENT29UaBcO+y+FiZBOKSFvohkm9W4Ibpbrpl5vhczN/Ljh7msh6tlZE+Zk5a
JJp3w0b3OYFLzitL5oaBDCL7O4YOKbXhAt7qfel8F8qjnTMZvuvi+P93CAIoqXDAXatwWWdzjAIP
2WiAt8tYl0ikpg6uMXZTOLRAAM4wdJZAtxO1BnSrOT3rKpL2qqaBNz5sS8spZd2H+GuhxaxKxjFv
T1wZ/S4a2Jni/Kme2soH5Z1zQUkx5eBKeyejw72U6GdRbSOKHMyMFTZnx6aG9NUuCSZMJriVH+4n
55sMwy5nj2rEQO3462UYiwfkaBJXYvWsreLgU2YN+HPJTTX0JtwvjNVIjJtqxTB/pe6+TWacU7XT
k68YBhGv/+ccwN+38yr3zKidD/LTWMbwFaL+PjBgYBJCeURjEdrpIl/79qlMS66xJ5iHvyKjbd0b
lvdZUVxqG0IrgKoJRtOiPZzoZfxZgsoDwNik3hMcx+UsGvwSUJ1rDNKxtKwyyZceU17xkk+TNVyJ
Ch+bbiOgxDnF/HFK1niTvd9nIFITkL+g0zh+/FLDg+HyBAxJ1JKXKd5XKWmgm2pFn3+rxM2rAJ5z
ohj4k+9QGoODjjpy4DO//zW8vErrMmgmostNNG+NbVjflRp4ev0uSvSvdQY1Y3wWiSqFcW5A5jxJ
jG4wRtev/KF6YzIYP0SlzTWYDlqAXVduKiDLfYctZQcmA/1/Efp0Z9JCp6GAjPjk8k5JztNxT8O7
7K9B+krliLW1ueVESRWrEAJYFF92PRs4Dg2ssyKiQxedRRoLWIK3X/aXQ5ivMTyyC20JsLfT4L5b
DXzC/sxfKHjoUO7irBhhQ5WmulxrDS64l//wj8QIJ5BXGK0rwmxZQweI3JzYBaFBnrx0HGw1LG+4
g2SG/nwMG87zEp7rwYBhD3/vRNs/teCV2zOIFgiB3VT+kp/VNArGL+EtXaXRqoSdaqjlU7OUkJGS
/jgxmwkNpIgH8zK8qhAkJ8QEFl9pFAe9wm2eYnUhMl8TFgJVwndsuzcRuDJeQEcTVNOwsjD89MeZ
tb1L4iDrf8b33QYJnhquXI6ipfnJf+3045A+8YUcxZ8shVkCOaiBzCcwPEZjPa0Ss6k20df5mXbR
v9FhOFqrdAZwtRzVvzEumYNwwfjXBWAzElhjqRf1iN6fgQA+k6CfKwjPbH6WNje4SjF0pJ38a2Ss
G13CH9Ib03v4kp7e9sYGUo3FK+A16R4ag9+KcFdBUaUOs1VlGdPB05/u8otdyr/ThZSFmwCSuR4w
01YkCrdRG24+AMSIayl4Y+6VDziSA7eayBBSYqBWKdM1j5o4P2mEmgQyDM+KvZDB9CI/dgUTOUjN
zIgGpjnG3Zykjo9KGYmH34Jipp0oEeoF7aF7QXQmNHRE/7w1TBSlsaXp/HyKAZX88oQdBbGy2r/f
I0w0rPNnwqF2MtSx2wl5XeLbc95/puWxx1NPGrIX/yaS8skWdFKsvzVXHA2LT9cDQtjyfyAb0ckC
QRNpimA6CYXE7iMVaaQgZGS0S8UEjN/TlshtxQdMYp0/LKPNa7W6RHxUm6Wn6en2sI/0mF4KsVCz
6O6jDq/KZL8w3SGjMZRHuiXzhw6CZeIhs/hwv0ktdl/W/uPKD01s09KTDiqLDs2BryeqFO8XIAP1
vD0EHK4jKj0ya+lJ/yWl7lGUTuKkd0suRmkREdj+AtkKS5QN1ynAVD24bR+/S28FkVtJWfXb+f9n
f5AMFYvkuZvX4YIwJQL6IFmVpbTmQzIIYXkLMa5uUArlMHnmIeSLYHDhzgWfDbN12zWNjC33QJL8
9dusUk1fQhskM9ZpeUSWK8PiGidH2DjsXQk7pO1+SQUxb4VWGcqa4BQis/0kkrCsAShHgH48+GN9
+MtpelK7Ui1ARnViG7QNDhfx4RYBJH3SalJ9AdUbZO33PY43h0lklHL4+4QZf57ooNwtW6j2554i
DDUZbiEvk1YkCRa4M+qcMSfjd6QikBpZHbQYOmPNy00AjQqwRGk2Sebxqp2XaqrZa5fMKfJ8XL3g
Q4QAoNwoBpGd5zqAM1fMJIIYFpGpDJegjmwWrRGQd/pyRYWeRtrOtlF5snJPiiRKv2L7e+jQDeA2
QUZsUX/kh86IycoqwbPckK3Uh7J3QfDtFn4NbRQu/iEc0g4kjFzgiN13U2oAKNm2sa5QDO8wqFE8
qobhfGl7+781WEityc2zS+DX1VB3RETrX42MdcmzEiFK6RMh6WECjSreQU6iO607lH4BMEr2Z/30
Ud1d4Ku9HBqIP4nXSIw7ZPaCzfbsiltNWOtMdCNBTrubUxkUIu1DQlOCtrrB8cU2fgvAWRl56A0P
rH2A/KCMa4LyeenYK4lA/hfP4/lEeY7iIH8itRaEMmr/r3pOcwFqxxKuOvo/hcKScbqpIhgLHcjP
6o1FJAKmHlJ7RxdZFqf5jUMV06vxzQInDsGrDHuYokVhLR+rD8AJDv9YqmKrlFFvjt44C2B/3dVH
He/7QKE4OvtaTwNqc5y/h6BfZLKY1byl+jgVIPV2beqbZLmUn1BdzbAtxVxLuO06/L2TLs6l7rYZ
7wMKdeWt039tEyd+gE7MGhTRLL5HFjOLiB6v5GylKgubdc3OY9oyarM3z4iSTdcHz/R2/Sku5zc+
CGIes1SaIj2AxHQjS0eaNeod3IW+yfUDSETVOOXuG1OayPC5bD+a3Mx2DB+GKOZ9oSKMyBSLX2OX
uBOHjTYpWb4DkuJ/ErIDMcqBh+jrtZrN/s4BHs8W+iXc/IP4mdwr3ygLjehWDv+pTZgkcpbv7ICp
iC3O8+9x2XSi6HR+GHAJQeQ92CCNeOLDx79nZyPBj3ex+hZ51OboAJpOgGfrsTAWD40c9oi/YT6e
WnIlTWXjXFVCUpaN5PE34p8QqqfquyO2YI65s6GGrKl5inne8Vq0GbyKOrn2AU+nhP+cK7EgJZ6x
q+yjSHqMpKE7a90djbA/PyEqiT/S/FmXESybfsfC211EbNxBAZXnzzGSygPIE3dHThWOzCrn2chS
qpCG+0Y4TC3W8LNZw/+/Japfaa8ZhJuvc9ZAaXrId3rjEmKVuUc95S1zgfnuMypbLPrCwQq3W5Ap
1hF3vEZiaL//ffwSfjQHiUKIcQaMAyfi1N5P/OgrNPjo53xR6Rp4rz+JuXzyB685rhtBRpWRCqG6
7E/SsqjHH4QMPLPBJi6zz6IFsAqZ2xwFdpmLV63oRBfznNwpeFM9jf6KPGajGzDTOMc0gQvuHGx4
O52ByWxbN5mgTToYr5FCKKFV+x4ZVatMqj78Ix3H/4fhvydyKOGDzW4W2tNy2Z8caaNXdEQm0XAr
BB6KtN74I6PMAnzSToOnYEoJmbX4Z27zCeatanC28qv3yfQ7IJongzAe2RdOtJYvaCHm2nAiSfFS
6+1gHpMi5/YQ7YQmX7/DhSa4Yer7VkaEuEpoOq7tTWdAew0YJ8SVDrbFKmiQt9THEtVNYCsfr7KF
kUvZjg1EhBmjVpd7N0BwAAMfSeP1tzbKqZHZq6LsmixxFENbQNFFUFMgCb8I2N3KlnJRhDpypDTP
Xh3trnsNrqkdQEffEjoyQOSddSnjpBdkWQ3Dek4jIbm5s/zg09C5hKJWNPotxcZ3gSdE+1cQPfPD
lYw4LU4NhbiCKK5kvNhZMR9FIuYFcPiSAXNRqqv4w2FYI0vagkTQj6hofQReDI6nQnYRUrb+lc07
yz7M8a2bqK1PG0byzqnbx9Rl4Df1g2spn+1w8wCHhGbaplRBuh1BnKkA1GMHvOCFk1+/VfT+83GH
zjDa49TCTKIAwaelE+uqf+WPoh/yoXnin/bGkHL5GeDYBDnIZyDJATE8EUqqyYeLV1xwMTeHf9pQ
phaKiuA9o4OhTBZWhTgTpUKuRcncNIgr4vgelJoo5raUqpGSQUrGNW/eJynKbBQAYwlITd5MKj3m
qvmd1QJx+sZBMn71eCx3Crk7AVMqc3saKSYVIQX2awdDmcBo1eG/beRLrF71o/fdEY4ioVHOwg+9
SrN1kY6zd/Ek0y9oH1DGEnZ0PQD+x+hZnrWoS4xsRyW3bNiozxFF6pEWVJeY2VGLOQbqsNCyxwMz
gNdxi5xfINzPeajz/iCwJZHpfJhlPwem7+B8UbIrSiPBCrMLY5vhbWb1rfCoVSQCbfhw8ZXg9RWq
dEjdLLAu3SlVj9xT0GqV22yGntvlQshUmB1Dnuruc/rNNEf3mtMtopbEUiuFKpZ2PXGPjWqKGvtI
uvQwEejKSWG1DvWNYi1OEW5jUbWzk4bSQNaXUJuBAIIlWLnSbtRxZpoxZMu/3vmghf2rUKZwrt43
Y7obG1tOtWz8jVeB0eCctVSjF4jLtyIHF3s0n7bJA5xz3ZfQqmVMiEDoacqeLOm9lyCwcWh1dWm9
EymMxTjMmr2f8qqY5/1U9rB94ApSP+wwEoaLmss6FkZ5z8oQQDe0Ew8FfKrJ+w//DTim01tMavPL
JQVFRKz0nJSh5ODKRFbgmPu8FkOxzCATihUqusAAgbncL3UCiAzCRv6NY/0OoLn5N5oMUPkOh5pY
sBT1CA9bbxtXjr0JwzZnFeQ88cevsllgdm6ziiUdeK3kOsqaJ97zDEGILqG45bQeDqgi9BCNhl9h
5OR8lzbsQc/VRPBDixxeT7BVPGQNAbBOnChpaEhdFA219/vjIpZVfMTSDktQ0V/5KX3/RTpuWqYv
XWnMZD359vxYGyuZDY4Jb2vNdisX5OZ2YKN65uR4zhUjImzpNtp9XdepAyEyl2q1ka0dPNYNz7TU
yyeC8iG8vmNM4Zklms3tnwT2Gl5CiDVHETgwXJpiB9cgAyWx3L50vK24Lp3c3kxohhOkGAWbof7u
Rz4l1uGcwILjAR4LnoYAXbYnzM24mJrPOpHdBEGY5ZAuxRNrS3uAyXKDoYg4KGZ/iuECy5j269VH
0r6vqxEMq7Wk/fenbANKIdaIzmlf8yVs9L2W9xIZ2DXDCbnNiZDPcL9czA6OAjdLjDQb7BRbEYGD
EnGvkKosFrBepnu/KcmijK+9QRMLwfAmTIN32uhpokDEkZzW3wjt7OxH5XUJnEUycv0QWLEPXjju
QDe8EqvBg/CtN98II7JsZAMUIwp3F0t4sTDGiN6S4WaXIluqfpsSN7y594MCDVJXl2MpCzCIjy2s
ZzBOscbFzfbYivcuSTk72e9kRtGWSqUESL62NlNDp638a5yDROltpk+yD7jAx4KEofVBNaMsdnwd
ojspvJbtUo+71SpvOYNRp6YQ2zcmjT/g1RfegyHEYw78qNEI/gZgpCECix0YUa7wGpSrbtIEBUH1
agapvEcaQjvBv8rL7xGNgn/3tJU4XRIVoCIUKRZqFDUqxDn127oHm4tYpRbVoARXaIeRqoJDVrRT
euwoEXP+tzX5Qypf5nlpjby8Xjk3bnbqVSHlg7/NNrgPZGtCFfv1YitES0ViOLXe4MzobI34j1xU
aYZE+PwAnC9u92uc5Oqg4O0oTRpbQVK2UyNbx++Wc+aaNJXBJTrwizTaWfvU0NLdWGdGzly6OLpF
MUmRiJz8uw5PslzYj5vQaKgU7n9sbDPsIo25gkwPIFe5ou2a0SaMiNUxWvfHNMeqiWp7SFR+BDbr
3E2IXrwW4NFzTaFGwyYsHcaHVeoOPEJ6BYqOG+Tr8CcxRhRAMQZ3LbhDf7CZTJ6qAkYVmVmjkqvV
VSip2RuDEYmNf8HjH4Q+otlQtmyS6bvMMqPwZoc+mzDn5xmP/NZpydKl4mJcb6LZqFRrsnyEcZH3
m0g5O8ouirDgDhkMu6W2Q7zf/Dhk2y25P2ZPBvdHjDD7a/Nh7hQD1xxJlpkRP9rAjEKypQYPh91j
RyfqkH4+kaSILaHY+pXxIzi1uHiNWFp8iqDtrtQm9EdYwzWI4SJP7uA9zYt2Cz4J9TLmo6IJq4+v
YL/K6oTzq7EO1QCsTulElEhNbUkR1Z0+lecQhUKGQ2kIGP+cXN5smEk0uX1whWSHveh8WfnU/6Ft
SBEnGCkDaxvQaRCUxG3PgsG/kl7d0JDpwS6J/Qsr50wyehvC/XeXzxQScASXSf6JncMJqdo/Q/vh
EJhUW0cz+HfE8/7xtTvBQVdTtg1m9n4PKVrqblHZ+pqILM5wjmoIPRRqAEWpjcFDyH0ZWpo7gGwC
sgIA0D4cVLM64GurYFsgH/Nz+tF4TTVQaDnqOI2SAer5KxbYQbGNEBPNxDcdoKR3+bthqn8BjDcb
IE0qNtkJDTMwi9f7G8rV92FNnGDkE48tDOD+KdHkIT7uGxFjGf3IBmEzFL34X8Q27o6D5kEw1HaH
9PdzMR0zVKFWG+Z0b5A6wmKFF2aCHFsbcsEXWli/Fl0/TR0APZsdmW6Ipt2h24AKDnbQeiTmJQ0F
7hYsp27/OGn/oirUn/eu0WkpN9QHWCjUY13H562FqDnpkuAQkzON43XtuBICr/ntAM0T7X2GNBWq
WDSApBhUFX209/AhQ2/hE0rU8F8VUWg1G+Kk3Z17WUUARbjmjrLlnh5T3GDHECKzROR99PWT5ukC
XSFb8o+O40DnEhp/WUzPUoaBve7LmFUC10S46qlnu4BqFSYxrVIMqF5a9dIBUgxqK8zBBm6WBMnL
o5/IRavw49RElP7a6WcMg6GYxC0TiKMNeT1XvzLrdELrEZqHIlp7KXsLNIirfShMMDHs+rmKPxgK
sdaSBQ8M85D5bGSu0CIJVJyUqCN81Dnmv0jLz+bOC3InWdKDHr3FkekgPRbRkoHw0N6rGIBp/gG6
r2tvlPso6t3zU04i77NAsJhAGEmfuv4sA4n+hSYWUdxXkde3rWPMoqTffjYvc1KrUhaGkz2wAk72
ljpw3HhKkJy109zTgY9rJwc146bEl4LIWoFqKjFxx2sO7DiO5wmevJIa8g6PIPT5CvdcWtMDeb8w
0xc93+RU/wNcay+0bpqzVe/jJmJ5QbicFSCFDCJjJlIq6giAuqy2TheoFiXKfFKQvg4IYBIneFhD
mRlRfqrbn2mHmH+etQ4TWlAFrYCjkFpJjf5UJ35oZij7bwhaX4OiOgjNbLmEzs86S0/2YAtJCEhw
yliDuBNl34JSeEqhhYRKaWF8k70uigLZDFyTcjSrtNSSIeKO02IPxQrX/1VejMHO8BiVGNPt6QPZ
XQZYObV/GvrC1XfS0DbnZnIYc2jHs6uPWsuMGTKot0cbcdzFIPhDoS4L30K3OZJkouRJ7RQHbJuv
EK82Y2cnxVXbF3NPgzjj7vBFE9apJ5DKKgGPvck6WTCFW90GymXj8h7hxswyg3jBsDiV+ujcetnZ
dTljLSIvXXGuncEuMTJg+uaEECKy/LSdyvBE/wgR+6Ch+g4dGJTOqrWe7G3u+EvoLazpFQAE4C/h
wZEW7l381BWc3s8YRcvv9Dv1BCMaLN5EUU3ciUbCbtw7sx7gQ7x9awbGRTS4zhaHBOkN20cVOvbr
8gNXyaGB8UCpIZW66BaYWrp+r86Iu5H4WR/RC8n5c+TRtec/0LvnLNvgVGjL5Evanfsv1iP+ytfB
K3l/fqmLY8Qu2Ir1Y9H2Af5VZ1x9mmUfOwrr5eYhKbZxl3pSrp2FJ7l7sB4OSKEQUdwrowEt3JfG
kTHL631UsD/wYSBHfOlXnZufhmbB4K7FUpKKjGN9R/aWWvQsOnBR9quezNNpdk1jbh7ytQ2hUhhW
VNBwKyO5hCUdTI8nLDJCvHrR9+CeBtCFtxXMbmn+SAQS4W383o8brCTTdpLIpqx9DOvRlzEf9FnY
iYOboiItyOykBJmo2JJrHXgWNsAlhxqyjNM9y3yFgx2pt3OPiPgIUOfAdxpDGpteGbvdiGUtRMO1
9MhZUJOdERix8yIM8biIe/86DC3GUVgBm66RYMtwuHBZsnwjQJrg9I1K9F9c4E62iOc0kyVEvt4L
Xl/cQOb+HULVc3yOc9kxKvlCumxsz7EP9JW2WYDV0DcnEM7x4xMYWlj/hRLnL3PzevRfiWTdmmjg
IpoxGlaryFgaFHaoQNv6tzuVucwmBjHsjSExZDAq+YpI6lgeE2Lurbl97TEM23gO6FEOA7k7ZF4V
CFO7+EQNRyNdwZs/3FdtompM5k/y2IVRNkUW3n4TBCJLt5dnvBdbH7KBKY1MjUGMfWBosnYvLFeq
u6U+XirpvVXLMew3P9OvFxnQgfSC4JLhJkE0ikiKaSWWMLreMqREKUqrGhpGBYIujZdBFEtuzjuM
q2AsQSNY1U3Cb/Z77RXvfv0uDeeDpKYIJGXb9jzbH7DJiPcno0CLEO1RAHR6PqPH7msfeX0E6jHu
Vhxb69HFbbYYPnHYsLvUfVaYeR0IuO7d+lkCTDw1eddF+Et+thUBJsRrJ5lD/SabNcXi9tNAhuNt
6lrQLqx9ns2nqtG5sjUAVHsVWFqHtSh9EeKGvW1txo2hJsaBxQlmTq8ymNbDquerk4sOHyDpYkn9
Cnncx3Y0LL62+fUcd3blQPdAZTnKnNg2hkgOaxExzTg2SuC9N41rPUDSq9tV8a95Xdza8HYZTHZs
p1HzxCGvX3S/9cK+yCW3SSgByIB/3YjEmQEtI8NTQb/h8EjHqfIXnUaDAhQMsoXRHZqsnZk7CtCw
MDx2pFjW3RVUCBVVFX2EBkoeTorfi7yGC/qJ0QxWZVDY3i3kfAF+X87yQ236Ij4MP7oGvzcXQsKM
jYj1pUjMfDPLooJE1lmQgyBHiemfiRbSg/7zqpp8X3pVt1k2nTZcOeBrMjip9+Q3FkEMzP1BEDOU
sEI/LOwj6uc9dq4tp4v84oZj5t8ETw+yNDoRSyPMTUv9eMypVynXk5K54/toxXTExU15gnD0bIEJ
/rkboc8P9lIbsPidp+sRx/l/ZSKoCt0EFhVQINm0vIMfQIQwQ44hVSPGvaI0s2M+LiJOOxyOlcUD
ZYb1rEznNLnI30jtx8FoT9g23rQmsB63gsgQk5TnJMajaygV7y6o493pZIaT2P3fOTm5SC8ZwgJG
uKmZwUso/PM431si5TfaPPhQ/5LHND0fkEGEe+Ke5CtBuxQa7Vk+sK2Yw8pTb/fH8eI5UDi7HDQn
UkT22QmKdY1DpN3ZrxWTdEH6Qy/KhXGCwhDHH1TUsq5yCCVZz0fPsaSU4juQk2W94ZhdpYjMV/Uk
FKUxYA4K0kv8AyV/DaXSOuq5l3+kzTWip3WoXu2kpWJLTgm9vWfitxmDLwjFqJEHrrJdY2aEREop
BA3iYCkCUYpJTUtj35iZllAnyNKEFjO9+totJPexBbxdjcMNkp2R8BBXnLjkc/BlaiSg7DlvyC+H
ztLEGzrzFjg0cUDO2PU3jYtm7t1CHudQ1z4SACy4T/WydR25fFVohccjQm/tT4io/kpWHOUrUeLd
aY9QawjCmOAMX7/SY7S64q0C3mxueGs/OOcuHkGHXoo98ZrXwBnlZD70q1yFAauko8EWL6VX/V5F
Ul9SXofouMYj3v4vUsRkomjDujTgoUw76QtzSLlxLyCNuE92Io3uudopDUWfhe1/Z1cLYCGEb0wP
agRZtJvBGRkmXqOD7HPEDfXnYknH/eBmL26n3I9lq5xHWcTmpZbyyTYyNqlWJnl6s6NHGf+Uhc+N
9Vn/vf5N6m7HR71BrhvqQSpOU+4HXCi5h6WkNt4cazxtp9jEHZ8x8rfwshaI+TEPbCexE0FJZAvp
8DQv4Za4vsoXIlV4SsqElCdghcPrXpJKQ7xlYXws2ub72d4XBdnQlqfNdwMWp269xm+LaA5Sf3qY
5EV8/PVuMUkyU3l3+kGK9pAZa1rMfuZwQlwz2eqebnSVwC+4PstSHgvTTpHTiuEgBphWro2bFIbg
36avpVm897R1ba25o7dwtaSWN7hd9/M7qFFtXW7/DHs1ChsktBKoG3PN4psErYTZDrTNdIMxU7va
YRae9ECcTk8g5DUVq9RV4od15EvrQQNL29sgJuQtuu9ZjzIGzPKaXuOmqxgrWrN5h8Rw3JgfmmFI
S7NqT7RLSZ5hcuS2hbylkYtkT/yiD98Mbc5KduOD4DHJIyM2Yp6HStlCPYxsuGEl6gaUVdJ/FqiY
74SlbjIwr6efLgxHJs39WaHVRxTvDQ1VVqyq9NsOM/h6tKcP5QMdACtpTd5lzAeRI9P5+hVMpxEl
c4Mu1eBejZ1bZ7UPNbN4IP/JzBGRhSCT4An2AoiSc4mYPDvJ9Vn/LsRtDG1XaJYb/GFdHuFlFefn
jVn6jWwAbWIDYqzw72TCBQ1ig9ZVN1/JNGOFnc+5oAbBErga60E75ovvT0a/d/G7E+2ei4iT6/1L
o6M1iRmL2Kcn7hWFJcgsJLuzjbS/yzoFHDqurJB0Nu4hEei4wl6m0gjNNDnlU9UGUQSZBjhxtG67
9XB0hRJSwiPGjB3qtMUmvBCc4qXeEorQEV/CjZQyGgwXCofYjzQ+33CIHfyaqJKxKmREKKkbddnN
W1qSICY25+0SYnCE0H1V1Knd5kEfHwfL0AjeXPRjZ3fv/+wdY+SPfxwivw54UST2LjN/d1Dh1WpF
pIO1ldsuWDa2mVGYAvhKquJezm8/DspZgUqhYJN5hIDRhtAXaYenZy0c6W+FE1KTpT9dltzBEEKq
SvX/WZNZZh1CeZzHdTsL/jKi0a93ymyLzewZzG4uyYoBcbWYfmY+sr/BbBQPqR0y4MCoIymO/HEo
b9ZErXb/nz93LQT5/JUz+qF2+4xJwKU41N6k2hlwuyK+GldndWUuEJ3AeO2yJbgvPf/fObEot9+l
QXCmZBiyj5pQZZUpPyVOs9dgk/QRF/RrHIS63QRqtlLduiosehwAkep2vSzprhVVLa0/5khES6ZP
6m0sZrtar22wFxj8oFEv8nK0A4IrSTt7RsoXKT6SJKF223UpVqkVPbN8+0Qv1FX+XYKBIcOeuMH1
0C9yILFeEYcDumNrIuKDKeexj8pgNi9Xakvba//ZsEQEkBx8QWa3DfUz8Ma/VeeLBu6GFVeTBsHj
5RdPfAZd0ywTMvBjFchR71uP5AhQ4oHj4Glv1vvDiM4nYJ9TMnFj0Y0GUyUuJIxnApEAxKhnn28q
BFCzUDw9qbZMWb40hSU8lLGhOI2F6E7i8sWpLId1aPK/yM3Xa+lF7sYyT81B3o1Gd3DfVlXxw0y3
fC343zpCLFw8AkW8mtZ5mDhb/zv0io3wO7xalLP9kaSUppoR7VhK95mHNOUlAQIX/BuAe5TBe+aQ
s55D94/DcDiBb/lKWC/2bWGHNU56v8ihPXlOksmQ5499EIKlpgHt/EuLtuv+kgQnHsfHs3+d+kDB
9poBTZ7UYJz5nfQg45A1sJaMhxvIxDLz+VI01bDHhAiKUR8oZirgV4zyEugBt6ZlduqEWdvLrqc8
skKj0hIqNX+pJE0233jrRydzpx0/wDKnWecd/8kVLu5+ZlHVWWIJi/AgVRHpI1gykBLL2D7gSFp0
pWjTNWe1d3HwUA4WfIhPSitC+XURmXrrq9OPlZBQmRwin/p5GU4rbU2TB/ux00uRDoLC9w+bh89u
UU2torsYx3NeJHEpzmbNcomEANe0u8D89vhDLiQtv6qXcCA5SYJxcyvU7M8nyq+te9DQU2xw2FbD
fOQCdwwNQXeRZXn0X+BegVr4Vx8elwvE4Opz/C478hLYyXBRHPNJzbNVm3BtrJJzkwdYgdeai7tX
q8QFgioSCTywfBkeruI4XQ7sTok4j2QVo1pMRJJ+MUmImRGeIeTWoTieYbgrwkQ0uBQG5GOeD38R
eEunl7tpg21JPUkp/+ItQuL4csFAA4YODpCYapZv1JXZ9/1Cre4IzY6u0HsxH/UkClHF10oG2rao
Xu1j5+Abi+YSuPORmvCwy87iGDHlH/rrfPBNpl8EYqpfDXiGdA7EnqBqwJGvzKGTI1tGFQoJIba7
RfEdQDbTUWYzFVqVV6a771i1UsmnR0wbm0xreWbwqD5qmxX8L0V2MbgeUM1R+wjS42L83Shkc8rw
eBzGtM06AI9nD41iiDc4+1hlA/mcgVCNZ7F6ddHy8vD4QF0CJjlVedscJm5Wwq7LFvZ9AYwqJ97t
/eBmTNXqlQ3XU6SR7ivfbJ3Ad2tgXaUasjAyJbK+y79ovYik4sUG2N0PPY6X534b0lQJVQ53v82+
A4kMtq+rsVpWDF4JLfcMkykWQnZpgRjXSRfgni4o5qljeBe7IhP99esT+V2cGrCTCXh5xw3wI/zi
ABqGu4K0GsBb6m0yWvBoUi2q6v38oPf5ewYJM37Jo5+0xZsTTHMVdCzY4hIn30fayXCH21WzdBBQ
uDXl++HJlMvtm8rlwaPA0w7nzYPi487t3DKROymHhzO+BeuGSjfzKvUKHXJ1Wiin+hkPOpmhB1IL
eWRZAhJ/n7Pw0ugQwtGsBHuhjorkr40NL117P3kGKyx0bldlcT/9ZzWNlVOUvTT+l0Djj9pkhNcc
9ns8OZcx7Rrp9UmZ1NUPCL3WU4wPDcvDJUWDMGgujUTRUAAlk0TgcHYaN0PjFvKSaePX7MD5pv59
EWbc80voiPjn5B9t3+wnSFXvOVy/c7S182rjzu271US8TERg8IiTui8TlcQnLg958HXCqJpK0Npy
O4eWRZ4cRocFTNLxp3xzi1RlxCTkt3ivTewyLvyxHR1Snx5nygbjArF5eeVOKypnhiJBfhKmbuWP
cbfwDqejVossilIx5vxwp+XQkSWa7ARy9tWH0dFJ2rnwN0yxnS0Puw8BY2EPb9k5I8v8NY/B1Cux
MmPqWjUnnMU/YrkEhCzh9bc5aEYXGeaQSnacSJag1sPrZn+zXkUsHiKLv5l7gBjEMJVn71Os+zWn
8Wkq6Eumsrndq7AIENI+YJ8M3HF7jwuBdcDPHsEfCfjKNooVTDHk4z573yfNogTQzbM7V2d8xZIz
nZa+YOz9VHl2webg5yJJYz6VNn4HmtvpzSgW5jfwHUoxu+3OaHgNU1zZ7tYaZdcoonkqvVhnzQnA
V9vwT0g4UDmP37PHtlMH8QNXIPSw/JkaL9KOZ1Jcs2u0//pqRpDe+ZtbdfIYB8BEJMw2KkMjimIc
qjWMflOrpCNft5UkcJdsi6hL1i39aVvk7tfru7ATy9eqFj6ks6gPn4fI9YWkFGLVNmOXHac7GPZ5
I9JlYurAsBuqpcsX3tqGt/lNLaOiXIeRP2WFypQBSOnCZDb2314BEZhHygAdF1pcdIXg5rVtC8zl
3V0vUfOICF/OZH+sotuoCWHEZTJSP5Qea3ip1EMv3UN0IGBx6Z4I9SDCOO+5RUEz4TyT4LBLWqJd
T0+bCdl/zJoi8EGK++QAgU3CwHLpEL3lQwwdtxI+jE4MgMpJYNvTztwpPASU7aZThyCzgAY3BZqR
4ZvfL0zY2JdjIRSaMnukzDIL5sw0/yWtYWqJUdFqP/jH3INIkKQh9aT6M00EEG381L6wiYNAxguC
MZuuDz869DnWmOpiOlfBPMuNGkpRVl+6/Qlum9kGKSM7fTyEM3jMk8BhznDo1up+Fe0aN6lEgGqj
Gxa9nkDTSHDnz3/9bYuO9BiIBXIRkQQjVgYTjMSeP7mJHWU2anIPojvE2054cm7uFz0UPrwC2e6Q
hppJpwUgPwsxWufZF5L5gNRitrooF2zSxy+O9mxSoxK8K7dzag2x9lN0fe1ClqaSfQLmIxk22138
rlR57pv8EeUQQ/BUwFnM3PHsgabH+/N8yss7m9cY8JjhuJ/WeyL+Y0QlWxiUsMPQEXromn1LoLHZ
8iHNg2EAnucsSgcry/tdfcRSpmIftW5NWKg8vVKypbsnyPzRjrpT1RJ6N/5gPt+0/gI/EbbwnNrY
q4+UsqJYJsHB5C51TBAL3O5xBcweg37M1oOCGiL66MLVoiGZ+60b5vRC/XbUE772YNuLkvPt3+gb
82vByuiMKB6xSeYr2PPvWhuxq/7B2xxe/mbUu50Rykblxf7dOGlgDudjc+E5Ro/i6S5mm0loxcsc
t3VfdJVoS6Yy/jPNb564tpMgD4an6XyaGr1TofCAPxVwxoCGg+jdvlOXjUdNYCnzBxGhQJmRZbjM
/GYKs9dEbZI9SGjZ/5Y11WpoTvAGddf8WsZeQ26cKBACuP14vegcKq6OgZEC4gkiULYk9eTB40nm
E1W+AZvGx1OrRcyVTEfK4sD0mePY9C5J5gZOuUGBvfIOEFu7YOHY4ilPGGMsWJhnig7KSGD5wMDb
nLEOEe/5+yiR74MUuWX15t++OV/LwNanZwRUEOc/QOUrrGTExk1okD6ZM8NsL4gDQ9XJGbXcR089
YVnZ8l8PvWQMD1Hgp4YJV1QheWKqhAlPpOrU1/IKm3tLYMXBL9Q0SPn1QQYtksu17uXg2b5ak94L
UTsa2rQneXlMXTOzDNe8cylmXclPouH+OdSy/BwtrHXg37/OiVLVWAjRvvbqBxMl/MPdAJWoA08z
Uw9uUf4x6g7x+XwdiFk30RE8KmWaPGmZWsuRNhddkLp1bV5oICtthfbO0ePk0tfjiYJdrCIg0LeJ
j4gdycvc5o+abY4YtQTx3GNyyaZLybd5zD936s6wqCJAKOFa+gmTzCgmWpkJBjs/cUb0l0i+KzWF
W46VSwffMTD2f6yWRKURNdVIydAFylrF5nasLTp27vX0yLdSl6lMQrecvc+6AO4GMtsf3r3w7AU9
nhv00nbJokqWQFeXPoLHKtvIt8kAvuzbQgKsRuUQTySA2WEzhNIZG5HmEvRMuU7BMAGeE3g8+dzN
y84zfDipHzVoEfzM0Wq7rtWxqISQasE4ZX5laZX1TCU8rBhjZdmPRTPScxVWpQkIoYl/5XSadEcX
Ye7M2KaRr1wDYH7yVx2vGb5W4Ue6/KB0kqwFx3o3XTHoOiu03NEEjFI2zPhfy8/g6Q2LIKifU6/2
TGZQPWnNJR86k1JLKZwwUD9WETDc9JlsEhhWXXCg91v3f/GKQza44dmjm3WJR1+FHQYq/BcdxjDf
fWbW9NaVIqe/xra/9PZ2c9ToB29hQoYPE9lbUbx8KFizRx0Jkber63BP+zWApbtaJFlSJFfAQEzD
h7FNqsBok4WjPb+NdYhSeaSxGORNBZolyZ4JhGXdtkiNA2xN3STCIl89cRiw/y1uOhzlFFkrjKH+
4pmAVl1epxjHUwlcXdgxS4yxnUfxLmlHfA6owVpMYeaflgXDOmqyvFhUmLJOaYkumsxlpw+rEYDr
NDbQOWiejJ5IDlY7kxhwzvhopBXcrM5/XADoJ0qQWIDA66Fxg3jUDkix8Zif5pmCp62I3j+ArYTF
zBt0HEG8jVnMeusSImhRWpK6+SgXT1fy9XLuJ2+4HemW+TXrM+NBISvaUG8kIEYEtxb54TPaHtQL
auxDJn/8JhRUoXkS0huIK8hp/JPYle8C4hsptiX5sGhllWmNyDXcKwBdaGEqbCI2K9w1/vi1tyWt
SfSGFVYQ1qwzYbHZkKQZKxI9hWarHS0yNhUGjjnnmMSTFPNBWGA8EvUaKtCR5uo/QkOSZZJUAorY
ASkhn4vZz2zktdWnWr8XgMj03PmXYhcMUNdBT3wOkhxG1eFCZc9AE2ZFrvMQk8vageXuNSEVPAPg
teevw8ZSuLfKj0YSRnlV2rQWf27wwtMLwA2x/zQrLG5LY0SAAvWbVWVp21vLQuYeYve31lxfTcRF
Siw0vWnZf0ebegGhk1ciMoh73RkwB5Yvd8tf26ujCgm6sNIXL8ahIrszNje9r7PGkF4Lz2tq1Emn
G/+u4+qoS0Ns8l5OxbuAAr6mE0PVmpkJlW5sg9XgXH2zEW8jmkldkaU72HQCuRU8cQ3eCC/TN0Xo
V3nm6656Pd2H5gwkLnCXC16fEeIrfq2IohkkalxKdqX81BCpw7uGJMsj77IYD3O6rKq1vFoI2ge0
9L2MfL+rwjw8g19dGTqFMsjSij4GvluK6zeUcKp7KaNgLmBtQMQVRuZ9f+Qk25Nds7plhv8GhJEv
MqP/g90/EiMzkyl5ys3le6B+eMjqe8kEJLSi6qax5dL6L/Cxbqf8xd9qB19QSmRVrSvgRMbKbuUn
vPU6ZMf/visKmGQiTK/z4nQbYUTb+q8pLF6X2bGAUNk4pQ9uCJdAAWBye37qM9L7PV+acS5Ffmwf
Rd9LGfIuIAokwTiT/tb2BxxaTryOsDN7OiEtKwFJShK7CIPe/t79lwZyroJoNiniUYOo+6OqINQS
/KLnhx42ZRBXis3WzqnkYtybgRx8kNeMH+519rWZjYEAnOod9xahjXqPHh4yqPUQ3H62JQ2fZwEM
tZC3nBW0rECtM4OOaafyZKW05ZuqXztQpAI7OYl1I4HS5AqJXkqgMZKriqCf7rb7PmsYReH713Hm
y8MNedflf4wzS5Ha95ZSbcDpP7M9qS8MZUsBETceNJcy4C1rAbADFneeglk2I9Z9F4CESYpEzULA
MFFdvjfd4xHvAYtUUWIat7I0ZP3f7oJPeHC2JCxsiGbiwSPGlnslXUpgnmuRGSeEdn5meo5vnRRV
vjgbD8fis5aHU8Ha86cBP7MTHe1Ns8p/Owtgkw3oPVHvol07fpNbC7xDbkFGBTcQs4D06S0kVoFY
gc1gJBBOGDL5+QSdr0WIQ9bNVviMcGSfupxPBhN1IpQcnXaRO8Eq+4h3LIlULTHga+aqi3qj06UN
J9FPHU9bb2C/BVdrLCsWU1UoO81TqAQDR+z+ueiAx5+1qFY8/pEn2yFARAncxbyApE6swVSd43lW
xL9naWY7r1sH/4uvIPTDO8Gl9dwikpTLvO7dxHICt+4XfhKlUNDy/BGyMKF91nqw5kndWH5RCM3P
xhZ0DeqSjG5WkQLI/4bkmb9NB7BjixzWqFN0L9r5tAAYIm4zSrY0L94iwd5YTBIgEhnjKboihcMP
b2wKtOCAohw52+4Gv6bUaPf3th+9h2wOITReBENsGUU2jdMv3/GxxZIsf7EYzqqvrToRHRdmj+ag
NHrRiow/qrLUQm5JM9+nRhfQHJNOKHo79rnIIkep8V2dY+/M9OiMUEWiRUkm1YSo513iqEyVbdiw
4DH8jGkzgZ+3ybjKScthYeEny2cRcPRUbwUJRgO0hCUPkfrsQ/8odWQnxehAA6oxiVkmz2KGy19V
Mqqpe5g5/bsZSOhsh25eyzZn/xkOfrFMxf1z9wBqrxjhHVjdfPAh+f0+ov0HGaeuEQdqhjAVQZrQ
O/dtDhdkigNpe9luG8eYfET0OsYPvvo9sejbGt1p+wJi/4YJH4CegjXgVYu4zdxN1VNqQbQ8fxy4
kzLIpeY4HTjxu+CvT4EEugrdiTd2s83qzBNn3vJdNyeul+1pzTnuxBde/nsBBC/5jH/rWISe2YUP
kNKjQL/9uSCJRwz9FQWWTj3ed/LeX69jXf8FVYRYY6ys2VRACqz5ECJVwPCD4u3XAVuyIa+gSvuO
22dOnQRLabdIsGaBYNI6w0//ismkV84dKX233i3PXuZv2VpTf/u+4keaHeK2Uq4eJhRRqOtscwh+
wLjIqrEB/0v4KR9Sp8Wbomo7LSHXepTbKdgKBVyreWiWNQp9dA1TWF2jnqsYnHz4b4CiLiK5KO8t
JDdswewCLPQ0HgMRsGNwptMdeWvuPlgmsc6GyewdsOjDHP+dQ5gStRJpGIxyf9/oIrCENZWr4veA
PyZrEbFa0IWXDx/8JGpiYjb8Fwsx+hWW2SVFBqWg4QnSZ3ujXxiWwPXQIS9rcFpNv6Gyyjxuk0RS
8c7yPCEMHJjk8Fz2zVRSM2pz0rCJUuF+mC8FRGxPhvM4XIOjOQkUfE5HwhmOpoQ9R24ABxySaJiK
sez6Jows13462EWpx5l5UH4DixVtSBfbq7s9yizXC2sXZyAQ6ErjdMddgNa/TDAEe7XEQie3kYqy
1CJTxrr9rwicWu8SNqgcsT0aHpiLqxPmTl8H2KKGfrghC/5isXjV1PRIX3qURwj57x6aqxbFoTnv
pI9y8BscXg3DolEQ/zMnCQ/ao2joFg3yl/oWXgHnx0gAcr2MCUrzDLWwtcqPrEWr7yuSFQrGKESE
GHyzI8sZGBPaQrNcNOdfJsG1/vt1KB4ac2Uc8RYJzJLNvJDAkTanwI0br/x2dZaR7xW74N1/rc56
4pjz0t4idtFQgVZioR8Ik1e0BVMZlDa+dCuQGBXbn22wr+vufDiUnvThivGkrdiEXTMJVEGqm1cM
z2/3GqrdgGDHzfOEwkoeOAMOcOoVxz/gYmoduPxZVgClZCE2Ep/50+0kYGSfwvMc6igjYNS7NAbo
AqgjfuLd5/ybwUdG5419DjZuI7eMe2ddbxyXasPQiHEnIIaoodUDK/RrFAWWrMdElOrN2jhPEHKO
Wrv4+k3VyIueXNfZzvwaPr4Tze/g6OC5jFUHFPa4nHywShGVJk3Qt62nAYT2+J2kWGYCDEXYigmr
92vyOknvyiwo9zv3a478FMZi81Rp0VvSM1ykXg31wLsFQpr2u6ocLenlO0AraO1LR+zSUQ/1O3oS
QC35VBFW/sLBkzQmbxfk5KZi30OAffQOZ/5m6dNYdz17yRSrY/gv3HfEjQJeR2A6gwK7x9tn3DjY
o95HteWiMvx6CZ/EhMe1fWOnDdQsssDQvqGqPEgCc7yT16nIOImHi7SQwk2GqME+Ti/aR4jnJm3S
7UPTqh2D1E5V2S+Xt5C5y7gTcbYg+2473MuYcjNnp2VN2QIDEzVmNFA+96cDu5bYAkug8QvdXmvq
QEzu32F1Nhd6Kc+9uX+Qzjyu7QeWNW2WgiSF4Nl/QbTq1Cxl30tT06ZFP6Y8xTkHdunNsAfuPShh
q6zrkxjS6LWwvJoWq6NtpSCOez7Dhbcj4oQP7q+tO7qmg+ul1yK8E7GFZzaG4YVODVB49bnTF08x
Jvfb1ccouG2UFkwHalG7x7oG/lUa2X/sR/kNPCCF9XGq5oLeNGc6XTOPGr7FJz+xyni0zq4i7J94
zoLEhWcWmB/n5DNzPD/xXvpZRRtsKF/rWYRSIixdm8Q+a69tF8zk8rtWJIoTpLfxGzJiLwl65hI5
q3ub+wMtM+XoHRWY18O3VuCilZTTcHuB1O3gQhV0qqa68BcrPHz3bdsHfZjnsSKU6VR0OoeUwBL9
XtlGkUTPY/UAlo6LlVsPE1Evesao6IlUxAxIkpKhj2o6x8In6YQbOlQgAVV/oMEytj0w7LLXNPvE
+DhvyHTPUKYVvcTBa1DD/ln6uMdWX4DDuS1X8xm8GOHnIVZB/yi3DQUogTRiPJpO5gpvGn4GLEuS
C8f6nEXMov4M2ErsSturzrWhcy87+bVfW+44kDC/ZTL0KRCXLXI6XxgqlcU6RwPvPZ5cL9BvgUTd
Iwku5u6KxQ2fgf8iQ6TKpZzWEFhAcV4BAGhUkCoJ43WOG2pYs4zyOoLqOwpu3CjynyckgGv/tGwO
lELx/Ud93d4ns9Rjc/dDVCcs9YNCRjy7cpVzah8jwLOvMyt1Z4nsn3wybfcKW7m7PSTCbXfS6Gj/
fsTIwGhsgFj3fedGWHVmkRgvoZ51OZU/ApWj63/Ld98VoHEqNBjW/Sek79+4l3vTJxVgpZaKfZYC
W2NCVu6ufAWRwVv8H4U5s3dHRnidQz45fz11lF6A3r7R51I1PRIkiCU/UyyRGSnIZOvMhsqn/jlL
mX7VPWxgyAto79DV65Koe9Zn9TkoLC54ZDL1wpuyRIXKqHCmG0vFVyepmiACqldOjIJpKmmBOjb7
eEs3qGU6mRWFIpiYBHyX2/4CvqW4x4N11brRPe+CDAe9/FSyTRWOJi5nbwb2l5/4k96dE68fqXqT
hDYd0N3HhIYYNtr4q/DsTyLHD7OkQ1xdZuIcbx91OrJhlSwmc3YbAPS9Etv5ajOwWv8XfboTmeDL
xhgrRRApWFHeqjNijhtlJX5MmuWOIQG2ilBXdKrFY63+Y86HQ/gFjc8siv6QAFrKZWnQILjDG1H+
FQ2IrZoOge2qz2NWP7wK5kd8WLc4RVKuMANRlYtUE5UDkxMVn20kY/e3xTsAvJHk/bzXVUhRQw9D
813ie0DCVAzAsK66YMOzs+M6e/rita68LgYz+OQVSiLhya2e8rJVTEsbT/DdyDF38CYALhECoCO8
s2YeobMJPoQCDsH6pobm2oF39r7TXAgDLB6PELQp+k6/HuDV3SD60lH7emob/XG+emgrjnXovxHA
3DVJEnPtzxN4Dfe/dH9cfXpriFnt9Oj8kMz0B/iSPQwT3eXGnP2ZL3nIlET+NV9s7d5aSq/KA9SJ
Ywq1DsjN9Eb9Z3M7MwjOW0gOOZr0Ff/RKy+0bnrN70NTQVCCrEilFKc7Ppnfprn0t3CSI76B7GYl
r6j0MWZdk7weimojEwu8cUgbb7cuMreuGxti2ajEXg0vLmsSRZABahuaDe3uVIcuVmjvuazp+thi
lxHo8DFndsw3u9cUK6TCC7eGc2srjIHBXei+gVCNJDabzM4OiSGAZVvpV/X3d7W3hYMVqifYgsDo
6CaTfqLhJz81KT5xp0xbi7AInIS5FNs3MAhfIfKwA9FeD6Rce8MgynlRoukUousaqkhOG75x7dIB
wtYwEo+a7Nr6MWiXcxAbl0FmArRDpouDTUlU77AruI6HeZtvpHzQ+a8RsA3Z+i8TUtB3zpW25/Pk
5SqodeV1/L2HuCBbaE3K5xXnACCynEvd1gPmPPhg9iNwrvuw4sba8tBfHAhRmW2D+bM+iRBp8vrz
GeooxeH2BOsXRarwyPTtKZFc5rjfThLJZn+IoGTGwZLxuU75lI6VAXpaE0L9D0XYPsyEuHivk9vQ
5Sx2rGGDAYJ+xf5BnhF4PlmuNMcsoLeDM48jx8UXOPvJ+srt8eJKqhf2wN0pBAZLRIdZ/i4PBUrk
c5rH58F8OTWIqa/nhBJ32kWSzAV00jTCat/DmErlBA2GkqaGYdW6bBEjYDxrIIvebJzxhhZPfjyA
7pmCSLlSoM4G7JlVPX8lCIFHjuuPg2Q6OBjc9cW2HGIIYLliyPDixHayY699ud1cPahLmFqYgq+G
LbL+/aJI+EWRXx3ZwKF48apL7iHlzAlwpZTISy6d1K0sM4Gz1swhGh0vrNbGV+Xxobunonpg4mbL
yzD2Dx0awNmGTKgq10aeQHH5rscM+RdBESLt7v0GlwYltTvVN0KUnJ/JZXbFr76TpZU3jRScXCVg
+y+TjaEAHliyXus7aGdo72T/X8a2R+WK/uZzXMxhVPtOtmISgsmlzXl6DW7ohj8gM90h/CbzkgQI
Acb3WjNmZfAOvMp8plRubv8F0xX5Lx9goVyKiKynmif4qIxtjZcGwxHZJHAizsIEgJGrlBrandQ9
CznLdvbAYQQHH6ys4fbWmCaV8Q5AN3c1yJVMDBMOj7dqCge8L7EvbJIwWCeVoR+uEbpP/HQ7dAkS
Tt6wOqZ40EDr/oMLg5vAsDLzfajPkUel9IM9yNqofMuHZek7PHKBzk9nWLwgXvEAUVcIuUgOvY6g
t5p1nMSXdl+IXv8Dcr1mVlgBAxCCLRj+bu853xS8f0k8t/sKYskW4C6zWWfA4Z2QGtqZKWzAHQX9
xyowk03mvTgRIOGJl83WdUZT4STImfgz8j0adn/fbRfMgR9EbstTA1Qe01W3LdaCF2G6S5jV7Ud2
w5lcHmG+0B1GFHoBa7OEkO5pzKVEJo94EjpNXrDrYbXSzG3LfpAODYesdt0ZdyNvSmCY0eJluH6f
2jYDk1rpLXuEn3aEConj6vTAZ4EROMlfXhjhzQ/UVlkMhxKrWFHPpXhVS4lQgWOGerDq9/Wz2Yhr
ka9lMCz/PxnVJqCPtYlGCbTEqCvWlfmwxVWuauTFRnplOBmeznubtFdv5ZHpZEOtDu/0TbkZdrBE
yd6KbJWqIItAsb+cnKlHGZbghmtbTyBzUTy42X0gI465Yr82wPqidGKhfkQx4E1NCPLKiZKIvGi3
9Ix3rcz/tfjhSiippJDf2hvgQUOW28UAwpYv4UbhREjAypl0MerUtmpj81Uuc4Y2GL9wJdhDZC57
/WaBr3JZjby7nG788DJiPpdaAkTwZqQDOXCvubqI4NgFA1VUu44bFFdfKZnefUrdljw32ZkBIEce
K0NbfgWqeHtgS3QyaKqL2I6n0e70FHceHXoSAXGwEqfeGyZFkYVNwzPeuWCe6p345cHQsYVV91KM
voifPwk+/PxOioiioM3ka6EmrkGJqw/FGVLpmN+wCgrZVHC1NFrD/EgnRk2pOQOplns3x+/b75VT
TfC+4tQlynZIhMziNzvPkP4nu1XjWeIG1H+1fwbs4ZHdKO+xPwsDvc0zQiLnsuXj1z8VkhkYUzbi
qPq6+JPNTo/cioDIDIYk3D5X9SW3O5MVs7PfzWR6tJXE7RHUQ81CN6LMfQEjzQCSzaiLtB/QBnYJ
0/gMfty/qVEFFQlcNdhdDUeDFKwb2N28YdwphXmGqdgMyFlvIYqzOVMphTzF60TIP+ktqyJSCmpV
O7Fx6zUqkGIK6ymyLUALGErTh8Yo5H5JxidQvQ0lfeIJouB8zVdu1tdNQ1a4rZSbld9e8Gc+FREW
O5nlsLsPYwdHp+bjKJ+SIrLNI4CxuHfLHbmjPgUw/LIf7NnUUIWHfifIoEvuLgOALP7tSrjoWZjt
HtvaPLd2DMdnfKM+pfCWYVFeme2lCWGGTQATmRR+BpQgySeAdMBCcJG0GnY5dWggEliEFQ9aK6w+
bAE+KQMdm5cMh/CuLELX0fvN3cg49V70bR/1DBbG+0Y6wfAP7RgWKrbWrLZrY7Euk8AS+dz6OgAl
UqPaRWnSrTMozt7jEZVTjVEUnqHOEt0sN7/iA+cLqPM/EAvE2pt+qQQKBsPQXdHHE7lHMJkcq9EW
mUNktaF/99SZn5adglfFYzKqT0SupbegOSGH/L3c7N9TMW/7ac++kEQxiv+NXixVMLaQ2Ze6hlFQ
zzucXPFhpNtBHAXbvYK6YamDxOLIpwrN0CBJ5F6lPHBdlWeLZag4rgi5yeqFbL6P/ERLFf3rynQs
fUqhfpl/aDpXTFZ+yL9yO7XiMpbvlwYfoYiiQjalh9ThGBLDZAuxpgKrdCfFh32YxaLARHkgLTB1
7cBbqMXUbZS1AiGtKPhHF5BeppbiZuAiF83/TGO3mFPOCq8EtZiVvABl/1MBTSy7A7slba+8T21G
Yf9EkKOD5LVyXEG+315nei1u7stFZdyzr/V9w1XgoG8i7czkjixRnLlP4lWmLUUM0GGziys4XKjB
z0Tu+3txsp8UWQCyQ335BBnNvv8svRCeev23RDWWQRvgaWEOfh6xjbS53D7VQiKMtpS8ATaFJYhE
aBV9BY+0tk+nb9Dh41EBXJ6THwM+rmgUa3dB6SHqZPmYSpwwGlswprxshuBHczW3UfdvkCDOvb4P
0FA/dzRjT/EDTd7B3NyZkLqj2NNBDGUMk1en6fr7cGoHGaG2Rh/Iunho4CJ9Xk4N78lUPdNp+n6k
ikF84wlwDQ5vYeyyHnI1NksQ00bSsBG/sJoG0pt8tbzEI1bWYUBDeYvtzpre4Bhv6z5d/Ha5M9vA
8pvmGKsZpKNKAbdvXnIBCUkIkardJMI1q+XZQsD8bqw8Iq3DfOsR6Goy8vdQNFSGiTJj1eXqkLHo
gOBM0NYvE5SQXZmGGzDlGifpsvAJV6n/lusqd0BJAHR3j2YsR08f7JD7pX7I9msHMquDwcopRXVt
GlXGK5NJivE26WnjBpwRb4lYdXs8e3k+1yDP9X8utqjUak82fvA6jwOqryHhyt1RMLiwo8V72fBz
bK/L8Q5S+e9qSuhsWxJB+gG6PgKTwX70gZLy4DqNcMEBkqTY76Pd1E/nGLUdUnnv9Bvxzz3Iyayi
4piJuWmjP0PT8iS14B1/duUSVId97pdcmCEqA7BberWLPlNOXgoJjsG8JwfYU9flI61U2PmEKemx
Tdb6hljFEJGg2Zre7UMvezfc2SSV4sJFUHA3xevvpdcq8UP3KZKuFco7oNlKGlgOpQvsXazJfQPO
bhcnXXbsQcxkW6gHd2wSoiPflWY0ni7i4VFSoPrx+eUsfP2TttWuGHX6UXDu927Dq47syk/hJZ16
vCfVxQHqdw99oVOqRNEzCLa7V07DVYQA+BVHau5ea3qet/3pUUKKoFK5Hx7MorXGvcwcNNfMUjVe
cAtMvat8y58oOLbajSJ1G/prugjGwHO1rbJ4Cxnbpe1cIKCihcpsvN/GWzzr/S7pPpOKWDnJQzbD
SSfaxoNrONoE2p1ModiIh1rPF/Z91JeNi4wtPxNuQ9ZyuKjjIbuqaIK6XTwtEccWm0ZIhU3C5JqG
hMjH3N141pbufomCQReFsLNGIU47Hrs6j/GFFXVGeIkpfPBQ4eC0gTGC+qcq9Q/5F9omRB1x2eYd
C/Vf+dFmPXxfv/HQqpZtiKri2qwuFkFogqfBJgkUyRXqNjXY1TP+qROQZPfIf8usNKtrmHnXNHqy
yEyCWTEWUpqKUyuUoA0coRmPGjZvlvLdJ+USt+WtfR5znSt/vm24TYMoj2h9oReycu21rMxOF66Y
i1CXJh7WahClhC85DLF72S6cjah7zN05ooS35hErNAkfHFNX5Or5ciKA7e3hVdlOmV1KRU2IyIrO
bwDJOj9vVLZpmXAErW6uGF7yk460yo+iKmePswGiiEVWJk8knzSKeAbnpDg7tKDYN86hBNVByd25
Gy/TwJQtB1/JMkzCPMcYgmaioChodJL3x6saG7jN9yD6qCRrPUGyg/BfAkwCRKZRns8BHy6M8mKP
BUEWnJOY3vzCcCiChZ+de6lybDcjJjf1TLNyc2GcWl9eHLjS2XMZr8c1wdfrElNhiV9N1RBK4RHE
dtkb/d12nTqeQUaNn6cz2ZSyxglHCmd/F9W8ZaV6T+IYzi9gkQw1AB492BTgvAdzMIiFI6GWL/dy
ax6eKqQ3sgk5XqGFoCuAR10OZijVMkSoct6vIyjbd9RI5LUt50zTmY7gy3+dh3KbBbhsutACpN4A
/YqNRKpRamlfNX5WANKjFOsexpdaI2eprUvfaAOpEm6aqi5FAOSG8TFTjci3ymrcJ1wZVDf2bFfb
lUNXgTAlTWzXtzUjo+e/kYoIvkJQOnvJO86Y2Osqf4QDjc2fcfGA91ictFLU8U8SUCZ24Llor/qv
Zhf+Di+bWcNgpJCIvnMN0kpJCrvWtrR1/NzIEnlAZN4lelMEX04/HPol0A7J/MvM/nn0HW5+fZBK
GsjKjefmzgpWFlz7uDQ38bpfqUzA0fwAX8phCMx3sgpIP82uy5gufk6QkxChGkp8KgsSAjyDT6qS
cCC0RI3BCpwQJKH0pcuPHSerwDBGRay9KSRoAc0egR4To06e+f2KflVqdj1x1pna0vqNfF0Vrtfl
HorjfEaH+8W6hJ9YICT/yb4PXUbmY0YeBwC6XtVXDtpMqIq51GQseiOl/qEl2ubiRq5ylXjVudii
Kg/RtNxZE1thkH/e7umjC5y2TpYLx7zRJj5eYcf5iZjRi897nwrO7pyZNZFxwwUnU+nY3kPbwPHL
0HOMYqP73e6Tp/YWOrDOCi/gqBmj0QA8UYCTjjodKG04XKrmG/9Wwz8NtGKMiyK4kNWUr5bf7OwP
qTfGB0I2kbxnaFVU9WQBRdp9C61T7QsvJSzrVQR/sYkCGNnH8Cnpy7c4wI8YKOQ7t/Y3y4zEvqE5
6lBAWYUDhi73PJ7j/qU0d318pG+7RkGjdYkKEsMPNzOiXGvCgv4MXq3oKKD9yBgQIWQP6P6HEasz
J7LjSvzCOvpEPJhtLwdqTlf90zFDYPAtlstt02EjfMP1S7YPpkj21G+mmYtKLSpsAJOqXtwVBQtZ
wFGKmXCQTjqe6IYldZE1rDlOlUKksBK6Sddl7qmIhuRDml8RprVI3ONlh4YcqrYby9vlfMLjFFG7
hI9EMeM5ZEMZgrmeCCsjz2d/ueOIvzHGjxmk8ErYqyN2pVXuj1xVsgw/YdHjCRMPV1EUo6qA0hYl
neHiZIB68tEobJAxYgiPu+inPTyQG2v5BKJQUBnZLFSGZOuvsjiLAbZK5DkH3o5THIo9t29/vquK
6/op+XJnZtsZU/PDZpXA6S4fFkGp/2eMOnuxVj7KrprCd5zFhmKapqKlVK3VbsFCpTK74g4lr4x8
Fr74KEUPTZw8v8+susiQHZjy+hZvlAAVAuqRDc1Xci4XDSvYgtriiY3dnlGTtzGXYmUP7GXmZH2N
XVyeTisGIY3sFi22qEjoADKNvN/js1UAhFjRv0THjnocTFOaZaBMuikILd6fI1vnhq59tLMaVefs
s5WswAyJ7fJ51fOe1W8Kra4BtS5U+CfFAKRu/VVpnVKnBeve6BINbbqhJt2lm1ZRV/blpdD0zAYJ
Rbf4hwnJDpguVr3cUOyDRcZWsj5SY/k8HJoPsCixvJ/RMeWL3zUr8n2hYqJ338xk/N+ktA0uK69k
QOZZeCvKI7BhcKv8jHTm2dAjk+DnIrmxPiayVrIrua0sZv9k08CN65dVVyLH8rvXvQTidtKZRjIM
CD1DKq72euZj5gea/GgAvdQ9mAqyuFuWfJ0Pf9cKCmlBNyxw4sY0JjRuDwfnv1edhpc22woeCJmt
CZfDr0BY2MPKIpxs75EDF4E047iMNGehaHgpHR0f5zFZPaQwdO+8NkrcTAmNGeCz7qVsp96ltGrx
y/1+FZDnd2u3+muisXkAfkkUQQ4ivr9BYt9597eGrzu1bA0yMh6Da3/T/nvofBfeGkEcavr5lsGw
w0XUZmTusHWj9DBpjgMfdRk922BaiYGhamqZ2n5jXX8QaSbH5UQrQPeFObhQ+ouQ5cT0068wAuU4
2Rzf72ZlDCCRzkwrv1lCFbdiXEeRseKr8zxmLCJOGAKE7oAgFT/TBGVfRd/XBb0CeVI9BkWHvHGl
tqTFWdiQ3BAMZSue4H0nsLjuCX508eGbLTrDyffnP3yC4jj29aOn5d49JW4/UlXHMz0H4NCv9hSd
SZQbm5taJ+GpbQPFy62Gb22ITBGbnu+lgrOAxoREz6eWHioaMBAIx7JDKJq+4jyQxZdYnBjFOw93
Wb/k+fdreefG3YNLKj6zDTI3JFkWyFBE+fgvBDy2MCShkmcj7P/FYkrXVqv1KmUf0ifx8fyBAqc7
fCiztDww8gnD8TamLJ/Gc0ZPaGQ7Xdibq0bgzwetNG4/Q4XIEEOtXl8GEAua5i1LwlML7Ygd32UM
99FXrrgIkZT7aTuXDADTSooXpSdi157nyq+cr5obd1P0+UVQkj4y0wyjc93bzT6jxBtXmFVi3OLF
P2VEPd8nOSUoHwGuJjB1pfyVZY9kOB1gRieJgZP1AxOOumXtg+BgjVdx54i9YM/NCcGLHiVxhSXe
CCKRcHqGvnG9ON9riqtZmPVYmUxcqr3puAaCwZtJqSXp9GknxwrKm2iVDATNjA3TXh+IfOeZ/Wof
lgvY7/ZP6TCS1C4huLyMItztqc1hJjP/4naxRVtU6wLtN0QnVTAfjlxfXbIVEF4qzovzkmDf7jGx
Rw3O2tzGTfJ2rWvQyZLuq2wjSdLVhXZ1tQ+frXhIvZ3MY60ZcQMmS0bumTJ5QGHy9oD/ueE35uDV
u59XdD/ubzSWVPrHiRWktQM50t0ShOuTkTZ5cPOPFp3to7a1J/SX8BXhOvNn8+qR34x5NYBFTLHH
y0HwteHhJ6W6d6Z7SVQmO5a/YvsylQuXQG2F64up83A14mHqV2XteEz4T+7h5wsrSLL/Vs1DeyY1
cp+Rl9RyiwwHaLdEioJs3qsCGu7EcZtax+QF5H4hkrapYJnxuBWnyRSa28GeddsXeOPpQ0me/F58
NceoPl8ULR+LcFXx/qwHgfcREkm+Fia7Cj5OiStC0oPsiBghnEy+gqdo5Sb5Xj63mKIHTBKhCc2J
lljOTKQHcYUYZPt91wbDiYTlv2b2XOrJvI3V+zvmqlfBnl42W2PZD3J5lD+iE/mmxkOj3ubm/Xg+
vX4AhnIgnNqAGKQkTkJ/e33d7HZZjm0Ikx0YVg5qI828biSzoYoaNihTVVWeSKH8tJtpE4bZZq8K
epHpHVSv+TFwfbJoyBDdmgabyQ8MyhOxnfBeLZhfNpJUEMN+8wsDXdMnUihibNp2Rfovb8c+PtFV
52uvomb/Tu64KETkyaFFUtz7D19ib2+e2XkmK5uoAjDjsfl7PcAi6FHhl5l1YZN9uFGgD8Lfq8Yh
2KUddSOKpozmjP7wNcg+MdggQlUKozxAU/vWpVJUvh4IEm68oXhtPdyu7nd/0DnUdCDjua6yV5m/
41UNGH197+IgsauEOgJEV26JWpeo1YrEnRa8O6MyJqmVBYxW3aFZBTTTR3LkuWbHVbVfVbtHIhiO
K+2cpQuoxhuev+UCvU2AxJz6cCwKJL7AesIeyS2OSnsh6TSYA/xOXtUB6oxdOEvX+BZQzWW5rxMD
bUsL/pwfBB1rmOsIQbuUjpbTPoJBC2GxprPCSEvYNSWR1bWjJqkMLliMgRf0fquyjB4RmAyNcHMV
j1Kgs8ynHJG4O3IGH8AMUb5o5cnObyiYHqHD+wZhIjDC/00/EW8ibBpkbN9saS4QabZx5ri1kzoo
Ide1Sx5C9HpleVM3l1rXJTjuWp195vreXUC6sovaEQVDLNS9bnUW+rnVeHJPrX+I8h4LIHf65FZv
URYAaG0l6hhKWbmcsax5z57BETWfaEPVlbkrMOdzp5E9Ac5xKODhyMaUK93DYgA6yN6Pn5nBzOL6
LTZFxN5D1evoEcTpSY2zLq6tVRU74T1iM/h/oBuDMndgB4ybJPouSBoca7KuFXgiM65rQj1dEsgZ
RUbMdNf4hqo9QhbW9whiHjE0x9e1n/6qhvlPXIWT+vqkd+79zp2GFcUldFkN255TmjuNeb01CFZX
D983nRIENkjuY9Z1p6j17ytJhd2q6k107de5xViHbhl20doEQLLj0TvjZtXHxlKnEdGbNET61ARs
0g+kXIRieZ/AFDrDR3/D78rxb/g16g0yuhPIwvHoFKGziZnHZ34YGXn8ZMr+mOUmVQkEzI/f504X
TMAq7chVLkS69rfBjWdUMNZJ1mDzIOq5Rta68eeb9fAVizmAkNO+ZL2A6G4kKm34bFOxvrTOT3oi
Ydk3uUFwY86JmwkQMCKsO+vIgtIkEesx1sHzpqnrRtQmi07vi/WmgwguEEz1nULEF0un85/EZlxm
SfAnbKDl3KD5KKQmoJfdv4k8QU9uq1L8kadcwQd7bZly2/T6COsThdoKCdK0K1nFxXK1tM7Strfa
zgjQ+MhGK1GXWcRJpXpFVzyS9HYwoeg0aC8QoNm07k4lIaJcFflKx0FkcJk455CCCf/ePP0xjkEh
FgUW9VezzWJB8wfJg4wn1dOacjXwOQIr9a0q0ueN451he0AnraSaf0tEPMl3YJab3B9eotU82ahV
Qmqg8Wtfu84yrvBwtMx9Fe/kboernPTD3V0hQf8XEezUT4ocf9SqAqBvYPer8YoTeK232778NtDo
Ll0Lxl1nNvxaGNK77CijVe9MMdrZbGGeHqC2Kx2kbEGRUgh/YCUUkvm8YmjC20IGrgwB+xda4hEx
KmFXPBp0TsMoem+0wC3OKlEeAHx4EgcEAUaVfS80TQpXimFPIDYUEzQq1KNvxMs/0HfKu8A96aIe
KIGBRg7tOvwNPwYeuq8wj6igPW4PRS2e4BJS0K0Woj8bM+0DHcffzgiuerqSOB+okzukwi5E6/bo
ODswMEWIFhiIoZgo0KBHmzoA1l5MmpBRleyu377x7apNsUnEWEKmGU43kI6vor2X9XLFcrvZ00xF
IrK0R6RbmXgf9r8PR8vRMGZ5NN+Bag7FB9DEv5DjSs3q8A0fXzv9+yvN5q1otr3M3sfKbKMHEXqP
VwQ6RDd7cW1n/cnDuZBtE6FjqIhusAq4hYTJKTuHVwBRtVblWCdjC0/yLwY6B++EGnFAlK0yAX3W
mEJZzM882P+zvfM4xxsD1M1OENkFH+mhFlW4A20OfFbT7HAPLvTbkPsjV2qz9ABOiDhnM40lSBFT
7MamXu5EtMh3YcepXQyXFQcor8NGtHhO5l0V7wGxpw4teL0VGquxsWeuijXsLHjcf3S9pXR/rCkJ
RF94OWJMQmY+kmqyGEEUFJQxr5SBtqGw2p7c3RLH+Q8gb9yp33WQF7T5gj8tMgucAIElvOP02LI3
NmDmToCAVIglxXZeCoxj2yrwIvTEP1PuW8Lfcoy9FsxDhsUKNDY3Rc7Yt/5P5z1v0aFvtTzj2sc9
BVEhCvFeikGnU3thGWq1UJDFWMKKpv2Tx/reJc24DHATg8Hjvwxcm8YIUZpQxO/2WEBtcph3L4Xw
fs+wRsjhDH4haw8fWARzn3hi6TQlUEoUgiFnPfw2SHkotqzcxhrpJ421OQVXMJ9U7gwYC6NoBjgl
nj7c13JifdvVHQ2q/25cq6Fw0TC9OBljNml+l7mNiWxRHJWIXxBHp11RiOOE959XDnhLURsVY3K6
qhFlKP7QkOm5t1gUE/xRCDi3vloXeacsXcp8/4j3GEGqasH6iPLmPfaHKVyPWYsQyNhl94lIYT/l
PYBpUxYkBYDZvw3lGxQETrZUoepNljha4ym7hqAirpphZq3dq1rMebnhgonkjmpYFU0SOdlVyLLN
M+Z3jYPHYoH/wbsTbQ9/17XI/tHcoKxMb7/qr4u9wwvXNzqhUq+oz81RJWx/8bVOJHK7szTSkwXH
VYF6B+mgq0Tvv5QscYhyGTaLEuRiGF4+tdBJOxcrOxXJ0N8ygexfBaJCg+he07KXBlMSpi0nyeoi
uzQSRJToj0A5K2MrYu3MlbqbU8fQDv/Fw2Raw+z8UjUiZ1Cz+tCMP5DJH4YXXIBasg0Tg37YvE2Y
hkohkYdtBgOxRJIHRoce7ZfMp+UMULjo+gd0twd5jkwJxFxHfjlCDnzwSMr9VCYeBmOSiDJhVnWJ
QkCfTD94aTAaPvKYRwqrCvJ9P3Ay5wYvLQ8U2HiSvpm02pL2UTdBu3bBdD2UtFxWnEXL7n05BG7F
w5Z23ANgvFqJ4rrl4iB3WCbeit0OcQGOWev4A4WlBdmDmc89Hx2rvXjAubC/NiiSGvuvx7Vtb5G0
E9Ewrczy0OVvygDz2ZAsDK/NFvf8/wdsX6KMQ2KT45enc81nlRz/PRN26wOK0HgROf4yTI9TIviY
RjhCKaNqLza4DHULBGlYh7sJIDnxDIUp5HAQTdryaTAuLHakFq6Q7icIvqdJizJhcQKFSl+3tjbb
7Cdnw3NSJF84vn7IYIAEQh/R5RlIxCo2qCy2TlHH3/qlr3ynssSowk9l0UI6FlvU0z5nx6qBq05i
+Sj8POmBECR5wE8glnsfO7iGyK6YZD7yM/hbFHul+T8eWdScBUoSlhUe4/PyR+vLhS7NFfFoLEQ2
AKPyTSvatXTYZzqQFrd7OTwulKhEeDf/gWSkUWYWQOZO9t4SBE05Tcf+wyO/WsvDXbnDfshkiULR
AqzhpPbTYjXdLB34YZ2XwTlpewWwY4YjjZuESscpP8ca2Opa2ykWH/jGZ4UGNu7XAtugJ0EZa6EG
rKQ47q6q6C7TWNlKulug26VvGRpz+ZFGZcjbqtdLaWHzBcxCOf59e0poh/9+iDA3gVdVG/SdNzQH
QZzSUzbcAXZK+E8+g1QnvkZ2fA+jkADBtaiHNCKsEb+NQ8yOGhgOisZUmdCj3I3KRNvVg6JyEE2x
GB9rF+luwUSAN8IMrPiLpSNqjIX1k7b8tiZHdQpXIDyS/XDZ7TvNgs8gKl7a4aksAXW2OSo23s0i
34FKj7SNwtraAfqk6F6bIB1vsvuAQen/TpEK5E2wadoZiDwBXo9w79HgP2eR9DA4wUDXKe+lbXIv
dZnfBkgU3CJlWg+s/pmDrAllmNPj0itHB8Sptl6cPit+qwmJ8lGgSEdMSPVUI6FUsAVFoTMZM13H
UlAPzC7xfkeL6D1+Usw0xQxVCrXudL+YTXMLD9p6oIwHtO93WtInn1snG8v2UZPQEOjWXAGJCJEq
Of6VAy4gRgut1ttejtGrmERbPMwD6YWQ0FEe+GwtDbiAZUnkS0kTfBYZjl1INir0hlwO5oGUW/Pw
FiWvTgDdR8EWeXp2+SkWnUdmCSCxHTwLZZBjJzit5Km6xexW0kfHSFB3CXmnSRzh0Bwx2nBiDfBL
HqiW2G0tfYlW7T+NoHWnUUFKLAjOI26MQ4hRNVvrhcThdNIaM50OZFr29FdvTGUyZxCsFWc2BuWk
YL/FOv1iwcPpXT3EikB5jiH48i5xFHCLntAYM0vyt3fja1RfzYxOrT+03LGHBP/clKngTAKbU2mb
EFXhuTsU1Y2KdiciC3CdnktzU44mO+NS2xl16eTOyGCHk6vLVekpyzoFv4tYrTrAoT2D3lXsyFl2
ziXCRGiKRlZzR9x/utqBJMOpReZthZYytfFRsQkNFHGkqbDCcie5wyeEz3BWZUcDcn4hDN1gMZ04
ol2G5D/MuQyE4uJyy0t+50HX0N98IzyB0aLQUmBjDEZAzmIfMku3KR/lBAGHnWCeRFSVKOocQgpp
0QqbkJDA0v5PG5xqG8pKOPGGfoL45QUmzZBHcsBiPKl25gLJ7k8aSc/rLHz9TWnXpRpPXGVm8uKy
VYRWDN3IDty483M+S8UhikyRHC4uvdFZpp6g+eTLM+WjBOqa+64X1W8TOwT8pNG3P/3KF+zPYuZa
WZK0jcVW+KWPphoZdAWQrGV8po73SVut8Aflkh8VhZjEyNJ5wBN6Tns+cY6Z6cWgjvZhBiqcVeCk
WppdzgSvziU6y9vJAqKC1pSf2WEVT7Z4kY60Ou03EdVlQWAGIqapMjH7McETEsDxu2nM/tnwVWBX
ny+xpMCEHWOosA99aKUEFTdMz3f7MWaLLffrceZAqkCz0pxS9blYFXvY5e/T90o6a245+w8inYi4
q/wqFZyQ7jAHjyZjjp8x8ZUUzgI+s50SG1bze3487Qf4jAsvYyRnlbP587vfWsbiqpyGA8OcX0Vk
Mz2adRC0WKdEhQrM2Nlk10MNSMa5GVxBhkgN0h/mdYhqSrDMWrYdYrgp1jNYKulZxNHRpKZVnugN
WFsGqUjcxl6Omhxjv70i8X+8KmVpDTJFLoV8AFbsylAiMcOadr6GEBb21rOPs6M8b4rgh6aLEDxf
3o17GGs/tpekFF5kz5uXzl5Uhc98h7IPPTYpqV3L8AqxfC3j8iz2vfeEaTMt2CIBccbitHmFIWE6
Pfydm/DBmhTxF3eoX2aEZ07MYP3FEcJ9S9KWI0lxSw2tdvJTyDtiNwN5++fVI/2r8be98j7T65jI
DfVEgDUmxU2jJCTumiLJTkY2qcTwH9nXRbco2pfYqPz/l5mlElC+3skW7AL3J4wys163l1mJ+57K
YKQ0BSavZqkZoBan5YuAQAOOAEIxGeqDX4mwgL51cPI/TJLOVVQU1UNK3nmHjP3jz1ts3F5fWvjH
gmHjT6M8utP8OwFcKkznzQGEzzLRNtet1AvSzJMMRP2xiYRXxCdENEvg4o3Q0pIe8cEeF4G4Ilci
fApwyQvvgUau3h2lsC+L0iiFP8bT8t/xNqbG9yHTupSvvnCkjIgRJM1fdZRqTbmawGwqPsWLci8z
RY4gH5loR/FZ/otawNrs5qcA6rQY/qJUcw7ny15yCDaWDMDRJuhLiBpvXnOP8W9fv/le6GdxMAYV
cHySP4jmWh2xE6uLgFHDmo9CzC9m5ldodXmNn0pRbVchZCtN3Wz3wSpjcIqQ8zopDZ8sldtP9cNA
1rfv53X1KQzgfJ22R9ctrC627Fa9a/CXFUcWYJQlaWYqIH/8K+DZ8ZEPefC9s4fgw9k7JnrJW+nC
TG+A2OOBWIKHOop6xslf52wMT89x0mZyl2PwENi7trmI9y6MGgoy7ZovCvMvrcO2mDUuNlrmy/Zr
VaDKnV+Qp0kwpumeunu4lqEU8dxdRtdw/42BtSosR9DwZlLCS76i/A2g+Oga84MbF2v7UjdBmpwo
/rs16NdpZmfGtoIhzxKQIqq/EzsBKBUtclHa22TXKJ/aE7pGyj079Xw4KfYkSwJc0LpH2EmEv1ou
K+6CpohrqlOtYkCt6W7Tdsgf7yPn1CIO6QgAXRx+Yg/S6l30EFUK0rf+ugHIQIYwKlZgKRDuz2o0
955TSOYjwvj/8gLFXmeWos4Gq5RzCaltief0HdCPWce/4tJ6P3MwNTcxJu9LKQIiR7Id1IDsNs5D
/VhA+5D7G7OYee77CwSJTBMOacbiSUsXxmjY2ev/8H1MtZIEdvRnj5AphQsTSj1YrChb+63MQaaA
Fgxuk2pTrcNGXD55lfVRoOchOeP+ozAcPMBVhuU3K/0IZG10IISIiunPTvb1UPKMfni76DJer73T
xa9xWxA0V7tzCqTN1LJfHbpifASaGpVCRYXEJ4e+flus2w3ZEzialbVQIoanQ0RAaKxMX+/PZFUs
IVRXfD01heiQ1cpmyCYQf6zdESs2CI8fom1siPLrZy02BCOBsj8ndQnzIDqxW2lwYGDjgsin2LfR
YFWuYvncFzDADXEbtuPg4NUwSQ+KvEzSgE2fKEZyFLrpr44a+sy2e9Qgs8wptDM860kLE5v1uxY1
SL8Td17mNtG8/hUss8pQGFwGngzEcflRqpq5RgSo5xaA5ulvXoIMTIfaldGfZusOLdzEjndgQCjT
aWiYK3AAGfSorRAGmQEdIWZ/2U2JO/neLYIGs3dq/N0YwhiRcvDyH5LPO8Q4GDCrQrm5cmT3qONq
+8P+d5mRuFr/e8LS0HTqyqCm3bOwL4B/uImNcYwvuWP4hiQn/TF1/isbnD9VID2ERf/R47xR7Ex/
1iaXf89o5oh/hzSDlIfjxs6dt7T8RPEDgeeOv1+nA0HRfiVQotZxGcMNWoHPlhoyudUxiKursYPk
d/kq8WoicC3sjJiWEIIHH31J6nsVpVmaa1jRA+vo9saXWxmjtUJNgTWN1fDszpnuE1w3+RjpQTho
7o2Bx1DSoZO90kFk01GLBumBacQ2oVYPNm47b/m3FD6fCYLGSu1yMD7Yxw9P8hSMwcpwXT+0yR8n
iAtAbLA1k2ygk33i7PjMadQfZ4KtEov08ntp6aTPiaGyLnCb3R9dsk+LAmor4snM//yvmv+H1TvF
D9I22tJsQPS7GfKDeua4hyvlgMVHMXJkeUSsMV9y08WdBqXUC5vverTONf3Ta00dGAy64DPekt2m
gtH1DXRYpnBwXJKpQiqhcyHK/Ca9ye3mtV/yvQNhYERY2Z0hNkB1qBxwWhrCqS8N3fq7wWPdi4nP
fYfMZjTY7fR0Q7PDnm8z8cPn/P3colhuyfYKQGFSawRdCrtzc6EXfOT/Scf+E1bjFd73DEOZ1a99
recRg7dkiUis6XmADScKnxFZ4/FQ8813c9DdyEowAmNE0TBr5TM2Xk8/lEybyKhwS+EGcVncbnfi
PCvkltLPwpOkdzVmasf9sIkXdiE9XZty9Ou6d9MOiE9wbLer1F9HvINjjLZxf92jPPvMzx5F1oxE
YsMlyUyZT1dgx8cenSKw9hHTy6osAhQap1SA9ddA3ofYdvWiuXwHFqWtj3xBHTh6lHchY82/b20F
popLjarVdp+MW4OI0sevdFmiga+YOD2BZaQJKiIv/Lg0jSGp8PzDVXeE5T5yro7/UzAVS/bo2vib
tHEKvcTgJ5k7AW/Ttjx9w1Bi4Plrq0hd6B9qCp9MBsdzzL/rIjYysak/8fdkiZwynnhseKaBKpRc
RZ2cMOU5GyPIxGdmwLi8tY0a/LqTI5Ta7YesGAIzxaKTAN0OcA5UWydVOZb9J/lLzFgU/T4wTD+2
nOxKkVJYUbz5P/ZYGgG25IMvFAOrZeQT7Tymfzzk3J1wqbCccblfHBEk9k3TKa6rJl3PS45fq+ud
5R9K5WbipS3eKH1rlMeoQnC4JVYSj7sEJ4tn5QrgngiUnf6lVyofRO2aBDRv9A670aZuan3AS/i4
J6KyuhI2SiS9pKjAm8m/gmC14t0ywOdlQ12ZoGP1BMjhPjY1tForbQnigA1PWCiAjuYOjr8T/VCL
Mw+YUM3VZkZMiltokhAVVSjTUDep1Lo6yUr3gB8VFDzONGsFyoOkcyI1khPN8AGdDO+mg/Rg+cK1
6h4C/DUXT+RWO21pLBdW7IHYphSWJSJsf6TGO+LXfx00J/n+RPcb/ejhhamuUJx1ZzvxzqJQDYag
bVQRREj+IJA9PCynmAfecKF2oX+o3VOOkeRXYZ8URFAKIOddD8TmdNK3juvYKKn8+iJWVsg53NFu
OSvVWL6HfzGxSdlkV9UEwA2tOsd0ZJQYkULuL6puu+n/+BFtuDLWtNDjApC9h5gRZgMsPJBFt1M8
MRgnUhUSpc9scyudO7iSwSc1+FvbfYntHd8sgXDoAIWPyqMvjPWw1ZvivjO5YJJYyH74hGlBThkf
ZRlJmMYy4LmKmy2/6XsBtoPWk8R8rkEgzNVdu7tXL4yEYQtcK4zou+y8/7MrBvoppwnoAuF9L4Ga
3aRnzR3HklhlEVZPzNU4UcFoa0gjh7aagrAw8TcJPNf+YSLW8YHuvKtw2L6jo1c6rTo3TvkMIJbp
3QkGXSpZY8QHXOfcFT5hw3JG8dQuNcPx1r71vMMLCJzbkHLz4PcH/bc8LWxKMNMk3ind2CiQjQoG
yXmgljR5oTFrVENRd6WaqnT1XAt/t3o4iGnscuxcGM/3bxNWiMWEn8DXdLdfxowhxvy287X1L69k
Je8tzBVzaonQ5DjM2QF/kGfFrMjmLA/xKq24PMIU1RFw4egRGlsXcub5fSVMYCQuasZZFM/NFBhf
tdCbdgkA6LqY4ouQxnY0ST/2IsFG3s/QAttq5NJ7qJSEPd4rLjxoTrUXi/63aJRG+AhxqTd9qQ3w
yMRjyH7v+wd4mz20/yA2kM+JgIY3X9hoY1+O8xig7zHi7xYhiZXq70u0HOwfQNjcM4uJsQNz0Z8l
kdXLCNQdtSO+fTr1i8JjKZ5UUywkxnRzcbZeVb0MGKj6LJb9BZIUPN+7xXeItpmOy+lue5+eNCZ1
EwYS23WqDvoZ0iend2zC16gY7AWeDk9ZiXziKX7NFTpZzvangH6OPIAWG99HtjScsY6RaIfJSNWl
Au5UBDbzOxU9IK0kmXDCnTPSz5+LFsBr9e7Oei55+EsUBS3d7VcYwCaaAxM2v/WNFT2sX8kGU0aJ
I7CrMT6FBF/LilP11TJZ487/MwssFDeab710OCSSF1NlSDjEiQz3XndyqkdCO958uEHLyoD+iLwp
boN3N9xLYLNP6VfWJUHUI76MTzkNhsPm/Q0I1Ida45VHAAIV3PPVl3CzHBDj5SNMjRaRPq8Wo7VI
X3swJQQ2itIvHDYEF7ovzlK0VKlkC5jlxHSacBKf9wpZVv0QKpcxLd9BAJKhrc+Q2SA2OyN/OLY/
iGjiRqMiH7Pup8kswycIzu3McI3WZpkPAwXc+AfikG2P4851OdZJyBAgzTl1pCa63z+9zUCe2O1K
NZ5jAf4sSwR3DgtsqrQypSiR8OfZfYxJyPA4Vo9tRPLh+8dXMniapX1bfme1Y/suBCwDFiT/nVTW
YFx3meA1T9IFs38HI5KHnQ8pmi87AqaB/wPewyQxMyhz3Of5oFkeUUNBbs7MCJFxMp576xN3MEMU
hM8OFoiYBIlKLAee55avihE8e6qWFzy2/QijA+SPZ+IGD0cBlqIuu+bKrguJ6Da5AVMk4L+5UpW3
7X9pssXr1QkbazgYemnSgBPXqF4Ht5kSlkXJoilNYmde7IufXIyAbUPCxCZFfUp2/eRLGcOs3L6P
5j/XIMJ3LDk6K8o2QEzDpWXGUq8ftUloOtIAb/JW64dvQ1MWTEu7zSE0aP82KmTuN0AdcgDzY2TE
bFk+eEciKrXBmM56INRrvRPGhdpkikISdqOE3sGlHjRsAy25VK2OXZWjfTyT4AsOZYkGitiHeA5l
tgCcpRspXfncV4cfgQM4LPKeJebwglvwt9BP3iJqAygmF+SYMylf0+GoQ8CYbr0soZHRYFE8p1g2
Vbo1v5y/117JVb6sRR3EVBZyfX5KPfNnCGafPGuH8OW+EUUlvJma9bmr6nUM+y1h5R3harSVNSV1
6VgU+LoizWCNCgnP1TJ951JvEnvEUbEq/hu8DrIk70bIT/K0AiQrySJQPTaPnC6LCf7agqyMvLHB
0PuzDtYdTH6MPi47C5cjFtaLNcsRuHzVSvl+63Jwoz4o4r5RQ2TI4FWgu6DdQjSAxdKfhMYJDTrp
PUFdtZlpqbpWZNOAKd60df83WosyVecbrYdHv7StstjLT1nNXZS9rOwNEyTTQCZ9fIVJYSUh6mvf
7nWi8ZhOQVHmyTnC+L/+UdWTQMKAiPDQZKgMLAuJrssM8wBs5G5ig++9lu8iDgrKirueIMIq+XJC
0K8D6FRjf4shkGBtt06t5e/urSxGYUIsh339NfSrLu1g121DWEkPpBqKqmjlIT2FIP2k6h/P6Vyg
Z/YG+lnUNs0AUQJfOJCv/e82h2MqYMrUY+dJvvqswEGNBeW2+dI9gpqHT4Gqi+4hd882Tr9SUdwj
Nm8zJKQ+Lxa9jNKo2lRMs5RO/OUMrXTpPqt54La3dN05sYVBo2sbypNEiCq5yunkT5pZCxWK8rUj
EaOGizJuut7+udrBp55wwAkdggyOnjup2s50/ia+zssXnh5brBtW4jrL36q/VeadZm7YZeIuW5JU
H2O0UI4XxxONsJ2Bfzqr5u/dnqLJw0NcrVGO7SoiXd+LQP3E3JISABE8tTGBR7ezld17Nqq3a0PQ
NwdROc3i60nVLVTYpUHy6EyoArx1ni+jmP6H1g/EAeQLqFiOFel+dI1VUnhN5wTkyBEN30/QDkzl
RpyN04gbp2Hzi76cxlptHPYQT55F0g7VdT80jwbL+2wUXH6BY+eGNwDu46e9fVzoYUzuFR4cSHK4
CEYQTUVisHWwFXGkDieh59e2mbRWvZOA3hXTq5wTdTBvRhFiqRV0JNwi+w8HVQXnSblN2bHeksss
fgS29i0+hxOzAArar2cPfQ9DdZ6ntPQljBnt6UcKwdTjy/EPTGFoNYFbqUtH4z9bEDyujWZTTId0
sS/Si+iY7FAdI/vKgNhESNfZPYGlqx1CyflkHrNHlXV/PynLcFUIQH2nzpKhU9A9QYFDRgBtZTfA
RcaOhfX2Ae/ylfdpg9W3ZlqvawQM1MgIBDjSuV3yzaJPb4fWlDZlLwHR369YWP0wtF9OUG/M+lLi
NAmO3hOw5atCXmTw2lsoVrs0/i3Hf+j6mqWAeCVhU+vsnEdZ6zAoYSEddCNqa2Lnl1J8AAIScS0c
LPzwqNVyk6nXXI0SrheC/CoRUfdNNJqK6MEv1wbD5ax6f24XxYh21mNj3eHen7fsWNOdMgNOnnJW
WzeMxKrDQlW+JM/BIsWJX8Xl64InivijPe01JMqchU0Z27ZfzOVRnGGx5t79ids/YQm3RTTcxYQH
ywSNKAe1Go7WHz8j0ujI2oceq1qhXvJVMERjb/9UwmQKrLQmEDQ4Z26Ofe1k8BaZT6Kou3JhGpXw
T/WhRehbk2wKkOiKZzGAmjF2EUrye2GtJPjbByWuRsf2PSffc6+MvsS8110cxvqIei6tOowxSgZJ
ahok4xReC+0Qanys2TdreF0awHzz40iUuMC66xIwmoGa+badMuaTVInJbqQl5n2gW2OTAlvI6u5c
R4E7HAABMVjwQk4rqeoail6ZwDs+Vvudk90OzlRT1u6JGc53/SPwGrKWVTlZd9GfT8sKXmEHu32b
Sv8LjGSi8WkPLy0iTX7yqRoPZf1KKkYCNKHyCdZz+6yc5GpBqI+Gvh0AmVNmmP570oYIwky9TpDR
KE1lBMpqMHkDSu6NKP1gsU0Z3hvHMOYoeP2Ryxklr19dwU6j9/B9iDZa/pl6nPEddSVodLrDxJ40
kspDhVLjto2pzLN99V2o+CcIWwmMwHjHp+RbPdUaWgeA2rUEz2sjSPEgmPtm1niUQhfslSH6WL0R
thsqKZuRbS4Qf5+oMOfT42/F/sTrULketkGR8a2tOBNglN62kL7z1k5qvflPWsX2Sqdj01sO4FGn
DcXP1toeKQ8+V6cXwM6+qzw9q7J62aDdu1TTAnky+TY7HjGP7vfu+m57Zj8yD+uVJFoIw9YYVLBP
4IB/hWrt1sFgy85jH7tFrYitj/jzevEQOjGpyMrmpx8TZxgnddP1P4uY2tkyhytBpkNQnuAMMmTE
KjB54OGzrMKYie3RnMfrWyvQH7acAGf8lZGxhx024akBkK/OdFZ91h6Haw8Zea+bfU640oRjXU8G
0KBCNz3XGsSDq0fS58eu1iPBGjAbIUhHDNmbtky8Wu7X68C/JvoodYyUhNkr9fk/XII4tvVh4NzX
We/f+27T1Agurjk2FJLL30M6kKsSU2EtsLlFfw2eTJ5t0KzWOkqe++154HwXp7ZuqTV+PWhLbLBy
42414mnTRR42OOdY7uyJOyAwyirO9T75Z3LCIeY6qCku9CbJwUx4NHiaMrT7Of/nHrjOtqXiv87d
enpYy/EqIJUBLWsx9X9uF1LHo9OdPF4kRbjUgzjEr7sc05zNvlPPCt4aRNFCVgdg2uu4Ci+tEnVw
0EZ7R/xGAnFDrWbiGQsHd8h4LAXL8iFNRyQAyHfatClgAZmeliI4GtpE65QenQFbc+hAISuunzca
JqVvaXKM858F43xt9+DJ3u2+7FjTo+nXF9olkL2xuFJqOKPATfwWU9CvcIp1Nt8DwfiPVTHa+5N2
dV6mzEYYMWCBn+wVRbm1uZh1KGfMxF+zgjbLazhQXhp1LlhVtUI/oVvmFUv3UazFjBG8ZVBHvH3o
MP5Wcw6K0SpA4UZoHOvOGc3Iq8ng/BSda5ZgNxciaelOklrtVwOqC+0JOm7CXXqI2B9PUDrbBd4D
rblnWUU21GjC79BbOOybeshEk/2+g4HJm4XxXCH5/9sqVI7UPT2Uz9w+TfDdFLoKMbPxfkoPzTR4
tUcQYRqsIVX49ZBqFJfP/OZgavExkMDC1Zwj0z6I2dj79P0AtMCrG8W4q0gLUJYRkRd40Ek4aOtw
C2shRYZ1UDQu/dKpVUAhmEEsK8S3ZAumeiAD0kzIsAFuxTWn2h9A4JGxv+oRF9ST2YoMN2NH+dka
JLl8+4+SWCZ/fhi/EMomn50uifEahqgXddAwpqJkahni06LLeHHFNK0DHBR+096W2qskGw9bwNBe
+3v8fWM8CpAC1/tXqvgwOToe/7lZsa6jcbkvQgD33hctoOHEPSXFpKsSrPou+wOyWezmkvJ8s5gw
ndjXDwxAvOQJ8gfC/q0o9k0lPOY3ikELio8WWq/JSkS87c1AkRkpQ0E45wbhGu97AkE8smDT9eh4
9eg4SaCvYygMhfiZxP77y43nQvN83WY06rCi+EQ8nJWrKk9rYpcRzQhmkniYp6wUNLyoOGuVk7VQ
Nb3wXMP7FEn9Zi4UhU5Bp3K3RqUZdL7BMarbu2A3Ol/5erewJ2WR+2jGXoJWqiY/cljwEWPyV2WF
qRGH8XVDBN7t1izNuiKijIe9bIqLKC3qXjqU7EPvp/4j5oXVV2XDSh9Ehu0/YfNDTlJmmOrGwlvu
7nzfgRWh6T9PJyOoKUTUoWS5I5gdL4DEBHJAg5yuI2L9R6YRFMHHU9Pu+Zvi82lz+Z/V3Dd/lgxT
zJATtGsXIqDU4ICQuROemRyyTMQ/xUtZ2iXifp8C42hKw05WF49Uz7UpM5SLMWs9VFoYVka6vgj8
GK7Yz9pvmqtpn3I63Y/OJ1m2NikKAhfVgN2U4wK9ya4phSKPm7Vp9diXhuGJZMWW/kDC6SLF0QV4
CwE87f/ypzGFOqBQwq/CsBRvko/z2WRtknWvmx1yipXtSPH9hzx9RQs5WmFRM0eJTs+1wrDlDfuY
spCiUZ9Rou2rMTQheosmM7Ok3ynNh1meKCI2P58y0tBLTZLRFxmZnAIbc00gW4Jyjej71QVlgj+Q
tCxrGObvIcFAhY5UfLKZ5/9PUTrPOx3zQaQQkxTsw3oPolnIHtkGBLq18+VOugb5vkulI5xxUAPQ
TZjeOKGjAzcSmLZQ5W5NtoIuYaNwCdMwykfCQuF68ExgIN5MuPH7agHG9D9ORkhLp8Uaf1fmrvOE
Abjqlj9aNC3YCHMyXbEFfaTjm9y9aeP03Iy0Syo4tkIEzNm/PlryPkVbuVNJsZTVE2wsLoY1JiUm
MGbpymGjuqPVYHdAkY4ejnFBBnzb//8P/H75NsUCV9L37zE0vVRjLFEr3dfunNnzpY9p/vD+5+8k
Hs1fl5fEMI57qLuYTogikRUwb6ddQWhP/8CwZXxiwCZDJlEh1KC4pHI7+SncIJW15Sy+cy+G6wUm
cwRkUbT+vrd/fS3Uc8tuQABMk/zEb6OUG+AOC156q5N0SZOEpxi1L7hGxXfHDTzMwLKRgSWixtml
Z+FqFDmLj7D3If6uAy9WwDGpe2Ou5FO4619+JiNFtChML1Rp/j3IO1LyNnMuPdQG4WdCd+tcHgnn
/SYbIhoTNLiT3sHKSpnjNfPYZ4g1hkdN0IEo+Q0V7jVHRnGo5wCLyKd0BSL9tWX+G1RtUkzBx3fS
fsJ3UnIMvtiJxB1zO0wyUIdH2bSb9oISkSoGbU0xJ4xuJbgFzFQAV8JpSTwPalUlpwQRwEAX9SCG
d6qkibUJSl+D5CwvINR5rDy67plJzN60QrhlCzn+23gpSqgYl4CqVh68mF29KeNPT4/s8e7K5gkm
SJlOonF5GIiHzkM1cKmtlfA/hpTwzXNJ8ysiXEdXa2CBrGkLo3ZNUbG5KPv1vbYiw1iQOVB8c0Wl
2TooBP7yCwdOnm9lSjoYiRK04IRUpQAkqT2rsh+qB+FYsLlDtvUHXiEH9VMkvsRjptDreZIAp+Lo
xetXmbSYXXBHBeDRb5JmwdibKRPyufGNSA+CBt6NX3dxUSQT6v32HgEe6GlsgxK5mA9QM9Sumq1I
CrpRMvD73T0E1EKwLZivcKgBqC5vFW5mDh33EB+CkU74IqPkJa8bcE98ZC1mKmCyrNQpnARNhvyJ
vW2kVZDfGJGEx9qOfzdYLFp3fhzeoCE44WT8iddZIcV2/04oVsHRD1R2k0E/YabCmP1r1KQMWWp8
EybILZ64T7jTbzKA+0RIbUA7FgbFvmuk22eVDKMLtbnlKIUtVQiXj8oyNKj1xJz3ob1KiYErK7co
3bTt+jVd/NRpO73vXLIaFa6z2F2jrPEROlb1yABgA888MEjkmbNYLwng74PGXSqqOv4yg7bnWIzc
1z41UTBCl56xyoUpATgskK6YUroti2kf+5wpkXoWgMkAxtQN1fainqt5mgNQnhGjNgwS9uod9KWR
bzQprO/6zkTUiVKNXxKnpck8anh4Wo7dcVQwH70gODc11hPVAZSunZqNV7WSs+0BeAJy6qppaI0+
n02lWnsyorWFL0lbhYEXbsZB9P5v2QIv7sXhkqA7BzQEeEZS3mzlUPZKu4FjGnyek8uvCPH/XdZD
0O76Y1sI+HPtrbS3/w2ECdZgfprQyn619mtUhIqqzHmSEWCyeMhyZHXgSaQmkezkoKvgOZ6EwTdA
lsPyEtW9lQTz+bzK0L0Mr47CocQ/oD+jDPv4ur7s3sVL+q8zk4pnCBC3gUCUwYvOLcjKdErE1d0d
6qZbm8EFhjplzjRjK42Rlr5UZjTCE8nKHxv3LSQ1I7S4GghWKC2DKIGgHj0RshQs6pWA88gZwuhp
bw8k5phTD2LbQ5h0SUS4CnrG4ZHNI+H+8O3XVyXsw285Ojyqv85jDs/SscypsW9TBhgD9zFh7Aq/
gUwHIniSGUZ6v10CbOsDjQzbkdDEEqgRhBr1KlgyPOGyIpKh8Aa3fcUaw9aDbzpzk0jMi+AZqfdX
xhSLiVqcOffcFX+wKdqEW6o7HLUx0arA0Ykq5sGb57J8TuKK32KhMqrCChopI+gKZzq3sR9YVAbC
OtoTWwyCXx+Y7kD61Fjju2PupHCE9EchAPOUyRzpouKJXxz2VZWgdpuiLQvooTzah6cI46Pu9viV
TNp1gffypY29WvbOYXNvJ8GYJQ6IlMOjgE8YWel5WTglFytJwyZfiq8AfUtsky4PeHae+jGi+qGg
l5t3PryMMLqGnbN+c0fkZySkySo1E+Q9Nd0BspWOx53inm5odhLSjb9Gd+425/B8YrcjlHYuXCR7
UC41GpXevM7tMOxUB/P9MJvWRUDZRkMnczAQJCEoPABLW7RDOMd7V2y5DOyd1t0dIyLLKvKUWX9X
ndMz3xgely+r/lQdT+UUAKcQEMik0FvB3UW6KOqpXpy0mEoYrofLra6bBXPXbNDVN0VPMFYnlEsy
gLJL/8H6Jhu4m/hzBNaoktyRKQNIPxfTIX6Ghc2lRspMlAnVvI6Q/09QEIbjF83n/xnNLRFm+qOe
LS7pdpCXs25ndSAjptrUdWHYRg3W/Tv8cQqkv0ZOZ/tm22G64R5m2mtZrwsmVmCSPFtdUYVQ4xV9
Ypw35z4A/NMCACFpi5e9e3HhEipBaGCzw4xw0tSa55AGUDnht1cxXDtFvor72ESHxzaUhqRe2V9X
uDD4A3H6QukRnCyhpxj5oeCYOBogjJVuTIBgozs1t9I5UXDoGZt/cyr4iyY56s0gdjB8VRiwM3pG
YRjBJ/NrhYHlKkXUB+nzib+TAvZChf1eqG3BUhYl1tFnVdhi2CkQj30AvOoTRnlEH3l0NINhaRTV
mWw7BUi0cb+D/vmoRe/B/l/Iy5bAO1OdWwgYhb/TantpNgkgOLqOlneq3vhecl0yvq96DdPT4L9t
g3ev5cb0ARl+Xrfg9x7yNmhwvyZTcO2/Y0gQCE85EkZz9omG/nouyMsYahKzaTp2IQWaQftkVSvZ
G94J4k4QGG+9TacWRzuu4hIMAYtBm0a2lrp/um/TpuHIpVuScNQ8mXtO6xBNjSoIXQA2nmIPwi5X
4LLOSY+p8qe/i1PYVWTWxVGUeO4EIeo7i4+ok+XKKGxVZZFKe+nVT6mLbLHKddp6WYJJqA7T51qt
3S1bbMWueiJtRlBwrm3GzlzzFlkYNLc6i7cP7a9UaCzS7Tms6JKh6uIcsFVswkIKEplJtb1lah/I
PX2tzBw2SHa4Qf2Y5UM2DKEj99I3tfx6ooxOSrhGD6Nrzy6HJLDX7lDEMLVLfVs90OouJClJiRlP
BRmeUMipfUjqWLi0/I52aC7wZzoxw4vXKYvviGAKyrkRD6qhH1yYDn4MDP4r2x4jyfsQp5ADQmG0
UM326t7xTTw1plFitMhv7VSQwArNMwnHaBWyESfTbrOrOmDUaNKR4DQILNu5wv0349a9YI+0MXQw
0RAUIT1GXnMED4TL6hDvHR6LLZ6jHts38l0PvjRY8aapND9/YJeA4YhcSrnW4y4Inq9604v8JHLy
trADdq4vWTep4Rb/X9cz/nAETgI2KOT7QLotcz5TzO7T8RviYzw5CYHVBffRMk6vYyuCCdBHqlKG
YZ/oz9vE8iAmd+zerpwmrU9yzPpAwaX/gCidtjDqy2ForsYrK3k2ZSeGXgJ20lnBYHZOlSc6NBni
PVwwhcFo8tlnGn849PSYiU4Z6oFVAYJ5SaftBFaRctv3IPwkMTF1foMTfykbMMfeHapD9Rc3Agi3
ZX8rjm3LZGfn9UBMEQgBO0j32TdkMpiutgh3alYZBUXraq5E+jqSEj26UOUYrEc2c+2k6KGGsWdz
qZ2gWD9Q3wd3FZ6lkxsOz+hxcd4q2Uq0e1FtGWAa8juVIZqzVo/p4Qk3nbu9J8BlR065tuqz3UBO
6KpWJIt+lCiXgTTgSCjE57f4TzlSvRmuwddgVQDyzMLIKCfy1c4gFdD4234wxxkFtX6YTE+eH7It
a6WbMQs2NP7yG12MH2CEFNmS6gajxZ/wIrRTTSj8/ifVgvcaL231GtLEJAHUfks5IF8n+al4Kv1k
TL1PYKFn4QGjpjs6YwH3W8nPb/ZB+sSmFBMUL7YGfdKN3qacBlrUQWeMFv1l5r2JVWYNsQ67bho6
2H9/9tJkV9MtzYD2PyMMHOQ/HWYnGOR7Tqz2L0HSulC7rOi6LaVAqggPbKRkSlo7r2Ru+VsWWrhb
COPW2Oywq/QNJNJj2i7OWoQnj9W26SwX8+Suzw4AGJH0xfA5APh6NJiM/KF2KJ/hDoJWM+D89m1X
EzdVbhp4o7Rsdu2IxWbjVzJMU1LCbGFiC/uC7QF9b/vvksohE58we485GJRSmtXFYzT4PArS8QLM
gC2OeWm0AlAI4o1yfARxz3b8gGxx0sSamPL//SNE4FzYq7+Bvj0SFTl8ev6rdwBdk8c38fvqCkDR
yu2cVM9pOLbFx4J2OE7IU+/K42bM7gHkOKbU8q+Vnw4Znyk2ApGx5d9KeL9QW/fKu05KeYlFIiYT
DVLYLJ4TC7khB4ytJ4Bf/yyeeEmkuzFa05zWM0/xMkmgsid/ahpma0bCtmjZT9P3vqdsHqUEtAl+
BLh7AVSUR9h4lalWU2FNwfoCzKJ+UKqN0/FY4xgK7OaRxajHei72MyuAHsw02NAk2gxQp3F7u//O
txQ6yDQq05o7zxRKTXEk4G9NEYwiC2oH0u04w+qmqLnRyVFRWrX0nl4QlDe+JveDtkCk8r8s0Dcl
A6XmNUAWdKD+zGkK+0FBrFIfug1t591tszG7u+K7vdz0Mu5vq/Lc76iXLYnou93tfO6y0IQqHv0A
bvVH+ipiwWu/sMlmf1K2NP6P0dP1eWLiMW41m2f2hk1AgX5c3LxayMZffAh5IpGa0GN9tURgyjDg
HHi9rp+OVd8maDxA4FH7oy+7BTe12RETqqr+nOQdi3ArKh9fiy3UVIOhvIuhyp3lzrwJ92uIwxBT
p18Ao1209XdHQMEIkWJAoalWbYdlRHrGUwPjSJRstu2AnmNumMbK4Vgt52YSjZpSlD6f+JgAb3GZ
LhA42jq9u84iIfix4LXApS9oH224ItVZ+BNjIZKvFvOz4zHnEb9ypgtYxUY/eZKEC4pwSbi7gr5Y
ypV5CKpt5kLMQxbkaIxZmYvoMe8pXPMq7KmDkikCOkLh+9yvWYsy/V4iCQ1G8Ii7+uNu3tUyRVB8
hBfayUZ1d0dzuv3ebz26FnOFtgttIDBQFcSML0lZtc5Uw+4pnUZkubATyf3Z+0JpInQVqH1dzBSf
UNp9rT6+5zGI5nKNZdHyo/Gtu2l5dNM0GCbtgt14PmKHTuF1rXKdI9XEwN4cgEAuAJUQwM0+8vQv
DVr7wUo23i5097gpu7pPfpxL6wOrSaFY9+ZWGr81nkabM97LVkGZnMJo4MDUMm3FnpgT8lHp5i9H
/QgT+3WxrmfJlqF7cSCnQlVtRqwE/VDs9N3FNp7qHEvwc3wsjy24LSlYuMZjisLbaAPA0Df/tWc1
zapj6fLga3wbW1Qv71JrPlMC7/6g4MuudwVNy2myOnmyHZeRtOTzGNnGCbmpsftnPiy+ObneTZoe
GqW2x6TsPqZ6ew2FWxgQfiuGvGlSooRr/+1x4JwIePirz0b0j6LpcZOSmbsKw4FRq0Dm7IBHWvUO
TOzMfGiI/WLZToEa6CRPrn/kYN4w4mUSPpY/jK7+iCrVxzvOQx0GEgh+THYzjUjuD7Puwfa2Acr7
iA2CyBttvrePfhFhFUv4BJnkVCLfOFkSxHVWW12wxAd9QidxaSRIRM//V2QNX6i8/4iJzYLbP+Sx
fFI8PxCMEWcLbeEuJ3JJP9wUC61ictKqBDzi3tP+ftgxulQtTalIIJn6DbVrv2FbCqFpwYZMEVIy
bYx9ExGH63lE1C7mcfWm3fC7QjJqYvY1S3ekeIhwAtMGi1jbl71REqVz5iZHPOVugsYAhCUIZfp9
T2dkqF2MngNt5Czd+lnmPs4444o4NEz1Ls7hzrqYW6MSYCarOrdJhDCu9m5UdoSYDbyZykkwyztp
RUu+T8t0Z7AGkpUEKe7PJEcGcUKjYIJmC8emMJ2rB2vecgh1nQtAHbESGSR/JYbwxCoEAWdCFcap
3XxOgC9w2fzYddfltgKuZHCl9qcb+8SHoAzVg23Eg2xlmTfrktvo6w9Dr9xfsJaDN94l+Ap0xTiu
TPM5BbB/MAMsqpFWh/kFzE3jQNf3OwQ5+pnvWkvFSlocTWvd8RDLxSuHcJapWDkHJMQjNJ/gECg0
k6tHFjK7X0UmEHw5hU3HwCnTbbU6hm7AcX9grvzArGXZmWK+fQ1Sq0/zKw+l23PIFK9tHH9GIJAR
FK4TCwNdZQa3MsxcGv59GJdrs11iUWMssoPCoZA6rLZRlt1Q67ndhmwgiReuCVMtFgsUp/FzHx13
3fdHqnAIAOS+ksyNYNkX+o4HGBaKF73PjQCG+aTKIEbdmYnHdqwJWonOPCx/9ifXF1ASlOcInriu
EhdNkLScgNoclMBWg7p6uVsmZoGHCJPE3TPDRMgN8MelMyQJAfOV0+oB4BbZOUShS6meCvwMhi1o
3FsC9loIliGU5Utpf+DjYohmza6wxMDgHkcXzXVoZouRNznah0u6MKatHwpRW1g9m2Kv5vyPg1g6
ns3DfaK1p3I3OJieqddCQelmATDcqYusI7jEv/UdEgKYz244augP8M+cZNhuKDWfWneATRhgg0Sy
rCRW5EugINcoL8Jd6fbGDTQozyD02+4h5hDdLiVfkFZlJ9JUVguWiiiSV1VyHbC7RKoNhPom6u/x
Tvi2ALB3Pk+Jsm+qdW3H2Ao4lR+fSFSJmAyFEPy8UPefRRWK7wCtWouwFskGTg7DGz2WD1hPL0FC
cFfgvPvx4M93gc5qblYahHd/muNPMZ5Bk7oG+XNHdYV+1VI7hRexz06xtp8jUySanK7NpDxESw/7
ZIXHLHKmqlA9ARTGKbp/3Swp0Iz87AACImvLRnx2VIJG8ZoDJF3psAv5fmNwYrbe7J/K4npLqaNo
tcGuH/a+a6ZUnuO58LQi1bYzSdx5Zk3Gk/xoQmqtoryc7UQJhL6NZ9JPA2EElowmATLLG9bgHfw3
E7lvWw5IpJ3IqnPTVfKPUFBhmJra2SJqCE67BGT/rtLzjGAmKVRM1o75IBVc9dufvEPhKpYJyFQR
scvfK4a+ABXUp6t5sL2Vs7V02EMx6oXXfu2cEh/W4twyIWsUkdagp55BSwRrzZIT9aAHQQgs2R75
EdI8vhUF6IOSfIGowUJJ53YH0KJ65vTJlSFvujHVnp8Px9DgG71PoyX5im8rA+7HAilXRHFFwqRO
8TdZje5FxmNnnEE32DR1/oIhSD+BVOw66hPO0FwNGKLL3WvVD8deUi821s08EUngCyY2fiVw4Xi2
X2WnmsfuN/f1+lrkWqprtLU0VPtCRLWyV82k0i/jSR1qQcc47Dijg1x6GtrrNKNaZiQOunjKx2IE
EGSN0YVg8zhPsnAfRvVmfzWxfUfbPrNl9QFC7JLzS2uozmJRE3g1sl7M2D5FrMwvycF5zAoTJyEZ
whTM5OEPhIJCKUkvCChWKL3FI8Ew2GQfxmJ7rgvB1csg1GIc2NUfVTWIsYefWT9bkCVTIZ8Lj5G0
pq2MOw6A0V9F048TzjvIfLLg8NBdw3se+p3///MKwKUHH0LDId/KU2a4AsJad/XZ8goHNKS0BGXu
fm3oqiqdK1tceEfz/or4JoDfqFZHbM1IL1CzEqTIVpnCoQGnO0GjBZ4KPvO14vOc+AOQKSAHKCgP
VIVf5Wt1fin7Oxv3cbtInAHTnkaQpVu9BO53OTlp2cbINHpusn3RDjb31gOalQ+hkQwZD4zac+h8
pD1duyis/Xtw4TK+R1902iDgS2usob+JUqebLPtz4jOC6fFs3bxCGBFuHQySFa9+Uvw475nzHzUV
Xx2P7UFnxqBqNyfcvlJU6IFtJa5J88MFswpEYg+WieV9YO7tR+7QRyOdF6+1TBWvsVL735SJip11
3nE7SVWtr6FJDd45LKKTElC5Wa/7CzaTDKsD6eYugH7s8DHXBDDpGifUPBojJT0v5nq+K+PTHtNT
xd2eBCQ49K2JrztEiTF9rjvJPuneABm3Y1SoD2WfTwFiFVxHrlX7Q7GZ0ZZv0ofLX78W98SM8L7f
0OunSDF376Hk0lpumVoAOeDqbEIZHYqR9vG7iQaIgCVCYBUD6YsxZUg6wShJH44yFLHFl0K2G5Jg
zRMkYTE6PjLBSxo2J1aB41a96XtHJxL9UTIuQ/KpJ6or0Jep/EnBngofJl+Chgc2P6E7M4Zvjsbc
QIAsdYV9NPRp/amg3huL16qJl9+ACUzpsh/2NmzRHJiFyDqV31pW9DWM4/EC1vhBttAzxz6WZUp2
3xWOwy8Nv4r5t+c7kat2vyHx5w34N3J3F4PcfAZcUuBy/6e8X3go5ioya402Pm5qm204RcJjGbqw
JCByWA7gaOG7uVRGB1D3lUFgxmfon56WYXuf93hD9wwlDEjjBrbG6CrpPddsTs3jWwaZy4vpfL0+
Xe4NkRd9gN9heoS6JDMMH0hHB7KNEvcekVOdEH0bGSZzjNexbXCSGhKCJ1EfNz0HeFHr8zq8WHmG
EKmKvmgffQ4xIATzVBzzdyvYYDHkDHfxv3FReJgXZssj4W8x8JnYWYAYbODsPv9p6dI9m7c+x+yA
2BjtqYZS74ng5peXPGkhlexZJVF/P4eCmIAG2LmDlLV0siIXnH5Ncuna2USniJrFL/nbKhzh5irc
c/gX/pWuiDxmZcobc/TWjJdsvaS7p2keqjrd213K5qR+7HUy+w6B4neQFdi+VESTeKOM2rBSSk9y
3l8DF7cjyub8er1L6JBv/htD6gXcWCt0POvv+2KNDysalNC60DOxeSqT2bUckJee/7oIksLJ0bsV
gLjbBsWL0VJcaZSYriS3g8zRXgzquaPAODk8uDhdCeO4h/o/SlEf6EcROd1UGErtC3qkTz+JFeVK
U8n7eFXFlqbjRVEz5vbvgCwxiuqawmifcxJYkqL61AHY1bDMYfScvn3DXoQ+FHwrlZx2bE6KtyoJ
FyJGMwh8e/iVWm21jSTZr+8bS9T0mRQQXAV7Y6VcxZKrDFm/hywQ28mLPBiq1FeGONPmp6pgJ9F5
SMUNxWhuKzYrfARLiakadXHZZy5shG1ge65zoF09sAhBJ11x6A2VlHOgjRvDlTa2sn4nGABHS7SX
55A7GA3wGJi/mDoM+rE4Gx3r8JgRf8XdN5/uVlkwSF4sFtWp3gpD0AznEZz4OaT77TmQRUnXwYUh
mcigp6LhpmEHzokEGytbuBS1PDSckDxqme4WjbvQvqxU0ev+PRflqFSpP8CHf3rHRo4onfOfUeaw
4eBpzP8q0aH08p3x4/4S+u4bLr5FeY5c/aPguy/ubBlyCsCDNGvfugpyFRAz1fglmllpwV8wPZZt
VlVXE5tNNs1g0a2LZ3tDxpuIQ/bn45adNR/3V2Dn31HLdWuphgpcS+dReOOAnErK+N7rOu7PFWyI
MXZtxValqEiL4iSjZ+xbB/TPr4hs3amee0IS3rec7GAYUngA8uTQD+FdBYdtkrr32Pja7Gi5dqA8
8REM2vqv7XnVl+g8JUPVsWi9F4y9/Ex+pHzB5fY9slHVJmU8PrU6c/Li+two7CBb4xHW70Q7MKxA
9bNxlpK11obL3nR7UMhCnO3NaOPozX9dNABU37ZILRufu6H25rDeT8rLkFqAcg8yffJyer9rNIiS
DYZ2IY++Izb6rB872ivhimwb+pp69CKY+/uPs0q0iPFngYgntCVj8pilbrtUwMKGIZ5v1NmkeAVQ
wxRFzjeEYgcRAPATkS7eCgJWifuGXRj+XnOxGDx8lGkyNFqBCFLM5LW4axPZxvcUaNyrI9m9iyF1
f4wRytMK1YIYNCbWNRlWc5rAAcp+Ytd+upJ29sxqVqGSBPePoIeB1kTZ20dOffbbSsSaVDWtR2eB
eBvTE22J+zXbkEox3PdjBph8wUuEnLMghLAMxKeeKcgeuhhWfDEw7A5OnRu8rCc9goaSOzPT76yC
3oUYzt60wKP5xLEuJnYZ8aJz5HC4kScTTOtqoqKC8RnFwZ4V7LjQTVLzs7MU2EzA/dHAUwgMmbaa
1P4Aobc5LOU4SG5tI3dwjf0B3lJsemuMOY6VEbvZG6/8UOH85hZ/xNOOXgORikeyrJBb9hXOty7a
/bbYQFZ7EKQpkWVbVqxgSJFepXbY93oMsmJ7X2ZdCGFnB48KhCfDNHqCLGB9X4HYII+WHkt4aPQ9
BA2WXHgJXN7hhJYbsTAZbc5Vx7DqMpjbVxIsnVWBf8am7WSdyHQebpmd2AbUpgQWbVpoEZR8MWun
GANC6REGVZ7eBgFNS4w32rl5zCHR77CNeul/c2zZc3Zlk9ssdZYwxN7ahPgCA7k8dIF1plGy1cxS
F3A/smK7pHL1Mvl81RBhrReRpK5DJO67LfcQPmBV3R378cpW7+K9IFYaIZhcbAJkM6z4TWSV0mez
KKob1JQ2r1hXkSsJ+9XFA3H5nbKhDDJ/1onXNUL0RSpvYXbKuMjgBmIVSzTx4SyR9KmL1Ianq70+
sH7OGPwkvuxldmXU5/B95jCjmlQODdtrOxU6CCooJRPiAURvAeckeKimWdrstvQYGKgI9PwXS9RO
2086aANshn84EdFXJgjmsIICiyC4v2kxtnYj66C9z2PpIAmStpHT7/SAX1eytmP1AoxJaWD29fLm
UKt4W4sZ+o3Hgx1uq77sOXiFGzSuv05ckDx/IDNHNifo5MyZ4L4T0AVZBo/v3p0otiG4lxaT035l
UuYy7ZIoH4ovqdLQYYDC1MbAhy4fqV5LIs4meWJ7gEXqNR99tSsDhjS+1lMRwd/Big9KntBP5Hso
pAo5N9KJhPxYzng+Tskn7288O1/Y6sAoRvLWbCfn+uOlcJeCIDwKuc8PM5uARpXdlUv2d87z73iF
R1EW08B6WyNLGT86EOHOTvvgtAAQ37THpa8nN9zuFI1wfAGX2WVsCw9ox7j1WrlfkfkYC9KyD+Ux
Oi/gEmE9yA9bI0ng/bSm7Qmt+L6/MsKFuXUXHiUaC+P6XQs9L534bmr0r5axgV2N77V5Bzasjp8B
lRVinn7vvBCJZgGMP6npOvFPOrXGMu79sJAzv9LCeSoycbzPPAZ66V2ac0ja85+RDTza/+YTh/8s
muwhQzTtBg+Znmv4UatXtWOEp0OVacAzk5fKn/qLXqQroN9wHizER8JIguXk9eaSWvEPnI5tQi3V
RuzZAWh3iMlEOEHfYjsLtuSmgoNNYJ5qr9teu+DFE+FjpDMzhcGpFIRXKCwkdkJy+m/7CrJDxa6j
6KzoJsVOMVL37gzIL3MDFJtItyQPI9kjjXJ3chjiPY441YgxWnAzQE4eI7EmWCS95R4fWUj3C+mH
+FU6UVmN/DndY7eyKhYJC/nHAJUeJWYty9XdoDlRkMB3vc78TtlFHt1DKTL23+BcwA4an4BmQHEL
lPq+4savCwsNPWNpy+UbttfBkIQ5UuTwBa0w1OFPXnO0l62CQK7LTcJTkVspE42Q69wu2CxSpm31
2gsvtXpuXwGCCIk6aqA1QrtarkDU9y5WAJSyZhkO4FDh2BPKsyixAsMEOpH8wF38EwYcXcsQthKR
LJtiuKwl7JmFNBYMpLuavKNGF5hrL9lD3Az+qbmPwFTu4ZE7UvwY00OYj3j43UvsHN+q8k4zJyO9
gPgHjVuvPyFSQpIj4akTH9ZtZiuY37xOEAlk24ZGOztwLSWKEtTDxJO2R0PhpDPVNvEw+4Kk1ORn
5pc38TJrSxvZzeZ9dynuwZw+1VvIg8vf9oFYshtKR8InOwE4zpLDJrfych7RsWUT32oxThdAMaNK
+F07ejuPBkn8aDHmRej/RfV+YVzekVFYChLWcsIgnIUDVPlhQ4jaHpDb5uTUYy94/69C5NGRurG3
lPGx38mfE57mVFCAkzrXIMBK5PgcWzBkFc0n54eX/fsMZ1GBz+3p54xBPf180ph4+ZLvkO9wwP1X
i+Xn3nO49qZkPcdLxvTX0ni1bbIEnzRLIYD6ZFgzDWZM6zI5AYbdE8IqYXruomvxmekcYKzjolzq
IxJEzA7Ke0kZvGNo/Yq6nZn37CHo2218Pvd4Wq4KeIaRg/dvJUWz6OWNyYyyP7lJi0hZ272guD4g
RLkbQuz9W1yQrvM83LFuWLrIvwEhtXXiWJHLvpr6lBYoOq4LijHp3G4lJQrX9e3BGvRWcu2ZfZVV
vRHp5jv8gyaM3ZcfQnQxO0Z4QJWugtJ5LC56Db5Nz82qPZLhg/iD9N25jmyVEUzGEJPt0zZy4yv8
8eIE7gzh8KocxTZRXlBSsY/dDZZYJ0yFobasbod7HcHsMxLG72jrd1ZqiZRE9IDHHZC4b9txV8B4
6rxqyRy6sOvZsG/4yRK4kNmRZZvjrgCdcT0p08NDPW5RTk5+REbhkEpehu802D1pMM6A/dhSLd2B
HUj6b++SPGj+hzssQOZCuYLT8UDc0UnJIli7VbPzP/ICM4nQ0tZhOK5Qy+TTnQDupiTqjB1wSuTE
IOXOEKVTSLriqQMyN8u+Fc3yaId3nM0kTlkxt03beE/RgW7sc+/ADGoFpUc/MKLsKfANecI/SRC3
pXxwZ8RW/TH1+0BApBpcp8l8UVhd0Qf+gYa08R4OOUq5SR1oBVw0J7sA8TbSdQLJilMTSuioAlg7
rM74vGWLFMtkWXTc1xh3tQb65K7v/32ZVHF0apKCuBLbDCreZmfY1BFdLI7cgj02L+BWjcbdK9GO
xE0gjSjSsF5i1gM4l3a7+OkcI2KOuH88twIj31skXvbZsLzFGezhAAuYVnW0Lvj7QuENf31Az0Je
CP3SKnkAuYoq8Ylp6KNrRE9A6svtaSkknpX+aH8THHHwBwCpilw8/Cr7hLs/3DAWUD0lJU0iymNn
OaV2Hd6rDAePCRf9CBgcbQ82UNyQ6ll8pINmp/Kni8o0a7kyn0mlq4Kikl9zeTr0lAF4cnzwGvJA
q3rVTQoUbCl+TRlaoB6tmr5juGiVHkVm82giBpyVCv0M/Yfyjguh9+BOKgRW9ZmfEaYGYDP4z+53
6p0LOAr/+fXEPzRAs+2ys9b0/oxm0cUhvwheQneXInW3RsTYJamQmte+1/b53GyxN7xfQacycpYM
DNjWs7CnTyug0speP3gHJT6tiru1BZoBwyyK3MIY33gYVWE656zzjU07rG5mkm9fjI1ugM7onBDN
3U2FlZfyVTXK7T1LW2iiROanvr2niST4cpzyEMoQQbyrVWpeddD295wtRp6LUy5Dss8O3JwLmhV4
IS7cXOSDxDt3FR//kAxZZRyb2L69f6Ik0ccjJ25+4pyQJxeTf7NvwGwD0057Hl1o8IvTZE6cy/3s
98nFEHmqrKCg7i3LtsXq6sabJLSuABuCFMcPhA5FG3ZN0j59ygKUOAAokze3iXk32ekB1tUJxgYU
EyjluPs+FSixOdFLsDVd1sxl72gCNXTFUWCL9DN7LuhcWxygpej8rPtwC7wqbkecxOV+lHDVjjMS
J7hw5kHhucqmMAlYdysu5E1y7a1dOoAb9rMfG6oXLsEub5gG/LhwCYMoELcxAwRRk1ZLSiG1froh
PE85kSdczrdgMvtpQEj2ODWcNlhnSNQ40lewhx/Rhvto10NSshUMR9jdEH+4AKaiA54rD9SaNCv7
z2gonuk9Z4LcTzhkWXGUL6WHrWiJ1J2+WTy2/pKwewoUlh2rFJjQwIsv4YDctuv2fQ+O83xsu8O6
k3U/4O0SAJln1t9Gq1crTcyJ5dR4jjfERbVEn0ix1Q60CYWDmGwv/JNpm//6IampSRasJEBygGyw
LD9yUEmokIoH9mAxuesNe3Fa4fAjnNk21BUgRdnrTUlKxRMAKqZLgahdypqSdJOHnStvGJZWkUK7
psuWzn9MvOjlpCYVRAA/BgRSNIzVK4pM4xEnglvAcSPYT0EF7nZzUhDL5avRR9A5KM9+7JJpPJHM
mX+L4KJcZe6qSzWnuclxWdZh7yYTdeAT+Vp+8lnpTTKLv6w62VaFKB6LXUd00iK2oYzAy3wvNdg0
FVh5jj7CZHNdDFvudAGX1oUGs2RiFylOyI6mBsO8zdW2xrnFoRQ8VfInCNgYG0jJnHBXFRrE4TJZ
y3tfGWK+i4STFqDq+om6oxpYcHx9XAGp/L9hJtQQNABgK/3AR6JTjWLPARIz54sXqmmY11lR5c2e
4zPa9buo/Z5arX8L2bPkdf3pgMZ62J8BaC7gDZIjkgAUh3t0SoTzkK4UfCvageH6rjX1lviOTXVy
6QASb9wxuKosW8468rxl4758I1FG7haRLvUxPe0BISOlm1vBcNpkVoTHnshYA8ihSKdPqAiTAVqL
1PxHzokM9wrfAQ7xCTlwoMiyQ78jv8856gykAOqnepCJFrCRo0QmhOKyKsubTfqQXVl4CPZJ+XhB
bO4v1NJ03d/lZjyPc3HjHJPjP4v35fjxs2OWV+nd2kQEW67F8p9CDjfZZw5Z3/+6ak9wO17gVQCh
KEcFjgtdV9GweChsGg2bSgXEL2tXN/6kiN6KosnHWKLOwXegUdMGYCDalm0qeBUMXMVQPmyaJMRX
pft5iT0eycWaFNdSWCV5IdM4krj3o2VpEhSwH3oyBm/xuUKLktTmekK/S3fJ50S0iDEiTC3WrCQv
+/AflWUPNIhEAiYLLJqSqfhYyCUcC4ZfdJMCgn2J+eahwZbqZUrrgw65eT2MJ9PnwXOZq2uu2EKv
5uKpUNbWWmtTF7jCyoUgR4DNR0UUqOqOdaKRD0JcDNNbhu+pgdlM+xjHuyBuHtLkpKV5QsKRlFM9
gEvw+d2wSe2Eivj67yN5vDHecfSUFESCU2l0wc2zRkuEn+5S3wJKxnxYpzorpts6Gqzqg5wWhB46
d4IWNtsmEBFlkHx+S6kJV7zCazwzUJs2AMDxksRuwdirGep+vwvqNVGw0RnwIUTeY013KDoxCYG7
fPm2+388sqMs8e0A3AFAijs5udim/hPfUN8rL9VqWqVQZHNcaIbtea+hGpPtp2BnrGHSUytIkusD
Gs+XeD0sSrmQUY7EllAA3CZkEwbsunn6mYNh2/sOO1bc9sf5bdKa7A7ZfraULJH2Use9BmC6RClz
WnQZF7gr9+gLMUkfChxiwT3ECLPrzMSguCk1POEx/Fcgbu4Pk/J0l7X5K9aNlClY4Dp8L5hMiMOL
lwf1djAanyIfPIpCEO9MISL63lx64BQRR1ZvwfYjm2ig+bZte77kqeWmIeMh/1SDOsgfyG+kvzt0
I3on57KlyMSo+jMXFCdKXxiztCmV4R20JOuXIl3gCsMi4EPTsuJtxQvbk3Iu3kri7RvLmeDGNsn2
tAR2cC6aT+Xth62vu9l6baSYLg8h7ZArfjNcGQ6PL7Lm8uRuDaB0EVYbakXHw1d0fKfmJoqZ4Xds
dJtN5tJTpwpTEMqkLS2lbYEAXDgP4TKCk1AP0m8UBPFmtlR/3c+YHh3d3ihg/I0RAWmUk0eYTSpn
oJqCPJtlokJK7MJmPQQzrDrqbbWF3XXwa8AF5B7H0rUh2pxWnI29Xy+5nTwfyL4TNpg1ml74JY0O
qNd2p3ViNJcYgrUd5d16iQRnfTy2akOmcKoI+3e88XnD19r2KOOxs4mOtsgXBPe9EsF+igGEEGgQ
1fjU2I0tFSeKUsfhAoQcyu2JfRmXENdQ1jJGynQFEbfxtGzE4OJMBsWcSnQvU2KlaH/wzj38JZe4
7f/hwmcaRVxOlSA4NP8NBcooT21ZjABzH81MRmnVJepj3j2+gSlZah8XqhMRhPdD+U4hQ7FAfQM8
11EOR/13w0GGdBpB8z5vL2VFkZt3Tww12fLWAdhwGMLVHdceTqJIqi+n8j0zdAQtUL3XtWoJqIpX
nAda/LzsQrZt0AZwy3VGzbeaxTlwlbH9qJ/+hODYZ1UVhovlEnoqnbN3mEciCws2cs3hwkJ3B9Lo
qLSqskW8K88pyjh4oB8q5313A1o5BsgwqqmzYOWxgY+Uosj7zhPXXR3Pd5Crnwe5+6WbZ5lp2WNj
n4KJpE20D+ZYL9napIvF8GQvungPTg+fVTfMsuZ+S2k+aupWGrUFPwBwEnYNNFADZ2ErhGucH+IK
IgS74lNS29qxTbDCORxb9zTtsj6HtaqsRB06hmjun46oHE+wDOH8NnKi4IZNaoXWtuY78tVOqQH+
x//DupLX6VGd6PLpEPjut6SG6Tu9+Tz3onEcPtjiqpzNQ5mYpc7qgxCCKPLYClKRgPKyOc79LRn5
gUwMtbArQkxmse59Rgy5R6bETQ75ntiBxPamxnRSZn/ck85LYfSwjIlgRI99O1p87EYiN4Ig8zdI
v5e6eEJkyo5NfU15gScaQFfHLF/aCL5o5HXCZF3Rm3C/xg0k/imOrYiqMYE0DBV7rB5ti2dkT/Ju
WY3p38UCYjFW4Pz73Ylq6jyTetoxeyRPvdAWA5tnsElNt5cpf5CC6wODl4otxBl2yvKOSXFhWzc4
Obw0ISkEGXtMT/KEihifSEpLCbIFAyNhnU6/yOu8qXx9eFwdf/xE8eGviFZTT2HKC4L/XbXEmlxS
MWRh8q6EmrrzlMkQnyRBPG3/CT0vGUL6Bwd7lMHRP1T+J4vC5EgHgslQaMHduU150HvgwVdy5t+3
XBS6U/uBWqhfpXqA8TWma9ozJNGrErHvurC8UUJM388j4uqYD8HUqIj/IV+o8SNHn7xqg0wS7DER
IBHWacAfKB0QvhBrhunqWOWR3V8zLYPRyuxoklcpTjZsGbQLX17x67HN/cZxQlY8i3W023H3QY8A
sj1iGyRmHkBxRaXAzjt3Bh+VRdJxxpyvss58hMej/+TVttvA8Ri6Ivzkx4YdJNmB60vH5u97ohAh
1BBVLbJOABZfWojRx+xXLHPREN0DnBLo6whFd0xRefVv2rq5k1/edmf28zG7uGX7fwk2utAvQt4D
3hN2YWgmQefERKkzx3CQHMJrUAqvyH2VLrMPEcJoCxHb1cSznPbTNcaUi6DGwEF7gpnwCzFCT8PH
wOtpKDpZY6xhUo24n1+AIal8zH+UxF5+ndcP6pAqSr50fFypQZaGDP3raMUjUI1ymiBh3Jz0GVUa
SWtrk+jNbry005uaeU4CpiblYZLVsgq0YXs3g1/2TzmXACxjcpJufJodLmq52FyAaRwYidMJBSJe
mu3CxTZg/RYC8V8GcfYD/LbqwPsXZd9KNu6ITjGS87VTWYv6VoYrQmv3pQZxWBbQyqhpNopzFrng
4sBXg45Tj96DFlmaWZixJ6FknZN0JrTXJ7IsqWgwq6GH6/nhbbKI0XDCySdhU9WExXdhyDZy/La1
y9lEqoaMsmqAnhQsqZ99Rtx7m6mbFy1gWothFN0Dpmb/V1OkXc7zQoJfuNvuFX7TrWi28GKTWZp3
EBN6EALurKUJyET/dZUQhV1a2kNKlIEKX6ywKVMAQ9/XYZ92evWcIHKZrFHQ4MbVf+wZWvCBeXia
4kqep2A6I/x1YMajss/svq214bmMikm2hPcXUb7F1884EgxZ0/pKaENKiV4RMUwHcyEyYGEbmKGt
TPvts8QXj9Vhsy5yorBYuqLbp2W2KlV3JRn0StHscE+8is6vGyEx45psVUMBT2IT+1m+5E36mkxw
NgWrKHzV6Fq6kGCxrurZ8YEkPnowg9sqrJ0YvGrI5oYuw34kZuUbN2Cqmo/lwGuwFoRUVrDkLk9i
Smgf9Fib+mtzTm+VTzHOnnkmJo41RYU+gIoNAjzMrc5BB065lCbwd7tGz82BizahBJP//nXNqyYh
DXwdoUs0GuVFv6BVAbFuW2sbSpRfQPinF5bmQ9uQAR8JspcSmF2++lfWkJDy79rpF05m2epljabk
CmlSqWewNRYJd498ifhJ21NnGSg6N0xvji+HVnkf9zLX34wy5X54IA2kJDKSk7Vj6EIfElw5rej8
HzaHGuSjIn6Aecf6FXgipkLOj1AOKtW4eRJ1dVtTdYoiuWR9e/UXwR+85aJaNL78XtMQTNebn2sh
kHHQAMXWjSxVeV4YduOfmUBmKALXdbhf5Q4qpnrhR9PceI9AoHV6Jgo4xOnZjZ4XvguSwODpt+WE
NT85E8mRcyN3v7K7Ayzm2bKPDaO6FUCb3bIgKNQ3nRpIzgk84aN2K8O+AIkSaVdt7q7DHytb/66W
s3VSVa2DHsQPqK/dyBoQEO6lV+xH2USDsb0BbZcojug1HpONdHJTzXPdQw77lgkj8TqeVlAMXLgk
zYbMwsSW0Nryw5WFuYugF9Skz3UYjoJRPvYc53QUufaQmicL1JEuNwYQGw2KWbc6IB87t/PjFbUc
JfR0w8uZ4o5ie+D2nyLFDnl0iew6H3tuAXwfuWvYlbe8VfTV6rK/mkN0S1OiPdr7OlDjv/bTjzxE
Ujuj6TJUivC0o9QUm76YpVJSbaJOSieVvhNdlczUhzhE5XrU5fkHliFEnHDkrrbT/dDfIC2CH6qx
7Tedt1ZxOhEhJ/FDNA2IptFUcuWWFPGOUL9z9zR2LSkNgiBSdZ/l7x7GirE0Hx2jBq2RWITnRbIs
zGbhTh6/mGtkdmRho1Ci6TlV/EMZB6Pk1vq1G7cOEuOxo5j40JtXxxM461RPFeC0/3DCQT1G1F5i
Tz2Cwi5q3E8xzOBLV620pHII/BWZNuD3ueuuzy1ah1vofQAjHDYmsWfhg81vyBm+NlMGq8YQ5T69
Aob9SvILmsM9Z4/0aFeJ1KADqP9BlfhDeoR+pP9X6jekNC78tVm0dOuJ7y1uTx0wJIqtTZQjz49a
0xL8/FBUUoZmEreDyatRPPFeWOG2OvE5nTLhouslfVEcX6eEqNSM+JDiZOngx/6NOFo/HbIYGoSL
NdZ6b+bD8vETBw5ZyHuK6W5VDJBTVYiTas0HCkzGF5EyF0O9Dl6sltIQfFdTl2eVDDc8y8uNR07a
epcsiugdFOaX2kfJU7jSBhCKK/eakp/0cZzckwys5zRL5i9GjvnNDkFpHW0DtehbIlv6w02C09Y9
US7+GcUTkPUK6aajUrIDX030UMOwucqbAXzBCEzRe7kGXT5nmAkk/kMqfgEZN80isYH8D1GBtTC+
QbxXNcxIzNtf/VH996m8wr5XavzB2HfPgWHaISpgtdTtfD19IMplIN+TM76X451+vYVGKGQr96LM
lA3/ElxABkJLFQnJieoqJdO2ElOk3OK6T/8TqNPDO8xU18UOJXGbfNqn8hLm8AW4jytAwc9RCe+V
4jTH4krh7oy+7UM6R0QP7taeqrlcyn/PiQMWcOb6+7FXjJ1nNxf6U+mZI+9biYxzLqcHGpPQD/qw
Sd1YPNEuii2uLebFnUBjEVG5h4PVlatNrslsAg4HvBmNnKTVilnE68qHqEQdGCxrQAe6CmYPoHto
EZI6cBVSr8GAoK0jB9swGP9RmJZo1QpAb56qV/MJyiqAPeI8wwxly6a4mrSqlfriqqY6Y+s2b5D/
wz1atddUAJGBzPBb6uFdQUr+EPTHitUM/tZWG+kMHpZGstMQ46PqFED7u7DxGKCcZRgenpQ21pYM
PMl7ELFWEbGRegTxmGWSUnDA42XISHL8Mt8I0v1J/r9mABAHeQOByaVbUAdIVVWiyQdthQyLe6X8
Qgx22M4pLQJssJU8sdqXhHXI2wB4JsIpgIbAc84eZ6+J804Li2GOpN7OywLPn9oZesCcO0QQ6e4i
IRTctfbDceYDq8udKhVWpXIkFc4P+DRIbeSxegV6CjOg5S/Wbcpc19A+jBGI+Xq4ILC2ZxijGof0
9LrGLXvFICqlSVUK5x2w6cNaFvKCaI2hsk5UTUwb7nb4/8hoG/ggACykpIUiwWTyAnlGaAJnADRq
hO/Y4XHcTnRWRutuMeel9f8Xtt2SHjcd826Ew2Y1ae3s9XxBYo6G+43e2ISo9IJtq9d63FDUmwuA
EQtNV7zG4TtBj8XA7omyoGH5H8FuO8Vr21TBLm41UxVz8GdpcTIXoS9jw0l3arQKdwDi4hpA5OZC
dmsYPmhn4hdJpbgjTimMu7pogdEx0dKH4EYms4EOLYjutIsnseyb2OaVpOc0ioefpH88o94hulKr
yd2Kj0jZVem8PUFB57HZ8XlGPOdrnEjWZz+nylcI1Zhp1jYarFMg+/79fz7MLYugw/MwtL+cvtri
WV1zopp5MWSwjEqIiT/j3w2Fdn0J6OK+OxGKAtO13PJww9MGuNYMU8OjRitUs7QVZ/Znxm6uxKmA
AhEd64/E19oHRVXV7XsuZf7dqpW7jvJkalhZuEPd1OEo06hX0jZNRs2JmCffpWwJjbkyzxWWirbf
XX8YJ1ZForMXv7gmA6VXuHaJ3ALr69igdo1NzyIwhyR2bU5bWIQ4BwZiva7bAThQ02beQgg2BeDQ
Qbm1sO8BSb9hSxHzHQLyzPKByXN42BaMqhNm9arXnt1BbkCZHT5AUCabYuLd/HHyGV5VZnAXFdas
Yy5YOg+H77njw9HIXDjWg3gEDjTuYaMPAJjAHJvUS0FpGpxfkLuWy1TxJ6dgl6M9s2LajW9tOE/s
d2NBjwHvUMeAsDh2GET6QTTmKyBLKXCr48rOp7db3bbEKRhq2p2Ft++W6TIvGSXRRtzVJ0g1NVYi
K09XqxLOitrQfaIgpsXkVm5/cYFcgq7ILI6ALni85KBxsmFs8/HIKpqoyQj299pgYz21jBmLrSdH
LGakJUbf+OKxVoVrKS/K2v8gwiHZbWtanCr7bTxW2sSkaTcqH5tKVP+gI8AmOgLC6y/KSEHptufG
4w7K7cnECXyAxNUaa0pYrwS5kXpal0x6kt/6wQ+/9pjtIi5P6W3sCJbDSPoL7IkSrJY4b2zakCHM
H81jv/733C04pHGWJKp38qYzyi63jVO0O9g0+iilbYDweIj53Da0vXBIi4GZy2CACLuOG1y3RikW
bCbUlbzh42CU8eU+pG19wTMQrW9AFrl5f1zaRs1SOewqAhTCttjrbTiZunOsSD9flAPTtnDKCbYV
txUV6mQghmLn9A/ro0lIu4nvZfcobtF0IM4wMNjWAGMcrzaR0zMcdXMTnLaZ4q63rjzOa2WQ7/EL
M55iiRImUvqhWOlj9YSHcOYp/A7BbaHSbenmp6MEbUGtzI5qX6nVjAfKY0kVnedI87atpF9b4o7o
3GRPvTk5gp71SbGoBHnCgKEL3cPA8yYPXLU4ZBHLPUh6kL7nnaB9wctBB3GxRth6Z/vQ/J17JcaD
ofeOeTT3P6B63KoNI1i/RE3KdZchw4KfnhRDymeKQDEW+c6Qd+UahBPDINlI+eo5Yj4lr1gBmgab
I8+XiVVUOOMf6Brw5lI8bBHrGODqLycBU7B8E+WfsGe5JdKuKI95xy2IvhXZheagMsGKtG+CSZIu
6zuUQ4CUG8uFlJ7V5aKMYFRz9Cm2F/NsJQVGqBv85NXowuKh1yLV2c9TdtpLnt63ao86Zxln5z8v
4/frn6q9mD7g63rJpn1XaX6saAKC0LrIcyKp16ObJwrpxhd9PCmB0hnWN7NBL7zSJTUUo8soOtzV
yeAQGaNrug97PFA7QPWvt9vcOy8nhddJPs5MNDFEHnOrWosm3f5a++PkHzY/cyBY0YAA+HSPoaS6
sLMrsuRmMzRLR3P1ZmegdB+xoq+c1S6/PqRuGfIMgqjyxm3vQrVgiE5JzZx+vC9TKM4wZ7WT9TKA
ATDvfrB1pUSia6g+PYXUZtGwKV0uYTjpp/c3NEY6GOlxBUoAUrIbBUFnVyu14eiOH3S6Zg70KYyv
Gxwj0AQWJ3FfAuvcw3HjaAw1AQdl9z3OM6WU+b6JbrGpbPYmfIg8Mbl7bUvEMgmMv3PEvcmdFA0Y
f4V6sDX5dIpEoMBt9PRl8WiI4HbIzOjyl2Gw0M5qD8WNMeLY5TJ9kjW6JQ7o3VqKtu2NUQdKXYMj
j3mDUvHa9dHsn783+jTCpp8EqL4Nn31amBoaEyL6O58Lpy4drSdVEC00IJ3gsfH+REF6Qw45zdK8
955pHJCiJ8Yba1h2ofdcZ+8L8IchaNfUt1/PQ0g/8lR65mbV/XzYp6Sj5xko6+stVA8CnbPuliCZ
10dv1LbihnB/0FMW8MB2wKE/r2DEeRtlsYZtaOrSLhLEY9pPI2+K7pFgGXgQbx8FbWm1s7kffz2B
HQKLrtyUcFoRRfQgH4q2OhasoUfoc+TBalXK5/xDHH673CQkrxnBPRioo8k4u+WkPfqJ6BNj0rpQ
RO3rsxFN05fu3My2pM666adOniJdwWz1auQ/BNR/VkjDgn3KrB4IwIoYSML6cP0xpRjDGEsBfJ4t
tt9IENsqjb3g6yda8ZoktYbjfMdJjuJ6qx/JuFcHdI7kWcazJ2MjNprvAHoS2sXYVq2isJVcqo4h
wOhQCb8O4I2JhHnKfGnoDkV+rEGkwAbdV6+tZapcFMDtNY/Bn/UFhMm56okG7raKiEX+/WpT+fo5
N0GHDa/QV9MPgIA3Txi7wJSGfeNmP1FR6ybfjp/mdWDKDZzYmJkxGukxfpZvEHslvzAEmmgdjlAa
JNkSOhl5upjMMXigbVepbLZIIc4vd0BU/CVoGurch7K87xBfGkNCUflmwRRBxEO8SYQZgmeArPmF
0j6R2ahtro/m2KNcqIg7sZIAaXoC2u197kMLT59KSqW2ymX/5R0AOVcbT0KoMzLvIzVirLEsN5Rd
Uv/0npWnPFmInOsMQfAFGgEJv9VyYaM3HxMnaJDRY0IMj0uivvKBPsVm0vkOQ2XfcRUIdFOHJux7
hSpkwO25Kdi6jBwq3ZYNJAN8UelIEhy39+QM2DL+/HAxacKGYA16f/1eCz6t0j1BrL+I2bwBvJct
PZiTjm18sTS8j8m0l5RH5tcnz+j79GamWuQhwxBUgZmp0x1hHxHrH1l3CFquNllrlJdDmMlIP+Lx
E7/vD9Asb/HxydLuLrvcd0/tnV9KyHIPFJJL/W+X46noTyxAzaBoaQ2hEL3Lba4FxsBqNpw2P9AL
XStlaJVWLnzfkGJk6eNrIxthZp3VKOofkw+xT/Rm1TP20ojiPCO0V1k8J6LPpGuycXLL+nc4UEhN
mJs9uAwm23y4cudEPS5Xdcs8qgLSlKYrCjHhkl8Yi3AK2Ovx6nlOVnFeDjZZDHkDCrqDef9DPS8n
K4mc1lo2TRItqi7Xu/sf+YCaYOQU1vH/48WaprXX+yTRLiZefmaEop9ZCutFX9GcbB23P0ZT1XTu
/mQF89hRQC5s9zilu+Z4HBbCa58xJzvdBa31kb6QG7Ka3uayKBr/zwKc7yEyqEcBPaCcxLexCjsD
/LTS3wkyaIN1T7py0AmJ8JfQJyksW8lIsGcptBng449Gli7M5GCv/SynDhG8vd7LchnAz6bB07tj
bImhHsH5HrwfVlT6xhq6C+9esy5PQCFgBY85cW4cjr5tAU6TK+g+tkB/jrCH4Gcsq+awkIR3V/US
v21M8gJje3g/KdYrcGpBdJWkY8K10uhp0nYQ9jDIHXoyRElhnBGSEIRFaCCJBD5Qc7RvJj1z4qIX
p/+MuodQcFFRjolz1Qhp/WbHQ7UzmV6n5TSgZNyGVQwpplez9BND5t0Vzd7cAY3230/3p3tV6wpm
tk7rwSrOPm1mt0lao5lD3+rLJUgD6RJBm6Jvh4MlpvGipjTKczP7a48Sh9cENxpGcZ4nMgMQMs1g
wAMW5AukputvLY2NUoRXTGgm6e5UUnxQ2HL99p5ER+SaKf8e0qV4WYJzlvzQ3XwayUAYu28SJ3vW
jfbwTmYO/Y0WKM9TSBvfFqK/XbSmRcVLm+8dSq54QYE7FOK5kYl1FM1SrGi8RF9r8tVQfwotRL2W
35m8PVtci/SCrcHC+UkM1laZRFZcRa3BFHKa6x5A7soNfYzMMobyfbz6vfcN5avi9x7eva6vpfYM
kWdaFptchSjxpq9wtZPY2uP0S+6EpuIlhu0dTLmXm1Z7JMYZPL5rs9MiJZF3M+ZcTivK9UXlGn7H
Y+sH03hhcySlmnfoCe11jsW+eUM2EhUONffbe5chJth6gFm3aS2zMPTGGe6qBBCTUV8810P228vn
t3WCKXjz39uZlaYBI4uH93mW9XDF0+eA/Evi72/sAy+ITGGSCPCgPljCRl/2sw3MWtrNaU2lkt76
A6B2Gg3cRJwZmnzMRiYjUcvrKP2OL0XYQyO3oEN+z8MPlVPYuih0tr1rqr+wPSdq3RkYuDZ4S6L6
Vw6L87uci/NiKDj7it8FLiEN3nd7DsAeshkFc0MKD7V5IdauBGcUEAzRcM3kDLY0DM7kKEJmaXo0
ileSr9z/OTFWZw92gmJxcDu/WAuI9lMKfsBvttF9kDBFlwgQz97TZSJqC2t+2uqogO7ovQELYzNS
0LeR48BZS5ZHxfGJ1dBY1/+yoZL5/Tq1M1vVsTxnha1ZM2s8CkSmfP6PXY4csjx+Y0S7ZjsE8tCp
2nNsBPQ61NIGgJ1Wq86bXkCX9xiXWMVmSvnsD24/JJgh0FSpTPQC2hXmTZDGwV1YLFoGUMxb9nP/
HZXz47i3+0IlTvj+B6l/1vp7AHaRP8bUNKzByQzTzDTCjEuYiMuFIxRSRdADSm39bSlYpdHMJS85
qjLtrFSlEdQv21Ez+YHYWnYXz4tPVRXUWIEYpBClUfN+L5zUNEJMqHDbztMY4uCc9kr9+/jT8C7X
OLE491VSTXAuR22E+LNKo1MGTw6amRMzhFfXIxhiw7PFUEQih8xx69cZfjDHUo3vuAcFvJV0sPfB
eT6xYZo7xuly9+6y7pG/bfQrnA87g/ZVoNQImltmq3dIP+SNL9eA5nchn8AuqO7lEUCXUqkYmpw2
frQP2SqW8JJval/JunCQpixWd6QnlTFggFCbQ+E5oFwOB1iY1B8uj/SukZcoHZppfZs922uBauAb
FHghgjXBWJfw4HEpFO2ubrYMxs4pwOT6KY3s1gejywBzcx/dtaXRR5p+7LD4f6jO/st23U7IUovs
YK3DpMZKtYKc2N5ENj/AMm+6NDeOKm0zQCco5eaV1HMWfWos89YuBG91cosoZzV90MKQUxqK3aa5
1EscDEP3vwAHQgcBlT+jcHTe0b8SCe0HSSUYBCguok76jbTH5xfQrxi74ktOER1L2QscATmg2TOG
W3ayEWdU/10TTKqSKtWD2jjF59J3c8JarVQjuwnU5Msss/59wCt53wFngYFGcPmOAAcY21vPWRYJ
mwSDLrJjjUhxf4uJnj29HU7sjTvegdnaUzNpc5esLQ4FUkAP0YRj90LD2ZXxVyLMc1+114BMrIli
n8P75JmhU5xvICF7XeJ9a5G2DnfV1v0AgLjbSW1GEQWjzKQt6QYRgFBeBkzMDk4iAIQ4rAuki/sT
T5itcZYv0omfHUwGJnMxgA0+NHzfTfriMzJLGLlaGkGfynaoeIgm686iDPIWI0pvAOjO1QrkjioE
MeBj9JAWW1jA9Hmfh/+1q+9HEn6tcvxc7ez3pLV++qPUYJkD2fEoC1RmVPtk2sINr03B/xh+Jxrt
zkvV/AtRoqx73lnpLo468t1IvfF9rOr7/TWrCilqTee3h7Qpx9K1qb7tXx11x2p4LjHqUVStkHqf
/Z0knuctxZklMw/qmk5dCBSpUKlCIn2WFv6Henkg5uP8Q0n1WShkyvT4yV15ayWcVp0wynPdqXgI
Jc9u0rmvW09oFOJG9vYR5JbK0l/sUPlK6MBSCdk6eKjd77k0X8t+leYs9vzbWguta+uZza53SNVJ
xga26gID/+/LyhcNkfEh+8mu5idi3aKXfReuy7GXe1+dcacM/030QCzDVxSfGpp7zvpEEv8K9XJc
wfP6B/r+/9ngFuOj0AsTuO25dvZ/ssDsU3t36Kyq/6OmlmPh5cv+exzoVJ7/bhhdct6HdiabHfWe
fNRGOi1LAKMvrF6f+TfbKE/Cx3fEcWvhesiMIsk+N7lASZN095k9dOOv4rLVUk4sPOPXgjm75Lh7
wglk/ha+Y6jb2k9uzGASKJiP9e9H2EACykqeTLYa/7niit6RPRffuztFf53POVfgat4Y2uGQpxSW
DIj/9mC+zq4cYBWhM7dX0iPOyLp9gkB90lxkwoCJqiqRVndlD0OdmwkDbw2lccSpu3qWjbIpfOcz
D+ldxPRdveekAQh5HeQemdGbMI9+lYM9CbDwYHyiWWJj26SyK5u+hY3zY6FJFdIa0kXHRuHFudTB
PhjcaqsSUNbYlLNU8WDywhPDw886eZbzeDLwQBXMw9CRnnQ7F1eJB1zcHGm6JNE5qoy3vM4R0Eep
sy2CNqeMD38+0FpymsLV0KWfHQ/6nKS2YGCwJcDhA6PREK0dhwZEYZiH0XATWsnZWM+WhadNUG61
kdghaAwbggZFj+m6SllP00S8q1zyda8LmekUpFeWY3DjNOBD+nXaA10x5VJjDXFO06KRikqIxByI
ZgPBVnTzpDzOrfHqFa1KvOBPFs1FhwrE9cXSLpEGluHKNs9MthNB8qlHhuw41lmjl6tjQLblIRb1
pL0AB107Bf4Sy3GRCuyJXTzbTozD/WYXhy1YUvEGanalYOysH+87shR1tUVP6TvBWyXG3FtADSsW
7xwjvXnKEGn70VtpHwAwfSw59Jke52YZnmsrUsFM3H7/GaMR1RvHzBx/kPMJv13CekP0mIm+UnvC
VzZvGDkAQPqpyYuLUqh5W0BVYC3WQUqsZW/loRCkvj97/DFytm81MdVJ56dRHJ6fO7AiMucd2k7z
YU7r7YFuc6+aM/Yba2K4QQl16XpM00F7s13+LOfVE2dr68HNSpAXLXjODfdcKlo8u90lE+gdKZlt
ZKxyY99ktkz3O8SEWSy0Vq3KGa3CIWby9avAVAhospoP4yv46QcPEZJ+S6dWkU5nAv9/PsV+OhUu
psk43ybu0xDC+0bqgC++87iJ4HXf5U5jJNnjGc4119D3VdM7ksJmpnJaysvBQat9FnGTJxe9w+Qk
QsQEdo3Bewd+5hkhatLUbFQyL864XZWMWSjivFUsjtSZTwF05faOMGAusLQyMnOfEOVTnuhoGFJE
F9ad1Ev9F+Cnm3OkbkXC5WRFAWig1MVEgq8tIOIrbDODsp5bbkNmHJKuQDnU6mW14+ipzMDj4rQk
Emfbciuk/4M5RRbfSBQC9hUqKTLBceaDJ+IR0EdaEsXMZ1l1jw8ROwk3HfaTEI2On/HUvHPmj8H3
Lw0SIHji6WpZcj5LfIX6OLARn9Q2tkjoJgVprVhNWOk1n1OJcCrmow1u78tisdhtrRg0tYuq03Kf
+c/XTFg3uLwoto3UqPCCgX51OPcnC4LGjvedZHj8IjnfuFydk6TTnYB/cnchTpSHWy4L1/kHuh1Z
l5Yi5abDDdqeR6V1q83fljEV1jhC+mPSZfzrPihzL5ZJwR2aRY+gDmLfAWmYzUwDBfu9Od5D+0tA
6p2kwRi6ARpaVGS5v6GpH/Y1X3u/lZkMCYQ3w3479bfLLixchjFp1TyOECrGlF8/UrSiWYo2tFhl
e+dvIWBrLcUkObJNYrOtrSJ6jgmKJ+qaCcd0IP1LwZTH0RJxKXxZtkQQ7vxNw0oNn7hAcZhE6yZF
edddxHN3N/naPwDIZUcPo05GAo7OlgspY95oaDpoXBllDh0EJOzXP6Ks6SI8gCIESDkp8ngk0mwG
wD8ewJq7MLoB9l0MMcAP/7RJt7URwP1FKFu6B0maFqPb2sfx8sgEzZkXKsT8gVsbIVaI4oU/+KKi
OZB+fyd9hKfjxNSuVke9TSrgdKj3Q8eeYUIc6MYGX3LXJOkJ5WknmzkjjZci7EBU09Kyjrdz6XH5
Vhl7G+kmdBvmGKATCbWGCtCi0y6cPABiAQLSLcA3yXoNdEWLw2p9B9BnVp9eHwd3q8XXd5NPJEBO
5sA7Ck7FsVHFiSDrVBctLwUfQ8LxOFbqX3KWIOyI0n1JNJVzp3sRnJTMFdCFpnHvHfDyP0EBV88K
5XJ7+WUrN9989hVnFppyXjDMxpeUsWL5HbWpEfek4xkpRLAClnCZFWdDXhrZ8gexQEWEKC0fh9pJ
frQo0r7K/FKC7raPk/adnOPs477ITFKUvR/2Yhc5SdkKZOmX4wu/CxHHoM0T+eKGEgoEB8CXpUzQ
2PSVRU4SZ/+JrnWRC9mptCFA7rNiebzu/iLEeZ1XSgERPlZSglBMWeZMfvPPfS3phSLj44jIzr9P
SEobZ6Z0ZtGUBY6fbS5hChyNta7QE2QUOvSDgNiK8TLdIkYj1GzFhALZFxDJNfhk3725SigS29d0
vwohCEDszg5VnL58OKRreJcNTuUD5/VGSYLShp6H+Qh8EEgxTGySCBIu4nCCGX8a+lqly1q7prPa
QyS0+jSrE+e04o7kuSo9ONr3BjxnSqFI+guF4b3QhD3puUtD/c2bPafCEt90qQN52+LwScSKeCnq
4REP4uX1YTImV8k+DcAW/wZ/nxiprAS64gaAtoHy5PMhKOCSE3scUjV5qn41QGRfHuIQJ6Bbg7lJ
4aHmh/T6QLhYtzjE31uwMDu/cRnIiit1Vdhsa/TvhtsIO6TWdoNTGiQRZfFaX/JwYKFUQ+MQ2iz0
qLXVSTyE/vX6UrOadoev+KVVJ+r4w0AV7l9qMk/0QSFcxAxfljBeRDeNz5/x14ORAu0mF2rndpcc
IRdg5Wb3fx+k9wAiustMUqDkq30JhIZrWhLNWTOYaEGcMiwSMr0uv31clA8/z3RIHJkRPzMRbIX1
AoFq77KiMv5pkH9UB81WB5Z6+W0eDBkp11xFFCLQgAeFXvnMsyrG1GqgF2ZvAFttDEZ+auoXHhda
9xLL9I8LKmUEP1xn5KJJCtzvKWs59pWnB1Z361arBqNi1fUzmVsaByt/Fm420rLCExawytRim0lA
Z+BsUC+TS3Db9V70wLw99+Xpj9epemlntdBAVKZamip9aagZRGJ3GbWg/5LCW2Yngc6DFnBUV4UU
doyZlH1NIE4y4X97F0mKYnD6uU3Why6Q2L6h9h/ITTevPFU8bOE6GhrglC3bP175tB1aqBHy9rHG
f4eEh/zBE4QO1CRnjtOk6nERK+HGhxatoI5RwbGL7X/e/ZoKLtbyxpCCre6LrNrb7+9wiEGcdTcA
H+GqNP+BESVj5otKIYhfayBvrEBXLxTSbe13SNOHbiyGWdNS1ACrqjeH5XZ30zIgdqD6BYXU+Vq6
JRmkseUEenwx3eyJfiQfO9hw+3nla97xPq2Do4YzRr846zax0XvTChonSrVGZEHFZTj24UhNN/gt
bCezwL+s0WOXEmHfAzDOs+gD9Y+c1AEY9JFy5Gki4L1RyZU0DRsdB7nScz0DdhKc1saLu1FYxqs8
JkFRTlbUtoUDTxP5tFL6uH9rWVWlkarCX2fxiwhl9YpJHxppeLusqeIoJv/8eHWv0HFM2OZeEuSc
Z8s3v0exZswXCx9TCgN37jMHQ5iR+m/LaTsbrtnlqvQ5W41Be6ftGukeKELkobERp+o+XTlLeWAp
mB2LYD7ipNurPRUFs7Bj2xbh6iT1MS6pryacXlrRe8YZc9rB3q+s4tzCfLVfglAKCIslCHtPIzoS
+q3kmF0azNeHmqThgX8HI036kcroeMvjk53VMJah17ihvxXd8A9WcJCKbumiKBruVZD7uZmW34BF
7WgbS0aqNzPbfJgnqf24GUkaWB9l+WeH9xu1DgcZJPts76vcUAIpmAps0sLeuF+hlyTDsYPQjefz
c8KCWR1s7XWay1L0MktX13YN139eCm4RGpgPa9osIwXcxMl7v7jTBuc13RBuSszzpprCqU3AAvm5
NoCentX4luTxS3ZnsXiNcmbyO0a5J2r1HiQw679LuEwrpU1jNfI/yzE8ipY0lU7DiI/jXiv/NDoT
OQVRiRLZT3JnjKUEisdF5U1fqHg9/2LFrG9J0A9UTqm27q26DatR5HtkRrcryxSZX65UiL+i4uBM
AyVLh2oqF+Gn2bIpdMDclXlP1iR51kvi1MobjNoarjtFphKkCPAdQQ08VH8BJdzleg+g8ApIXCuM
r7WxKoApYLjEP3RfWy37fRzu3Qni32b9AKDp43/SYI7aJSywY6/Iw5TiGVzxS3xT/XoJgNgG+grL
dat6pAu8WVnfdhPc8lCoA9gE1+sWnYNmFGxRc+k9ykDIbTeBAzJyH+wi6h+YXJf3KC//zPOxKeIl
GsL8sThkuPo2RojBker0TDJ+MA31wOS/F6MrzCI7Qn4Zc+ulgKfyesYXiek+a7ETBZAPBm5QptRA
5NCOnXEIAvZHtmib+ldvkTWSAYoHcQ5Xl44sK+Xhgsg+gR0bH1Qq/l0JRO2zRqVLJqQ2dcjnJp6u
/gA5HWxwdflJXrFtCj1sFD2OpnuWeACV+sDmBODSjLxdGXpyiBFn+Ci4xkG4z80eTSTwV25l50Nq
YwiE9JxSWSqmxL7eGXpzRjB8+/JggKckcC52IkmyOK/j7OtbiRaasMX8EyM3PTCUhzn5GsCbEPu7
qnlwDEHBbzU0KpEHmSZfzwatAk1QTJQE7sneQFfSxHJuhp2GEIcr3A1a1pXzZ21BH2SWX+ZoaFm9
B6fcVtrwMQBofQywn3/dsPk4tCp26d4NTU4nG81CdKsDCuIYl4a/VDaSjz51yMH3/rg+ZmhyAGVZ
+MLs5uJpdMawgt01Lfcd/FzCJZsvzjTpDgggWys6oXdrF1zGD+2mUDDw6940oPlVkUBFKuhvw5jE
lIFe73ItXpYaWqEe9jdDdazsG/QKa051zHsLLPEXVOIWZvNAsjnXLqo/58VRG/DWDU/SexTKFSrz
dkAHaJhBQBbOSqmlY5ISkd6jQ56otLaw5bT26XB3jNJNCwoDJAIMo8L9E3Pj69O188HJr2ri08AS
VvSta+5Nejzi38UGqZwnV34Vc8ACkN64I9BtxLN8eXNivSVVhEkTDHOFSpU/VCLf8LGPzzDzkxWC
5n2aHuqkpyKZiRWzOuRCRJjp56w7RG6Zzmjhuf4RAXPzRqmVoG1uhcfewhh1liaGceRooXSi/cik
Evv7WhlZGVWcAmYvQ65yRgCTm78iR2U5kQ8XPaUk0ZmBoW4roP6Y51hKKHYy4l1KBGU41/3mgTND
Birz1M/qddFSghep9x03biSr9+7Jw+RTQ/1RRjNYrwIc24uuxhIcG3tu/3Pwwie4IYvZSGI1Ft6D
ayH4nWg4PeDx0Pyz0FjSWBwTAJqdD70zy98BmAZ3ngWJiur0tWcZ1fThroksjOJjGeF7RLGXyuYD
dTCOzfR1sa0STwQbAFGX/wb/h16PPbXXRFVtjMDrYwNz2HfMyQW3czL4xEIRoRP1B1+2vToyRNGJ
UV71wOR24vDCEtDwPCRovWwqiyqZQjhI+DG6rtCMomEZ4qMKePvnISWa5ZuSMNXdTJ3bmC5LafKt
WqiwHn7sivAwAyQi5+Xxr0OmkV7e94SEtjviw/xeZQe09zvQPjVEpkNCoiGUIVUSidh8adbzqBO+
OOkt97ySy7DVkuRoGQeSUrTyv2qyNpAbUil5n/qGn9OAaS/+Ad2x6DXAqL2qR+PENleGdNfE4Elr
2Xgg5EySey/nFkqEtBN1a8x8zU83sF894TAhbkfKZszShHWEktY89NJ9Fw07+PS/g1FgoC3wG4YH
VJrKALFQSOb4tTQYk9hVlf1mHhdSAdIQIX1gVrzY5qftenC0Jk+WsAaCQXdH6Zq+T8yqtS1bW72Y
BC0MrEUCRjdgMj/IN+J8ehw31lGbtvGYChOdL1X71QPh3yVU9F7d/dqNHb/qBRKe3VyeIcrQOnEO
NSWtV6tvkko6eLDxaCxV9L7AH0jYqSN6Gq/ydd1rns18MwPZ8r8Dq4M1Ipiiv0D/XBg2t29yr4DJ
C4GdWemdqNyLB+sylt2QVr0FT2xnB0r5I7y58OLC6wdJ9okAondpaHfQLRl3gAZMAFzK31tdpSAk
H4UpSWY7wcDj8xGxNO7P+9VVnkKzXeiWbSJka+BMlK/bTbb6js7eWn9lvUk5Bz9AWryVBKH6s4FG
MfiI1QGD6U+b018aNnC2OuCLrHtNwrcDzZ+zrqxRsqjJorpkTuR5RsgODYFY3oy5L15R9Zoxwihk
yeE0qLlhnaeOSbvQ/8kzPuTWIKRlhirKcDJ/GX6le38ltcUK3sxL9Kf/4SRcvbwOucafqG3G2wcl
eB6sOPCcTQ3wR9huCXIIW9gOW+bKElYE7yIRS/M0MVcia4eMiwqClAQ89hj3DGX8fKtY6g0akM04
JucFzMN46E/5PDcWMoKhDJutD4q80UVXPJ0rFAM5QKk4Rg3eLqmAffjdFd5AEa4zGO6Fe+I11Hom
1Fpa+AIBdvYGEb2x1xVEUgytYZw5nQCEbcOJXCyn0Agu3ez05uGOnEk7rRBb3Vst1m7weylPfiQT
d8RzXjZ9d9nJlqvTaDHJGoIwNCENGAAglV29HX7gXDHLobOUxOWhlz6rr8krX7n+1yUj2bA78bfn
xb3/Vhx+Z7TkwgnH608kIPSo2nkjRBmgCrBh7qENZO5TtoyPtjMbLOgl3XrvTRu4+TjjmQeZBGvc
0nz3Qg6sg2aFFGjyy/XQMITYZD4XlhsekGmJNxKl7VahQhC4mSYcP6iBJbflMje+UFJiKMRypz14
D9zYot7FjYJ427X6pwc41cy5We3Br2hsMip0m/gmEFM6JhVdonqrjUd4e2DSVhdDfGIhRwhC2Bub
fdwrr2CzVcuXXlBb1z9jOSnQR+rI0UXqZth3Bv6KPx2n1MEMlA+gZePSeGfMRS3rmb9qA66OEiD0
MhMeL1ud2wEGmAIhlhvgnSo7AmTmMPhKoPBtAJctrwfbwxocuVJe0doMFdY/bJQfLN9YVKTF22ym
ah8Fimm2aSzNeNppvuhrq86/QF9nsx40eUquCxlWemYqqThiwe4I4duw9JFCZlCO8RRMcWhlwKM8
/6oAGx/0GzpSH4x+0qULR+VE7ngkiGFRC9Y9WwVkbdmYh9rJfDLkbJGpm8dO3elEKHC5EXqZBrAy
oPfrkK0/mWEjjuoQdRw7C/uDd1qOXAtzPi2Mk4HKLBhNLxagqRRse5ks6IQeDvuRoGU9EezkpHJw
KWv6PsX+T3ZxcrSsBzW5tBbkLTuP0jdD/xcOI9x29zAvAuVwYA5fQAHCFY1MezK7S4fxwv6v6Eny
+8kq1ojYkCa8zm6V2sWS8gZoCoIWhuNmGIvhA7ABzxTIyyVEI3p6mHtGf+1Arx0nSZI2CwdDKwWi
QQwS6uWEIRbPIGvThCJQ17o9JYjB1FRCTfpBldo6Cmvet1QgRQemjfLs3GylNETPhKg4CdCFwK0C
lbMOmyTGmuy3kwFoDYiCMSWQ7fY5VBhAyiL2mpqzw3z4X2odMr/MRw+6sOt4a6PjxJJUwWWkEvK8
cdpXSgwmWp1T5eV4AngGxGczSCltvzbFTA7hpkKB34LqyNone7bcqJX9DR6v3vmXlrV+Lp2FmeCy
Z/DtPTqgWxZFBHZYyKNYkQkE/yU5TchpsnrNZMiTcZ446/sHlw2z/6oM0dXuEqVidhK+ZHaRQBuJ
SBhuXkbb5eGo3twb+t1QImXTiqCRbmd3YR4wqRxCrAqX0kETVeMewU7qRqLSIQLVohrfsd6iK1K3
ABR6WSj/W4yJQwDJr+mfkMug9IcFZgjdmF1iQj1k3v9ERcYinE7pT0i/CcWfAX1dbHSUwp8WovQp
foUdDPkQtqnkwFUpMe47J85SdOsFBV6K2aY6fEizTETsw37gRZ+r84rO+SiPKy8Ck9+3q7iGIZi9
goCpk+PZjmKgalfLn0Mj0G2m4VpqRCf7gp6x3C+syJdgrc3hUpTP3YSfIPXtioqOLmhxnauppkOw
EI0utMIjKQpiKNd3SU1x08ssKPaXrbv6NNi9nR1kXPChid6TwpRXhVOtwnjqGs5xwWtGFFwQTDYv
HbzaVUZrnxdL6EU4xFDURNqHwufmicx8kJyRExMJ3CiZliBVoUMo/AU+pa1WdETbTDx2Z81Mxwuf
f/kj2fFGLSSZ3LESLcIkst4mP/naMaRqaHWwmtowPFigY2I3JjD0PrS3xzoW6MYqh8IrXkJWwEkd
2xf98w57nTnXgvhXyY79ZWhoadjdB9GKM+0ApKUPc9pFWHS1Wy8jZHUPZSZBrW4teJet/tu/oiQF
1CHR6VVlO9Io07542LOZHuNordoGYFQBpnSBXvvgtR9kWwkh3PS+h1JW3vSww99LjSh+8a7TpgOe
rRaNfPf7DCywZ6rex4memmg8rN6Z1Q3whWWaGcOZseXA7cT9TpFowb9lR3N45SLbGLg/ohrWnX/Z
CkB1qezi8wLweMzfQeDrIrIjVf3dQ9T6nShCkDTIOtzZx5J4VHDwK29hFO0RcgtyL7OYAbbMHts7
9dcoyZQMa0UXEnEMR7hnA3El6Wer8Dklag3F0sG0YzTF6yAvwggWsTpdQN2LJFZxs9uaLC3NBaBh
QFAIuyZUi4ypETu9jT3qN/fY/WRxNY73kK4ejvATcCuhyy8nS6aBN4vH1xr/J6diLY4UhIimriRn
eGB5+StBoIVPJA3/tJewhCqe2SVP9JFxHqINQo9f/6yFnALoUOfLnqo6geMGfz4PwuGj1Pe72Fig
s/DwygRbVNDz3g4ChxG46KUAICIt+keGNxCUhJv6ul9f54hWdtVc4Hr24fsCM62mGbvwxGf9UpjP
Y8v8V6WWGgV3tmT0gqZbNBFRkWCrYaroei3yfaIVkuo853+YDnxGv7fe28ofqERk/JrrVLDqRHIq
udF7TWbmBffgMP2n6gOxnvePRIYcDUYubClZ9okn7joJqCxIZDuJIhKbRGmSB8ZCU24e3OyqxOCk
zrBBOoqLUPjgZ+UHwPdaAr0IpHbiU+aJQz050TovB50n5dI6TQmqTsKPxSVKJ0gkdJDi6KL2owpd
fLb5x8xlY8NDZjWZm0UbugsANkwTxD564NrsahwmmGkJpIEy0wLEXPn7urGkjFdfjc6jHiYMk0b5
U+/UuPJH7tVI+XMMnnNGgJxEhYjSN7JpHV9j1arsesgo48yHESzxOySTWHSWatm9/7UEHvGSLlgv
yulBOBYp1IN0rfcESzv4kkLUfvMJKw+RiMIHaOQ7PJpO9Xh5C3m98NwFnk05nPWwM7rDRx/dPNbU
++u+NiSJq82HQ/S9edTUNmr72S1u5LFkJAnob1o+ZrnkuvgsOCBQ+pnaPkaEOE2kwix1px8Xcb8/
rf1Ywuvc9bxdp7WIiIGsxACFB4bTJqt6Oyscag9QgCOLUuoOOoF5cFCDt7vOWyNpajetYZ1oGFLx
/py7lVtcFzgyBRE6KksHVTuG9Vcf8atd1KabF0uhuAelYIuo3aZZ1hf9hU9qKCLxmdIFer2hEnBC
Dg37+KYQmMljp0qRtRBgrKy9MrTU93K5tQqIg6zhhxbeelhePVi1ygJ8YpYJ0WPkeNzOXLPhSSuW
n/BUpOeL78vTtkly3qsACA09gzoFMx4PyyV7aw7d9jSNYKLuj6mFS9OGqljyjK5GtJSXV1mtIGQI
izc62PXeWK2jk3vyyzaB2E+S92dxNTpeAiybrj9ohEiiUxfzxZV9nmUq8658tcitJmcE+k7LEzXb
fz+E3hmkcKiute47V3Rm8krWJLwnWP2H7QfnVzmspEpoT+N54DkDy12c1mJr3pZB16ZtKcz0wMzI
uM8Vq1hABJe3iZw9oWdm3H9P9YSWMTxBDVT4Dmm3tOS/pEe6LR8LcoGipPn4qJv4VsKN/g58Gh48
qqCvG6TBgjGrWsNbV3YVxXYYBgozqTZ73wpvUzT/0iEO4sHcCxp5cSsHPXrPBQgjeiJWJnlc1+4x
86C2LKjkBQL2EuLjPJahq0UXfOY9k2K6V4tGPPbFzAhi3Lf96QkI4B7X/E1X2iAkJ6nv2df3fulR
70+ZHnfXAXA3Tt1y1AVpNDTUClyLGP4hnltfDmxwicb+T6RB30/+ZtqmBw4XCkvTEAD8hLAU8Us3
FVuNwlvSD+EzBOq7cT1CU+MmEbOo0DAG0hskWqZFmDiixmORbLD1uLJOODIB6fjgEd7vNFnBq6Jy
3dzM43qNr+aXv3YZ/IqAUz55/65BrlxtoOdLGaF0wdDdJFbBh/hduSsF1hN47q2pzYa3I98x8Wrb
YnbzxHw5e6iSEMfBp4g1YFEAMBPIxIREgb5mNLvD2K8n3N85K9J7GfwZAq0cfEqORobr9K6xNNyn
rbCueglr5DJ6CtiOMKmp5Sth+zmsEL8B6uB6JXN5HtuUxwydfGVyPdORjPU5EpRH5dxno2AQMIJB
TcaNJpgFSZCiPTEzdmQI6aVVjGuwKoNRngMYKZwdcAZWut/X3I8DiO/ZwYSXOFpV3v/lGGYGI+TB
HCJbHfzH1yVWPkVEaQ3pwOUjR2LEqawdCCzJ2WNFAQdmLB5EOdwYrtZBIeGco+EadpggYKIvxzkm
Z4iviTzMjAaU7qs5paXnc7KrEZ7b69d6mD+Wt9n1k2pL8qMm2UJZrt7OIcK88uzeeJC2VyDNIDVb
dCdavHbOlLHVKWzgu7OEIYKTFTXo8xhTK28+ww563+/lmp431rXKct8FUtYF0VVgtv3TbcaH7WRd
AEAnyjabdYpLqttCUW/gStkuyR04H/xD9fBdzn4/7dxNAq3ZlstJJBhrB7fTjcGTBZhQsLjt1suI
DcZiC0oUgMNmRuztOMcjuf1WKlhDFS+aJJk1t9OlKmoGp6wLeAvl+lOGA/4jYFnjN79WK3lvM2Hh
254HrQJ6YptmU5MWvJBXxsa4r/+4gPCF/9K50j8GqaY0srr2F8V3Kg5Y6wqw0q5v6RlGcj2eCU5Q
w35EMSQiUgr1SzgsfSS7Sel7zbnfMXpY2klZpqSLtrsP4dfDk4wrLbsmOny+6QuZBrXoTO455aOP
VbooLQfF25HqfRKRdm9DrSb3I2ahUhS2Pn3RB/LSvQDzY+uxlUJAcDIvDz9/DSaOsTtNCG/OGqoP
6B/16l56jZrvn5UrVjpiyi+qeG4R5/+0OeS0SPCGaA5IZ/5gXtTGcGb+RQ2X+mQ7KTI48sBsBbsH
F6IfczS4rteMv6WcgoR/BxXPTZir7Z+rWzuRTeRT7rtvQOvj1yiRH+eWz1QJQCWPGxdJaX4z3w4l
1TJlpDsoMujoH8HG/CxpMUTHiZ8aCKDZIpAhXecZKtUERACzCcnsMxFDAdKN9pAGH2VuJGX26ESE
fVYG1M1W2zRRDNiOIswZ8s9VSLGIea8231gJ1VGjE6BiNSVXxFitTObKXi5pKj7KeEtUjx0p2X2O
xVCyFXJfNEk27hUhbU6ehHrEi+zLpuU4+PnQGVphbpNRpoug5tvnflKL/j+OsxpeKMmB0GYpxBYu
sbfrU30PYRc8E1PCa3f9VvLT9vQYUZnYPrQCT4QYtMEumBpHdQt9S6EmZtOfDjX0hghgV4kqkT7Y
tfqgQx3Tbwao/uF9uH82yVTh0iNIbMsiNT6T5KfuYrSt6/t4yoxQ3jJuCgj3NmxAx0v4DfoHpQst
Q5yQmHyGGwLDgbmroENqwFtpZoMXVaX8ZzPx078Gy9jgdjj74MZB7K25AvAqWo93znnETHaCOHTf
7+a13IXY2pRj7zKkjH1pqK22a1Z2h8t99cT1H+kcx4q4V2UXt1PyYxL6wDxslgZK/99LU/MH1yjf
8dWT9UP4NnjEC+dZJyV8tfOkTkxQsf/ywY642+NzZWDO31yh3Ft2dxXJ81jmh4LL7TFlKyJdmU+b
VGyNiaIGkDYToBJZ8Ubz4LHv019kAp3iO3w78hXGay4C1+AqmYwUrrNdf7byRxVxocE9QV9j6I82
v7+dQli5WrzZk4wCs+YIoy5fVxHF6yBw+g3Ci9y3g+OqaMzRW6IybdhXCWp4QvcMPximQ3JaVuum
6jqc/3mf0NWdTTe3yB3YuIaEiBhkFb5+3y6WTlRsvL35Pp5pD1qQRJnNBkGEd5n3oVrGaJonlqwH
4T30giG/M3HcJYFtdxWToqC521f7jE7Ncp0/6ZTZnmrmiPBopbyS2KQ+7tuEzuvK1XxZiPY3P9l6
hlvf+HpaknDV6xn/lycIN+5KXbsnOMhDw7WGtK01Jw9Zw+kGimH04SrJCEEViMKgLWJymyQ7ru3B
pcbkNp989Uer+ehlc1erGFBiD9YJ7lRkggu3kCXTEltaNiCVl6qaLFry6aKLtDmqWFNWJ0NF87G8
hV+NRFRxAazwlvBiRuenhPC9ScFO/Gy02+6kSAhsMxnwGy7DC/xyF4l8zJhltEqgQM2njDkCvD6+
ZT5six1dwv4y5zXan8v7aRYrmDTdzscqRgl5iqDJ1K01QeWC+lZMNbPCrrbz/d852rh3H8ZwE7z1
rAuyxaPmVNiY0fIDfGVrGAHJj4DY/oSclMYRN2AJEv5tzes7427c+3Ej3ukmifYIKbRPcvmZlulz
SQILXreEM9IWGHl6p1HrePTG3pE7c7KCdoHb4SFH8H8/lASw7VMkI2QckS/qvGBVbg+kLCajMneH
9Kg9iq+KaE6HPJKnVo3r46/CNNivYB6+3Nh3UwZMQU1v2P/JmeaVashWFM9RyoLmzvcWdbee7A6z
k+ZNmhSkszVe6Dbs1l2XaQOaUvXbmqu7G2VoBMfbmt+gvg3gHKAE4zlKnBA0rBogjE8AesNgQhSA
Ho8gHC7uC4LRi1XpnKYPvOTgvvrCdBh4sqSfR+ih0K+o0xbhjFrpjp9ieLg23HJ5DHeICxyDy9Fq
YxeIJH/zO3rOdayGyeMjgwfsldUo+20jKHbNnQn8UHMqgxlkWTflE8l40wuKgpmmd8tOzhWB/b8H
2VAyRQRtVkzNWZcRLZ0c65znNzRJ+u+BZwv8qpS8kViVKCOISHotKDNECn5GT3AkqAWvpThiljfm
ZtACxduiYFcoBo8ZOqD21QQ1/AUOToImZNzBafthAjSY5y9A/Kzl3Ak/Itrp1JzCxm4CeWQ/JWVJ
XRxedV5kJEVB8i4n/WJ1eZ4yI/TvSHbOKoNLnSg+n02su+WhZzf82CVtWSuUzd1zL5GSCfM3eQW/
g/sH8at9W21UHAj/6rkLNEH1oJRWJH78udHFuoopq5+lnEbPiaX9glrnlE1G/wvT7rTxv9DKJr19
G3COUqz+stvkUArvTjoPjuCETkI5IlbdRQWbLxxnfkffi5FQfUjILC1pKfXHVdpJuZw9gnl8PhaB
jFDe5Om3lVeCdPD6nvjy8tFpfVskj8mfnlyfjd2GKI9rNYfqanQil+Z6AmuRwa/HA+n+C/+h0wXV
D/8HpzsoCO0oXJLijPANz81D1wPVsopIrwrXxQv5/KDx9PwZVEcqMIpHM8Ep7uDFgOvI3MUwhUZ4
8gw7RBnXCtLP0h+GDyOJ3I56ZhKN5cX281fJUz0Wm13DAIEvb0nruk5DO+K4KoQlKqNoe1Jj4Znp
hrCu2KcFYu2QYN9KajWSBpz0KGfau3k6ouSw59FvQTvzw4vUbx1/kiigBWCAtYrHFxg0V4yqnyE4
uNJjrYnwax6WZHi7x+dL6VmySwbHidN7ttzN5kiZlOz7QPAb0rtDEuADC9sQorV/W9/lJwltwjka
1yiZoT1ILMkU1yQSd4a+zkyMalE3di1bgehTxF3FOEmFKmE6w0wbv5XPkSwyYNPaiqlVSWAL+SQ4
ccLEKGnpj/KIpuuj1I/HyQzuEUQ0kWXyxuc2QPbbOik4+LxazaZjE9Q0qZVmGsBYgjHVvE//VhPB
hdtO03AdUrpbHomnDNUyKwpt6Xi7iGa+r7Cf22r3/rlX0b7zXGK2KvIWnxpU1V8D76ef4ZZBhLMX
EDnnHlxYGpks0C8ga1fy/17AE2Yly9TS8hY45Mw73pz4UC9x5vxrzOnyUQjGIOgi8XXng/G/r0wn
6KPK5oCLGOrsaqIpQdXsajG970UbS03AgCxchHEe3BZSEpmrx5Xa0p3vAxodoUJZwBc1YeAgKDSM
wN1cfud2QHSb6GrZZ8jUj2pIQjqRVUZdhVbTsDCohsmjpBIJVz7wlWHDKYJDU8r+5R72Gw6TZqi7
cbgjeNro46PbiJdt/2OoEoK4Mdru8/9cmpSE9dyJ9Uaj6sxhsehXXaNOmmeo3prEuecxvndHVXa8
11lPBWt3TnTPdK/j5YGoOthvhboawmGPryCvBp/HqOdp2ID5LKU9RpzsGS6d/fZgQGn2IfBQ6So7
sktB72bXMJ+Bx98Wpz90kJj5vJUf3XHDDNRN+HLCaeCS7OaBtwOXtvPdwTalaVEfkobXGL0nyt0A
WhbuS8vT6C9cuFBHzErR/BBFr/NYv4QyLSaX/vhwTOlSyfL6qfQM8cbRFVn5sonKAoiOkOOMU8CI
qGTZFrFglpCmV4kUG8ms2gFtdWwDcp4rxlnswV+pc+C4VpAIqiWd+Br0Up5zzoEDpGvSuYSohFmZ
d1UdTQYTS+JLAn+m6bg9jlW8x/nJwRiRM7pZrCUKBb8wtFu+35nfwrACBkbXsSlWSnFhQ690e3ds
bOpUsr3HXlW/kQ1OvwbN6jIUgYZguU3yBgcH3qrfGh2yay4cYn4805823x0R9exLES4CeSleN/4Q
p+EY2TqMiwxDwxnfthgNKGDf5xo4Q/WgnVj7TLh9q6DNKRC1qXDwEbfGy4nsjaZe91VTavAG8LQn
kIin7yebVgFieuW5xnHrFQzD58wfRnXEW/LTLdIFW5pi/BMcZdiRWxOBeYxeTScAerF6sFkdX5jw
raK4sGOKXL20PhCJGon675ZSlG+2ljHztJYfsfLtwpgQemYYn+RJSL5UqJtp42+6lKuYFTqJDsp9
O/NHvYP15QxNkNBxHTmeiXB3TcPb2tvbuVpp6k0qsOe159iZg6cCHwo8ljrrBhEiJ44I2dCiJfd1
6EJl16n26JQ27WUU3rpWnT0XDNvZuUX1ISJDJv3wbrAKPaSHobitAMtWyA58XGUF67c2PE14tZv/
22KAZgFbEQAHTU9j0UxoAEX3Lmz9ArC3jfSNzKuLASdH/w1Z+Q990YZA7VJaZ9O+mf7GmLOp4eOA
wDV8JGMfeLNIYRWtahZEiBGi0uMQdvKBqQBbWQHbS+3S7Z6IUB6aUEOg8cMHjlma65X65m9rY2Dj
V0AlyGXrQcCyNt/qDQvHU8Gf9Wb5Wahm7douJV7s1dRvj5tTBKKhZwJSoUnKNvMDvcyGX5HE7CnR
j/O9lw+5Deg2r0TMN3py8d8b9BG0+C4fo+nkflJWyZOv3+yiCA0ZneogstbLoCi388k6fcv3LYf5
lVLTKoo3dNOGLRYYX/zCyprknTBOb3sWCkDt9hIZJF7l3CazdreHwrJYRoPgz6VfIbHk6StAoPr4
ZtkjGu1TKck7bIBzAgrU661bUYpI3JuXNRSkMr6RC0gYtvQH3FqhgmNDjL4EZutF14Hj0QZY5Pqh
QYwqWz7Dj3bVLMArFUPD2zJV7pAAYILB3GWGVTt55782FKY9DKHRDxjnF//L/qs1UEFUNMBcMk/j
TyLE30HIQfESbCgl9t4WypZ3VtObHGm4Be9Vrp5dzzU3DiBbfxmtIoudhJm/pnzFY+oiLE8uavwA
Yj6f87g+oyhEM6DVTSJkAUJPcqrnow3x+IsiFk69RY4/+Gg+Kit5lbtObt2+h3E65gJXQOhWZbfB
iMYEjuCSKV6plaEHIBavWgtdV2qIMv8CPNpLjTn875tXhZLFQ+0xPAVYUeJ+kXii5xh+w127gDWl
W7MTVnnC3I1Ns+41D/qQRAk8mGEvs/HTLr3l2HR9EKc5JFUAwPDGdU+VWCsYaks3biP0wZLfYbI6
J12KOCpsP3L4zqC6l4/XYOqU+jRlJEq2rDxO06IkENcqHzuy8eUzAwYrFqJYiOqCl+4zm+/Y9mm5
UpS4zzCsOMGlYWMBKzfGJDf4m69GaK8Sb0MV/AT0bBuTqLgAGt9t2RBeYmDujOA602UmLS5wDeOK
pgOdy3TFW/HsruwGq1K77gbxmYD2jaMfcZaT2KpcwoNqDX3BJP9ABDWJTCJ8xfFsKEPjP+IWIYrc
rS5Gs/NhU4b/zHLaHUJXlXW8G8SeWIifc7bDiujD6ZHCGk36dNB7x1cqnOSxh715jM8qSk27JFiS
Hd+pIqHsfJBfZtc1+oQSfBhcM68FW+m6wzOOgygUWPpTyugKXyx4gp/8/wodcCGQ0Ytgdz2Of+/c
yZW5h0aBPqRvCyhl05RNbsiJQlILbFv+9nBARMsLhPEnYBKwAWDy5S3A8YoPUrCOjGNr3MHuCWIw
00CyOXYSUxGN1R7dEEpt7SrSg5LaNS83tF5aTFyiJuPJkS7PiykTth3+6ncaNj2Ia0OZY/mi75dG
kc0wa5yE8MqQaJ1KjmphScJBlIw6mgsjGAarWtY49DW+bOwyiaT8uW+XsBLDpaAXQr4F6DD7dpSe
xA0fy5A6sqIaFDWY2v6F7Ws1dlRoPDjoCSMc2dLxgMUvXdd7fQ4yAIx/3a7cAq4qwe94R+r4ZcRu
6SqVyIgnTmps/OGtbR8YfieFzjREBSQSFHqLRaa9tA5UH3OhsiS3yO67vkk37CQLDVDpuHKBO2xC
pymAHGC+xkJw5+L9RBI3k9IRzVN3CnRIv++7DhBoDjkRIDIUhoTnCGOlTduNq7apNYCvF96XpacS
X1VYh1+wfs0NBzW0KHidRlZkHoBB5JIuFw5BsfPP09yEgWzAMqV6xvpREcp73uV4zt1JduJRofvU
tvpRZgUvoybp6dy3QHy1cZ+vin/pAkmeR96Htji569aSrPQeP3neGSpiJvs4VJ8F221sXJXWB17u
vQJlgWxPSCLQp9c+nDxJpyW62kyNxuI1YyjHvLUBXCYDVwcIisFDyW1Nbx5Uf7HWAkMrDtCXsSZ9
LaLlQLO4Yb3xKMGbki14rnNAWRpOxyciFmaeb9Loq9cfAJNUgFDgkA5Doj14Cgu8RLp45NLLEpM3
8ikNCzbZHXM2XVcNLEjASTSsP98jnykEoktU03GtjRzF13DTIBavhxSxxmNQYzcgMZd2M8ptJFXE
qD5h1p7NJnmXyj+JT2kTWZK3V95azxaP7RSu3ZG/JGDc2gZzLa8D1WQe/IQ6wUSzdt7vWUvle3Yp
gpqe+D+sjMPYRXOaV5SQidJWVCWYazB6Gp5Fpbz1sUB8lY9UoEGi2VR3G6opwywWo4guZxsSFZgX
32oPBysBZFO3kLmwq3RmikDbRmTRi+Dp3isnF5wOXLRG5dlabWrWaFsDm7b5dggIlOjZSqIqbyzR
bfUFO1jJhPrtzZOMkN2Ft6F4Rxf0qqf6OppDOfjRjavh6tOUxjtzVsmd71AehBF87AXtJ3fj5w3w
K1GdHDON0JB//ms6/ROO+oXoCqWDgsaRVBIMVA7Xob01kn9DpdN6qNYH3m3KTWX/Kj4V4hiNd0OB
Iras0zC1Yy+HSEvGCgyNcLg3RZSTtv4WKOkSdudYf8gdfJ0uw/moQZ5hLk3cdQekyHBxWfyrmJcn
XxaKs5SgrpCCFOwj5nWQ8TmwQz1gWoaBqy0M3zMl0ObOa9hv0hBXIQJrgCcnFLEVOyueK/apcbFk
ZmopN9faUCxLbvdnBeX0mkr8yqNhm2rs5F+LmzcQKiPL1Mcjc31EUt/SEOewqrTQvBm1+DYt4aXb
W+2IiuUdUtWzsamZMqcvYRAM7a9FwH/PHUloc1QBMi3u87x0bIwDiSauCI6gdJUB8U6+VextJ0rl
OOBINr9J5P/5JqK9uOFP0w1daV3UyHDLNgIhXnE7+WshqZPnM/aDtAfKWaPwPn0Wt4fabKB/jAzA
2c165jfD2GFfH7CbqXQku1h08xBLCxGRJjapQI2+qThOG62i7uKYK4xOwAFBP78+ddEaPmSQUCfo
LD3MtdQPJSkrxgPC18hQldWLo8ZPB1HeXU+GVONt4TP21Anr7nx/co0ZEdWQ6ufH2S5iUrdFRh6r
nwBkY+NHaWuFHdFSGqV5WOpfOD3DuPa9213WnI5vE9M71bDHhi30d+BRzPkoR+xL/+oZc4RU4PrU
F5sZJ9cLVgkwEHKj7rCetEzSwYKtvNfQHhyLSDttfrwEwKE0pomS9ZRRZxEIEV5kFCRI+tNx+m1b
toUmfqjOQCm0CK+vJyiFN44HwPT7E0NkCnd0USjVFlPNd/DPHzhgjUeVdaopSBcagq3jkcSYpShl
9R8JMvWb55Fgl4+9pr5KHyirw3mg5NwLOjknzPibklfaFgSsiOrdsiYwQ/ZInVjtluVYAJ9AJT/T
zZktUqwSRPZPeugiLe73pCT0ceZx7t/nVTlFLDSvSkNZjkBwMYPNvyplOvCtwpJGX5oijdMXs3SY
pVLlBK/60F4bu3Wc6jo5jh4RKdYMD2a/OIOMF+zeAyL8sn69HjlrWqVPvUQGCAxqOuyJpfH/RXhT
w2JynM1YA8gjsoDCus7+j5sEqyluL3yIBNcaFPpVjkzl+TERi+2J/B8teE5M5MxZEzaXBhgeDUL6
XLqy/+Co1V+dJjnmwmAOlzJBfHdbhWpFIFmZCkE4kLwREKSmNIGwG7k98Ipv77735Gn/gX5yaNrZ
Mfal8qRLOk4uJglynWhGq1ewFWywbcjOfEi3Xb+hwL3/XzCNAonnK/TuuNJWcG+u93kofdly8+Fd
lJ+OLWDOHv542A2VJxeZMjDvIIdDuBu04wM5pV1V+48Z+Wbv2O742/hQROVaLkyWDmTT7DQ2whCT
vpwZQQ7d5beYdTcsblY4RHQnLWBlV6bP4LYvoxazLnOLanAehCJepOSdZ68gbXYqlZwbueVxNq33
rSalWHbUClEGJuln27PuhbA8TWnahxMLrCpbNWxoDlbwCaau9Ehprk5E4XikBF7H5JJy31cywhtI
Ycyf39GuM9EFc/K3+TwGCK6mobMbcKGNRzBlSMlvbnUbUyfZrIPf1J2qssP5ifpvvaohAHdXImjp
AJW7AQ69NTuNpY87g6FjfqMObEP+iXoGIONjtvGE8DjDZ4n3S/3R8fJc/lCq8tQcNE8yVGdaqG0r
Ovk8MzaGlvKQ5HMLgff6T3/zPSNQkwLA0/Wshe6FCOHoJRDJzYBWTBEdVixkIwt3cXccrJ/zOSe/
4D9Pj0LxgDvBDmjHs3vXit/ZbUalZs9DkxO8h9rlnG/q8c0dSHcAHONn4NxglDH6IKhK6/ytpEiH
z+cGRPCfPZw350Grd1GDQVM8caMx+ezbNZHb+nhs5pu/DX6+i58HpbYVkiL6o9M6iXfIvFbgpwgU
WU5LibKdoeAZNWIaOMvfZg/tu6jANNVs5oO+72xLz5n0mKEQXrVYgE1HlkoAqaw2MUBc+Nl1UWMj
puQ5C6Y6fL9vAd72Om7EOcMcAdQI3KaWw2BznI1uYrNR+QibDwkhcBwWpFhdThLBGsoGDJVyL7ok
aExukxpeAwhHrWw+WFpsJUvAJfPKtW+dcQzKj3HOfMtwhSLBRotZvk52O2tEFy61bDPgCW+QQDdm
yOUmultNSI/dgXBttbIy0gJkscwrlZR4WMilMF82BCvH2PjRoPDsgXeXPD07GEU5yjSO3HeU8IBs
ighus4+bvB6r1lTe6BDoyN303XR4nm+x5JOOP3hITNjOasR1t+ktUTFg4Som7N49E0+CmpUw2OtR
eobLFNb4fZBvjFL+8RlRtV9iDnhpVjiqagt42m5/YFiJrn35nC0KtxUd/YCVlS6j5JXHqHGhVfH4
f/ncrWIJ5jbf0TDeMPaN0rJXiz9fmSXzEVuDStNRc6pr4QILtcVbrAawiKjPk2j8ASPcoVSnbUW6
1+A1PHHTtHd90ADaaP3avTrh7GHVhgCHJ5UyyQRTjbhWdIDTxMX2ajvEteCJSfx+l/J1ruYobm2P
rflIXpjYNIiDg0oMOTRIEY4yNpKHI6P/UYR3Hi0cuI1uqUw3yX5ARbi1U83C597qtUgjtsmpb2tp
OdjOPVjzJ2IQGjl4ArdsjPnbSjy0c+YLKhXHeEIFHCF7n2W3soDsqpIoMD/AvL84odkyWSZB+QH6
jnWDVq2DfB1NjgHSxPCOaLkdtOHj3n8z4jzR/6cLcWdadAPpEULSaE21oZ9vCU+yWXsv6+/rlF46
i3uDi3pHrzqi/UwWdWpftqaE0RaKukNgwNlM8Cmw6kNz3nSnZAoZLi3WPjurQwUxKefEi1qP1Nwz
S+HK62ElGr28sFum7J985OVkeBd/kY2M3IdopiXliB5xy+8ihd4lxXIZuNsFBpySGgyKJAUrbBrn
pDwxwOPpZVoT5X0jwRCVF4ho0ikPOvhAmg/OWFH+IbzN9I+3HXStNdtuCe+nFYF8bdYxWYdRtCwr
ujFjcnBT96xrljLEVdrpJyPSf0V0J9MB7MY6pGD4x9G/2SAKLKV7Cf2OXfJTrTNX+UWhFbf0bBLo
IXZo2hYK+q1owJtGKyYt4b9gMgbMy/cj3bW51dfbES7O/17tgio8ID43m1J/Hu2dWtcemBqXRgSf
JaTotTVkCmRlnP8dcFpsdSxDTunlhBXCpZ/P3GCCkCkoHeAdW9hbZ6mAkl8HwzPeRNpsCIZp3kT8
SWIwaTxqicaI1pwlWCq3COLCEa7EGjYzndSRN8eNUUfmT9H8nL78cO3V2Dw4qN8z58aqtHNaAXwx
WrZMt6cN/MyJ2gZqt/zP6H5voEBW2ALEywNpfcR3vnehGzByfAkw+6K7yPOFyxTiAk9OPVuYsnvH
VknayirFtGD24S5VaKhHuQbIU/IPC/TGwsnZqWeBFFXONN/aYhdEUTRx3nWaDva8ESnTNsspvUuL
mUSaUlT3R++vEwwReX0PkUEqYfD50vVt8mNvz9D2zkw+3+Sv0tcE/i+02k/Wuo11JBqke2b+rcVO
lSqHWxRAj2f0yH+y0Qnb+oJWIbr5hkDY5unpThzXqsXARwmBLoCFbnbGSLcCgfV75hYpqAt05asx
bQzo7Z6Ax38YM6Qy+UbzlYRmyeNyfYfxhYNjwnc0O2VZPOje201a4RcSkJw27dxcGoj8JdKiO4B8
0ybQwd+O5cSBFl3/fA+jGsQcj8oCzSYYy+CspH/N9vDfjMvYs4eZ4JOlHBgcBG07cw6oRTpMXzOw
igJNWrVpoevNRh5PDhapBTPsD2UPb7vdrTQTJGYZSfFOS288hhg8sv4Am28DKZR1ec3AsGbB0fTG
hUYis4RMNI/bp8809H4tKi5VMn8W+uQ0uqiJEH7jEU3/AoS+gJ2WmuiJI+c29Y29WWmmn7yFYhT1
Z/p5ZISqIE9PrCrKb819FIeHqUFbmQVzKn9NSBj67MNp7rtFXgxvfKjBSpTlQAhJOqH/4h/J17mB
q6derC3R/VxV1Hc0DHeVLRqpSYThWYnEWHhDCT5eA0Pc9SuXZ9nA+6fJm/BgkXC6wPNwPpQo/kAY
x+LBEZRBdn2aycYaKjBmHJvVzQevaQHZRFum0Y8GSoeODfvDTlRLRse1G/LA++N45Fd789h8pcCC
Qa80zdt6p7UQeFEq4kutPPThc2rXdKAklo+SIDikKWDJgl6oGN4sL1xyLFZpfnU82xZidc8pxE6x
THmeqttEb2T62zGf377kuDAhxqJLUV/YvWIsCmR8p4X3S4DRvG/j9dzmjMlR7fL/Vqiu26GyBGQO
qKS+9r7l6uFdKFJWYRpGhFYGa+dhFICJ8iSJldGkl5CAu8DVY8fZyDMH+evdar1VmAYqbT6KagC0
8WYhNNVbKA78y1ri1fDxh8HAkshuQiWnvbCuCE6YW0B1yeazkJxdtNaiA0eh+F5vEXLCWdUgwNyr
ZA38AGDDBYcrAcMbk4m9JPOT4fFh0/XS2QueCRBpWwHBLBTj2kLRCQws39ZOj/HnYlAI9UIJQbVo
ps6WVX0aIlJ6zcbKlPWn3GF/qcsaqiM6tldqlT9QBpwK82qo/AYXV39ODOQLRexkxqKdx4WVeIys
An966ybANvcV4FW9YAMPA2631laeBdr7pgL9NRM9eMoGttOucKdL5UvRNI34TgxOoecb2V0Wzw3/
sk/UyVOfnADEnDZPry9cst8eseq2Bv8iJdhw6wWs8gvd4AKXmoOpQhNe1Gdn8tJPNSRl/+vNV1fX
beIPjEBZ7x5M3AWPtOjT3WQM7PesEIlLNgQJS78Sy3QWPX610vUTFa+ZSxjSPIKheymChx+yCNC+
gb9cJNIYmuH6QvMzevHQsbf27mXKDDoBKa087HiAKzu8IF/SF9oTIqJwwKss4XJhM6AjR6zQJe4c
qp9GSymAUK4olTDv0kpvlBY3mI43oSFuieqMjJsAC7tHmU7++yfAbLGVGpw4Tnc1UEq/SyCva8kT
uy0+bPrFJKIf3M1p/zRCjKraGLfjNv3qenDkJwLMyyqYCrt3bGmODbBrnDHx0jlvwzQ7A6bVaz4J
b+9hnzozJ+oN8QL4EOeYz1afygxBIeq6LymQGxrpo6L52OmZ5GXx1TW90VL39dU88IdAz1oI50E/
IQVac7eFYp4nRZhFPaxtQ9UAuZc7zNUPQqoo2N4ctTDDfpc8JWH5162F8jsOnAZp001L9m4PEtPy
MQ/Tn3PuPuwYlKr0KfsbVWcKj6fWcS2JoawzfnLduNs3+m2vLKU7KTJpMOACunT13FMEsjZke1kY
PLZ9qcY6jqwi3OjqNUlNFCX8npDVrTjETFuKH2LhEevOSel+56eMjTwEDM789N7BGAGZn1Jb2GNg
m2nvE0WmqO3hXYA6IFxH80qQWQYcD50uFQVwkj55pj7+nNk+l+VQz3m4ArCIgnIywT7WQu7W08wD
5YP2m20ENjJhOiqt7AYSsrtqnNnfKsp2F1ehs2KMSpOT9Vr7mWd01V0UePiZc0bIFJNNJXW35FDU
ueXoOb0E6GqIeSLGAPdRKMW06+oiayCbcIsNljsbc/rSf/kwy1VUWs9CRkkADJE0Ti0unA7ruaxm
Ovb2A7zfghU4Nkug9/RJTHU42IraDaNTrLqrGTjrvqTAbu7VrY+jMLrVbn0C9N4XnAy5ER+N2LNZ
CGGDXPt2Y6Zq97sbRIC4hhXiQjKgmyqW8PqvsrIEvS66yMHT7MzO7pkjb/yTze01CwWxfETDycLV
fbAaOyyOsSS1ekzPkv816ioRX7+7tNYIrx3Vn9XWDndH3i7o/aLotU+zzKpJ4mOZVhLZFNe8unvl
+HCuYkIBhjjimI0aZw3BEw6RDOERAdHFl0ddncLYl+iJzSpJbt1uRXSzO41tdfsKem7zD8fxPzv5
1IQWzLEP7sImnHehPfQbug9x1KhXg9aKBwbc48DeFj7648ji4E/Bfj18DWJNUd5k1UxfziN6YSbg
BXWVF91fHwNmOPmUwg+xQOC/8TONasUladBHvYswe2l7UkFpnFRUSIltTXfgl5SyfoGegD7PDBEQ
An14Hbh1VusuGdR8NXzrT4OOO6WgJvtAW0Qk6EF2o/g/du5UEhIZiYrt65NbOvl1XaJUuDcA3JMW
tp1JutemBTe0t8F9kcBm5YoooFAHg2nHjgQ+AsdVuZfhx72Gi1aQaiCx50uQKc9ZOmWAul5URPY3
Z4DOhUDlFCLd3KxJfSzAfCcW1TDYDA+fchCPkP6aRvvHkwH8C5OQwmRlkMH+e29act3mpnYX7AnA
PgQzzJ6kt6p/af5r9PlR+3pHu6uRzLGyKL7hd/9YkLdUeUojoB9ZcmR4uC+bDLOs5TjIdqXeDFkb
dfiTwVQ1NnG0Yy6f2hyhVsknh1vQcFRTVJ2wWLH8LZWRIwIZk32jj3PYkWePlLfeXlXE4f0BIuit
NNtuKl6o2FTmoIuOvAnKhleNHmIiQq7yBRXaw+TULMOy7HH5lnISj7De45aefnDD72Vpr/X+5gYN
ffqZiN4EOs5cSOTm3eJlaFZKH/etrISRxms79IStFdTVLBoPbkithxNwgvilD9vkoPFpMAQLgL1U
zrVt9nADG/6LU3lcmJ9nqdYFBsDv/N50Tw9C0+jHQAINKzTvPGRQ+HVQsFGPzIu2a5shML9GzuVd
EuGyhAYJGkJXTnP1rlHpPytaZFPhDpV3qOOpgohVCPLjbJEAQljlEozgXHmtyApGVOjDsvzmNyJl
utRXgkfsC2l9VVwWc7IKKAN9Cd2+oCMdcT0Y35FE6IvJztyll0x5ZxcoTd9q3+KuKhg54uvWpdzY
6KdEgPBo/RScqvrtuKegRHWxXxjC52CZQs5lPQ8SHFBNypCEYf31a95YJuk9cW/Xt5ep08A3vNRh
AEaNAZfJ8FRCYje35PjwBjjoHUi1IVQR3ClCXOkOH4E4MdeLJrwDNMlijHt/tdZFb+soXK72l0hj
8qizys1q6a8NfcBsH+mHMSS5MJf7R+AJMIFdOplx87fINC9SEdeSo+5z/CHo5BqQga8tmqChvmXC
BF0xTbQckWEupjfFBaTqsBfagCYfj+kL+hcjyBi3sHzce7LrUToSICP/9an/1r/CjwJP8U7L68ZS
h5fe3M3yJhiiqtSblk6KRQTt24+JZZolQZvotdtniZbWZhx+WSCqE4l+kk+L7u7ssOdtPkvyH5z2
SJoK5Zig760gToVVVRrkxTe1T/M66v4UJ++oAfgJptUa0I5726knhP0tatB4lT+MBoBM2dp9v9ct
G47jKHPmdqi1vIFkl4fSWDg1tgpuRTmYmt9lQo3UtY9q+xzPPtU5eTnmhb/MPdoi5yUHbjN+3XpH
pU3YzGqK1eOf/tKBLUn9RWrahD8prmHlWXeEG/4JQ7NJIDf/8i9edw1xwXULcbrD90/050oKnX93
Je6kbvyUew9zO7JBfbNXeEfGE696vf4pqqHuqFPgPL1VNiG7u5i+qELVWaF+hAiMj+7+qv6RJVj/
cD4Tt1RhjXN1+Lpu0C9129z3+WeaBgLdX89ec3k2hpM1208XE8nUPKXuhS6rjbBr3s5LBDiH/qXB
QJLUjV8gwtg/+qq6Hf/lLGdzYMl3A6qeQSRsdHysm6rF/qxyM4b43O/ih518kslEfVq1Se9Vmx+A
fQ6lSmU4U9vodQdsEbHqg+I6iR6dS4aE5EZiwH52mf/ReOUg4SiYW3cxM/ARRD6ff3eCwEeVquIG
2OqMpk0acXB0eAfem2bQoTmvfgpSLs+wyErG39w38tXr64A9Sj1LkXyfGYHAuLnEPc4FtBFKG7fn
zPPzbScQgeL87ptQMRm4NbLx545yV19dxBe5hu8xcq6lpaEdcBdjR/2euVlFXbC9GdswycJ3JQGw
YqoHlYYnLzP5JeRQfWqL3wgj8uTq6OV8nw8yIuqyGlhRYzM7Gp1WOjNk6A9jjaGH5OEuOiwbRDvH
iyssVClrd89XGX+UE/gSHChr7YiRoslj7rHzaju+iD8mkKBBwULOKGcXy2e0mCHX/jVfxX6uY6ht
nOC0VSacXvqKw05JOzgZKsb0l48ONwlfLKPitN1l0zyZk2gELDBKIw6YRhYGr3dWTRrkXuLFwn6h
h34ZFlXe/+etqcCMVS26zPuNM4oawRBn2HUt0YBzwDUBFu8ktj7c45wNem41B1Vjx33T7mYGkecK
1X03kapi/jGCgALAukm/GPXJsbVpb4+1RsISzL52Me3zwZuiqL2mwja1ziNGZEcb2zXVHhVPerTT
4fRvQoXWQIFSMmWZ8KTmN7HUZLkdsGx1nLyO2FTPNd4EZg/+RMmvZeP/n2xjX4ODAUnPeHWqkzTv
Eh4+v0MeQs4IAR4Hy2xBxIHWbBYyA5jEiQ6TrMMRHfNVKIK1J5JgEpwvRSaXrA7b+yZH8DyQ1n/W
4+Vn94/r8w3wH0Wx6HALJ34D8LDPUGTMjbwiB+ZeHCvTWJtqNvETjGZD9rQcIWgWduh3TfZvLGEI
cIrS6NApWuRz2NiPP7wcowFrexoq2Kn487ihN+przwVFKGV/qYhvI8ejqM9+KIrRFeTp0qP22XSy
FP7e0xg2gseu841+4O3GVBKN2cokAmHcV4nGNBDVfcz4rC93mVz40WIs9eKRdi6di/w8zxLyQb3p
OOKWxcDq6gcAxqB/KAtPgDgN5NukO4uaj8JhWjvrduXb+NNJ5oTbrUCpwQMgTyr7f9NAJ7TpNtS5
N5FF8Wt4QQNYFvd/bAVQskYQED+LBrONM1lx166yIfFxsLxOaL12nnV9wBmrcGTrKI3gwaJ2mY4R
Saa9RTiS9wR4xUIk4kK9DB3khMKLZv/WsH3lCG6tiNrNbIgwlHXrxnlNpKLFJen9RcxM4YJxEut5
fs+19AugO8Qx9Clvb4TKko14/eCAeDC/FJxR6nZrm7/RbFfH2O7v/M8WcmJGHIWsX9E9VB4B4Y6W
RmJepLfjkniObiHLveBJq7b/gqiGW3kreTHeuyULc/nHqWJeJsMfVDFtVRBdjjuFsz6954hjUhnY
GJnS1uRqlqXbyWqfgONi7Rhk/Icu+och3il5i5yhj/3XwuJ2vZcQ6pyJ363IaY0Xuo53k1I59+xy
gmwJUQD7DGd+gYcLp4wiaM633R9sME6E5JLdB0W1MaPpodD5Hql8turc/VLrHTAOLeloY/w8HWOG
hL2ZTuGmMHSkRbj5dJq8zkbWRxtjQQNnooRwO/WCBwTFAG1i9OEZ1Wykdn5H6Vx/Fo2tQ4THSwYO
+k/PZiXyksHqTRjHMhv1LxXAtSLqXvorUp307057JlmL3tBnzvdg0r5Z76/+OLputDWzPlHwZvsH
fDk74phuxV+E5ramLJCIhTb0MTOQVi5TT64t5OFTk8OwQntD/a4h3mbYHwvCfOC8YdnGSntxltQm
ku5U/19kKe6OSEVdA6PkR0Ymh9J6XCFWKZrXO+pN0d9T9+1JaCbXyriUs1/Mb6t4+iTrxWYPEJ1R
37bo/C+AOOewvHpdXxaUxOLKqb1J9XRwgtBPaQKMZxZmv+LiX2RU22CB3HR2eR9HSjQ/AgTpI3Z3
2L2EQZawS/Db6YliOlyrJGen8YhyYgKl+jI9gR0LGI+5CXE+RneKOTzqsfzM3kCFsrSpUz1G/GtG
di3mPIPLczCn5YeTudn3JOMcQNQblthlpwAl+3sc2IkoLWZiQJBf10LBQXLwnGeqyzCZzxI9rTB4
+6YtGdKXoOpOkwb0kGkadSYRsuSDckc+IfdCgGwCZhCIUwI5QVMxeTF5Y2Nod3ys2zOT1/snPNSK
8LmBaytJXQZC/CX7sRQLohPEpCB22HT4P6E6TtcRpSYhcqTCFuuqQsYqbZYK0IH0E+hpKBE2E4M+
XpastaSpvxH4hNxts9rSdDcMPyTUn8dcg6yfVbay3X4JEdFa1vwsv7pmEnsrQhp/FoxEB/SzHXze
QNfyTuxa1wDsfa99r1cCYKxaZYTAkoYta2KvV9dqcWN2dI+kxX+fQdADISw4YjLl/FpMHfKOuDxH
ed/ZYOjai2EhzJLokKalaIPAhx7XhI8wWpmKwIcAvZHF+p1RXqssWnmzvkr+Ym1/woeGsUS/j4ae
+wAB2QT/jORDVu7olN9AgH5Xj6IY/YBkO1pN+jqhQLa2vr5BnEPLT0k1/fYyhnqoE0J/VeY9fXt9
AzKS6FHgGQOcuSpTZoWyoFGJhDCl2iogAoMkvohyZMLyXJME55BrB7TnkpdcS2qAlDur/WLTruhg
Fu0BDTnSrppTa7zb6LA6rs8mwKh/+jU2rpv2eQ1b6DIf7hIRSVyg3jiOhdR5ZOt0NAIMDbHo8zTm
jNR+tQ6wJjTyu+1eozGMtAS6eMk+aRS4uVXVNy2m/mzTulCPekgGpbn1kMOOcjpXD9TWmY6FbHgR
BtjYFGoFtS+SakbBWGYJhccLM50+S75y4jAoVWCmDzRF5NyxdBkA93SEDCWKvbznjUzN1oTUocai
ALwAfqa2hUStVotnRDKo410R3atPdhnKI5vpds+ThXDdCt5G7J35iH0SCVrQs8EprnpJFKXZOq+A
89+e9+EPM/XxsQlnbKcMrxW2yJmXgbYb6OXuCeyx94KO/ypR+qzsynLxrZLd/DKrcLOV6VhS4qdR
FboSwjJ7VZ4Sb820PldCUJmTnAJ1WfITCYwOiypmhnYp9UHiBEd0VaNRQLymG+6AMbPZ17XVP0+M
/jkubkqNRuU8cDqfvb6aag/vh9VOAzGg30nnldahIw6pIS7xLu21zmCh3UiFgUuYBRgnSR+YZVe/
rUiPR5NbR9Dw+pmN80oyD96ykc7zAiSbNdonsUiUMnn+OBVlLYMFgH1TNWNmEsmE0tc+Rx9xiloS
Z1fqOq6fKnHLm8ACeJOYOQF27Y4B9b+GxLswiR+HyzsaU+QmHI7p1YB1z833X5+w1xUtE5iFZwQ9
KxrhY+VdZ6A7A/s7m7lGAfMfEkczl2XeelMi1JMTYW7hKI7FMwbtLtWoXzWDGlJgVbYYpmpBIdAq
Os0mXrNZDZ76cwEq54Xehlm6dQkkEWsSRCAFWAemaAR8bWN+337ml8gEWTRRZ2qdVBhiM8h6CwPj
6tvLpQiFlLbMWb0uId/j/mu3YnCyatiRSst5deNB28iqjnF6ICPt7RmkgIJYhVtCkSnRyMejpCLJ
+/B+aY2cChPrc9uN+7E20uNz5jSbKK1oK9vMjTlAmAV+/6kc7QFToRTf/Oh9teCojyLSM6NfHjg7
UJM2M5jmgXS76ufpnIdX4+y5Pv+0LIM/geJY+i6b7o3jvQqcGce+pQo7f3yTkdQS52/zfLCqwrpd
ap4iuRqOFFKKUYj5v1xhPp8ufB5+hxq4rXC08t0rKGHCybvF/fAupsDUwvNNw4+eQNctdZ4j4Lij
e9cvh9SNYOcXwSSOmeQkWDxolq1N1Y/ZplMQ/YaL8nAaBdrjXPlv37E8uYojloh3uK1iYWa5Pyu1
3aGsWPkhJX0yYBCo5THfl9f3b91uM7CwW20aYCbmaJEH9y4lHflmoeZfSIbsKCgCPbMvGA72OR2g
7HaLqz5IW3g5hRDdRHDlsQpVUPQNNQ/SnqZwTRG4W5vN9hsYg4Hzc+tW8O0OKFH9aJ6nN4e+SXLa
weAQTh5VrtfqVdv18npmGCH58sFBjSkpgQnfIMdt8nmvwOtI06xZwBe3CyRKGbaF9QmumNFMCBVV
R6zBvjKF+60l43Y6KReRQfT8bYUbZff+9ERXooJR0f3nyHwk7A6XHobfeGRto1gCTqZwcLqOtWgi
MJjC9xIIpGKLdZcoSHuD/VupkmyBM8iEpyA8PtndbmoantCc60sm1JvKnat4xDYTsHHdfK+GxpTg
XavpnnToL0uJUY5tzc3Twd8QSb2vpwlUytsiJ3UwoMSwK4RV+ggnu4PU7DV2c3VHAkE4xQeXPjE4
AHywmEKC+EJDnt3IIqyEI8r+Jl4A9UPVqEOHWepjnov8XWB/Ye5OQgPY8QVfLYOVKlZDjcu2QYbY
5FZ4N/xBJfauLxF8V/6780Zy9cPC/K7qux9sKq6cU7Pju1v3+xtQ//AeXetXrkv/IynzqWwPgzbu
sYCxh+GLPRp7o753iRuEQxS1qlqR51sbCm4nK3+1TYatgckZfW+KUoWAgqL9uYkwWuRw8TUPy1Be
8/wMJ+UcsHOZcJC1xpN5JVVzmPBc7Go6J26dPhfveK8kI9XYbxtMtdJ6BiEfmASH+S8y8/hPc80H
X7ca83adSMTx3dgoUrTuvapYNqLn5wDhq1+qqQCbuOwrfEo5jk12ZBiuteEGT2YOQuvVyldYkdfY
zHNLUjaMJ7cay2YLxywXvFu3BsEcj6mY3kaP57Ea7TQyKQ+9BlOgMOruX7LI96gyGTJWdjwXMK6v
klbvVAZ0U2LxP+LZDo1JlNF2PWZN9QvBveP4QLAPymrSuR5rwfhfNUJZWkzy3JlH/bWP4sMv45z/
+QOTpEZTcduk5l8LOYrT+ynoX7IlDhfIwOT25CBq+OFI961OOo9g9yvw8nR8PlBU4djR3SZ3dt3A
4R/3/idMv7IyrbZ7vRNk6vt5vyrIAHJZLiEJmCpkjTmrum3jsTvsAe2NEs0yGyJraFGn8oX9LDhs
VaubpRkElm7xFq603TP0JQZG8mUcNGGR4CFKAobWPO9IqHy/vKVgiZrkwQ3t4z7EvAY6ev1BE6ut
9ViOJkC/lBX3IwT/ZoHZ8gUOG64wlsIBBsBqJTIDcqje51ayWaLErPfzYRDT/4OQdegf238DsxV7
FA2przDmOVaw8aq3sH8hMD1ZNWv1jA5oEcTxnnrO8LyZNNOxbp1H4gV6+F4RhlQRdFxqy895WFzH
OY+H6+93vbwd2lP0WXosSHyP8zfMCRDVujVGEJcNrhPwvek5l18c2raodSUTa+INXmaqT7sNpY8A
O1wLdJ1AecSecgbtpjV43nnwRhfdQcGLWIae+VTLQUewZcMvVVI6hVXZ77Oh9p9twd0jB3PWa34D
9uHBWu49XwCQlMlSo9gUCHdN2q1hPI2+36a4CudhIjJfoD+0AYvvWL2zijU+TE6oaUQV1gzl50jg
at0poeYHAnBZTIzss4QPobhhar5WGy6Oo2WxoN332bTq2FOkCBrm0RX9vffaNyukMp0Hxdi76S4L
cmhj8Y7btBu5th+EoUJ3VgP7SNxL/r7U2UoBPRfAEW0p9sfXMSBSKQLHZs/iT6i4Tt+kQfSIcx8P
SfJQ5q0yRJ24njc1+uAYOPtJFFNCDK540o98bINez9PqpPU7Z3ZRriWjZwJqv9BM1pHcyO+4Jhmg
A/8xJLQnWiuwQL4xlgUwckcSKTXZPGxlsot6Xr2mG5v8xTe9x8Ss0kaFtY9Rw4Z6KbH9S5ozm7qA
X5CW7J4s+DKrOl/8dZigFZ05G4m29DjFTEgfG7S6bbncHaSH5y4RgpJz3Y//D0Xt5ZVR4VLVkB7e
P6t6rk8Nd0z4AMCKZPhCm6060/EY7SS4Uc8EFEgKF2MEdBseqPFBOusaC5/KjCEZMGnUQmtaEex2
+JMGEGyCQPQdKxtf+QFP9p0rH3Wce7fcFGPgygO3ccVOIysvGV5vct+oUvAIdBRBISsHGrZ2jTxc
SBlmbKshAcKOujMoOABNDxCrrAam6PmEubU2Sxpw4MDD7D6KeA9M94ahw7r3BlZhdn2+LeB5AVf+
kRrvTl0OA/JLQVlJng8CIfLt0OHAgw02FNDuRlUycp1nlOWF+5f6dUIYMzCehmmqJapW3oKJlpyR
ISVaAHnmOXXQq4LG/H/X1+ng6NejYZtbv+7mUgYi346+Dfc7eXF6kvKvM7XgytbY5s6lcCI0OZzb
jTL36Koa3BPkEX1yql0YRMMdCcCbB9OIrlQP4qW+BC1XY2TS+khPCP32XTEmOBc6ZxPKxj96qINL
7B0Ax4eMT6Y5kER4HD76iMEV7NVOnXDt/VkrbO748Xo4z03NI6sW0whzbOtbfe65qVb/j5qv2HX4
GGuGFe72uFBiFoNcMrn/uhPqGX7iiuCFV6hz0NKHZlJ8dEY59Udgj4FI3n6+DaXlHx1a0j5++diU
bdafZ7NWg8Wkvjm4gw0N0T1afpRdW2QP8Gx2u+qY86CA8ydwWPh2Ohv19ZJ+yrsZzjoXMwBnVuOR
ZfNB9U+miLlxTrPM/0kb7h0zlQA2Xm9zj3pCfBcjYVufn42k4h2LuwEuHi+cdtbtqBOleeE0z3aS
f73OWqSwQCYXTT+WB31ErWp4eA99lrb+wQjmaj8v5lwE+azwY77Yq1cmr7omXpV2q/I2BDw7CMTB
eUXUavs+uvCyJUfykcIVkFhLQ43D1TWp0WMVD2gwpNLD8XVSHqwFp61FNX5lOOUuym87oSnsA7LF
RA1WdKSXHFfUT61euAslDbdEDeHBE66YbuTO2WXvs2EAeH9JvFhXXfLxOlsj+MIPWDwTwL25kEgY
+b6/lGnzekJmvER3JMRMgHek3udfvyqu99x0lCTwCb74vZYgXViWbcoZBgScs3RF/ie0hudGPDYL
0VlohJHjs/nPYNASNoHI2jiQ6AzcW3mILwEfWoKMRaTA4ZXk8b0G0k2BfFjZBBhHPViApU81Isb8
/2W266HoiMbpBHnbXlRE6PlnANfflsgM/tlOgN25gOYGbJNehYZHFaMiDM+kfg6iO38+XWJGgndA
YUOZbwmNdqxBWIRGKz73z52zQa3Ag8rZgnchLEBYSfPHMTwA0KyggahFrXlSYFMgZ1fDn2+A47eA
zhkzMz+KPYQyAm2sVAwqSBnSvWfMyEai3ENeYJm9iqe0ML6mJYFh9gHKUbrkG8KDiBDFXg6/focw
VFT9jxLwjJh9jYD2fLqhGqO6xFQBG1JnVHSILPgL0QrUQka9YOqp4CmQTgYn+djZ+hz5RsrTa8Zv
z2GlxuFjFIKQWUAAbgSQHHnP6bl6guxCLXX+maKp8rMbEkk7Adp7ZhdkaqLEf9bGQ8G29DjPqh//
PiZITAgVdKe3HLkSaQVtUsMeAKjJofBKkMC9xEdpNXEHr7LvGYNj9+Rz3R/fHvOlgKLST9TPm7Ez
153EdbmzuPHm7qB6pOLgt7ThxkoJ8LHBdPPuAacBUUxx/KJLft9aG4IAXvfmm6x0iIZvw8bJkKWh
K1718GsD8dym6OAAugJ5wj0ukxOyibSQ6OkhAbwZknzbKZ0BwlcKCxC9aOD0eL3/1Ti28vgD1dRC
T+lvc9oikhX9UPwfWBU/3/Rtmm1B1vYMarUp//EUsJjT1B7RyjYCvepnFqMYx8Tr7IuSwEujfuV6
XzPB1+D45qFkQbE3EMohg8tNHgV82lX55lE9FJMo7ZFWaE8EkWXlzNP1vY5jvpbUaDYG2N6hrpbF
KtUqYpZkgYuyvZ5cV4W6qKSoS96JAuCO47qz8tZwdOAUdat4so0FBb2/GfYRf5hREKbuEqx+VnhV
QWNPPclS8mfg2AMkp3GFU1DSfwdxZ8qZi1+6aHPtO8jrEIrHd2Qy8K6Wg98aQfG7LwEp5DgjX00l
STPblNS9ehY+hcO6JSE/hLwmKJ2wtmWs1LUfR7rRlsTfBY7c5xMSQpBHEg2tqsKV+UsZCvNEqIbM
VsHMOHni8RiuE57Lj4I7HYgUzqfSXfJsnYBarBLtZZOO9Wu4HSOgQZlkCch1r6ovZszBhaotNNDm
ds/2JzWShmsL+YEYQ7PLe5RdmrK8zt+O5vHeENWOazVnq47aErxWn6X2hNB94iXjG3QnoHubjzZ2
iSWuKuoeBHyLd6roAhzZG5XLcezSYpB+zuvDC57dKz4wEoH4rgDib4oQ1Q9dzJEuxfX9e1nQGjbk
Zy/zGMWVSSg0+q6vGetSmV5CoO2rQdw4Ab6iIHSka9WnJZRzlFtiZTT628CKGGdad0KIiOXLwCY+
+rDK1nNV62vmjQVBiF7EJhW8Nkrnb0QkNTNlAiY8+q6cyBEptu0Uv7pS6tsqtZWYe3bx/NdW0DCJ
M4Pf7BYox+P8Lv8UZjQ7s/Opy19NEouHiQJougwIc1azqW6LB/Z8L87vcyDuzcqkjEfRea6tvZMO
tD92T2SrDXjM0xhKVQogQSbgvY9k27Sh3Lp+IM2L861bRtMOizEtnGNsPES/Y9+F5nP21sPRhT1+
RukNfU62y4+6+B8BNPnLj/BIhVN2KL/wt+BYvvWcfQrHsC8RFDsnib51nUF7D+v21wWCwWDU8fuJ
svl4JOxNC73DrCq9zQW28A4pkakDOSVxlK4LdRgiYGMoSdhIV+yn0HJBCbw2OrP3yMTn4zEUzl1W
HK3DlQG/T37FGR2wBrfk1lG/q0cY4D7+m/l+HhViUSa0+bojZtSMe4BwySBMzqLu3mIFZRI0P5Ar
vsNjwG6icLlO8hySMXqezydMjY3NBFlbkBWsWFamfMLhXEsay6Gtk4N06Hulg2YtrTZ75saJ8Jmj
4+nxV8M/oJzm0Qgx0E9hrYWuXEUxkPQxvD/sBkt90qN9S3wxyUSemh9qVLJqFYjMaxorlcQdQ+2L
PTrx/bejlj8tlPj1EaN5cDzg4BLAjTn9QD2KfaHeVu6vQ8xnQwNPJemzVW9QeFDkDlN+ULJ9wj73
WO/uEkLvoF3FjdXBmhea28tQBmuLMHk+c4u+9+231b9ShRYRWUW0xGHdWmDSTFNUKk0LEF3qO4Or
cO5buzZas04n+z2QkT2wtV90/XYxo2Jdn1z0lAeaoEGUxI44KLKFcQgFySkRcNjMNhEghpTupNUr
+DDlIBl/gGkP2sZIMtgBwelB4VhvikXV9By+sAzQRZHyIkYJtdj5esiCWYIzcxUWF+GL6OR79RlU
w/w1aiUkD84Xg9X+Ftga2dnWt0xlJ0JgHmZhPdZYfMDuW5PEAHpybN7nfJEkQbHQH+OXZdhg/aOT
GZ29S4d9m+2eP2D7LjAaZMUifLGqyQVJZMQD517XvHdZE9r8t55C/5AXB3OvTbp5aiBg375Rx/48
mTGRnvOx+VREgadKxS693Sc6o/tvsUS1O0+gYNt4rA6dRP/4v0rF1rKq3wwFm0UK7j4zoBk4ze3s
Bql7Nz1g3ttOKGyjOPQyW9K2XERCOduvOJ33Z5JBg25v1uuPotD8jvydmzTfOIpavXWQmyQLDE56
/qdbj7WPYTMye4wvqXm4098Td4YsjD8W+SyYW4wUgkMmB+b8NGlmmNuYJnHnYDgafUPN3xmTfDc/
t58ceTm0bB8TYCfUY6WZPKKX4mun7MaCUFVl3Lxgl9ILqsgLLsadvLjivriWsB/ExhMrzPTmhXhL
eAFFRepBb7kVOKqqKKiPEvAz93s6nKUu56Ro2tiqMBWdYoLn4p6j0MIF68885xJt/PTrmfgSIhLk
1vFnSq1zzHXCvwF6oQ2nLVfVH27WU1T1N7cT7z4p0C32efvKm7QGy7Ina/17r8XYaWpNtaW+lZEI
Wkkw/d4XDuqsGHleiwdz4BGffmOLtnXUV+fgoywhwSunE37QE0Zs9DVQFwGGBrvvaOFUSH4qr15+
7gNLbsRecj05TCw7jc7cTNUCkPhvxgJM6eyuyjd3pfPJXokovZ62Kqi+EsORfmTMu+Cf51yweeer
3CukPv6UZGsfJmuhxvIiUW3hcgJIMGYo2MYq4E5l1iZegUy+3wSM5FmhJD/7vxNbHa8KHaV2zypX
zqJm47fqJ9KFmU/qI7OXQhNR2MtFkKxmiLhhtsT1Mg3qq1UBrCYLP7bvpul+/3iHdj7MNZTN5kbG
C7e0bex332U+tAJZih3ZdIqv4J01CY3/OzKM41Ih9lVMHyAmu4zEHDoz+VwHYgsEuZQ2X9InO/cb
tQEgwpxUcKvsZIaSLrRNMVuWoF7zyDD7zOt3T4DoRu3/LuKXmBTSyCkRZpAMP6u8m1BXC6MV75gl
ukwwfkT/o0Zq6Yd+Ov4nf+wCPyKT3A8bIR4Ew2AsSFcEcMiiRUH37pHNwB6iPcfEJtFOQbaxuhn+
W31FWdt3SxBbetoFD0eIjDkz4opWdQcwxiT6x/tOdzGV5XEPhbnmyhqATG/MnG4GZzdEGIRjbIH5
MQyj74Y1gsRuFBXOGywIYCOrQhoAR9TxuDcnd/iBUNfRah/ajK0DY430CiVTgddwlpFusVmlOMzQ
0YnjpnQmTT6TEwBNSKrnK/JyzeBjr+3fEg+R2a/XvRsO0cFTVFWU7f7W4beD8AtnEHJpfa/eYp6w
7kc9cvWiOAeqFsFHnyexmudzscr39obgj4qRZDVU7gV61wMb3mxzV5FKySLWCfYp/LFlnL7J71ak
SLZJuN619Zv77ONxX04/v39DvPs7/ykFRF3UafAi2yYEVP7/+qyFifiUszN+mICR6ENxX05WB1Ft
X4CUymbKwYfhWHf6JrUPK3kTaIs57vYkZhQ3x7sO3KnExpDyP4Q9rJMc2WF7z6WWUHbW28NNWxwB
K+RvKeKCaoivW+PgnnDnDWfFWOQKgYK9bfgHfYBgetm2CWJahxi1nAeTIQVERmyFJF/OhZOsi3Yg
wZ28G3TZocEA2iKa6l/n4lPGwwwAotNS0hu3AsF19UaxyElBpaC6y2sWWnrMoKci9gsWTKF5IgpJ
5JZImwf9odvEcwdRyuaSvOrtlFY/uxXMr8Af0/L6SodbnaJX7lSuj8j6iisU+AHOnDM19i7+Dzpy
SpAWsZhP3jSH05VC+xOmmY/mWgSzPs8odrj0C/cZxzZ2KJParbMTqVFcREf8A8oxTU4mSM1njLxj
+c343gGNOmoYE73MZF/zMs/P+vZ/+fkOiawRHBj9HuQS7MFePfDVjUP7bSiMfSBQLr9N1aavi0ei
NyVX7OsaZgvfc76o5c7h5Z/bavXy0Dq4q5f6Uj1hpQQQcK0puzdhT0fV5bp8PA/s63+/puAq/L5c
ikZfMxfqFcQQyDn7Z3HSlBYd6BeAqpDfRQe/aWeRrO2+Fp7sWvcc96KTGbpjMZeDjyIS7QrvScRu
a0a03f84ECQCkflwfJnH99+NltyiVaoa8PmIfu0fsI5YaPW0fMo5LPpTamQGUX1INmunI3TQ1TDD
+vf240UvtXG9b8iLTU/0y6g96kkA60oX3ggFIqeS+1DxQfsY0oAhI0qqSmEF5jVNi+6nG2ud7aws
49MD2Vh/Gz5f7kCRCfWSlBEzA70UX9gHNxcvooucj7zq90n7iTOPmsT3fsCGKYbbM+mECvRYO8be
GTROpWfXa3JtpwBzCKlPZwCn6ZlopcmMtgiYDicQTzTBeAnWfR21pZpaFAid3UnHRSWFldFnijI7
tIeHMV6z4SQMl9csAHShsIGkmV4P8xaOe0LRHO59CLwGYfi6jUATwrPJOVufEtqMNXnRE++EzyQ9
ANpfuDRpHjJK81Yn0x+We9CjlFa/1vC/zAVhAcIhRa7AzGU1giGwj32faYKy9VHW8AE2dQqXJH/A
3hZ0cRkBOfYCem8E6KeBupSlIZc4qYdIZLZaf8dNWujZlhAat+mu5hWvKIo35KhJLoMKHDlhdAKe
LQx7+G2uvFAv60+Gw1l3K2DB2dWu8cbC7Xe4IbwdUIc4sEZ65nqmFHeoLTRCjajMVZHmvxykqLjZ
nuF1ZerwWa4HSUtt3UAI85NacrHQNcKlseQe3QL1ZzZpaJZ892Nh6eqy3VCoWm1RcyQmI6m4YcHg
2Jsm7uljDDskl7DjHDfn0mvo0BRV6gQ2BRKPME38Hh4QhuSxntRfVvHQAmImF5aKv573Sn5gxKMM
jXexBAX1DMgPcQ/3vB1v5gR0IY+7m77iXn6YvSrMxGfEQtnuiyhKFFQFohY+q6CEzq+5sTb1nJut
l68i2O9MafFdDZ0YKQUTWbT4E+Hh6aPQdmbYFPpaSSAgBid1pvZwLvog5YofAWbfo5Wt8d3BT172
VA9puDZ746e1aMb9mNre1ZbVOQhQK6HI8FgXQWor1L5iYg5+z6ZI5ET4JTFSDJxZsi6IeLmPJEKv
Ai7xitOp1waDAIj8gy37yj+bQqlmeGj+bPpwL+INlsMsUXlczXQlytqmYwqWj8Zc30aYKAQJpTds
/saKHtJVzUXe99j8k6jWLWqIeLtJMqO23hZeOB0sAFYlCigJbaXLvut/Yg6gQvDuV3f84MjjvEci
b1nw9oGZTQJTI0Z08ZdoqHL7wX2DRzLL50f/EoBTtlABSQUBqC/j8Jch4O34FvySDjwUCBFkwUTw
NMJxvsASlfwDqMhHoXxgBLD2x/6rnUMNLL3V9Bj5TvLpuDxuOHKNKmJKXWtolapXMcf7/e12cw6A
MVE7l9gny3hOtWk4E/tSjRa0/Dz+OhQ7xnPraOc5guuZhT0WApT+ra1c6DlctfLJjaOdvstTZ5LL
Go5ufOmZxWqv4eTHq1/IMxTRKe973HPXja1iBwZmCBYZgjKSkCe+9aJOvZS3cQiW9mBrdDoAnqDK
XrBA/iqKPGCkQAl5kmIWJig/Oquda3wzGG2VVVkydRAyw+6OSB8RFQ6fRl7EjjSgTKjO7vT0IYQ6
/vpXN2Ld4MkQNo0JCnTK7R/44TVtyduJOL/fOe/BFfk+k0YH9CIOoEIwzbzbY5vOAbqvF3z4YcRN
vwUoxQVPWkCuU9RG6ldFXzkXeyUczRx6zGcERGnhkNDZXtzb2sWjm0/kSikvHy/5O1SyFrU+VnOe
QTOZ5pCyNnd1QY3wxf+EG2lcany4X/zNmpoU/wFAXlmRgz9XNhkoF3SeSFp6Nsiiy14oMEVu00PV
TyPpwDozjCJom6EncuNjJMUbWtqi0OIhFGGHqxoz9XJG77QCuSIt3wSQfkG1/m3lcw5paUM789rK
cV8/QkORnD5z1ReyaWieI1MJcwY4XRjDI7e2uWZQGdHIk5BG97KKtw7qo/imAWbV8Hd51tRcHY/u
Xy+gcwUUcUG9jUJi0Uhc3yFVc/Iyf5GhmwO9SEueXroL7PbknNTcAiS1cznfm+zuy3OR3pvG9n4Y
6KHlvGSSoc84qysi0xw0XEmZ1RizEAwe0HFZYoRsFqCibPOPdxJlKzy1OzGU8tLK4az631D625ai
MoGQ8V9AfaSocJ1fbX8AHymIA/6aBbZ76dXH6kHtpOSgReCYRTZRph04Xsqzl/69H13bZ/IAfPRS
pWSZsraUQbOX7y99X7onb+D86QrvLZOdnI9uPpJGr82Pv/H2WJlT3IoLEniiPYDHWvQ0U27EMLMP
vv2b0bw1Z/GyjlFwG4ZhwltXeHPTGs3otG/IUyAZ6SAOTPSgIsrChaZWnovyAmNkm8VD80RSdfqL
wlWaMQfa7lFxPzKU3j2ZwNjIvp7S9QVk1qYe+5d6JUNsRqNh0We4Kr9woEMoaSySNqbDkUunv8k6
6iAjrFaHOSwQklO2pPeI7s8uXccOytLdaCCVnsok1haB+7F/Hr8SnTcCJlT8B7seyigeIRbFMflU
zpX+Zsu4PqpPg7u/tv1pwWX81r0wlm+YbwO79ffU25DBQO4A8BTRHna+vKyUSQivKGBzVIYlCGH5
5NbfNqMYuMwYMy+dMzxssXNMNSSkF3fsiAljFnhBLW/KC4rhuY7zBQFqIKxDPP7ZbhAZxvYJSyn0
cKSM48Qg3QS4tJQginz5m4zNmxy9GzzGOr6obgVJzCMh0GWgItLA5GbqAxLQv9taKLIuF8yV8USw
MSMaLkimiyr6aJPkzzArhZO2Uq5DxiWRaS1C+xwtGf3EeNYAGZniDJftLm90vd3lBmOcnJo4NXbG
SancC5CAU124rLp9IFXUUaoyXdG2dUk9w46fgvQoXesX2IlnEqcYymFm9XLCWnSwDxjqfY+wIj4M
LQ1/uvKJY4fuhaagGfzePmWYcTC0mOBs5NV8L9CqwHm+0AIw8EiHccWvKAqIz5ujYc+Owpj/VrVx
vIXl9e2dWmEXoiX4YUQxR9RnLLClroutLlIbRZeeRGJ9o8FuktpeIL+WoPYTw+WR18xImjyhX2zk
1CF00qOdBwmli3K1ChzxTczwTB+lypqKNi7WHMg37mCWLcOAy84qHzzjOwVYweYJeMdbeiU8iO9w
Fkx/wcydiblJUNR+C2440EjiOZ5D/UTsSZ3Kzrm6viSv3+QU299YsfOmWwM1AHHxSNhjX6aIe0zo
/ZUb+pXEO4vybpeFQBdFxdvP46NvmuHAHzWFboGx7Y9iuIg1HveWG2G/VOXc3geoO5uGkDmyth46
hgfTyBHlHKr1HfyFvFuvSmtuR2eMTwz5SWypN+OvTz8FgbgTcMkc1CFAawaqTYRGUFfrq8fKKDN9
tbDQAvgDHGcU+1lr2FYjQI5xX/qRyNrh6TzRggYoHA4PsvDuuW9r+x2h83Hqx70qTGSSgP9yEjAh
VOI3Ad95h3f5nUEh0sfSgzW/L5EEHbvRVYpxAOf6rw6pl8qQtAawfo8wKFRr0+f9Ajfw8Z9edBn+
jBAvIkaSA6zomMohpY5sT8JdTCzH3ffBk2wip1fCVY7FIGOPTizmrTfsOVm6knnAykTfKOElPnbp
5PtB5jx00lcEBbDTD4cTcHxyLstUENgfR5AAvpvMx6NTdRTy0UMvktwaTcYtRaJ5jRHYX1ej9but
IhqBXQ5x0MA5JId1N1wZ2FeOacV+hWNRzUYOBwEj/ca+olxq+op+7mDH8VdSmWBwF7t51vW55/wK
1eroxO8JgZfrY/Xirk9t33LTd0AbwHXulhHsLqWja3bOhkKB+1uDEovwfsyNbkIXWIEo0eO00Sog
F39kw+6cd15KCJkKccNGAKBmU4zt7TNQts9S0UAgvj1cXmGa0Mtsfk/nILRfeBj9sFxgkDx+A/eG
a2a83cZVwxvFNwrYQPxbrePyEeC+7EINZZnfPXscpF/ddzGxZZoAB2PW3Ej3VcmZB5rO13wYzg0+
amtG0lbX/6KED1bo0PhtJdeo6ZLw+mxeC/Ft0+SSeQMaRnzSKtTvcuyUFfAH7S0o0wRZUY56u4Ln
2WQjVUCbKC5BBmVtjmjePORjkLT+OayM1pqRFHByXT9bKU6oHMREjSQSDVjUVGdRxbYYQsiszb5k
u2afCU7ynal9hyIt78ffArk62FBw0/iVrX6ypoxBLWLm7Sjyx54qjzIev1+VeyHwR1gyoD9DecZD
gOLeH9bBU4DZSxUI19tNU/tN/YevfNK0Am9u5ZTN6HomdWpx8lW0O6WGL3djqlUKFFkw+rwmEOJc
xewO1CUYI1mQxs3ujcrdl/DEO0MXbyqBOv8JHnt58vVG/5xnyLPBx1OjcivA7SSf2EEuYJ+JmcMD
VeCH4Q9W4GAmeWQRBInYN/tcKUmwlN3qB8dnUYz5A4fTNjC6OcbsrhCdLea1zpwJPp2FmkTlMBSx
g1rGe8fKNoBBCFFaqcVuFJqcVKhg5swKAJecDzgqL7sHdn4v073aAw8Lu8jAqO06bd0qXZQL1zXg
pN9bZrEaFCufW/if1PRrJipxbwDRVFine2QUao1cq9FMTTG1RtZxyyft/sa+newj1u5aPV13lva7
bGaucvoTw560MEBEn9+Fx85dIAR10hG472o3pOCpo9x0lzZGRp70meQ54PRZ+cNpgR6kBfnp8SFO
3veGDtnm3rBe0hJczE2rUb///yueE0KiDlUPu7aEdJMdvqVUaTlVzvJ02kqocBhqvqAyOXjcrVs/
6wJzmXYGFbvU+Ygjnsg3ZhNjik+Uj0rcp1zrF/BjCKqxt4k0ulXL/XAA0v3kUtI0hTC5irkq5OhE
Ui9uzGSJvwNnR1A6l0U63EZb5uWx3eW76IPepe/6EEJo8C5zq/E1dzqW+XkHn7/L0RfKZnSymFUR
aGzCAbW+PloB4gzcjezW1wvSZy0zZoOHvi1CTMCTuJRQil5PS2fQZdojwXSdcJFPvuCLBlLCTHxp
o+CIuCbOK+r41gUCrrr7n+pydzdLxBQjFZTrr4uRSlp6wmAWoCgDWfAbqyKdzL6/9NWTAdRXldC5
8zsWGFPMsd9rSWMs8Iv6XNpgJ0Y+P0vaSmzZlt7r1LdErkbwfn+aL23YFJgWFnPzO9t0+BjMWq3E
5sS4jxyPWwodZ3ngZkmNaA/rTuQeqZbR3k/OgwzPiV3nSWfd44kBAQRhloNcbt/vYgwCcbD+x0pU
pMszqmVPEiEh+cqACY1MO+VoWt3KaY4IfYvnxlvtwwpfySGeJ+5ZrVFVqLDrjmjlBKx6bcc7fxSF
d5pFbmGKOT8TSnSTlySiQwkk1qzYme9ntFt9Yj1uCTdsUKrLkv0a0cKdGl5lUzk6GPbQTqyXgboG
Wj5cEaKGYibEwX82i8ePTG8BrIo6siToU1bQrFjY4RmHhdUDlIYfBc5De4iPtBsCqg8DthGWBxQf
ACCe64gBMDrr1qQQAWpm6WH/DQa4HycPpKNpSxlZqB0SsaMTjqZVMVxycdUa/beArMCdWJCPcXe6
ESkyW5Q/fDhe6vMOHieboA8AihOB8FyiMtWljgeZDs+WOeCMpCYz3i+NRPlneNGPLZy4C2+wxgFc
khnKT4arw7f33xh4X2Y/3710rKvPh3zUIv6xL8iHkjznOu3cNx1gXBPETYlG5ZEiZf3vBjyXgfd/
rFI7bUUuaAt4UkfazZuSDS0fU8OUNs6XF1X57zmfEFH4YDA5DN12SLbhA1WBlwMzxXU9DSobPlZg
ZxLPNRVKaBgFhCuy8+GauP4K6LdT0fM/iFTRYKNbM5bH+FjOwqFFBy14AkRbw84KeITeNqsoQ8Y7
lSFdYLID4J3nwXd2EJvD4z2jTS4rP+ULhSpPmyosile0GpufWGZKDZmhcUes/3iDXs485FkMAVh0
cRmoGjzcaBkEWs+g1hRnbHzlN1tTw/vjomSOJp+5tyLzBqlwRlouCVutIdAZ1up19g9uvOz8PL+q
jRM6xcpSIkoG1lpSkuoFo6mGuLMyVqWKC96gSd1fCrSB+EF61m+4OzGBLpfaHYeTRYqVDD5G/lrh
+cf1bnLA0ky8q30YF2VWjXV8h4SyTqzJOjRjRitYYLSWBPNmx8bw5sHYzp8xc3h4BS7ff3n2GfeZ
WXxB0hJskUDIeKZck777uy15t2SNPLTUCJ7MQDrITfsSXWRtxidqzZuDsd4hh91It2xySd3jsado
w/Fz0wJ92ydb5LII+gwJ2cHCJMDXjvt3j89iqpWqvrzlmCqTzEW82lcR7+UXp0gNaWW2ISBGlsX8
uCRUXse+lDVzH/JnUvwGhXbuyfqhE80Fc1wRwRRx6Rh3bfrf+eUpQPi3fltkoq8Z3iGxhAzaontD
02PnilfuJLSa/6N/crlWdmMw/f2NC5V576KCklihkhwJr74WbNeFYqnGHELYcs/o+h/mTpplIUb+
46Bs4bYumc14NnWgeCL+vU+lbqIXGpRHAjt4fUj5Qn4f84I/qXtm+SrbWP0FHUEkowrcJ0jTudh7
PNshtEayRSRI2pPYCq5euhc4G9gc4hFZ/f1XBOoT2xYL0gzJiXgM3NT86oZADHOMXCbS+oY6fBE8
KRz5Pa3YD90oINnbBhes41K1NhVmf3thtmoytG0ORQE3krH2q0Y1D1YDo4VDgMhIySMvLWpFVF5L
yuLWz9BvawCr8b9xYJYbKznS3/g+vdzwVHj0Xj6VrpjTiUTfsJH7r48iIzYncRyzhvwYANKyj23k
fYZUwMLWCAP1j0luaXGVJwqG0riDuM4CTQgKn7YaoHsf8Vs6Sz/9Y17PoM/Af7M8F7m5Xn7+uA+N
F8HfrJ5UP8/dSgJ0ceqi5zFkIORjzdyB2RFqVeLLaVkf3ltCWqmhC58HoivesDVMhZ1GEoyBaZF4
/40sOfFJkUBmAVGdirP6NCvUXXAJQzT3o81svX53qnWKQb5YKQWH9u0NxgxsUZvj1h4tAljub3M2
s2W4J2rgkhLa21vC5Z2SfvCw0zJskl2Nzk4LhkFLkhQv+t0/F2FZQGyUtOwMJ0Oefpof167O3cmF
Yp760dw0afs57eaN24JYwEtEDzH/dEWOS3u9idwfUuLfbqXjBgp/4B0QOTHcv5dKNz7o1fnsUf1o
Ao0K7Br2WTvi5gq2faTyyPhprsKLhMpKXv/qsVxjawBYAoDsF9WzKlmJXB9RModryQm5jNq0MDxI
92wE/w6XJQHUQvuk7X5wdhDAqujKa3CleCifwki8nXeA/MujzhSrb4vLfkPazF0bCPOe3Z+MENZ+
hDFr9x7Fi5hEe84tanGGaPw5RAWnog9MB1OFJf5+/qg0I3S0tsMAEy8FzcURijr/kHaDH4N1/gI3
PdaHNeucfTFiKW2GC0QiSwh/NRdV2Vi5l8LLynpPEW3xQR0po1xSoO9TDDE6f8fLXd5C8/DXmu9u
4jk46r7YtdfQZJY0nWlucBdmVOSACHEp/IDZW/kNaQmzSeG6GGny7iSZzed+E4kJm8aJMeBeS/Qb
pr5ogVAQ8hQyYhfOih6RcCI3dOpBnc0PeozRwWR7Gd6GX0kG5Ke67JTyEcmdqg99U41TXLEUF50r
g0Xc/IFCuXIR8B/DvrdVjjv56pRbJrCNZ0YKSKBCZFpX59Q/bRT1xZxvI2UBoylkPx7FKP/Ht4EE
lVgLwk+ud7ccCZY1jrlpx3YpzMekIzY7GT6c7kb3vRb3q+jby/MZVZ8oW7b16TMk7vhIpBwt2zNN
ag7E0XSrsJl/+vde+FGxO9kLVWBvTEsUNEdhScECaA0UzjqQlX0yZAWlrkfs2+7qumXwXbwzZGgZ
g72ee6E+NK2w2cx6kFW1FdRvw4KBAzOSOK750gSz4LJ4XbXgZc+lk24RqbEJlur+k+aA8xnZ6LSa
b30rYGc5FAc+WPGeGIeZmrUQHXegQ2V0BWQmVjy1G6OvBuUJteb1BQl+hTsrbX/jF/iHB7Fkn/YL
5E+UqlhueAVnFIQb6Q3JeJXwDINYnUAWt180L3K+3clSR2VkGc8kXTsGD+39DWxsKCPHh4LK5ziV
61WWr6aQygGSvAEsygfl4d+Q7g+9Bckms/GJfueDTT7i7upmMJcXInx9qTG7rNf9xdkyk823s29g
jGXetaLWNP+e4uE4RCsG4DkN3Mts4MjVeEQSxUBVhAtyM0rRhW5R3j+qxyuryCa4dy8jHa7mWUhd
IwfS+TzbHDrvh7UlmVi5Erq6Zy7hlycu2rySLo9NovA3ud+U9/xIRfJn3LWCWw/FZebQOjJ6XWdt
xsYySE4jtlMQRiPPS4WOWNbV7PpBwW7WBUiw82jSJySRn0cC8TgAeRcdX/UjaqHKdKq+WZC4XAYM
2Hl7JwYDJDMhuJRayEyEGMoBaT5aG2AlCVAfy7Dzo+BaQXOuMEnz3sGC1ZbT5UowhuYbxXpEb62I
kneRlG0S9Jsefq7LC367/8wlOsK0kwTbHuMMY3Uz7t+k06+CPTv2aCzZYZ9oKbOFqZ9FoTylZCPK
v0QWSQY4dzqomHnnS+zUiXTvPvzYl5Lb8dP+B/HPocjeKJ48F7Hnx6EjvYBRv0WbSf5DS9E/rleZ
z7Ra326dwbH1wNM2Thatz0XwKmJIslJMYwGTzButEyczd13xPi+VDRDbJ9b6Ov4UjofT3wxUWki8
Wqn5Tp+TWYpVmSf9oIK8dfVCDAPpRYzx8LHUzPGx4RZT8vV8yKi5rze7qF+I/YA4m3SMTp0irBYg
b071kdVyDX+dFmkmkth07jG2yITGLNGV7CTHyeheSUgrz6KxQ24eRjwVc3yKmVzVy6BK61cATuw/
zRmGz2OXsKU5h2qfZrMf7jt0JilUhS19cqK4U18RHNsONjJuoERj8c5Jv1SlcFN9zD/mOp4AqykP
gmceLrgRuCOAPkANay3Ym3mCNBocxu0tIjAloK+qDOxRnyDmtCUnodCuMN1cFM0FJCiykHrLRFT9
kWUvQ5xCExvvWJC/U7Fs+Lzbr9JAtrr5oMqDSYThClR3lK0y/O4ASeX1GjIxiiOeg8ivYKOONhDP
HVO3oDCMEpyT0K2UqKBxSMBpBCSthjiUh3mFwM8FyVSCJUkOVU7YDdrPaaRKRM4RgoQ7AoxuRlYX
8QuY4Sn/rfanr5f1NtRtZCApBkTz7oPmQM/UI4LIBIhF8ORgyLBXHpgddnWtD23NfM0kelFBotgs
ilngkuTRF1E8Qp++q3uvmTTzYXuBYFp2Dv2Svy+QvFQAyLjSoNEyuBzaYNi5hoZZC2NQiVxHyM8z
A6ER2cMBCIsBunbWOudFBFaPHVIjNGWItjUENbzJgcDJrWoSYRNg6V53me6h2oW2pp1Qs/DTaYqt
Kq/79N4NrdA4UY2NCM44KwnfVNsQ+px3wzPEU2Zih+E09Ug0eFR1/RnmYe/4Pfbsf6bKxXI38BZ4
6rFyytPbwEHY9GkbBlaHhJh4bJiO33rFVh7vY0m8KQuypB7GVlAFt6wSsBdihQZ1bsoFYlbfQADy
c1fAs3BOhYeRrw4yuBu/s9ww9KtfRpGigIY8LpLnAD3BK7QUKwi9eTSW/9123erAr+Pa1u2PlldY
FPid1AJ5uWabQGyzqiLfM2QELs/O5fgYre6JofTexWf7+MB3lIw/KGF28q86drKpoB/Ees7O/fG1
oNZ3QCOUTRp/K/qWZr5oCD3+Gdgt6YIMGhxxT37Gv68pa6YATmxp6ZngrZusrYl+5V67224bvk4d
Il9h91Dzj1r6ueSmTANik9ajeJNW9a75Ck9hcWiEk7l5V6dYSP9YpyqqVObU3IznpY9sVfx9nDIC
jrmQl7iqHgSVZNIDcNkXogAXkPrHoKeuFi/eK6KnLOCCyEG8A7ZulNcK3KAZOeD5IUYcHIiOAsus
3L8GxulyVAbmjxlsF6qpXpfuGIFqKux4TzUtw/ZiPsOyXQcF9dEw0k7U3sPpRRwlpGP5wQTFzn1z
IfYnYJbHpcqh21d0Q2tmvcPQ2v4JnQNuMxrnEWcG/qabQz9u9+AI0dJxTnQFn2HWKnUoYBFhG/bv
YV4qGjtfwNpf7M3Ov8WIju6HI0913LNLyuzrlD+iQyuZg5xB5di6QVMHjBvBF0D1xwkgK+4wd8/f
nC09mW7LAd7wpQ1ZCca0Kim2Eg8eQpckct0XsXYT+7RwSxVbcwaToe2Ygckg1aSxXg7LtONlTah0
bl/xINdAxc4ufpUHksFj5KZFVKdCb6HbB04Rs7sDuQMHRyzF4S3zJhNCZ+/372+IKzmGXJGGRgOQ
VaUX0TIg0cX60Djf4hDRecyR89Rnd7WmESBlLKp3gx1zH28SVnlT1hjDwLsag7gz2s//qdWolUiO
JWU9oO1waA9V7aZG3gZlardmvaBg/ThW15kmHDk5jOIkPSucgKN0WyYiV6hAY2AEULQzEGLbOC+h
BKpczhlroVlXzd5CEPXoq7f/ZiZXoWlc+BmEki+HibNCbCXVDo5HkjaXoGJ/DjUqMIBkeZtSJfzF
LREAoX9l6c3wpbo5RV7nkk2up7yIdda4HV0L35Rl73VcXyqBBmXCew0uD6IqIbT5ZbppwEymExnz
/6e3WGMAfWSu+WELGC7PnackUwOuFkGXyxv6+va6fKOaMtJmyEt5Kr5mmSVgRiPKfcG9FikgHF7X
eecdLMwTG7pSOrTvnBDHbeNDxfLAgvYI3F3GK1FwvvpweqU4AbKRTWicrNt2QfISso5PAFbIRKzw
bEz29fr4xthLZK78oDgCVsRXFnyBKcXSefoE5dhbJL50zua0lggSlglgNEj/8ek3ceTK5e560/1H
zpphUew0EyJtj2IJXpAJLLubdmPLpc2D3DQKYeRgzK7IwgPJe3u8MWH265yLwKmKbkLmu2UQHD4t
6lOZbyqHM5K0OeytIWJQnAS1AzhecVj8hA3tWkgQoA062wSTWkxlKffm4tWbBXDE9sviJLTy4Wgy
fA6vtXMqzRtAGqmPOzz5EjXTmb3a3Dk5X/5JyZRhoFLMGw3LEOh8r7QrB6swIyRlj7U5tXX59IFR
0yPww5gksC1/MvmeZ87iRpMgu4Qt80GA5NOBPEdn2AKLThXgYcDmKzEihEUp/zZCPV6Tz90ev2uY
legQqmZGhhDH07/O3aMdWLp24WfbeRkpodc8pgwOtLN2MFKJcP7RXgIBdl+Y34X10Upz+x9eWYzn
/sSGpCzFAovRN3NM8A6IQ6Xl6gx4fX8kkhwuoCLcmpd2eUEvhSt+oSwiCL5Deo0GYV9jVZWSY+u9
pINT1GliK1SiRVKBvPX9kg4nZQNtyVzuQmQBz1izdYvJe4R7EvXMXpe1b4+we1dBgX/O+84BBkmM
Vxz4qO/ufZw5vWmybfvlzjdaJdPhzME9mr6VGPs+vbpkO7bZj3Z7lmChIbbml7SPeASAm78nPVAV
y7ut5YIJUc8HIqpKMbLAB8Z8/QwFRZJXAKoIMdoPDxqEIREbVCH2PC1aBTCxqcKR7NHP9eMueCLT
csxwd7f6QuTWngY0w8AjUZmGusipWD5G89Tam2xwwDrtPjHOq60psqhv7zh6DM0orjWtVVcyU2Bb
uTfLVBOYSMSVNLWjUwHvDuidYHNlWHJwXbTdoRvVncX/stKrsYsAJk87HJhzPJ0zm8fyssWFoX7s
4GQeb0REeuO91Ezx88pVlCZgJ870OyTkh+L3KzxWbfFsynWNvW+xB/F6Pe2SbZOTD2prG3/kp0By
6jy7B6M3yfepEBp6zZbZlLfuECU/ZSu2P6U2JxDWIWFhDK9QXfgckjUc4S03rMwxSAyeD4WdyCpg
3wPfE8uiS07nCAEq1cLGI3r/fot8mmeiylUZW10ZDjgGu2eICmm+wdR3eIevt0KACqlAg/EzglJV
ZQfDT5iVR+JPKX1cA+Z/NQdfL+mu/bD+/D/8AN4yEsLmFyjpnO3H1z0QtuptQYHhlAo8vLil+Nl+
u9a0PaoOsmyFvhUTQBB5FRKnnWerAgRDnxusgimR0I0NNuvCWx4A0mEcby5Zn0TGASALYiW48KGS
OZfktM6sQEqlhR7wjYtit2Ppm3Piccsez6AYVmmCwWS0r3hDBG0RauWP6TXZc/DJfTRdx62TAKje
58MXgFjhhxuL5uUDD/O3uTG2/ETccMumF+bXDORiIhjkuFmYsAGiPQrS6LbwJELWYZkdtnnpWjtz
lNCipHkiSO2Sn4sHl5NqjBf9Fkm4++g4RwkH7JvsGn5/izKJbrTM4MTMEkfrB+lGuts9wIx/DqLH
f9fkwn9bhT/XAQiQJ/i7efgugBLkK01CKKXcnZy1DCJoc2V8IqkwsiLj3d4PzSkROdJehRcQq9t2
mHsUtXDx/BRnQii9R+L2OGmmzovWUDQsX/w2+d+cjF4XZ1GIJCmzHcS2jT6p+rywm/thjuYlUVxM
2asgEgahv7AxfyfGvHXcHfrmzHxUUZIW65vJQMpI3pKnTPF8ds2ag2A476F9qxQC/Ngvl5HxlP4q
rsrGXYVzFK8TrqHsXyy37TJV8pqwlNGh8t/S5nGD+f0imZAf2ArpofPosqmz8gks8jEqE0BiwJ6l
zpFSGGQPafYDMIhhC+jdRoSGVfo9Yr07ZA4XhVjzRWiDHyOy5ADzm/nxcN6e2xoUe8UQNPYLSFlE
dcozliuWieWAmvnt2nvYvL7xIHF/89CsMfWyhXitOSV18IBGAq9PdkZKRvyTOy5UuYzIOaTOD6nd
UGyVsMkloj8A9Z9Sx/CAz15gs4Sk8TeldG4Y0wy3rO8jQvnyeMqAiwK7TQ/cWbZHBCfOQGS1wirN
6I53VI4zMI9U1MZ3y3gBRAPxNVUcTimHodKhGVf4hDv3IjgY8Y1DBFiGm81avVvd4xlQeNJa5u5K
y/i28SI7/X6MOUe6xIGw5UqmP+ecpGSsDOYLH7S7s0pCZVGQ8G+4SvyxNIcY2BTW7GPp/uUNAHv8
kNAvtPpJveiTi5aPMIWaTbnoqGjf/2ccT/nzXbZEBZRHkcJ478GK1qk+j2wHehmuBgJQ/2ZOGD8/
nIEI97XYzoiSUB0DptCSJ6Mqd3JRE4UlU83pyyeDkagvZ8/ccGkMcPHuRPFJQIF5SkvrCId/yYhz
K/HfNvFuDaQklLs6ISsUm6Rgq4qBlJe5osHGoBGDPpH7S5pKvVlVFFfzDm+swvHwDjwqXtH+b0ug
JiXy6Jjr8NblKUv3qtf3oARYe7rp2pAskBX/VCAn8kn033agIjjLDpY55g9M88GhRd//nl+VDwxt
l2JAwak3dFNU8Zdfo773f6gILglhOKqox6oEbQ0j9oVCvBNwO1gVwflNfSC8NeoMCAtghN7IVn5Q
ci5qVSEEvgtW+0YXzWzTX09rxsOF2ZK+11A4Csb+RYyddkFr9M+KiHERxMj1evwrfW/ugCsQt0/y
X2DXF7NliAEcVa+Qvq+l57VbKBoomvi6AKcE03kDCHDcF3RnC0OcPeUi6FPw4FNK15Y5xwNkZruy
BBABBJjigHstTz6AJLWqH0a+hH+IIlEBsiYagZZmXxqRLDmuMRsdGf/jDg1RqYfr5Jg7GxhvYu5O
bLIp8MBiba5y4kLsEc3dWPujdQ5FK/oH8im4x+K7aRKxb6qJZU89fePovjilhhkM5fAgCTgvF3P0
XpDyivXWct4um+HNCRgiXUsDXbP8MelLFKsN4hoTvUbD6JLZP4Gd6POBqUbRgq7NITQYE8otH79K
baH5TXrP9a2TQATf+hemU+qVxdeJJBfANh7Z8j3FZaf2nEESUtvpxOZotYUJEVxvfawD95j6onwz
L3/R0mlHG5nP7uIh5QfBcO9TFtAYKJcItP/F+gg0DRKQMUP7BOTqRF2yoYCpHkC9HdU8HozVOVga
DPAt+D3YXG9k4xV+1SCx1vu8rnXPeYeEXVptWNpE/kqyni7+3xffpOD7mK1EswzOX7bl+bwZv77F
LGifiSbKX/WhAL6cSK8p04ZwMxEjM534LAAkW6YzkYMXPTNJ3NvReM76FWB0kJXeTCLwVgVWpBX0
giNQDYGz1xg8b/oF2ebPkkp6nfi6y5VkWD//WY1rsKpYyfQSR7AJNP9Ny59iZa40H0gBlRgjvEHu
WmntW2kPx0+OQlt9mI+v9FUbp8jZH1+R2T/J2nqof+jK01xp5C+OldEEeOmgum8vYfdhzbvdZhz9
VyHC2HS0mBdToAV13sJ7DXGA/pF4DpuIcQAW/+6W9338UTFGO0Opij0AxWZwwW2ac+6cIlY63Zw9
xQClkuEHQbrR+dtbTf2DTWfQnGlCIO/fg4Mdlk9GNzjVOdDhoZVL2/Scc6F6gnuusu+1x0+qN8SA
JCw76E6em5kdIdZdVtYbasMdMy2j1NahHUo1eMowdhtVQybzbLL8zzqIMMU+gX/iqDjOWrxL4pgc
uWekMrh4UZ+5B/qfi9gax7Ax5WSA7yl6BhSz2GiiWxLkM3JYgmAxOF6CVh41YycIZ+K1y1rep/Xo
LuSW92ObVHt5IwTpUKqHfmRukXK5Z71eIpu7BSvpyIl8Er8dzpFTVH9PJD7fXtpbbsHn6blV0MAP
1QBcVEYPkJPAe5AEBR9NlKd5K46zBh+/+rX2atjRDC/vF08iefMQUcz0MgJf0VCRa13C33HlaO6F
H8DIjtpfNOkfw39wqNPJgUAGV0X5IcaHdX1oKngvirc7Vy8mrO/j5xU1ImPorV+e8VT+QUQ0A6PM
0EZ4EcNQSP6HOu61sCDZpEk0CULC2PO5M0nxO3gbX34hG2xGHGFhXssnJrOlGYZ7RIarcIk1bxAv
o1kMBk8VET5ofUtpBvDilSdOl7S6dFZm2Ad5CDk0COYwEYqW0Ax6OJ+vbQ19i3InZ5tapzOPvnsj
JRg3xzwRPDsuiaH8XyT/1chN5Tvh4AfTMlgQnXyWNxG5HeEphqPAXGbNoiaskYdpqeMQEHvVBwRk
QWoj4PF3TKvfK8X+VXd6oJLXeAIvzEi6+DcRqxDqMcoNkOzIxU8jSqrk2F8F3mMM1zwafcM7vdyO
JtT4gzCV+MOTPRdjQx2t7EVwNZGZzi5FXUxBZ4HkK/fkhSIpJZQl0cBlpONa8BuabYdL07MCmIeJ
JJ5XeftQ+e3sXsgTnKCDLhyLEtgYx/xqFO/uBJ7U1J/uIawUzubmEZTb0QJ15lTdBrgEzCqf2bvi
AGCk/zxwM7vZvsdzPaUAvS6WTCT+ardjP/h7cnCB2oBsHeyGAlOFUK4cn6rZxApxgYtOsNs/eXs0
PovI7flGN9C8cOD/EYQgZK1TTUV/1aElRCv33N/l3y40zNF/42f2L0+pJoyY0HgMWxZULBihqBj/
MXTziPr+ybNUCtRKP2JHVDafqDJmqZDItjS2hsdCPJwau5u7Bh/OIZ/qskVxluvIPwl6JnRbr/wA
g54E7qfxxSDO9WLjcngpyTzMMjODiyYhzgwR/whXT3A20P48LXCUAUJAnX+n+gpFxSf6sa9XQdlB
fg8yxe7DGXhaH3Rhl50z/Lo1btULYrwYXbt0wph7m410rNhOfv/SkkRIqL5JgVHrOcSDrGsp4lek
YA32giLbJwE+txuvwtoBbN134gmulTJDihzZprBsl3uKxNiA3uxyKPr/bklLXY0GQ7N9blKViZrl
BX2KHayX1iKpaBj/E65ADa1Kg9cD3+M6Ya786sfmD6/3hwUAxZu9lraZhGZIdbkzz96C5mWscdmd
EWwegU9QnPaZL58RTcJhKqsI2+2kxcW1ENfP9+NCGB3L41LJbWuSLX3qkKHMd98B6OU5SrmvkkAJ
y/vQZGcfjb2U5JMiCoIvx2S++61ZCwWVF1SpgbGZK/tNfgfBIFwXQUUIL6QEF/8YUwyPCP0mraw2
HIFWF4nE8Y3I591Gfw3Hjexfa6aXFkJV2j38NLieDTakBswqhpiomaSbEAvaWnmoMc/BIQ/eVBjd
hiTCBGbnYKYvlMzVV8S7xAozSDHO9YXd3L7T8p/8F47QyNuIhGIjpWbJ9F2Duy15BLkwIzbRMLLp
Glq+M0iNLgKzbKUlg32nOCv0aOet4WkyXF02eIR2JEgeTIgnDcq0+U5OBvX5hAP2HDf9g7XL3y3J
MRg8m73E/1wFuvHamViKqj5ix5UmZc75xcwV7RinVCraCdVu0XVkvP6tN1jBp5e+cOs9yEj+Oynd
yJySUYRrLnusVpGgbe5P6Lq5b9OREt5TwbxT3ykAt13f/7bTAssSGwIBByZO+Ub/ND6Rh+jr5/uK
4F6s+F4Si02SC/8+B5zutolOS2V7TfMGKDYKJzH+Vac/l/5RGrQC2K1+Ilun3sgtIWjeKIdZCk6x
Ylktrnx200LvhCGwsvs+rPSrwuaVKjVwvS5l9tE+JaOx6QVbaonVp4rYsR3H1V/st1ip0hAs84Qv
K4KIBwTyHiaQJ4G5YZXoTbsy75eMk+nyu/zwiK4vaGVNEbj0dhbRoFzjEoxJZxWfGKDKlSMLEZ/B
i7VIWUBT35iyZ18IJWGGnO0yHNgyH6LAxbSrqJr4BdTJXabeXnLDgh2KUQCbpK897rl7EHXXyU3L
gSsKmdoT+TLsZEoBChF9M/06Ks6YH71uYebmay2tUTLphzjDYRmqdb264icG2YMpR1Hxq8zbHg/Z
HLK3pBG5riYQc4Fi/rn05mdWP0M9LQu96/P7cStMzGEdZi95n9U+OGChlhA6obqzWEK8aB62cTWA
g4uolvuIwRpIHwA53EHB5KrW7juxtGqUdDX5mhMymaP1TVlNjhjY2UPApEG75JPvcXAwOPWoO9mp
7hnb58FRdS54GpfjGyRiBjlEDAWVDORJ6F5lCUCPL6A6A2B67TTibGiDRDxftGR8otgH8qM78BCg
kakJzh9t7qwgtD4Ru2i9UlfRLOQuBsNeC4zQZxgDkAJBB6CPm+4Ggtzz7mxcxapspXJIrKcaTMYw
5ww1XhSrBsqTZ2GoTd1O0KQYfCg6PIvURk82UiPgkqM4a5XA6SIvBbpKVVSDjuLK/vSqXvsF3uIK
g/EOph22UuYuR0l5Ns/9o3j+7ypBlf4LRqLXTnKZHTYhuls9Jh5kEKptetCxRvokTmdwaaX9Np9d
Ocff+WlLFaT29h1kiSwPZ6JTU895Oyt8S/LijfCdV/irGl0wLCPBlw8sgO2dDptaglJbOQ70tfbg
IjRFVLurSHPMUq++BGEWhgKcPJvTMjsEyb2XU8Au6E/1NDoR35r/z1Ner2vbkgtHepzTUrMo2LXK
bkpBV1B4mbeM7l6OYA+mBmCq2TvWZKaDzIRfGVUmQ9sksjutqbSH6qb2X6FY5rtTonDUPb/Vokcq
XtcWo+k172ggPx2Aypa+KSzvPsyHUVUcBRPoQYjBK1txn6pITjVT0ICywNXpNNkF224yV0VXMKjq
zj8mNgfxJqjuek0pwQz72EP/rNLCOmEKU0HDN7XUv46s/BcK0AEsLZ2st58BGCALqdbBtHbjbn1T
SQBL3jKewYqtBz5l19QDCdkpt+htX2bSnRJ2cTKiYZxzq2kzrYbweUpWFHG7mWKlIYQFK3p0wXpT
HWCC2XasmQFtIRHGG51LwPX2ppMCxzVIknktL4jm9T+q3UOn0CSbwXwULKp+B4A0596uyBGdZdoi
rWkBdam0JgW4LtWN8cXpSC8vz1S35yE5Jr9P/rs7dGLt9k6FL8sjMbFfN1issULv9b3ZtbAaKgKg
rC8VKasePyYKt9k0YKasaHm6/X0RMvAZ7Ov7lJ38k4Sqzm2heIam9RhFbtRXxMmgqMx7G1XAhY9a
riIA6MnCBn468Ev9uUTRBoty13nXocMs9olljoUBh7Zjl+/hI7h8BpmMq0pvjQd8bd+UWpktZ7q2
1y8+VYkcex2mxIqQyV/D3ButUOO6Sbh1lYzPnNOPKJZwujhWYrVucKGjhS3IfJD9deT1fDSdbZ15
s++NBTockOhcCICNxmQuc48AZ2ZBErgbQaDo9F5gPNxRFEGhtFLJtMcCuc9F9PzrqNVxogvsVMwz
/QOJXPqgvKEFrUXu+wFJ3p9QO7tqZs516q1ELgShhy+mo0lZ+K9UqnXuEihA4MwWb9/gpcJ5L11v
87EeDZORYDdZulf8hYDYLKS3K+Gdx1Kw49TixvialQLiU1bfYRtJUYDFi4ceUlpod0QVnvY8OK3U
9XJcvE05hidatGHb/7sRxGNPCReZplMtJUvmb9xOJ+OZgJQ80JDmRjjl4jAzrsG7nGr0QrA4kFXu
ih3nbFYu4y/+nNaMjn/8JQ0DJk22tnYt6PmFGsiiMvL45JX6ZEqRIJri3mI3hioRVC9wXgovWOo5
2Cs3sxgTSH2DVJYuiBEpi+bfm4HWp4e3AVBtwL4loLJljwabsYEqNWK1gihJOumwwxyUVTqy6aFD
d0xVsqMvMj8aMG57hMXmYmX/rHievFzUL58fO8xMvJibPYfHU3d+L2akzyWCTOsP1BF/i3bfeGMx
9twJThZirOB3g7P0IlbvR5Bqa9k1Scx2lY25VbaPV2pLt33y3SE2moBr7xarGabbUiKJDqUM3UL3
mYa6feb364Yf+Zm2irlVSjF0/60+3JR3rxggl+uP7jJBWzKkMcVoU2gwyKj7Bly3OH62dxeyoHBJ
eqfE9VAYgRl70PG3sByPfath7XMjYEAP7ZMekFSbME9ltoK4FPLZ0oq1rBe8ANHuPlApK5uR0LZy
2ixtPHvPPJenMVXJqXs4IpiZbD7DwKixThbJfhk9xFfzKlnu3QbPN2W2xhrobO2/B3rtB4LTp+v0
ITKIK8J33Sul+VsX5VpngufQ8171PtnxOs6szZqDyiJFxJP0Azh5BT+Jy3PxoF1QXYh1IvaaPSzq
EOGsy8gUXe/8NZhj6DE4U8/45jaCsueVZyAajYh6mDRUTfAZseT/9WxETmi9RccbJTrsK0nG3I3x
Atve81I89mPSBeJUUmuwf2xIK4qFMqM+zBJopQIZf/j2X87lthrvab0E4gYeZi8qgkcQfcNyklgh
7uDeiOaaioq0ARlTE9KxrpDx9XU/fzRW9t8mNHlsgQoY0oOQCCuVY1u8uo5FVQ+D1Fu+MpobxAVt
odes1mFUANiHd7P+0LYCzTTED7jWepOONffsVxEh4c6ZTouzhqHsQDI8j+OUPnCQvgSC00IKqe2t
PZLfkClgTtmDdtEtTluUIkD+b7RNa/lq04qgvO1qJR3HnhjDRlDoQSMYAwMlS0VXl9M7LAVDfTIH
u3S8gfhXwMOifaSF56nbvtz1nhlZHYMi9lMh1bxoCsTTc3UvLUmd+CyH3fQHM5MyWPdJwjtuSXFH
LadNWjD1Jor4k5SVkM5v+zx/RTvtEynOR3akI5URCsRjuwxg4HP5UDM5YOvKXXY9i2EWiTd0yG3c
4miYgSodPyT08BbAqOuKP/ghN6vI/nelX059vOwGfjsgUygvMV69xHgUHU8ddGqCtczEVMUmILjT
rYreF03HttPTIR9nOIE+6yzCKK/udASfdyYr4LLG0aQBNEBPy5p0T0olJ04mx1OSm9XGkybX/4Ct
9AyXkz/zZjyUuj7H3QiIY579WuRMLaZ3BFk8py7N1LnT1Wazl0gJ7YnkugZuJSUzVCsUP1lcxVJk
Rx5OJ8FKm3n9VNHdZzNeHYsr7IPnxOOBTjyjBSHk/FMjd2lQ8ffpvhfsHV6RS/ghuYq62NENoCKJ
IvJ2FcZU/LeIOmLDfBaSDhVSqdKx38oM2k9AhT3HEeYklTmKulpBbRcqBApB2sPnoeldzl398lT3
ekqWAeqBgtz1T4I5cuJRSsGeyJVgamKggNVd3KHEfL6cH8+/N5HrPhefgAaCM0AHMvN/LF5F3FgA
N/6bVwUL7wodu8+gAveQVuaBTRJPG2WREboR/waJs7QAm4AqwSL/r0qik58ecLuQlT06zdXY/K86
lYb4JfaNB4wJZ6GRut1huar7Y/71EcV+EuJ49237Q/LdgYpckc+qWjcVctRnYmMr5fc41+HzjeQ7
MSV8Haghdi4oEAocODrBBrKTT1v6u4ZDiJyPNkcm6BNFVv+HgQGfrtNll6IHo82BfxcJNw2lZWbe
BnVGgz8OmSmFv5kJGX65V4qpMQUnvU2otbD89jb+eH6BmcLnZLbuGD3OkPz9NLmb/mtiLuF5BWKe
aacfJ+MwDi2Z0ctz1NWbtSSgXWf79VGAEncBUgT+MtroBTlb0RHyGkRfnEyP4D8+un+NLw0LlzI8
VYNB4q7eg7OBAtuE/VPBRm+JVWH899t0SSM7b9Pub+YBn/Pc7eb0owtiZ4BQoONbAIVRRFef8RGs
Mk4TuZYCBFTjCQZhhYj+ONKUT1bQbUNEY5jvzYEQHvNlI0C5vQ9npHOxhTB+I+AzoFasAhoQeT3y
rtGLsVzvXz74Cw6CJE2YaKboCegIimcilHneV45TILbIYpy1ecrcSnIyt/La9Gz28UMG7NkXG1C/
enFWRZgIpS9Db6xx411q+sI0eTibpd5wWUVad4cehUu+q9hePvMGeLAJV/DukfalgvS76BKaOnFu
8WrUQWR9tP9cyI7A08kiMM0ndcvH3ObpmAn0d4E9BfiILw1GDPJdo66ib5WS9hR3lZ5bD1BWjlIA
Tx/VzJ7i11U5HF2xmVWnRXCr/q5sEd3b499FxRb/3KsZPbj0iYHiI6t3fYECOWW0Q+lgHJ75cfVR
1ROH5kp+WxUJ8eudxGATKYTGnZ5z8OPQWBePcQL7xg5EjLHtQhJ2yZGqTXvBum15VM/PdDYHgSqh
XcSBNO2YirmU7N4DVWASEQEzf2tIx1onEYqwDwXdxQGrMerQn6Oh+5EkpOwPdsQpmtlOVjDo0asx
OoQwmU7TtEIFo5CfHggCNXrrFyJruCgNRmWl1ZRsz6z3XHq69StJjKh2mdHbGKWi+hzKlv73qubx
P3PdGUh+GPgyBZPr//DNP824WvZ0o2xOWjgvgAS9TAwxcBGEjwAPqvU9MCd6pB6VVFwadF7uREUO
WCjIyci9xaXGLH4Ra55QyCbJabmEPO6oRadREVcywd7A7ZLIAiKRjEEsIpkQ6dIrnfnVrDGARG49
lRMkU8LvMqYNVE57wAwge57+Mva5XaOTL/EDMBrtIDmuXeTkkLC9+YjtysSCftACmf+RuusE/Ga4
gF90tkV05Ol/yXd7PBU0mAMmNJw0DOEPsuvTRuy+3icwK3cwWXsY729RBBnuZRtzvVGc5enKORMW
qYFKaB0MNwcHljijvlsVG/JVSmVcM/IC2ulItAR1QQHEN57aG7qZapcy4V78pcX63sFxLEE96XHx
DPEybI1nV8T3lb7UZ2rrOlT0obSzeUye4zdrbpmutazcZdOLmm14cQk7HLAHpNO59N14JDCK4kYJ
VQLfU3qqdS7bOH0Z0BKjeP9/UdEdhamFgTNN1142zJeUaMF6AUKt2Yd+PgghzYYLgZz1tDTGDXUY
yAsC6ss81a4r2Nh6XrGf288Bw/D/GUcKToqruKrWqG1O0tKvXRy/fHnqTQw/RyUuIzQRz0X4wh3f
KK5YioaStRnp6novhln+j/FacRJd+AQpSSwnLpke/AHL9ip0UexLbWHvkcYPP4EtNQkXBs4xkr/x
nR7xxOwt7pcNckbwmVsrLlSCCTwFRVu/2HvUoYnJDxC3eMO4TmezhXX49yJa0/R2iM943se8y8lZ
ljbNxIakV6GPQ1cbnE+In6ffjWhHZo0ZSxUE5Iyfsht/k/B8F91MQFRIYBzton60VTIQKOFbsdRU
50DKZSIySK4r5ZLE7SvP7oGVj3WeVTKnJ1RNjXfKW2jpvji1W2ue57gq9DfvE8eTyBXNUhVqriUH
Pupg6A77FYGvxWzKxcYjx/Oq58hg+dt6UhZveGIsA5JLnkWfS1Sh3UkM9WmYRA+n+QV2KKrebqzE
hYB7GJXw0GtwsgR69TxuNVO0JjJnDM/3xI+d71Waa+ahla2n+NK43rDnPn+ApO741u1EJ0wqFNKr
xGvisENLWp3Q8Nj0YK864xgO8/oXut+hXrb3Cvq3kxfswmMLzQrLPkr7zDkCAhBbDBPmGfflDH7I
Ge1uA2GGzPrt5YhqwRjDNyBNvbXk2xUhArGjhfY7EdUGKBs4YYCxB2rVs7eAMV5RfEGnzocHNUAi
pGphylBSeK7izk5NLeR+byUw/PEWqoBgGUIJeNpYOfZ+1TyQAi7SbQ8qXPmvyLNJAAy0829Sn1Sw
sCjiJQ+V58gW0pREatUydcGKKAEe/DIgZgYWIXrRb6uaOIsVg6UFg+s1l3vYwUkRtI/z8+AYTHhY
aIpS+K1Wg0ncj/wVsmfQGysGsSSHK1IHCtF2h3xs4mv95p5XUlsmg2uEyCEx1KOTy2FwJ5ufSKTF
cs7+G2W4QKQGaZnC1luezBnPQ8wT0lW7tqZU1k2gIUXFZHlSxrVukaX2GMr7LXFND4T+4X/MlqkH
itzwbODub1qzSE26rzAWfeJlyBqSR+qPMf1B7Cf/Buou8rx/7QdtOUfL9CDm5DLtuEnWfnpvPKFP
jbQlmBuHHX76mQIIjUpfUK8A633luj9MeIMwg4UJ7UnYOFZNj26NO/4BZ0/l+YVzDwmbm0cMAB9Q
i08zFh9/MtbiDFIE0vG1KNScDLtXk2i6q7CUobkOTq+lIBSnPNxYWMv9ewgEsPSHRrHL7/7jyIJ5
jrUTe15+rqZdi6xStCVlM8qIJ0bkqDQi5K0rd93NCusN84TgpVu2/IapxXHqSlat5b98dXfp8ExA
plwoRlMnpe13kzUwdo4qfv/wt9xhsBxfQFrgxMVIJ+YEdklBKj3QOBp+1+bgwB2FC8TF8ax8gBEA
/S51UnHpCvdakEp2txmhT4saINbDUZ1CIVN9AcmXbbPt1v714x0q5zBnWC9REBI7Pa8HnEvg2Eyo
KKr7E23uPA/J0ZgG9F2M0oIpr3o4WM3juFQacWJ4z06G6LxlPovzGmb4AUht1oBfQIIj9/fHoe9d
NAgyBydutqDT0R2byP/Aksfr7mN/e8kZ0kD2aw5PRxp25Alvsmz/snCIpmt9lcFjLjrrfN7c2+MH
5Dc0Wfm9A0s6/amkiGaiHzby43lsCFp+kJA8UaK/Knhz/D5Eihgc4lbdEWzmkuONf6hacY3CTh2O
ANnw+cX2C2L3Bg6jrKXZKGnFgeYU5fFZc2LEr1WeHjRbq5UyhrgBregJ7AqOwCL8QRm72dhw7Iow
jBca+eFHFt6ZmsFi/WzC+XoaAIxeEhGTOznOyrLlLLqdBmNVzDoZHlHmSq1c6aUStfVNtTPYLCcC
xKqSCx/rFT5c/YAz1v6WtfsQFV8f0467N3f/TEdBF0nEwsELT70zaANYavEf43kgtLt5w5tk+nAV
Rw6gncRHA3rd0IEqYRHAe6DFrJ4GNq8jJ8DTgYaMJ669w7gxT3YrbMrqZaqjCKhc9A8mtJnunMSC
igkwxrPEslAWvDARelZRU+Hypi0bB8TKtz83NF170ZGrz3hCbVdjoKWrWuy4fK7cDs8MBZp5fdTa
TnE9L8BQFPJEhTIT2HgWxDPkhsk7KiSCivt4Ib1evM9gshuNvb5k0O3BS5aA5B8TyDls+7JsXkyE
J1RWbLKPEJwog3CvWrQh4OcSTkqcCF27+KwOwI5d43q79mXIn/onMxv+cu8mLyg6scr8QOrLb1jZ
St6p7i+stEumKZjBze/uspKTOtjtoyK8PxT8cbJL3njL6g+FlgFTUE5IeA01GUtB90+8HcVE7LJ1
EjWFK9OJquF7SoMLa7kFIv2VnO1JDliTdpUTBR8JOBbCmFQU6drZPw8VDSnrwzZsfInh8hvjvKEz
5zgj48MJjAGvtSWvXSXCViAq84v7Imqpbb4U1psg02qC879FudyPp1XKFSyGbWuTKVl81QZ27bf4
RhPiBNqbRjIUWO0dMVo4VqG4T0Jrf8+ckBbFMQzqimggHbesat9Zne7n/en0+soWJRELGMqkMFK5
Q2ZPQHf4uIQdXO2UIiZN2nd7ToBLnIrpE8My9ihV6qoXxTqLR14mosOGfSct9fRu//hd7FgrAYZf
429zggInDDre7PdHmz88y5YbUmpUxuQdnESsCCa1wB2vTrs/Q/V35eSZqAEHLcOqrdX8WhoZP4yQ
H8mCILTcXPnNd5vkFdY/XV4psfJYC09VDwblT4lt037+T9zDF28IBRbck/oblYhf1OvdsC4W9O1X
SlywHtSWIREqxf3avv2Au43RUqYmv+JOQ3asvCFK7PdwSpdhBk16l4xmE043jVDj589rjnRsDb2H
MvAbJo9kTER99IL1AC2vwMlGx8IXnISk3KjH6EhFaYmuhK9gc7DOjQe+w2bwyYQAJOe31rqC8iPX
jsUDSFpvA5iDTiImrPfVckPsW6cUmMzAf1keHLw6pQd+NwtxLb5T1vVadcWJkZ0vASvcAH5dDFBz
4Plaqrrzw0xDujAJ4pT8EDmJJSu4kolCiC3VA6lGeCyFwhWQmaD0ZWFjOlC4rFQWG3+c69Cndm0i
bEbDlKHcSHfGklin7OAHIyQpmL5hEjOfp5ex0vPA+oeCdlxJJ0si9JqOEXyOWxzVhKxTGv8/qE6h
TbvEL06hCuCKA63k7VDLd39Y0aUXmixRNc6ZR3rWlJvc4XxjJJWsaJX0c/GD0MXIAKUYplEGAqH2
rxjUTH2xGIjrDJQvqXAy2rlL9KIuZC4XCLqrPX+OmlMppUyfQU81tDAs5GyrwBn24Xsz1K+5YkuF
C78RmNMrzY9GwvW4HAXC9hPN0Nv4ypRa8cc7PuvGdEuPvYi/rIAFpjDWbWo2g4ZA4Uo5U8wPwSuN
gX5AxXtLvPNYWlzY/z3t9vTQ/8O2A/Wovk/svLaKTDrNaQt5xK/s9XgvTVRWTlKV3gkQ4mX1k19q
yDotQp3flDr1FW6+yGe26OlIm7YUq/CTeq5bMDWuKWCGZm1EeIXAxsq1b8VeclxLrrqx4++dqrF4
177pUYwsHa6oyrCrAVn0NpnOpn3nbnMjjgJMtU9zeZtFRWDoWK7+GCP0Y4eV437Wf/bamFts57Y8
nUa99p2DwQWgmPkFhvOk22g7hswtoiZqVOGXOFLGZ6LUhuSKWHLt/pLs+9NAMC+lpM4a3JZ2yj74
v03EUJLQdfgsXwAoc/p8jJZtbjFgikfRJS/GZ0F31sNAkvQ5HcSU3NLo1kzOk0xbGLXdGzk773Gg
xg2LDwi/YiW3hHTp6aLfe51pMjO/CWVJlZ70/iM9hiKQwFnjxyR+BnqqTJTGtPlN//1/mDlY+qq+
Y2mPI8YcIRAt9mwYYkH65QkdOfuGN7aPski5irJPg0/y/QQZFonz0jkxQPKwQ3bil7JZtksqW/W8
npcP8seX7eZ1pkB5x+lBTMp6vkfjwVC0BYw2Hw6H+eKk+FH6sQAhZm2tWgOui0TrJJ7/NXpyjvxz
Po7YWJhPG0JzbxmQX1qtOjxso4clvUD8H2vsC2SAm8qeyDZUNgK80ZdqcGOKHUf0lJ7oLB32v4dr
MafkYbaPoLLW00xJ24p38usrsFiDN6pxnT9rCoUGnfC0JgyvnZpeDv3vbUkFLvZjQgdRZVNlgslF
Jz+wPbM8VJADHL4ZI21QDQ1IDFDKHloEhlADk+xBxAiE5iyYuWp2cgH9SpIWHrL0gJbtKtNf6Tau
TQmAUf5QcvFYcOXsTX+lEmurVam7QvdbR1Xen1sE/TyXCHXvPK2K7sl/16C0GKbYL7cY8ZTUByqa
WFM1FnVjbncSToUNN1mDGxCWuRQwoirkdUklaSYIskuA67SkuyocYCEoLFE3TUaVAlNNF9ih8s9c
zMY9iPNWRoQORcL5sFbbIo4ToiSYZ05PCpAmpLmSVbwxClphiNvrzWDMG5kt7+wrK8NQu8x6DdVj
TzMQHL7jCLwnScPbxt8d8Iw7AdDNb+VBZfqVbaok+KynMvyPtKYDidAg7r9gxf0axZTS6bTvHzHJ
n0BvJ5mnb3brTAGT2z8Z98YnQcrmCum/zOx5R/2DQfHPTpFfFBkhFmItCTkTCKbv8TXzZytvHTVX
XizVeHLJUvsPsT2q8tHrtWxpGb7sTEv4XAOi20GFVoAixJOfdSqQ0diUlhTatWx06Ov3bKujuS3O
rih6hZ1iStvcon6pZ84xbEihqSC7gXxAvFSQwg/9F21bVlxedDjTvapEWzcqc+a/ox/C1V/NFs2E
Eo7lffhMtWRqSEictpawbbbxQ9EabvvfetCPKb2qpZe7qihZw3mAwU6+S+hJiqi+WI9wCU/j1pKo
j/pXiNFbRhu+1VadPdymwlha0LDW1MnZN8he8x5LYoJfZqkTslzeExdDD1YAr8o0loSs0h8oJ7hH
vbonsD1k7VOqCKkeywxLcenVfn12dEp0WIrltFUFGgbTKeDAQS5cci9pMMns8ARw9fXzdFmMM68L
aXWek6V28IQKGcNm3p0y4BUF3rjNijeOp7KG405QjVdNUZVdVJI04SGUITGjOiEnZ+/Ei6C0TvUR
fA+KBz/7fY6AmlacRGVnzgZgmTc71/TxlXVRTcq390DEfFt7F14YQVMXXHenTrAV6xLa7OuxuidJ
zfijQsul5JS91k+a/GTLtOpJcaoJivssZ0fG/i4ww7k57SmZ2/FWbZfURPuH1aTBk6W8yUzDdkcx
lv9k7ZWTan8vuGp75g2UWsP5d8OVFoj1Cz0hGCUczJTWYOcFMsKORTmpKMdyOrg9dnNM+BpP580H
haPUf7Dm0sphNWDw6f1X6kbIBBqnNjZpNn1t2kotGjl2CwOgku3konYJlfwPbA1TtpTPuVAFwJXn
yPeeXCa+V25ZaU8vmzCHWVyFuevDvrhOJkwxrF5z/5m1FZ8avLxIYM+ZIxmpp3RA3xKIPI4zI1Kd
LLeWY7frzEIQQEhjFmmxRbvvDrjRrL7G6XQTkWk17P/UZ1A8a6rSdy9/dSNNtjugrk6vDvsvBdLr
ZYNHewKbLOZK3RtsCXLHmbMswW34VI99yvzfNeBRXfZMu/C59ft3tckz+2/thKZ4bKV7FwLw9nT/
b7T68Z6K1vY+KtEW9J1DxVD0MUX0/Rm/CuxpoB5zO8vSCJwSLeqjuIPTBVRvfHBZV9fz1AXeE9QU
+ytSgUupxHILp9kxl+Uz6pyIflecY/drLQEMWF6xo5ljpavr/QJxcKXrKBGu4p6t49zf8+wi/7ks
YuAvhKlJK9K3PO/AyP6kdybeyXUjn+u2lwU9usCkvjakT9H0ITaf6Xy5RPL2RjdqtaIp/pSrYSc4
cFFFZKz60aQiySlAYXdE5viHHiaN+K3hIakO7QiiqtxMSGqKT8BedPp3yCh4gldu4Lqo8mIhs5qo
riFnVFgO2LFX4K/I5AvNbVdiAc7uwnJmYAcxQ0tO1ggfRM7ZdpT7ngN9TJ7HeTL4OkLw9kLqR521
iPXO7FKJ4FfjxXb9gIyb4OtAed6H138twimqZ2FtkMH8bSfqlIvmx15xTH7WffvlEV/HBDNToAuS
m+D53e0keCKKvuKYzRc702rjJ0pNjiseoXixnt/XL7vlSrZj2ORlEgfLVsKMgHQwN7elMdICaYfB
0jgeCf/0TR6I+VV3vM0pbm5RLfgjYH0gShKs5Jnqgk7GCt3SV7yDi7X6vdn3WKoXIaIS/KeniVBK
Sr31bX3pOqIn6Nb9uKatCp50X1usmRMrTtUbXTujENLBW0OkALvvIOMASjz18ZDNasMmrEwLlvfj
avFvx3QkLmJnkuHhBGDvaxXMhIgSxNTCmUCESTrCHBLlzwC5c7/dQ70zNY7ftklhXFtboLR5/UnB
oYTUGXg6KojUapHedHCRgFBhN6oaLNxbqi4PX+6suA2+UCkxJRJ4Z8yXmfnyisS41RdR/lid7gf9
4IpA/nG2kiDudaBSmj6wznb7enNQwNjrlCXGrIbo/wt7BHkKs/ru9bHUQul9vYZ6nTMRRru8kd7n
Y8z0HBBCXUiaC+p94oHg/FdCsJSxEXZTOiuVNu+hwjtQX7891yBXjDRovp/QTR/nJD4UTk1/aVsi
Qs0PFkxTNhTR09F6sU5sRh+zjKJk47Fs0DrDKOxMA1tMTOf7YjIPKwvUmfgw+e0PSCdghP95zpFA
JHG365Q+dF6iky5WikrGPT68NZQ5SY00Dc2Omma+oBcxFS5LhUxWcj2z67vHoz6d38R4cvP7hHzb
kp+HxZ0gobw1p7w5jjpZI/qI602Ymn7e2WYC0MUkUTaQ8MnVu3zVv2Qenu/jwc5P5dzn8WVKQZOK
XOGBRZayrDOqIHDlCFFzM/SAbflt6laMptWG1sDr4J7+9OuOhLj67W4XNfl5bj6xFRkes2fsAXYw
iK2WJZVcDOFTRF02jWPtgAHEUVMwj1CRrjXfH5eUSeZ1Sh/LSM5qOzMTWanEuJMIodNYvbIugAed
UVFJa37KGouvicfwgmNh/FWg/3W2Z2QFFJmLPLvj3KVQpZdpO0xWSA+PTycnX2F/8owBJNZfL3br
MbWEcn1q1BARV7i209khMHHaAjqZbBbLA7viPHjtjZpm4V9BMqF0+jGk2/yMoyhRBlcYT5bPu8Mi
Nid2HP+Low7hzvM/xXQPy36GcIVBUv8A34e2quTCVlMQJ0ZcaZqqiSu/qyhqaZUsEaQLaumbDxYz
FKIm3L8m2xevGVvCeSdLMa17Fnr2LuRnUXcUTf4L+JNn8GnSKVWPYP8lp1p/XObodIV0rsfk5bp0
WPAq8gFWgBEQJEhRe4BGfuGqhtkGJAjRVMtPwJ5ckFJgwVdTEsSJc2XvvFLMzKqFF5U+Pso3GyOT
2XtxMB/J9YyWX38Z7zGfbPpgfM7DgHXJMDR8y2IM2/vIUiiH/dzlEoJs00owa6eC+eDNEV+OxBH5
9STIYKmeMFogGj8cCv6FtjPXfxInvZEmBTR63HmVP/k7+SDIModgkqpAuGlIthYTvo+VXj/vbD+a
8ep6nsBn5VZBrPuXDnuPWXGBbWA8wpk68XL178VlMr6mr0VQr8DJJtbxjM0yJEH651aIKl3ung0Q
a51p2uoswvJsDMvcvGEwgyHM6HGWUrUz40JIOCWHeKz3Ny9UD8x/GKthtPTNNn3+TNy/n21T72eq
q+RUpQ8nRcC7jDwwGv04qBE0cm+Kmg1wKwkEevzbqBUa64KE5kQf1OPiz6dh7sd48JKNRH39zIq/
0eXWmIQV7Izen5+RshQ/GOLAIU4qPr/9qIrL4FAvWyjUmDxr1Vx3dTUzTw9dPaez3egZ3IdUJKs7
CjDaU7Q+FTuE5EiujfOXhHUZzmuQw5NKRDHY+zdxheXc19IIiq1rCUSFkBT0O3a2OkgbP74K27kg
4icoKcNeRbI/8iMWrah83jNwjVPgJqJ5F3u8Kz/KBHrana1EP8ByZrg1i4bwdUzR1EWybIafR3BF
iwEnrN9/5cAw6t7un3ITRVvC5e/r8fPTXftiC2QvCIHvX2swpScsHika+CcfUcucCI7ozmxpm0k9
+vOU7BLRNitZ7IgXynjagCPm+53NLsGL+CN7vjjLMmwjPNPkvmvMj7Qf8C7q5c/mDd1oAizWqd6d
+Z8BKCJUdZa95MdGIbLu+6Yt8vkE0vY05Z1YtGxa9sVRbaShxo/2hWhcgNlkkFF+XJEoC+BBpsnv
ssW/ZHQVwlNXaZIgZMMQM8ARr4PBQzv3fL/81E37ZRYKBLt4SeGRbbVhBA0u1AGxfYfzWIhExfln
mZaQv2/diltMhj9OjvKZC6iA1LeIGa/Gm9/9xpuyF4JsM3KGXsycZG8sR6rs0cB1egNx72E1B0H6
Z6L8Mupx6LeHdMv0+c2qHzo/ceZGNd5mlAobn0GpYrGfKW0p85qnhmNiJMKWK7j5qJqgYlgkeFyz
Si4j5NjNrdYqp0bZmUj5clLgFfP+mQ+F7TwUXnH7XF69muZlZosfGDrdzfgK6imRNsqDekvY8bwY
UTeFkRI58fvwELkTVjQqZScTiv+hS1wIwGVoqbZLhdwS5XvtnQO+phAanuO1nXuoOciYicmWMbqk
6OvKWoiqsatq/bHPNP273X+metjOenc2S5H6bgM8W8IkVRc0kG9JfHUtFdf+PSry+1vwqwEOUop9
fbq07RuIV+w3ACDiKMlMfZ9FoQXZ3k36njsBplA5DFuP9ZEqdAoOvEUA8nH6P1k2rIwE+HqE+Af7
MHBorKuVYNx690tEbw9ucLeNhsIM9kVElKX0ELnCA91+De/SyWdKtnU7KJng1Rkr4SN1vZcM2HAP
jzA9X56JNZClT2QZbHOxzAdIqyo4NQ/edHEFDM4dz4DvHHD17yJajqaEkWwNNu00V51JdtxyYSaW
7L7DRj4YvoyXhrtL1oFTu1iW3rjMy3B1tvfQpvGT+pByz++Jjqw/o+kP7gWAQDXsxAqyGRP+r4Rc
UKZz9RpJP1xs/t14ReLIW4r0xB9FikWu0sqyV2TqZbjh4ERC/wr83ivAjDOG3ODXn1ZxWP9bYyag
wSG5TVsV/9s7P2iEH7RaNK1Lif4MvWEiT6azWBtdXoyvcN2yRkkXIhJ2UDtYAFm5DGslljcWVXWx
N35KuKUsCKL1IRMw7XFvxPd/ZTQW8xoWYv9MK5h+V6IeNwbLvir3KV6XYpfTXggBg27vDx2VX96q
nm07KQVlG29NDn/akjp74dQIGkVvitfwE1hG18TdYb9JRhyMt2UH7lrqwEi5JlHWfZMCYXDxPq9q
JywgAeZvsXRYvhuUsPlnBa8FVlmgDbWoZQMhskqFe9xpdB5EXyf7hIBqEnX52vwopr1o3YgmRFP+
ulasl/mmPsTeTIN5tI76DwLHDZWzKBwsZeYINoRFbSIjWmvAnB2gA6VQaz4JQ6yA7PhwaBrRz/rS
dvfCKbWuZubdpYaw/D+3H+euPRy6bcqMAwaA9x1KRDrDr7bTCxOXMRXhdJUmUiiqBEAT2MBdAu5Q
ltYyLT+EA/Pj+bRMalh56pHbH3mgcm8weKOokKczL41GukM9PKKAW/C9Yhr9g/8Tv8uaholeOBKE
X6tfuxMOzBBrjCoZ4kyjUu9e/GxwTyjA0VWe8fY1C56ILcTtdPtu8ACDwKUN8fYpjqI1TRS8q5hj
efJvrS5Z3wqv6R8ndkz20LsghTRTVyIc810Csvhgwh4weySpCnCGxnbwTXvYK97+f1OTj1Z0CAOg
nZvTR3Jc1A7XqwLnuL8M+sFMhjT00SbGe7O5TlSf2/g+k064IQWhq+OyaHAvW0mq8YQq+4RZDmXP
iiXfDQt0OKb6zS+UVXvbIPq2DutkTsMQGTXUaRHUY5AuhcBjmXvcr0lBbQDpW5njwG/6FobTPdzB
o2ne/Uf8AZURnQi4LHBNz04KLckL9nXHcQYyUcLt0NRlmjlcXKFC/S7qdEaltvGXPcprmzoaWHfj
aA9Fc0d1eE0wUURluLVLFUHCjeasxErjzxOSCBze5l0ogH3icAwMHhXAE6oQAbPb8A4zeo1HAyJ9
B2wCGfpQSmv1nZptke6eAFx3cFNqI8scsEmN4tmgInBrVxaZVZnW/+S76Ay4y5FzMnY/uPFezWOy
+ypJYEB9l7lfuk615IIyKER2uoc/8IXvIVquzcbqz9Rj5oN2iTcW7CG9nOclxm41zkknk4lZ/7MP
ZL5vcNkti54EJ8Jz2g+PzLXid1FyoG/fVIm9fn1vV2lC5/Fh8smcBcixaHdOpKCM9JTMyaWc4dOV
bOn3cZoraZ9+bsJQ6o5rFWyciwNrnLV5/4mwnCRO/AUItGYtHqRkpeaLFyMjSS/JIYFg9pmeuqsC
X+Voz7vzkz/uHxZ909cui5qf4mRwxeleaAUnUGhhP+fG7mQlm5VqMk0GNw0DGKtGhoL1bZWgUIbF
f6ul5IATv2AJUglplKEvY7weqF3yOrxXPUNC+ADxYh2XKq1Ak+iLR8u4VAtRCET6xh8wAzVKJyB/
+oaYih7nnDV6AgcECj+wJRLPmtb0oQ4lbN2N7iFfiSWZ/anQkDc93GhvCfZLox0goWZb18d6Pxa1
zutIcYRykRByB9/QU/HGzgluppimrctqplKSMYufCjDb68j7jMRtTj49e9YNqYZCKr6NYsAINH17
FZ63bR7t2zvs7XkYPJAbMR9VkygX6+zH5UkXSr+NCyO088+sD8Nzi89UdVam7Rq6NeOZTConPI87
TlQmej56EDoMA7voOWBac/CSiS8yiKvIy6dQHL8p8k1CdC8KkKalkF6qu0tyVSw4r5aLZq6rmWNH
npowWzt1j1YwsNEqV5zgM50ZM3IlaC1EgiKhPbJiwr0s5JAaPHo9p0JDmW6cXD7Ku34TBmhezN3T
bRHvdqDk85ii1+xCCYSKwvHJhfzsIT9fGdhJZI48EhgQkOTARUd1unuxp6aRlcfTl5YYA7SzIzYi
mphFRep1pqJtCgi9ih9HMRpKD+yU5V66kWBHK3THfdvwtq+9psEgRhyiLyPoQj5Q4ySy5wDKK30+
cShi3wDZD0I9671pEI+bm8yUPz8qR/Mca1zaFAOqd8FyNO0hfxiP84IVuZO+5ETvRa0Ghdh/gJKE
vAmvqAA3rkgdr6wcdFAUhx2l6IWD2mG8pcDAFCrpzweKmrch0/B/6WikG5K0mkSrctmdPKo3Fjki
M8jkA16fpUC4dUZObQbQD/dsoZC0QXoDOtfMBbuaOhAmI0x4KIngPrch8kWzwk7C7z9HskNPzn7K
ePAVD40SpwLPq3h3IPLLnMFRTYcz6jVhH/ZpaTd5xXPpmj6G5avjE5erxK2ozY/Jj4qAgRIgfZEz
5I9ERVW5kj/cclPEU8GXJmG8W6JCe9ltOvZGh3hkzHZgEff0Ncj4n90qBSuVv3siOPA+j9pfdwIq
O3JOCzSUXX7Wj1Yj6s0zm2ajjLq8J1S3CyrrXPwaWvtaaCRv8Y979U3rc4D3WzVU8Mm3cSLCsMj0
T43YPzHctJKTYkYXV6Wq/oFiwIzssZgO8JKFqfibpcsPBa26rTBze70r4VNz5v8ZOfskcm40ZLZv
QNGDm8Tafi3oR1CxcAcaxioDwUxYM9eKBdCKjBcD7vSyUGN9fuZIBu43GOCqaivdT2Np4TG9lS4U
p16otFYZcn1Ol4ZEkWjowYkw7KLpx8aYcAz57Ml2hrEdB6ncIj3Efp8abc4T5zwh70si8bcIxZjm
9fCtg6y0xmrarcdzz0RzRF1GgrKmKBu5Mnl2zLkCVeRdzXgtFZ1OsUFr92L0XvlFrPK4rnlmn4XB
L4XN3KvlZsbvvvC7WHwc4+ADfn/Ba8P0AQAHHabaUYz+Fwthd2TtOtbocrghwafBvQDfBVHpcBjz
p8/sD1IVT7NZp52xo4PZ2kw2msUqvTld6raOL3haTCpkHzhiShKh1J2dxzJh0iypHJzcYd6rZMvg
blTMwXtECu1tXouIjwrkRCHVEozJkx0UlpHQilUTq+MnseEHr45FlRzzSP/AM0IPdIEbm3qrVOZT
XZ2ZYfOhAQhLBbzCBnbhaWiK39V+Lj31P7jnrHsbXrzsj0hm8IDqRh86ZJ2BzaTQd+eVcsd03XsJ
zagQaaOzRF1JlsFer7zqjLu1fA/qYTuMSx8K1+LKhbsr96gnHVN+VAwrp9kngkMTUcmOyXIxVCJ8
5YsjsElSbpPlERRleo2p1gxWBCl9zAYgefhIwswHoX5FsCz8/rjUkzSrumgYFRnMXB1YIV7g0haP
rtyxEE1rV0Wh9T+uhLErvUcs7U57zW1bNIYQD55xhKwLRPAv7y6eok0AnhNFheddLG+xlw4f+ZOi
qIAWxQEvDGo1kJx21d+9WSC7Pndhleb6snReECybJh3aab8UonVdiXKKANIS9QvYuyrSwAsxbOal
/9EWuT3S7RPekF9Wvz1aEywl0ubYsbk+MTnbO527lKsAdi3N+wDn2QlsOOaYTYE6pA9wkiUV+fHT
vnDWyiuhN4CaMcngWjpEdHf2tBhUVk119kCXUVi6hN3arBDdi2Nxc+ffZZ4BwA2wmIXwROzP2yj3
ptoop6NRmTUeL/UvRP/qeLS/cZlUDPrWXEz8Ya2c8JfA+1NmZ06zhrwv0tIXH37AsC4awDHYWM/y
AX4Q3Wjsieg+clrL6Zn0H69GrSqf8noTPpAGEF8ZvEwG5JCCa3AG7NY0EoCNIXFmG0WNgYtH54ue
winzbR2g5qyM8SxdUAzYcNsVw1dNuEF3CEQUNKjOqhwLHzCsuUf9hptLpTSbRpK3XoWM4obBlHLB
9Kee7GSpNu8+zYGX+OX178zcx1bUgPLhJnaNuTHViyL0UAWKTIzFqICfEYYQu5ptyjcKTrHmSpA7
tZaOjrjTUvO8qfd4nzJGSItJ4cgYN5jmB0K4/eOy6oUoQvaF5Gu/10+18nhC0eXkPlLgdSgbMgEC
UMbCHUTa3nkVsUmfV1yI9IU99phs1LjPSAiQewe/CNHeX/5KjCJ/KlcN6Twqmn4sO9HnsBDR727m
AjacHd1QV9LHx4sbul5pG2RVL+GZ20YDb6PztMHVY95/5v2wpPbarB7pyk6xB2UAsTTQD8/iaRQg
XKuODgm3UbQ2W9NkbuZ5RhsMRLjPXYcvFuqCxHy+UIQDTJCFWNLs9+CZ9Sd/J06NZ7rzjr8Nie1D
UbQvO8UtUUhxu4ccKemhTuRxL9dmcsrj5NP101eWAnkBT6YfXV//SJqTX8D/8obOYMbQ6S4ERMHo
Gjxjuv0itI0B8nBw2Im+py0xEf7QUTmfAxsL0sEdgeEoQ8bE2UzSj6VZyjSxmovCRFDrRVmJm2fT
wMpVH8399vXjHjHaovClO8e8BHf5F5G48eXndD8EC91Ly+VNpgR5iKXV5BD+YIo/YrwCjKhwz8qZ
K1xwvM5tg49zY7KKYYo/xFWmL6kIFWnt9s8DsWp/lLT7dRGxLhbQYciq/zwrg9or2gsV1zMapj53
jw7GwcU5pH4/yVoC1QYlYfFT6lAa7kCY/khNHzMgCFlNSVbWuxdS02DNlHtC7eZtpuw5eCPTnNdH
QNVG8ds8pLZNzzVFqY7MUOMzI4DFCt536fA+MRg8lvwQMKncm9RKCNg66+uA/Hnwwl28mKIQfcji
gq0CdTqIMvP5tQck62EbtYuMm+TZJ3pIvTolgLg55ZXUXVn5cLKwi5bxVNsp+lgc1rNBeTEx94Bx
WUYAj3L/DDKEgIAwQH0GD/8h9tnuwsYwo1IeN4BEM+Y4kz8oXIthfs80S2M5NRFWo1k4TaMxXiVa
g3XQvmhUgKgC3bsnMzygrw3O7hM/rWJjAkqjX7WRrgU1KitIPcgRZHMhXeDaDnWjMCtiQnycKIwO
0KYOYircz24Ebj8U/6k5QF0i9ll4Borri0rfThAUopPzWhLBXg0lrRug3qFejFIQQOKRflwVaKXL
dKl1xs11orvebu2y/1vJ3OTvdXemnHFxNadfBH2NdRzw69Fl4KmSe8QWSN8BRU+S28eOObYW6GLK
Vx6v1lB+naA6/LbbQE7zXkNopssyZA7ZvaiwCnXfel9feYKVbL/QBAfBar7s6cQgBaT2rBVceEIZ
60hfuWvU1gqIKfnc1iKjQO1CdupjYkwiNrAldkPKa5dYdPJ31y36pU+LPEO2AkBPV3f8W3QsPjtK
Xur6UatngY5+J5pm3tTmh1wJ5SJFsl/WIEux8iFOYB73M6mye1nPOPK9mQ/mhklUa5lD1W0r2TZ5
96tfOi6gJEvxzWiJbIXSccDBUprnHDx+DaANAxWCr9k0H8CPFhnjDRTR0p/dYKFpIArpBKP3TMBA
LFbPmVXoyUgMO2YsOizUeHg5to4T3aTsyArm+YaSEQd3QBWUEQb5AsLxOzzpx7QJHI+eITlErv//
FkFa4af9xnRlEQM5oPH+iy7FIB9ESFD0QfENW+i8zEcf6hE5wVMCzYe4tIikFzSPEWTwCcIQnIx7
BA4gNBLsnyXm7Rk4gkGD8M9EiQCBULBJ5w9Fr81yZS9PLhXjHqOSQZxzg1TTlbhzHBMcrzGbVzBN
CKtYxWF3h+lliAlTx8lZdjp6zzOq6608p23cN9n9pmkpi7JTrjqYZ0hxHknndc7mbwZZ0M7qYAp3
2dBTDnf8OJ8s6d+qjDLD05ped7nbalIi+3xtBPXj0rG+SuLRXqk9oCQg+7FUvOtnxpnI79Hd3DA5
nC3umLzx/9VUZ5XvgBzBneg7VzK39JNRI/xP+ZjNzzd8I6b7lL2jOF7nnFbzto6iPjg5HDhTm1/7
w5cqsqMYLmQP60dOgnvolUt8ZNIMxh2BghOKjD2/DEkbxveU9EAGGv+d2sriESy4nmswQIUfeEWQ
eukn/NiHn+Gm+PXyx2KNYGEx3YmXgtPuG9g8S0z7nQjzoDBRAaAapY0J2NKOA+Z9tmaoyG3ajSKU
GT3KOO0xx4/rRsHsQ5hWaOuvLdmeV8ox7WHI7e9jAfmY5+FkDta+lzXwNe9MvqyMZ/qGbMNpZSNq
fnL779vMRA9yW1mtd9GgRBLCPOpupiTfsw0GYnVXiYx0iCIqw8iSK8TkpvvBVYf76Bt2aQDOTAnQ
AcHnR4id8TFXXaHocjFjb0/ZYINTxZB4fneZVlkFSjen95OadcM5G9BQz6R39D2HuQABKcHXBgsX
judNCGv8EEIPzYEueNYg7fIa8r7ZhD2Xejn0EPxCeRsq1Gle0pxcoebrSSnqeA8K4C/Lm9584vPr
Gwas8Cdzl9WDqukNWJtbH0OXhxy503lZiTYC0u0HqxTmv2IxLAOBCPGsPqQaRW+T6Asav+cfIj43
MUPPf3Si44d5Qihcl9EzbS/sBjIqDEiRmu4j4gQywpbGYAS6AGuVdA6UFJNP3eZ8y5WxR0mRp7A+
N+1rbDH8dzi5tsF1VG+Iiaduf3cTWf7xJk1E8UU6Rw6eVr/F5RMsSBTNy6VexypbtQZPcFQexfOs
JOVx3TOpGnQxxvBiT62txzj0WVFr9yKHCxk7BL6qaqFSV91MyKdGMozbYno9Gn3ORYH9rQ52MfIt
l7z1njZsSO9wA42WpPt5BinkRCQhXg3DCVao8KRnpJ5fAy979TNOK1ZMcRYbqU+yMcQnb79lUsut
QwiFcsDpsXzCDaBcFOcG9DRrY35BqIMx3Mxsds7WQyLVAkJpUohZ3k4UxQHXGKQhK0cz4oGi1c8h
MQMnAQSWV9JVYXmParaecOGfTTghLOjSRoZun+u1a8g71z/HicgQdGEi/0Kq55CmnPppHQwL1UIN
+qh1YW5mWUtpOLaaOGNvn8MzGk7exrIoxMR1U7GCB2eNvuzD0XOvogMeugj4iWRzeRnjnyplJwcW
OKDc75sCO+QUrhd4cyoKCHbEDFfFPdRoOPZxhhZS2Rp3ZO/hg8Az5an9U5ekYyo//qr+WPsxQ/7E
Rk6/6uJ3BcbMCcVqMl9Y1Wav3wYau543G2LA6GzOfLTTwspAFTOa+diT7K5fX8xdjrWCWkVFR1C4
9F/R3Lh92D1Bg76aY+gj5FNORlSSuqTMN9SlAZHX1W3SsJ0gtPs5uR0XjJ8QDkWtzjGrQUpfpZ1p
BbVVMhXgu6RuhuedkAerQWj8LHiZYI6K0E9EMEYDscFEXtG4IMNpYyiEYL69FFliY/k4CVhoJLRG
FMQjQfud9fUubmssoDhwmtQihsXTBmQQswvobMEOtEFSX34u2WNb9batXWK+CbZRrqxjx2LeBYeQ
0JEQZaT8ExHiljV7bsgW8NFFwP+OB5ogYxClNaNEFCgfyYwRNh3KL25HjtGABPtShVsUZFgEEQsR
x8fYkAsypdMbK997MdwqgbDEvWfgoeZYZIdwV1ssLVvt202H18A/uTn5JjVg7rudZwTejBaHmDf+
Lfs7MNF+/k3oPpNAcKPgAwEKeJu63KwMoljH/q2vtEOgwDEzd1zJGdArqJAu0ztNp+u9T4uaAeuo
7lJ2VMNWtdHDIq9+bpiYxQkvtbQ1jj9sqTtLLCOBNDdiKm0iuVayUJn/KDer85UbKA1CLVCWmYQB
3a36eOdMLUGnhP4INI9+Y7GdV14rxWI2cprr89C0tD0IU7kWJ1hDxQ1/y8SozuAEhhRwZPRxb7ef
du8p2wuZ5KkCHmLuzLdQyg0bYEat5W2S/xi7nJLu0jMx9DOf5/CCkMLYnP4Ryni4OJGnL4lp+SlI
iQ9AWZMhh7ZF1jKjyAvRfckguj1BHzNE8AxK/UmxoAtGTjGNn6W7YqA9eOdA9NzERgKVff5Lq2fp
0w4kdDbrG1kDqJFM9emZh+s6lM1Ph98wSTH0A3w7dYlWDoaVdzOuse3rHQ9LoZ/JtZrzss5PGzPI
ssHz++WQDAJmhilwwFungYh0Lbjv3JioryBPQwzWpDBKQRob7JFXW01rKE7hSzRKK7jvDzgPqhhT
Fx4eDz1S09KqAg7ZRV/URrfTNGurYW/l0njY4ZYXZh6KyNOuOK5q4peHdQYjmf6CFeNjXeqSEnsF
7FivrNTu0JcaQ2ZfJlFDcADCwLdhcOMtXv+KaLkHRp69l1SYOySq11Wm7pt0ZWOFGBDMpjrlOeuU
u/fCaLHDciyuqyRcSlN5nuEErmDlY1pYoGl0NDEMh+6yOq8bxDgwo/7Nhcxr4V7GXm9TB3JKT3sU
AvTLgXGTFXN6yWTrgsXtToDhde98+SRMApRUi33emdiCypv5+Mx1vMytzrv+sST2YrjWhQpfgjTn
Qvf9hiYrDb1aZ6MtRAuPXXsucG7O1+TUlI4fSlBaoaMrhcelDCpDW6o7YEk0xpmf5NlLuSkzRom4
XvLihQkiqH1ORBsreubChN4iwxNi9ZDpoJPC/2bM869IxJ3t+FPPLGRQzCqG7K0qooPEMj6HoN9i
bc19FAZmjyf/P3qyXl7br6b16NCCakdaP2jKhTOkFJUlDYTjOXx+wbmEizODsXRPYQTjDpBAep5I
ze4VfgdvUN01CF8BNj3lZ7cjzi+/0RyqdAZzwTzFDvaOza4M7Xq4xLBZalts8EtVPUT3ybwnCZid
RNYV+SKWr/HYbKXW6pMtA+fBiH2PwMRv00r5X0s3bwzVsmNY3SALROGGyd4rsHDvn9kNTyRt3e9j
3ODr81WzWK8+z0uJTVOfbAkCw6sjPr++oorhtu2A6QODwsy/Jh4GXbo8Mc44tNeeZeogM1X5Pw5n
cyUSHvHcvogGnNBT7ouHCIA5rGCMTnN6ps2DzMUHgLNzyKEuJRNFFS9ig1jQkjCa6b2gEM17jkis
5w9sQ4ViU3YAu0NjhJIH7iR2hDe43fsQlANTMGReSOUXESfYh+jWGm8GFPAcJjpbuoP6B1WOSH0U
pMmE2ajvuvkC3zaP3lw4RnsJHljj4kMYmx+sqlyO3ml/nd6FCc83r7k3JY6JdTiQpSQGvJDQAzNQ
ydUGiSEY8CPC3zv9WO742P5AdGff3RRWi2TMXDJvqVhSDTmgfgP0A5msJQelUn5QjHYh/dSH95Qn
LA3ZMzKw75izuaIgusGo4wcEatnPN6hFP2SELaq+EZQIgUs6o3AOYcCvA0v/b/aSrcljSnUrKlLQ
VHNyuGQ+AmWnbe6NXqiDWv05CUa5kZ/k31LObvK7/nGLJV4JEcy5Ad85xCmYiyZmfkuOSO3t0ZUk
+1F13iobLb827pQ/C3h4aIgqmhaGWIEF3MsuWBtEdmLt0Djyf9G6EKFcJx7RIgOEpXe/AbYMzY9o
vv+E/a2HfvLNRw7i4RzFNFfX7kkT3eqycA8TQWp7PAlEoXXbDfzLuGCUGYOYNTmayPiKQAvI2JPV
+8nMYxvO2arV74P1l+nVxiIIhYmfqFD2yYVXck71+4wTR2Cfh/+OA0KjPfpkbfnRLiR9sQWNFi7e
TEi/6v7unb/PH7nJ8rSjQR4h/+vEotLkAgmkY3YM83CdkMPIsNJa3BuiEL7jEngpzvA71U7yYKyY
h2wV0O6+BS36oXVVTQAmUzpl812ZbtKUjQrL1CcPA+V0kgctjUl5RStdmgta42ObzyLLLSsgEely
vTsIQacqQcm/SHZfDhxWtqGVoYFUaQ15NjDo9TTI07zVabbx1oevArr8QfqQIONLAJsv+JlVCfza
w9zaoV0VY6l5n4M7uXu0NuBcWOre/Soxf18TFVbUY6Vq7qLXcqB48kKgY2b/JkydcOXVIHnS9NP0
AyjI3JCyY3Nau9zk+yqUF604GS9puaiV21+iPhrpH4TBmjfQpsCIjmsezdIo6dldsiT//Ua2pXRV
68J9mUrnIrx7lZ7jL8iFHc2Gi6QvuQ0hEqrRWmWwf3WkNgyGVpTApd5IUIZZDxxasNdJQs3Ikso8
7XR/DKXTSy7m6DBzwVg87bYO4C7WKgniBKBEyfXGwTlewARoHga6w4loMOHHYwUd/d4/ww8Ktv+W
/E7LCh34e2nLstSaSVpvcw9rLvdxFOrSbGTfA7rEEk2b9db4fl6U0FVRDdoe4lMnIIuCeOOpZ/6E
5Vn6gQWvfbJTrLWmZaECsrzIZGsnTCSJAudImaa0ZHzGMFu3ncamZG221ohBynHdqwPvWQq5c0ow
qgM8uKiHNBlRshhAzZ+ZdWY3IGjk8iLYFcrDyXG64VWlWEtgOsjMe9m0c+ctEyr4jP01fNhhBQcS
k5bdrK59pdFwC39SElunDw1NPRgBwp/yWUVNUjTJxeclIhHYcru7oLmk4UMXh0ML67nYYFtZtTg+
XsYKVzpvwplqewycEeG3jClYwvRCbZRNkS5fNPty6+aOX+PCBuCpXrt5LDDF2bmqQPgep7v3gTFr
rNiDMSRC177Ynz0wFXg7V8Z2KhttAGurTsiGqnsivpQvqzDaK4Ce3rCwWP//hlPTAXMjejtdWxZp
Fi/T8WHUBkqjfLnwR/SnbdIH7DI71FWOnW1qFMjuKuIi3F7yKRvdjQJsLPJQmKZZ1TbRiqFO3mRs
9ge09SAkR12XwO9+PP1/CO9hWDlvR6dGhkilHGYLRjEyN7jH+3Yk6EO3oPFgPPlqJPL1Uv2LY9HC
zeLzM4FLWPVJb+1EEuIX1GoEVkPEM3fK1jnBPnc6fr2mS2Xpm2Ntxw4N5XlpLlrOVa8gOIyEEd+k
aLExlqhK1yfGyfavCxwCsjAvbdNjCOOGKQCimogFSzTpCLZY/qNtdXYyDMlM4hdr+o1S0r/Y9z1J
H6/CLiuUexOQHkfQyvgzePwIe5+xWmnoDT4t9Km0sor27PgqpugxBhpuqhumgnhA10g0bOM50Uly
h/6//YRVzyLvOPzzEvoo+BInNeZd5jjY/yjdo1bSxJvI3fkxqA+cbd6Yi+7ejUOkY1cEouaFI3p9
HjAlINpSgLz7nMSdNmxgryNzNRJqKzNCKcvU3TRorvnJq4GlQYWYwpbUrBR1f2hNPSbqvgkCPMy8
D89AJXdXV/b4BfB86GMJgJPu1aBN9VNKNZR830/9at6y3BXqg/To8e+9LWcykL8dE76EwMTvBHg4
kWLZibsyLHkNxE7U5qMVhunreiLRAODvzYue9v+/z/xxQKXhT7uztezatRo0FdcggNi13PNOtk/b
xqNLmXgJMvrtiFvbkPuuT2ivDeDxZkL5+VN3V7zhP4U8jonVI4D6RDJfkFE8NLVmBPZ3txQ9HAQ0
ghOTbFZdi4Jn7Se9/3tupds30QlNeaDS4Xeeq4wFP65GK989Yw0N1UskiqMu+rqqTYWq1MAq7Mqn
rDJr3eYJFG1aG7ct6h6CilEF1W2UoIQlvfGRM/iFxnaFTNk98i7fxkbheT6xU2+6gnBNzU2eVPnJ
nrfgGaG+dqOsXVf5i4zrmv8wY21n9hIpEcN0Dr/gLgDWjJMY2KiXNciPIiX/yhnrcKComVsrZQT+
lk2DjEl84wlQ0P+r8G2kJUZ6+JS3Ddyql4toZ8xNGaciDR1HgpRl6QNaSamHuQv4xNHlzRYZZ3yZ
z6F/HhStA3b1Q54wQh2qnNT77nmlrj2+LRJTHCx4BX0ZqKBlHerQaMNFBeY1TQREV8r7ImIrxocL
LRHfmnafGX4LjzITDk78z9Se1R1lA+PgJFUpZIBkobNqkaGj48Lbgju0agEf7socE7tK5AxWII94
T2gxGtMrdjrVWAzH7X/Bz6iuxqKHcDlEfDrPwvgyNHm4Uo/TmTy1JrDNLsk5qNWVUKO3dyEiJ8ZS
EeGoKSp8ia8Ra7swhsB7tJn/sDfl443rUWv4JFfG+hbU7K9Vzj+waZcjLskHe+2B+kY9Gyo0nUPh
mlWGbvul+K0YRrS8KLiZQxkrAgAOF0jPjn9ETZlrX2v/E2nJl5D2MBtPGei40c2/ZbGl9d7GuCQM
8CSr2mVgUwShpRBysFU1SSPLp2CsJRkpdp3sb+Yi8TByTjHhzA2y/hDgwOwDohNkc0KmuFXpOemx
1ilZRafHUmb38yCMkCxcNzE6Tq1BE0Z+9t+OJLlgAfnwh/CJQ1UpToMs37H7aYZAKf4h3K+CtBZ4
KXFLja84/vJxLhX2d6SaOCR3Me2ZzYk+XH1oPVzZU7zL0LyM7Y4QDTW2QBtam5LH4cegWIzZGgHx
w5KzIDLwbpCxOHph4DTKa42j4OyXqVwygPM8wggM+O37igxGui2Hy2Aov8WWbE56Twih+NSMcDVi
nJxnZqvntGzxpduzQkCHeTZGyCK0uQY16u273SQ56VX4idSY9r0L1T+r6Jbh4saq8w1mQAW66gzo
ieBdahC42KpCGwTwF1wYHuO/vaflJet3yuVqdRJuHf7g0587J8gA6lLCWypAoQ7j9+gy514CY23Z
Sz4B/2gwbNL0c52jVF9LcKptO6Q8vhly402p7haxHCfquWNA3YwvasTq/+z6IWWYSPS8e0+sX8bk
DYUFndbX3LgVl9VDTZ+6Cy4zJjCu4h0f2UMt5WmvXSDRxo1iI6NSlYw8epLrf4TUwCue+GU2ryTO
HHOmUu4HIhz/G6URxEuKSIy2Y0J+FkVGLBIxEvXnix1TqlnAl8LXH5es1mU8hDvVe7XyXwD4/tmO
VolbS+At+ppaikhpA7lYanzoU+bCfmT7VmlpfQOceSJ+EAcvLURWyF24mtTRQvPNkEJKUKIn0zsW
Yq1VGryE8vfH3Fo06VQWGy5r1oyU20uX+Bt6Y/FbgPxCFugPNkQKGQtlCgeRrpzIRy1Y2WM6uU2t
HX6322u5WezqNHsyC880nmzl5oxiK/2+r6ul6S+DnnmUSDJ+EN0hgORarr1Tk0W3gfAssd8uLFE/
dFs9MoUdZq23nFYZcuyE0JCYFfnPG5VmHBnQ2cVaGGY2865tpUwZKlgmgUahYjBUZwm9l+VdkJ3T
8m2yCdLBaVy0OEgEyoaAHtqowlIoZX9gzMC0msmkueGRbl5Ahi4TH3YfG7chCO6yzDH18r+sNjwb
ou2sqOFfv7d9ry1RNyFns6kKhNNJoK8UaiTyweKV928c6j2w0qtghSoRys/cGzXqK4BVHjz1GfuJ
Hzq39zH0kEERVIk1zdLCMB1s75fbAO2jIzx2e4XWRo9Lr9s+iOLUyHq0kjDHF69sdBuC7Mxch7aO
qXjLf2+pTzcqU1vcbZ9XKi0ujmKqEPvFC0pmadMFWt9yl1k+R8WbmTXCY00mXQy/4t+8lB5x0Loh
WqNIXIM806+OGxZxUZZJ61XjHIp6gb0+7AY+QzFk82NOZL5v2wURlNAzRnMNPE/VlywQ4+wkQQUd
QCcAGAd+H+PoyaTjRxVcb0lvYnIuexFRf7T12kqt5y7kFW3AQXrEA9p4H1uvXS9IXnSXMhs4aevf
fpROXKsPCBQMlAANiHtRFojFsCU48IZFvD9aBbU5xSiLTuVPrntMx7VOztLSO6ffl+7iTV9Cdv+H
MSyrokqoE89lMSEbVVXsERYDpF7kpct4KnkTuI6G0n1uKUkn7qrTQx2hHf6PWPVit88I6EIZmIr2
fHwXFJdhbRaLjj+1Wf/PnUcdMPCU8/sib3d6hzRF0rVWQ9tLIErb9Vyi6keVNzWePgj8GjJztKiD
HI51dSbq5sS1oTTT/6dnlDgoeSpO3ymQ6vEw9jbJaCXe3fZmBSqSrlcdaa2L1DbVfGPwPyUMc/d3
u+ksuSZhsIqla9Ume4EyyDiU9U+o1jlT0QYROZRXOEybId3X6jQUuzO31U4muOskZPBSqxQYD5hB
GylEtttPAtoWfbZq1SASB0gteOYAEiAYOIoDs22oGGOo7DjKVqg8gkPSz0EebpTgMdiW1jfYnCy0
LIAq4fCh4cdTZdfoGCk/alcHTo56aXlgF416ZPqWJmTvGEU4MxhehzqsORmD+cEf5YaIYzLe3hbX
RPT5VE+w/rlpCSf+sokdNppKkNVQng+1Jbe2rpygc3Z1xJp2HjY8wtTEwhKbpjlGVp9thD9LVvid
sOWyfeRRTaQAbZsKqxBxycKxaqZJL6OwRJpM2jZZT0BR7C++CjYlgK33X0Ut17gT04UAelZm/pGi
jV+oERM7t5OXyakWcQPziURRdIDu1WnRLzeK+ca6N7mLxoSUZxDZtvY0UOygcQO9CwYBKk9kYQ8o
blRt87hKU1c1PaNpwMr+G06KzvTk6IES9llbyVLqhspUeSXptUGC+UZ8kVewhMtr5QQAmN5pVI33
T/EJF5W3Qtq00udSObAS5Gc6xrxTBRmBiPDSxV18W6qsY3puQe4oelcCh1pk2HcfEJlV0ffdPglM
X9plf2z/HOeKavavMFdRZHwbjvKQWq+ekR4UDfa+gunuhYOrveTKyf2C8e/1xqzZBzszZXNI4S98
+kl46iVvomCkioBuKa99DlTvJYkDIllVgyBz0Y9T9QoVPjLobpt9joHv28S3jNp9vos1PKFk/GpV
lce6vV2koasysBY+sbCDRFN0PK7lrGa9KEShITFft+6+VM2oMc5q0n3pxHf6StbqtsDfZv5Lz4bc
bbCjXfmfAeNnT/ZN9D7QwE28FyJjApRnGzr72rUMKpYIZr79OctK7g1XDNubhHXM2AZdkc93QTDg
nCgyZUHEz9IpTI4yoRxVV1J4BRWWOgIRCgtIrR76J8ipTpne+jLiZzzUq3y5kZCggL1BTq9AICef
/td7E+V4RbywVP603fx9qkGlDd5pTK0JrxqnRlnLE3QcMZ8AcTob8K8jz4lq6X+C30HHyx+AcPNn
4NKu50dTxMRtQnQJbqfjIhTEXYDzrgjXYGv4flOsA4MPp4hCMkb6mwAo3fcCUlLC7NquJJegkqLL
eX23HOeh7+h/MHes10gJvr/H/C4eCsXiynBDV2sjHO6xnIbrjMay3LgB0FYcgSDkUgrSOb2qtKei
c90TiCCIcya/in11kVUD9lLy6j0aKQJoBzMFpVmbNBboJrf7QF25PhdzmMeVta21bXrOjPKa2VmL
VMmX8nrY470Zniri+Q/NM263aANrGC56/ZaoMj7xGJ0RcP2/OH7ZqiAZPdRrj5sEvA+dWE56aLWl
N7fVkuFAOWQRHFd8+kUCQETUscA+lkvS91pQ52uGfDf/fxqphL90lJxg5r8Sc29rLpEMXlgZWgGD
zTCpceriDg35MvpnJcVC5dwoYFsFVVwD9GZ6gvKM4yXA8ZIItvn3zvU2MdFW0PBhavEI7UQC4foN
JrcML74fJEvUrKTcQ/8cu48NQd2YuiaWLUKjysOn8KLu2Ol8xN3rIkHoBmbemYHpnstdM2xg/n6v
QoyWBN6JD+0Z7ki+OR+CiIgkvmtv4uFegx6WOn64PJI/T7jjeXzdL5Ex9DEl/PDqia1a2OnMPSLM
BJwzz+8zG50p/CLoSVm8LHCkeY1ZfPZ/ljnEpP5G+x6aIzNAUoNGX6q9fPuqhED1N+gMoWwUuc+h
tzJDE09tjjq6ZD733D3ak96EQVwIP/BqDZli+lfZuu9Su0OETrx94zJpUVRcoKE6xjhaZGYS/HSf
t7XHfHFZplewZgyK0vtEmrG/Bg82x6m67sEXr0mVoFFHu+CE+0CFCoLRF+wisvyyYDURa/WZGBFO
bDJHqjM4vc0ahX401Y+n2wHwOjWQYhRt6TdAMEQujLQxmEYQB/2SOOvqiu/9CIGa1VfL+PnPJDqz
lSreMj7BOPU9zyMqjl8YifyHK9ZOO4qtfvEVgpPisR/0kqFledmzBRd9SU0cODT3cuVJxTwQTAHf
AA1zkXs53A3FZ8E4o8qt9nvBdrgFwcOnwfipmoVDcRjFjE9yrxs9qNfjGf49hGIBb41k7agS8Ah/
Twfmqj2cEQinKKToXlWhmqEr7ASotX7llvU9n+tFkH3FLoMaqLd/IMeLv49qx4TiioPuAE93MOL6
V4c5BThDBn0kvgU40qfYeEsDqW3jRJFe0vLf+XPZtapVAlc+PFDNPr5byttDlaLqX8DC91uOQWax
nbmG7QrrV3CxELXD5Dx9Mq99Wa7Kid3t+wcdnb6HqAWbSwMiP53wIzeUuZyzYslzDq5LB6NqAeWo
TQlp9WQm0+gpeLhl48nYtNnxTzinmm9o9BeOkJQQ31VqbN/thmbIg9EkxAc0GbYdoLcsB5Pv5dzP
rwaHGzb1yxBOqBlaEMgPhNlw2Ta7tJk/4Wfmc71Z/8tYf1YAe/Gx93OvNLGBKpmZNtc0mONBUfsi
JIDgF25JAnSedYn8uKfFlJOCi+SsSO7gJY84/7EqWU7LoLztjF3AsmwHg2GbTsV+d+blOKfn/l2T
0tdfyHXMa6JZ9g0HzhRDJU14+kGOdDXQGXSf2RKcICwM17IBrH9rnB6AfskiirsiQUrd7kcRmVRS
4dkfREZ33QvrxpERjwT29J5ZL/JlcjhhRQL85G5btmUTQg8G1+P04mYAcHzcTLdHGhcpF4wpDcvs
6LF+FZAU6UNLa62ax2c60mb5edZgDtxcUTianMYkmEZpuMAl920zS8Nt5oo+OrCFfDpzEZWOIEwH
1xO77QMfhgZm8s5vfeY0Y9+SiKJXiiMpWchnL2uO1rg4fVWpXqhta6nZSYAxoVDtck7jTZ8cfIV0
NPH3Fdl5M7d4/K/D9xiTUBYJpzwSTf/7EvbrQz2KHbCWxVFKT8rjaoVdEh319YuNkbndwvO8U6av
ysmZJPDyLOx4fen0iUu1hyze8wJDEagz0zCqDr823KwDLihGeOKMphkc9dqaeqJkFB4XUErJfesb
r/T3zoOueCXBXs1oGUNLKOgIxEAcvuCHIprvq3lqPiECMJUbGIV3VjOg+y7RxhakVFJTenttxT5a
ssMHis98ZBXoNg9TthHw3JezTfiRkli4SY+PdKqw8q9OS4M90SZkRyGIIEre3RVWiRJlEvngjA5Q
sVS87HdVgsFWCEMYvGQcmtwxfAOydqJAnMnUd5POTd65Tfhk3Ws3lgcjUBn05OK9E24CaoqSatdV
OPR3fq1Jev4YdwGeR3iJ9PsaYwhghJHvJvVBXvoFuH4chBz0E27dqaTd0kIaqbnrNidHX4WGxubE
SIctzngiASeGnBRT+qrCRtqNjuoLU4wgHfHgLhPBmhKRM8sLOD2hm4txoFDcAkO/qskI3ZK/tULs
15yoMEDXWCaSnCrVzQu49ID/L5inmcpT4owhGWSXz47KNsBCeagOBD1PGfyc3m7iggMQCoaFT7aG
NhmpLZwNin1wAc3aiM6LA//zEX0P5wFsmAeuUPEBpzNClA6UypLzBQ+XjBTWblr3jiItO2+PYBhw
eOFVpMCE2OAsDyqnJle7WYidtJ+wgLKHwQ+Rj7QpkNyPaqmP1EzsOgJ6lyjAFeYwDgH94AZLqh/I
K1hWVCl8o7/4JdiMAAPlhL8lKZ47Yizk7EhnEtkQ7LtA1LTYcDVNmSNdNWu7XjwYtnyp+MNySQxJ
/hV0UihGJjVfG+g4sVyIbZfnOOnozoyqfkTRvc+0w5lrd9Fb2y85b84xm8RYh409TmrPiLVlVTnn
aBsFAW8SGpwdYwlGbvuCziPEtfIXuZXm9tIYWSGry09UhC+jMIGcLTGN+HeegMulXZCnBM8xHCOT
grRsN7zc/vQtq2HBuYhc+nZwjJgYpDm/FSwOrL8cPMzs9rIWE3Jn6b126AKLHJ1MNzi5coPZSMca
uwrWBwSHZeZtv278OtAhAyFVAYB791aTUj7evGIqyMwVc1WFlX+r6bHGr+HEAemTPA7LthmTvSpo
xGBATymNc0nQs7uXrUFOkz76eunsIf+ozgj3drkWeuqaBCRjqSmIHXUF1k5U41PkbnYYAMcRv9eH
Ue6TNIHgMEtRcDM4TCxIAjA7A7lMqO5v/nwooO0S02GRN5zVZYRfLC5al0OpRppWJrY3xL4oU+ot
liwfMnV3x7FUgUjX8X9jbZBKKwlwyPs5sGwDk3oTxFvU6GYZjH7JQ84J4RYQtl4Vg5N4RMCCoUdQ
hAKtnowWxvlPcec5aJ1+R0YULsTAKsK13z/+e5hP0iYS3wghQs6B3GiakwGJzFbyvhapC0WuQBH5
1yYlLXI8CNCO51tBh6UxOYq0rkyL182C7g51KcIHPhlZhSLt0KsLIAzgDFRjOMcggdukBvdfwHB9
eq7oaBuHHc874iC3XyKP2tT24vun8mKD2EJW18cROrbQwHlEEM2lfmmEgTCO/fkEZ0OwcO1yOpgJ
hZLLy07iGSjsfjCktpzY+Z2ldepR5osgC7NdJgsEqtjLwkQTChqG/IXV1iqgVfAJSJc8WpcU7xFt
D0AkiOAd7BFVHvU5yRddnIqxBmG6chD3OkU9ZRanSUPvLzQvU4sx9g1JswugV2VzezvOrCS/qDE+
+hjfB9NIc+xUM7J+9HKlkZ5URkB+5i1AG+tq0olzazc6ubOZiB6L0n/o3KU1WyLG+CAYYveYZi+9
lvTTve0OEck1E6TgVeY5KDxBvWALGXh1Oe/3GGxpoKCMRgjoE2LrKqldi//UbovxF2Xvyr6d0H29
6Ihae63mzhXL+tIAAzClKT1kULjQQFs43c02ELvFMsOXVks4bIYHlr3UcEHVRG184x+b4W2lnuPC
rHv4wgHfFz6ths4SaP47LdDdyrjBy2qmVjjjMMJrTXrax83wb01j2H8HPkM53r4BglbPjz2+z3WG
S9om5RsxWZtUUy6f1F3yZ3T9ouOJk4kXV9ulWo0Aj9jVni7smE8a/CYi6DtPqb389bxg3+ylkF1I
RfPg0ckQftLlRYQ7NUyiYidp7I74N3K6DO8DbMsPBJgj1EJMHV9yBC5blZTNYXX3suo0pDpaxaOl
jMO3wEJ326WoN7Dr5miMeXif/JathsV+LLimLYQR4jAebRdPx+ePUAE9ACjOoODLCBhodZBNDPlO
3N4suGS+o6kKdbq8Fr8xr3YdgE+XMiafWrClsXQ/nSoT/cYm1PHo284fwv89bAXLs/+WtYr3Fl9b
+kBNBi7cpWjjwXc/JUXhTLMl3jWYQbaRdzlQHOwkL0n1I6uIjekFz9BrLaoLzdjTHkvt1CWXZ2Ff
bK7s7k8n8V8CfeT/3R0gH/B8WtA8ridb001RVCaeXhO57z+i5UgsMXWaYqatUUTINAH0tow42I8k
TFbZq3N2iPcPuRg+iHJLuey/G9nybykDj7LQKC37e3fXk4qaESryNChMgQdasCiUmJSwuT9jAGTp
5iQXenloWeo5BinqK7WciczhIQIsTy9kBtLDl6B8c51cOYDVaFIN1UwPB96vPZR9Q8ZXyVU78U2i
NYaMDTkbPHwnPvYgf1GKbzvUvrGFE3Pnqb6YDQsPwOLwt6SQPP0DXmvIdXskB490QJN7yF/jVorX
q0+ZapJeIG1aAoTmJrtkRhCZ7h8tC/S1n49hLge8gTooYx/oDOmq93HnBSfEqLoQETO88Xfk3QWX
71L0xtKwVcCW3pDEl8UrmtHtVPwXE4syk58pgKqGcP0T/J+FzLTbyB7cGm118DgUPBzjQfyn30wx
oPUVKx1ArsVevioXc8tz/jewIlPCOeUGu0dcfiHFZfkmuaRZtQ8ksgzr21m1IPhNr6UKgntJ9a2w
dfTUzZUMQUibMk60y3Fea5IWj/ueEZk9LhSLJqdER7d1reJ1n8xgmffqmvfxFhCaJR4PGGnTTmvU
WRZnGK6ALPnsZPFLiP7ZuR0hXxLaZvQveDJt/7dEWZJDDw8jSzmBcglv2qaXlJZaEs8fzi5y00jl
eTzN305CYoDI7aYrE3M3JEHgJw5VMPavn27pFEqNGeVDVWs5tZMyogbC56cS4G4eioY8yGj/Uz1/
G3V8u8nR/UD92FLV9jpWRB/3M8FW8OLgZN5/nXvdSQ/9Dq4JViJHMYNai/HpXJr5mlSCgHpmCR5z
MprSJ078yQyW0dipEhiX9/2pzkCeDBH7kbDAlzUV9lcLTNXxFDdOHJTcrcprQ2H2+IzDjNKO5Tfa
IBrc3hGd82rJHBNOwzT9gdXzJldj0KEv8a89nUH2Tqaca6XtT8HOCH1VUrZWmsRQBe/UpiJzbom3
u9Az0JwMTUSgCS+r4JXMyok02yyjS8SbihEGU4DovsV5F2wMG0NcQoE/+xQZ9BVPVG9R/03WeuqW
1ixnj6bdxh9wY04R1HDqWFZT2mSZEs5yX9UHCT5UDZLcz3cEPReLkYF+S7UU7ar6fvhhBBeTBJ4W
uGnDikY5Xh8BeO9BlCNbsTB8xIl5/GhcxmfAzuf/JM1S3/KOq2qVUfwPFirpRMMD4ftiQZTLzEFm
n0UcPHkNkogavtWolqZg8Ixmwd5aFHoRPPR/Mf1b+ARXK77GvFK0R/C5iDw3x+iK/lzGa87LLzMK
Ytpi+h4Do2ar/GGUXeKaLXrBs7E8UOgJfL6+d1jGs7u6vydGLF0udZ/RJ982RkFnb0/4GAJnDOS8
i3l2haXNTnVRVCgpeDrhfBatEC1fVuZGw6vx8pN80BnvPLttDysXTg5dcGPNZbDtfWoAhgCItLwW
TMZHz3CniEwqq0rGHJRKhoXXN5ao0qMPA+wuHkDAiim7VD8eolYPpswj6oICNr8bpi0sZvzuw6PO
Qw2oFUBhWy9htRuJTpDXwIiP4xlYkpsUKGyKAsGhqrwkUzf1x+DHsHIb80FJE+9RQkidxapDaEZy
3AhanfaDaPVgp3f6uRjg5UOcr6UxnN7jV30O5BpNr5dWuGpvVN0HThNTlma+xik0w/epZvQlV0HI
vnNoOaSPzWU6N2teKZWqSP60brFgnZg7kX5X+ftc7L6X/K7Eu62Uznrp7Jm+MH3RgxzOWBfwOb8U
JAWj1iFskoijyDxerzFD4NI4H/iLV0IS8wpOJOZgZGhgxF+NuXrpEo2qBsYq/qbDz/c8nK0YLRj3
bFyYYwbUsD9jFIGQZoVoP0t5M7RhcNMkFhUnhcf+WAnTX69C4Av/6gCxPeuf82VxfpFCuF6ofxGL
fgb8LBPfRwxViU2LPKTRXYgayLiFp6JRSB/v+0SozS0DPBP5V19eOJvmHtfeV58xBSkhB1tfnBWm
7y8aPIhokoyGk7J+1iJXZlOZpEF4XM8oK9R8AZFvYLGwwjioroYDKNCHpDyVjnhyBesGdG5DHE49
NW4EH/ao+c19YTNjiB579RTroXxTisc4IsO2Y5dZ98J6XY8PQ+YzYp/4Hb9mQhFH9gS5bupxMPgI
8owCbmBS1FGIvKNt+LlKiHD41aSrHzOjCokMQdv3CSWYpu7f39Z2new2L7hxuyTNw8LFGu/F7Xok
ZmKkQMbWVGiQ9Lz8fyCKjfbo+9ZSnnJ0qHmUV9au1eDdeHDKKxlgdyjfxUPqkYuFzeZU3h2brsYv
pPEW2FYwDpbqhPV53y7I+XUVI6IyXP97yw6V6FHIPKMlbdA9iuFjKbyy4SCQU8XHbc96pMmFHjXF
L6TuUYBveNo7vXSW1Ix+1vBO6OUTD8MynBC7PHtP3dW9wL+iA8SE3Ja4q6+wwg/ZTTWdQ0VAnrRk
cZX8tU29ArohHi9rFB4tbqDOXbG/9j9qaXfSxCoo9tmaUJX00QffS5os8aaErjfuMO0r++ZNmuRA
5DXh6FILfAu98KAix31Rnlabz4zZTWoZkwnFswiyO8DmIrWmwrbJQayGmSXJFGCqFUwoKo6QBuwq
rzgp6usbDDcJIqGJuMY+uGVn7jruUHItXvonTSHLXSv7iRfmyvN2JggukeU/7f1T1v0CBNBTZRB8
Rb4O+jJPQLpbTRaeT1cPat60DecCLy2G2GrPXu2zS0MRJvbaL6yIqPdC9MqL8vaFV9RPP9I/Af9R
Gk5YdqkCHnQlkyWyGJM5YmcVnzcv03VZYxnJcMfngd96NWZb7ylDtVVp5X8CE27SeNeOxUmpbJl/
ihtz+gI7xeYYCsUJQRmu3/jXU3mMCCeHEprsP8IooKiHeXi+GnS30d0OwajA04HpVdxfP+MF4FHD
6lgSQxpK18KzZroYVg4Iq3Y461COXJlWVBs61swPN2ubIw39bgGFz2EmlcaTch2bX2nMgh70duKU
+zfT9k2wO/x2l0CWUY9vMcCgs1cRFCejHXPPiR1w977ItIstKt5C2ZSxYmy3NsOdgd1LJnNA8Wxc
emalhECcehS1WvUyclNb0uy+pr7GY12/vtRyCqTs1w5N9ZL+G6LrFY/OOx8JyKNA7rtT30BDg3ht
6tA8UT+ZUFroZQiYfqopcJoHpb4GA2IkJkjWCP2yZxOF2E4UbrZGhHrUTWgIkPRmmKbKQ2Ff91sg
GazNSJmFWUyZ3IhUPpU4OfOL3w8zt/wMx47ayPNji660L04ohpJcCWP4+ro+bylyf8Yhl13VpVjq
SSK6kKyYOzv6do7tDZ5KJp1jn98GADh76qr+iDzd0IRsX+XWtUAvJh3mgsEtPY319jkCcY6nhTjV
b0FPJ6JCpyD4bjPNkfYBiFawQC7XpCZEyHxu0OBJReCc+yuV8Ga/UHin2Q0Ua9qoAaesJMAW+qXA
Zf2YC6ZsTeIdv5tVjYsYRk7lRVwdv2IXYFLNQE2cr0ve9ln+H/HFTPjlgm3wwSq3Lj2YS9ITZ6hf
W1q5byezbVbQDuH+nZlZDUg9NF4RwPMuJCT4p5DS24wOAjva23UyO/tDL+jvvjzHWU7FIG3aqtkV
vkP6wTuJL1txwP4N+rMZNxPZhqM8Oyyr3rywRn2vtBP+hU3butmWRAfgh8CaKD+P95ISoUxIq5oS
Tf7ez2dAfQUcCgMrL9ONIslJLazJdk8GuIsYNENKQk39Uqks6f6N8wYgTa7+05feuxM9czhHcKXQ
Sh1YUkbrdl8oxMayGk1TqC/qkP232JmOtmSqIMPCf40FuwsdhR7Hjx1KLdefGZUGzLl4AkXJyyFc
kgPgx6TTwO22SvJWta5vhMLESV4VGUiky3JP7wqnD0ABz06FArnYtRGFOFCzWY90CuuRog8KiTo6
hM78bCCiakUWfRy924wt7y2L/sibYGhK2jTKeINcvaJDesCBUBpXFi3sYx+M4ZMRx+V+Airxporh
DwoKrvyRa47Qh+BpSNG/P1s0nt07A/fdWP66AcjHumfn6xMFEeUVnDWzNa2ej0OKzA0tDN/5gLe/
AiRAg80e30WG0DGcvPeJCAAkx3gHEX884lbaWU1qYafQhzxGVxKLP3Q5w13rLbV3Y+mFtpiDXDCx
RYZzCMXs4Od6V34ZPm7K+Any5SmoEUVKDr6v/+fW2KajPLGsGgMveKPyXS3VzXSbz2FymZm8MKND
AgxQagn8TpIFEsD/q7sVBfDiZ3hIwe8Ib8FsaqcD1XcWfSZPwRJU0g1YcfByr2gzcUCUmNtlPZRf
j0iJ1B3GQvqoqCn59liGAeIHg7vu3QnMJSfY6ww021a0F4zwpgFw6iYMgQZReMjCD/42dFcW202m
/FnGh0ih7hXD5s4EOd8RxwKM5eIHXHTJOwYCsLtS80PJr4o9ZWzNluuoyZ/68FF47oBlXrbdBEGO
4OpolQzYZ5sbwFeaaI7mipgb2OLPfodKDfcMQzfNeydcOXAP6RJsbk0DtyCDjlN/s3f385z5pkIq
6gG7xKFOpfc7f92UPejIMub38wKY2Rr71A9KnAFyheMxT2zrEsVVaJ8l+q7KYw207x4v2RtYmye5
rTvaSeATc3h4jEKDh7TMTnpozZzTmKGq5USaNqZZ+8CyoM3VxZKj/ZObDCbui/5GSiGvnJuOAdEr
jEYlu/4kwyMIfcUdETncGhHkfsVUZSlmcNbATal4SqvkPNiQuJKGkcZiKgjVZgcg9Pdy8JkIuQPB
a8G6ml8itww+zJUVIp9H5J5AlAmYaT2/GNy+YApJnEQuzbT8Dx2hI4rOOzyJ4+0/tVirGN6hQtyc
TKSH7HeneAoDQ/5SEzfMlDI+eVNAlgRqx7agViRetp3Nup8qR0leVu8DxkTMh9TTrzN8LNofAg1v
H1wDDWgh5sVf1ZyiSw+J46UxOE0VKtqhXrjT2iKLL3AGp18rNmDg2dnnLmGKyi1vlNi+rJ5uOH1X
7AWHraZaZ1KVEuS13RWuVDt8yeYKQpkFiH3QPROuU7+adWzlB06oPECSgzdpehb61qHqOxJek02T
vaPmaX0+UEBznj46IVsp0fJI1W+0kiRTKSpUMHUzVYv2KmT34Tw2RGmXe+ctTjJ9e1t3MTASm6pk
LrqhCLOSH4LgUoLSIKxsCdeQgc6lTPykvPa9zXCRtsGRpLZnezAzCZMUxlsEi99No2NHlnbVFaCJ
pF7HgNMybTUB9oRP/3u8YOYJDsdYk8WF3wnSFdDHCZ6yVu+l7mQegbpvKdkQ2e1i/613cmLy32cu
o24jmfmRSo1j4cFYBxj7IxSBuGDP/iSRBb1y1ifQXLro6+XnXtHtLqy9U5zZ6vlhTeZa44tgMnej
tFYmQjHgkZXNDtffFyU7i0JwFYeogHZznOVAniJXNL95X04+DuK3R1Vnxtn/S8V/ALbSwu1oFUm5
sdbJbX836AudTORBQxn70qTv5E8ZycbPHwBbKej5aq1TgVKWvxKbGH5RFipOwPIj/EzEGUoR5vVq
kV7LZXN15+vzStW5tg3CvTz7cbLWPcBCH4JOZRmDloPOKP85+c4Xnd6hd8zFlVczH/6QmroJl4Ah
DEjbtwJ44Qu53nFKEMrQCzd5wlHvqKC/nHU0zZXBN8zmxb958V+2l/DF85hjh1L7fgjoBfUTTExt
g0Ux0j/oLuIBZGJ+AoQ/pcDGzv8o2h4yE2KOsszoykRnlSVzKIkiP5byWNhm4jvGIzNMcYfp4JSb
uw0ZWoKsLx+EafBSEO8HYeI+CCED8TqebiPYsgojF14JuAcI6+7BiU2hy0E603ElF7RbKKpSr/qp
1kye6xYw0W+iDvyubozjFWD5kbZqyV7GKEiIxeyYiI6UJueORnLDg3KnJHKqyKtcOO+w70/1OGPK
QB8qhnQF+PtDfN8LRmGYKNw8eojyD7Vwm82Z+FtFe63XyKU0A1eHmO6ZgRrrjv49H47PbQh9HwX7
4XsLbS727egyAIRZkEszXRYqHfKPBz7024wSysBDq+WJXdDFzUS2Xjj4XaHc0KEaSFT8agb0ZLVe
y3P/5MNGj+SB+czO1w18II324OxicUJfmb1s/Bp0tKhWoeK8CBj+Lm/S1FfzuN0tod02worTn4RM
13FVM4uYnp1eMPxxUeblY7bmArT3bq96NU/guDXj8GxPZhSqd1dAUn9eYO5h3bDCfj80uhfQH/G/
5scdbRUOx+Qo4E0JkI4EmxVepUJaqW7xUZ+TqXM5yGeYQYlkpzy/NTAe4ji+uXmXuQG7vjLY8sad
kGc3OigQAPl09Z9s47hdbdLW60JcAJZLkyip7Z3XHKd/bGd9y2eGMKJ5VX2QHLweqxEEtClSOw78
Yo005iwPPk6fEV/hW3hOXJ3QirMb3FqOD6DtJbhhSFtDDOXy4724A3M4aoCf93dEc9dT29X2RkhO
EBwycE1mni7orWNqte0Zw0ULaM08U0H5Wsicmex/gEc5hQZqUxXQyVoSKbr9+s7k4ni7HOnjcP4X
eI/uhtLNfRZ1BdjMAqOuNd8lGES/b50wyy/+SmtTrXCpeQobWsbI4SEjQhLPldye8DFkFSbNDDcG
6IEsJNwm3dPOlqEfeMZYClo3qzItWsFayXb9CbQ0YNAhOPFmRvwMDr2dhJ5/8nWCzvzf448+NZie
bI9/5/P5hg9Ubf8/eUHgIBMLfT0kR1P73hY12oe+kRH0TQJOMn0EmzFsYPh2mVf1OVBmxDqcQZps
PRqI8/e+pggt54sBWGVGGYCn3F8iIFVezI19a8Wye2rIqXsTXQRgJRckvf33yG9OkMQtCSKswMi9
YPR0XpnUuhoRIS9uLG/8mBsb0Z0vkZbq6OZFmxohcO6s9P/junydLUf8YaqLCra8+JG1SSi6SWxn
R028L9/i/dtSiKnLjVoQ0J/hnKBATQWiEo6ADkcPqZG6TuAvx8kqdC/qeI5ytMuk2Mj3XIqoIEVQ
aG0Vi6UCsjF7+5k2MiT1m2TV2y68mEhaJNmAydg2yIe1r0dSA6dXA5WfG050RuJNQP6DzIrizCDV
1AgDk8qWlbRDcGQLmQNkknIe1pjz5GxHNhpLGUCTFAOmACPVW6GwGZ4Lv7JaMKv3jqzClSNlM/ny
6RZhj5Aci7PpM49HxG+gPLjgMrKVD5uzgxcSVLvSkV7Oywok0Fe/PKXDK/zJ5RErAYInyFErmf1B
6KgOaeQ0zNPywdGDjOj3ng02IrJ7OaIBfzSOO7l+ssld9DUk0UTCdB1dRXCc/EGCVR2b7Jfu1Y8Z
dlnW2Zf09JlFHpeThq+bQ5pxh2DA2tE1Qih/VNgMtUIpxvunF7Duo6sv0AfGn9midihJP2aFF7a9
YPptVhDtJMD3P1KvAFM37i/KGKJtllMCyEjzSSLJoAzLhldDNqeSB4xf37Wf+iaJQmdm/a8nNCtU
9OBx4wRFM5ZmXe8AviRwpMiC0yQZFJdfa6hgSKtBCQC1DCsBT3O2vxN8Rru0MyUlghwSEq7+2IXZ
u2p/rY6b7dHcG8eWc+0jr6gI+qWyF2OidNOJ6GSFXljV1mmB1cCMb+BzEXh5WqPqdrscHGW2ID3B
zFiER2ootu9csijyTwDZij9Do6+eVdqqi88uk0ChHd6JMjSSmTAJ3ljo7g3zF+pQ/c0TR37tIyuL
Qj3ecYs1bcAOIeRycACXFRBUs3fnqYKph45qehgIZNUm/8VK2YRvUqenmIcePMGh2G/gfUBPZyty
oSrIYo7Samon1+NYPa3hibkUnW4w72VHcLYwd/8ZQq2FPhtg3XQc5vfOEDv4Krp94o/x9a7kYpky
k1vQA6Hpcgy5s6qlsM/TZa7WeTJBbOK1jJ/iTUfTzv1CZaSI0AsLFgmZKsZcHe4RhG5iQo9W4nus
aE93xOFkV6fqBxkYgZnZdG9WJ+B7pfP9fg8lI90FCQcwPryGVwq6qrPmWhduiuITKEHlzR1F6LSp
BZCu9ShOK3pUb7E4Ydq102C1HYMS5vSCc75aEUy59i2CUEtpXU1VRTGR/1C7IOV5XfXhYipc9vYp
g7Qq7vUq97JTRqhVWGGncQ5CjsK4q4BWCS+Nu7wP1HivX24lL6s4uRjKtqX19IBgua0Ylqqlt5iV
3tzR4jDtZ8rdhq1hGf4wCT1wdp1gkeFEpgnupC5b42eap1C4965/vR7ou3ybTwUFA02uB8ErVojY
Q7EkX4Vc4zK1CDhuEgKC2iaFkyGSM83MBWH+uDOzGjr1tEmn0IS8vH+ECCMhmaCMLy+nonEB4qwf
+gk549wPn4QcJVF6S5Dy5NWJ8Q31Hs5DFGqfWEHtAfIcwD5uHcq9MNPjYXaeRNQaQH/NvCLbS/7i
/6wuF+yNwdWmRGK8ox/htYujDskk9U3qAjIrhRKNN/4ch4/QSi/lncIODj+NF4vnZxniYQWIW+9X
uRGLfw3zdgnDf0qmAhDNTVGNgQKlqNIVfsphyeeD1LdSZRNR157zXP7H2CVhi1dNIvaMIXsSEavw
yJ+VMFuWS/6BnMcUs/z8FBlXOzwT4JCcD1wdAX6z+s62wkl9fvDHoWrcOUHMBqDmTrcw5Kod8vkX
72xe4JXuzFCXhd7T61FZDm1U+3bpRFXg+9XranuGz2IYC5UcPFNWzWAPoQRxiwGEHALD/4OkLA7I
4RCCODnV+7YSfSc4FWzmx823ugvqDwQge5tIQof46qhPO4/ZCPdZVBwdTzaPs/aoixu0h+3kDhPB
qIfJ3BrLS4cBdTxgmK9wHvpnIcrnoV9jvb/Ixx5gP7ipn4hXZIbBpo/Izzweug1biSUHer9rG5Gi
mEEG7OUKu4Ob4osnlyVKM6f1CLuUx8bn3wHl8YgemqwmHPkEDkxd1hMsy952t5WaNFrCdwgd4zap
Ih7TfeB+YCYIbc6UAn6pBbKEu6FR1VHtds2Hb0QNEA52A/2iKiRTDcDOa63gSE5tG8StxlPdslxc
v+11a+WmigrvV3Fq9pLcwsOCsWgEIapHSI78adTlq76mRQ/1m9s+x2P5S0eJ9KD/sRNoekyIjJlc
BUTzzPEYHBWm890dkh+apeAEWEzNrfJpyPAAlVSJBI9ovdsuoI55BpjXvra2bZWLc+RXr4AecKim
9BpngqR4HfC9FIa6QdyHDUTGmN6+PCxHw+vXOriRxLXg5HwJe9HQh6t5Cu/Ul9MFTD6a2+Uvw2Jh
uzXJrWn1ITMdowInswPui5rs7b6g7cxAwl5ELNSoqsCq6SrztQIQhlYgUREhsX0VfVNZUlVVxGeG
bpVfpYA6zpjMopv3ZD8ttCSNy5+Hh55x1HyXmE4SrXSIXFhl6Qtl2s20Gcqs1DxwiDMsXVhWgllr
fFnKeiClxPSoqwQd4HmOP0/OQsu9lSZZ0mEqHShukbSMI1vbNuN/NO2piYem5m+Van5q6wFmKfTp
wI7pttXMqRG6VuDjrhlj7wbjEtLx4U3x7N/K+AXbJeSmrhBVEsglre/ZScZZZF9ZFtaxJmZQKo6R
9qSUNp9Ys0kYUoFoBugGut8ZYu8X7Yb4k3bLNltZOFOqn7f4DP+sJ4TH8V15is/5a/vZigxxf1fS
wUtZjbOYMM/JBgKq0KST36SQkpXzMD9NPisDAaGy2oOuTrH+I4hk5f2Eiv2KdHA2mvj1fXVdIRIh
Ql+h5p6u7OM5IgDgRdr5rAkAXqA8IoA57D/9YpofcomLZtpoAiEFC5kfg7V2F+hyaAcrwSpOQc+W
Rg6hHfe8kcC24TCabd+v9jn/SWhjB0Mp3VvjI9qIz65oLo9IkCPvEpFaNO8xSqQ0R9S6ifz+yuy8
vOU5//gua8aGtcmfGYkNYy/GmSV7y5yhMpTfXN+I//11HZXpjl9mk3b7p19MIh6L4ZuUk63oxPh2
loU6SG2JGSWdidXnkHp2kUld9J04u9d98RJ6W15cSvps/cFmMGiTh3QnPlUIuksZY0nNXiPICtaY
wUUMxmJL5C7ARnglJEulvhmBCvA5R1tzmuSixvg2Sm1DXKru44L1q+vvOTFu+cCdw2OarGvgt3gl
/EBWhC0xUKZ3dptmHkGHp9vN+x0/SIpcL2SbAJlDilcq9BnAZlrHqCYg+W58YGPO8KHzzbOUiCQ9
CO4MlpxhInZ1YVwcp5zikllcTEQf0FgPnRW+4ErLjI0lqjYt76yvaCc/H51+P27mosslwMWzPnyE
FDfd84VVMPlL9VoXHKQxW4IhX1UhmYtg47vIIH4wHE8vRKSID+V4FYNFyVFKvtAcVA7+B7uy8qwC
yIrlEGBHckQE+Ie6PeVJmGcthW6ntF+0itylWPxcE09+etvg3bpg+BmqietPs3JGIg9aramYZeWy
Gyq7yDPhhKwaSRA6kq6RDp3KRZ4c1Ri+snsFHLXUIbUPAFi0az5L0WHxooEauGJF3/EORodqCfR0
i397tddrAEAozwdkgs8kycAM1HQa2LldA2fRfhY/8L3X1DWP7+ralGYxDjjccVoHp4TJAI2xSA7Z
QqB4GL7PkjvmZ5OT2SKxzN9onrEH9CoiNa7o7albxSqqZZbu9FfWbxwS5SR9LySfwnA0vPWe4bOe
EUkGkS7IfZa7aUT+IXoKOQObQ8X6/QEnAU2nni8Zb4lYU9MAAeoxNELzluEMh8C5HfIo5na1RFtK
xJ5Jcl9++Qjoocv+2vF4yB2sBibNArsfxAxCVe4wk7YAPmw0lXQlXxG+ycvI+DgmNWzBAy7SGVi+
fvFHZEXnhIQWrA+w2xZhyPP61wokUbMuKGKIGHwNrxoIPHAuQ2/FAOf1cFQX7ps/Sp7Ax/v8uMxI
Fhy9Jp7d+WOt2Zeb6pzBsCA7uhKYYT/mrzHXmLJQjkHJm3hknJ+jKP3IoE42JDvquUmc5r/CbNZi
aBgwdo5FAQ7HaA0eV2jp0qr3/L1pZN5I3U/D47rzprSOM79wySsGip3bpo2fF9JMQv7KnBKk66va
2iyftf07OTulp+mcRREx8Y+nmoca9wFbV87UfyykjJvfRwAL7sg1C0zB32UsERsTvozJ5BQYNM/b
a10AzAmDsaSCpPvZbVdJJj0lB8pWLRDmBBq7obn/aXMOiWgdIY26IQT8bMz6Fwnu/vr1RLXDmB4b
7V9+Kajjnr4nuajwzw7+3D1ZgRzCBr8dUz1j7tuXH2jxEX2tPUx7dP+TUaggY2+JU3Tpf7vqnV0p
1BVVaWWDCiOtypSVy3jf8WvNpe3XP6NE9jyyxOkGAq85YbE7AJ7CyP02g9fUb+I2CTFZmQzADzqz
LS2gTlpVzIBDx7dLY/M3rXqPRof+LQt03PGfxybtiN7q3lxCzZCfttXsxKqk4MzOBf9CEME3IelD
NOSuubNKQef4WcCZDzXTBHYUZ3ahaZO9rbSEn/Qk90Ov/snSvU+PUDhh7cGDw4/uE0eSoqT0H+25
ZhKa+du7/bKHGpJunO/86y7mSyUzZZ4fIEc0eUjMu+uUQsRKhp4uxBsTD73CLP80Bh+WWGioaNvo
ewTytko1EboxkF6HALzyd2GNWRmjyW0ZVXyMh2HCJJ2Xx5K0oSaA8PH9lFzD4AZQ7FSVGpadzDZs
P2u4jOcriYtPBcjKbcErijAHnY4SV5AXD4cavttVqNlomX8W+IAhLosgUZs5IFCZlcCyDoovnzoP
h59BsFhUsah8vYrhJYwoH2Ntudg1rUbHVxi5tDHLyyVwef8yMjnclbfNif9/k+i82uuN82Nai8/i
JmQhMDfi8GHharl2srkioI3QPJD36w5mB0e+hvuxhwOwfoDjCS/fTL1hLh2T8Qdg4KHDux3OlL7J
sXMtucGh7RtHkDQpkcIIYvCCNybUyhQlCIV4j71G19MQPbhtJwOcfQqamrKcGRq5Maevqck0QheN
BkqcgnlOErDtXQXSwRhIXCfIqFZHUNdP1JnVI45qIAYKpG+jD6q9jtDCkL8A5S55gb8KVAfR+05R
rZSUL+yAGpL2AJO2rNICQGnLFtPH3lBkFyGw/LVt8S8GLEmT0df3ns9gQop4aKFcCc1gSe+1laGo
mQsWxRS1IdGO8U3PVqVU51mn332tE92ShHNLU8Ap6d2p7nFSDctRnMYL5NgIeaETsAbZCKoX5KLC
AQ+oQPvTffpqBlZyMh7EQWIjRsNIy9ByyFI8vQvYPcFzDd8kaImS625f4GBNzKaKHr1PX39JVOgw
ngOa9obLieiKN7faoOqb77JHCuKy6kar5dLHg4fEIG/7CxGV5vMbNweHhQCKUpJpmsk3pcT8psfu
UaxC0dxwJQcSHZJt0XXP3Bi2uX3Ti7IN3wCO0PdykP+DToyAacVmBsuaiQFT/lNl33I5E+6295so
LLLJbkI1vQcjpYsy1ZSOgopA8DxmgUHwWEXusqf9TU8a3rv+ftvqLvTdcuCAi+GPwjA03rvjeyZ2
t+KqtKznHyRWZJ5nXEc0nrnyde3kWyU6kF1F3WLHew2ATNx81USUiA4ZxvHIMByLBenRedrq+cpR
hVIh5hku8sjeNCougVmIIwuh5vaH2PCXbVoOcHvj3zfYhfdSB/Rr+NFAv3L4mHTgKLtBs0I309dG
RGNzE9eh77amfDWTDVOiJe7vcv91xGTiKfn/Bs5Qs6HyYsRhKDZnp5wxcISPcdAxi5CtV8rZSlAW
KUdRNyZj+oKJ0p8daUmZ6fXQbD8++/8bYBIBHZOlH7KUH5Uva4ep3YDPdpu5mRnEeADjt92jDPfn
9KMxg5uo/MliAJWWXVbZH9LypvaR9sKODvZcRz++4HyktxJAu7ljAldOp6muVpCcb5IiUN9nHM+/
1h9pEZNdJ+6oAJFscVRIo/abhrjpdI+z2M4l10bi9RjTOO3QWCu7zy0ciA6U2UmGuo9KkDWU4lsd
xIRqlck7IK5U/LWuCBUXvCjJf82XBhqlZvYcmnCR8r0a/RR3COWT9YGALQdD3pn6JKLiWMNDmpHz
J5Pl/UF2cbe35jq0hZOZgdn5ymXXpRFhmJVWgAprso6SWI3CUlcODjnYUQJ95tqX9krPODE4MXJm
AcmwGjl2qJGMCD4Ahtdk/UuU2iz3hZOtFJODVfEIc+R4JLp6INfwGD3oXR7PDqAqczGaVfZVe53p
ls842quhkiNCxnkMFmWwNlFCHPpnNuAcqOerOjpd84j1S97o+L3HR9cZGFzDDDTOpeV+P9vgzN8n
hIYJMird00Z5TikE/xWMjs93IFM2Lbz3Lvq0qBL2UdqORsDpiZymUCFPaRcltky35DJwutCrb4aG
6igjbClRGURF0na3SicyiDlB7wUmQr62vZ96B8WW+vHBD0/UvgCcekFfij+zk8r5oE6/+GWPWxmu
dyoStsNXcRFC9fyR9Xa4pzujjQ4fzbhSWhU8ILqanPy2cxP2w5i7lKg9zBIA8AskbIjNXUCBP3dU
WZ6NP9UyXDi6syHSGWXCQLWAQ17QySIENAa02DbSuFwOSUXokEEadCSDhUtkbaXixziA5j7DV0wG
k79vxBb7Ie3YBlvZNOzMXFEQia8GpQqzZQbmhDsOrSbtgKMZHNUyEDvUxnRQ1VauNTJ4B0vO7onY
XK50aMIDdF3/oeQmWZXSR+EVzKc4DvR3BK8BXoZrJUNOyJDuW6pNzJnL8MElSl8FmU0MpnYUtWHE
zTnJxoBu09uWRbpJWsrbO6Ypn5EPte/mLv647OQftzkLWRzqoHROTdpfKK/ONxUKLtjK7N/JsRT6
6WHFvEoh4+fGQfP4C61fSk29331GvekaoMk4hNg3Pmx9HtTEnQe3s9hSb1zQG6liVucSDXkuCYJz
QZnoNxMaZnf45ckfWUnoIlfKRkOrxZYjawJH/SLG+0KAA3jLKtkXzo9xzUDx1nk9DfaQOuG2Dd0u
O5DN4ACZxDhIybt2efK5SfOZOZoF5z+MYZXKrfIU67E6t5nkbnwtZJ8XjycI0ao7P4R/BZGWQaku
MbFgGrBbQaYR1K9Rr5N0DRez8BfbGwnv6LMvTAewAzJxgD4OY2b9OywGVZcspKMkkeTILAZ7P54L
r/KCJZHxGi/dhMIWG9FnOK8ACUhbeM1m56Ja9nlVfCB6ACkkiUi4ZKlrA42AQuUvk67ZlhVDEVUG
bfgcpFMYN/zSnT513i6FbMB6cH07AIBbmZgv59DtHFe70KGhCtBvD/C0+jjk7Ea1WJ1Y3J5cmd4n
gvPX3ohjLOIRJTkug91DcRad+6RAHduFUAZ5CsgtQn8ILu7FLQUxh0yl6dLKRLPv6QrFF/3MbBy3
AdHJ6bONCwmlDN3AmFTkLwD65f45yl0+jgAD+1Bhw5Ux/3gwIwCcnNzDP9eLzmKxyGm6SmXPP/kW
Upn8NeUVex5Vuke7+ukDWUQy88/ec1dHfZR4M4tcMvEUrexP8WUIIXMcAV0XbFDFGcjTLo2or2hz
nR0Q9OJIZd/rbfwwUKfzcySyjn6pvxUgI5YPSJo+dh8DTNBWSq8iLAiCEHSG0Z1LxpEJJ5o/7xJ3
Kx9cw8ITo7cjfTegOE6A2aSF6ZjCx20CoWdvYyBhy/Ova9hXcgc4e7UDm8PDzJtHYo6VwxP28OAg
y+gtgajqMbAmZVuvV5Hz22LiAKEvU/KQr5BfigdJpgMQ5n4F+1a2kk87HVCztWe+y049bmn4bs0A
JGnG45ib6Qb+W1zeGqbwHzUpyyGmPSWaSQEJOOtBRA/gS0y2iwzxUizxMMsKtZXHMfLPYXcN2Mim
X0vVwVL0SusdEuVzcXjs17LDUrI1VzixetJgYd7LhMdpBeTATyIhd7mbVSYe44CzKscJXOiIWqoN
kjVK9LqDv+VL685UJ1E0TuDIH/YtGtFTuMa44+5+hq3KlQIlAGDMl04vX50D2tqu5nFW1wZ3Oozj
DgoIjfYfvFHVeobD7zpTmbjJ4kb9BEXd6Pfbfui+Se9zYE2aK6+JxMeB5NRf9dqHi/ZeGLhl22ZE
xzucmIdwsHG32qLClh2hfFedcXyyV5SJJLYVbqqe3g7jrsEVuzxLp4+D7SGeZCT0tOWEwuCO5aaV
QMX8o/xYhn5zb1YOnz62uylDWnhqXHnPA9MSPu8OP0OjlDQ3UCdxPdiTH7QBU/fKpMjfss+D9Uet
AW38jGFJ1qGQCQJltgkBabHN8PQV/ncZ93QBAhX0xB8BmGlU4lBFGejnVXnzdHVbz0UacAFkoOQX
KQl8p3khB5gWbt3DQFRjSX0VMvrMf9+kroBxIRtIkk879V3Rpn0e8vq/2P/0zDb+AAEIg4EfLsaD
7vqj8N3UD6FWEdzDbC3fH0TpFogXMPeIatxmK+89EJ7S8xzDaoarDMfHUf3YWPA6+dRFuWaPu/TX
P8rxYWg+5eEp988c237coJ9Bki/+lpsY+bNaJJ0UOgw3g/yRj35XsgMqm0w4aOQ2g4I817J9WTyP
jQCkg4KMJNeYkPdD2BjRK1THSNH6jf2sCYO1skWhvoiG1rVN97vzX6T/x4R4MMTsnSnKPLregvcj
QDdcH8MblYwYFEy02jeVsh5tPHA3uKgQEQfYk8mDJR7cEulzatGEGue+peKP4qhXvWWwVkEuxRAX
ytQn8IzgbWu4wtie4CTyWymVMWwl0c4qIJHdAOFNODVgZkr9EOj4bW4y+rNfhQ3CNyKWho3S90We
6o123VuUlJHOWnhRWuDogiRcN4ivmwWfhBDJg1gucbzMo8Z/SyCuJ1USvC4JvTMw6EqOBjvteu41
/vM5KFhQAQ9ip/vwjvErZdOkvOuglA3dewgQslwuka+OTpvCE9AkVvsavYM4A0w0Z/D0R53c6VS0
8Rc/24fBLEyUwPyT58K7ITS6ZrS6k3U0E0mvwInXm1ae8rGTV1gh2TMoKqd8SwEQpyAiZq5WjFQr
MjVohRAIeWROHF2T54x7RLPjXLaK9oIZjlhGBl/i+K6eR0VVcmFB6+C98nJvtm3s0TOQCfi9eOMG
T2C1RifHiGdsB09uiVfZpjnkz9k5usrdnCFVcz0Vc2IOrkR0bke2KipTCn/qlVtfDEsGhaPtysCM
06VM6uOEKGCtDmH9yC98SoeyhFsdO+bD2LrEnSBVZcgHvEWmMc8UDptMI7z8dyVXebBHnAq5bTos
xnZeVwqevbqccyy50jBwYbqG4aIbPGD8S7OiYfynORKHlOC0i3EzZOZvX21MF2O1nSc0eTnlDayK
v2PJ5aOtLhncG4YbQWBNa7P8E6nLFVjTKk94+e4n6bjG3gVX+q5xu6FF2zZOYR4rmJn6K8IJx+Kg
LAJ6DO2HP55gu1cb/XZbl3pgj/RX7jvEWLfsW6yvUUsxl23YmlGrf7TRXMM11gOvZgyL75TNcqGQ
x/MrRPOTNPGuwUt6CZriSK3Cwt4iy9AmDPvNFP0Our3Rn5BboOwCKw3P/lD4PTwhJ7Fs9+kH0ex2
dVqbTmPhW2W19jyFPHndAseIr5cZsHA3/iK6EmdqQmA3tH9mbyReAmfES3ul+DWLkQgLHXOMD0MI
vVY8eh8379YKyLO1w1sMAkHrYYS2cJvWzTpuiAmRFFkjGp3jqvkMUNJgczxxbivODH26nX3CnyWH
R82lTF2kRlFzv5UBNxZoHS3G3eptHwvtkRjwC/LmEg6chqhwcYAsflVWJgr/krSwKXqzpjTo5kE8
QAiXjRafm8qg9dnGKnwONhR3jrJA1nzCQ3ucSAWzktfkJQFiYuHzzwybEEeuO7vZKhf2E79N2F6J
1vhBa86jsLlHsc9nw9oQWX1cNSuptm4XwYwR9TkR56Mjs5FPNI6R46Cwv0Q+qHlFGGgDQ4JXClLO
GB5zjXUu6tvqoiEP4GoSyk3nYfzFe5GYr8eO8wuxzcwxWnhy54JD9QzsJitHTfR4zh0aztCLFytX
HTFuOem2G/rYW7rHIVYILFCwRo+6SSwWCD/Re+zmAwZ7hzck6aGqTYhX2ItL7VoE0UyuM4FaqExX
7rW1T+MzOdcye4KN3DFB4RSiWNP4TIBc94lyA4morBpAwVsn+Im+dt1h4+Tc/8WxQ6Kodi+yJ6xz
K1k2CJ9Afk0xOm+doy7xzRLqHpy8fq41wG79XD2oHQ+0i3pwXlhcmxzRqENLsFRE6oOyNa7EHYp0
k2eeewBabGFQByAdAwXo9r8q2MGbi3e2v94uGBKk7gFsCKk3TWl7udqQXvA+weStZiLk4C4iqf+D
3KI1I8JR+kyj7TfCWImgxTl6Rd6J88ADbNlkmE13TSRxsbTR3L9aq8R9tPJ1Dj+ZPpBMtIafmWne
zY/UbeWp01lIfnetKwkS2oZcrokEiqMpxRo3QP0EeBmtVZ3mZySu9dWXN8OM6ZEbhCA4KqpF+TLA
iNAHnccSXB0KXd72F6wUaWUxr6oIONei/yMGlrKuXzWSyl+bEizLOnNDOLKlr0hypNVWWl62zoHG
L74Pnm25tycIMW56MwiOq52i/oEdUVundlFMq2aZJB8gOr4/ndKGpaQf8ZeR3Wq204M+xBIDP7sX
UfHQIQy3TpD7k+1BSgfAVffw02hjw8Ou1e08yFFxqjRDA9/H5WzW3R6hD4XJncnL/fzGdRZytOlA
kRaHxRsE1bHA8cZBve27W7P2qSgBEq5dxi+HAUACHSO5ulhi2iY98eCU98ctrhVCcwoWab7qhvF7
4gTJarHOxXqxjVM5gDAETcYotTWI7Dg9snNDbC5bOJDkN4Spl1rkB1KuUjYXIr6I0YW55SfvDHcp
7MBdnXyYg3HM4umhqWah8/WZMTIuW3IBH1l5IZvK/x4pleIqQIG39mDPqAsWrr/JZlXkz/me4UpZ
OymY78AmGMnDNrfBTS93+CRB16AQtQvSwh03Fj8grSBE0xuWI7Hp+dOTiHoT16q0IZIscgnkjvGu
82ahOghjHuaIN+5S/VeX6/QO3ZCQODcd/6IdCpQb4IEt5LMI+2K9ALwYcBVqM6iVDAufTMTYFQd2
CoCCJtsjvacDNbHB1he668WH3nTQWBzuRz6SRjeWkfAXDyqHVNoGSHusq9cDnZbxRGjklaN4Oe5h
4upJxQh1lf0/cInquGTtRJjJ6mDZQLZ/+ygUjWeoNN8rT366GuDZTi0foCb4xns0cPiKZnDTgzsg
qJU29FZyEenOHLfTOlfPdO2aLyt+52o6Fg7AyM1lQtgFkWhXBHB3Sq3rVp3rWEypcVQGbw5kpqcF
eXDQ0FLlCNs6abWkdZ015NBl+V9LFHtsVjFWcd8w48kGa4/Wcl3/ROQtl1h2AT2RE70nxSJvzM9j
ZVFsT/34MpqUrBO/CYsEcOm/5CKlIm9i7+3CY9wO9gCA3US2nGQz/t0HkAK/D5C53HDDWVikkqNf
PjmbvREi5Via/413eWebT/NRkpybHVLn3EvABYo/6E/aXNRqEiUbiPtqygXCKf9Nlm3kohEIGz5C
3cqJilEODN6BN/M0bTqQLwCkhG+8+xN6HshPBoV7F9qHWwiFyQ4sa8TI/iiqf2Fay49VqdXQlu8a
MclDyQEjZDc48H9F4hak6zg1rFbXHROJjxy/MuXCV3CLEX89YL0DlpXD/n8kMLPHXuehkuDus0hw
+gfOZROFOtAeN3HHAJ/WpgC+tjEtJJ1+uudWJmchOvtNAD15STYmG12PCAgT/bUe7Jvhyl15oVFk
mprmycUFn4Z5T2auWihG5kap+i4MuVQeYoJkDkU9CB/joiJnDDjNIGxIsjrI+9adDjGWfzKq29PR
0T3yh+jeaJ8dYpEQMPIldr3kOnpIZ5RXNAceq6QwKWutNHz/4556PFIs8EAEDNM9L7d26/hnThnh
t/lCl+niqBG/3je2FbzGQVVKMO7rWaBWAnIsWJEqTbTlsRMJTT4+qGW2YR+eAH6isOGIKyMrcieg
g7a0RGzD1Zf3amQgZLmdOcQkmdmLfoUQKht2Q8SolhZLKbbCYX+Fn2zZNu4Lt9CKiRFDMB/stLfu
2/JIQ/Yda6KzMrU0c/KpYpBfZqOfGLPaGhCTdFJc8vlH9aP6vZT/UulRB+5Td4/6amRNP5oH0uYw
G8ItOvEwbLnmBWn4eqj2EUdk76eeY4sG+HS47m5M2u+bJv8U7mSpIHKPIpxwkM6IqahS6XdT08Vp
Zys3OMfA/UCezbtKxoU0nwf0YElQZ05Rm9JvIrPQrXsBP0PvXJWlgVBNOHxG+nhIUDAQjzbYY/bP
yD7lNOMvn2fr3J5qOTBS/+82wRhqg++NBJs0p1BTXcB70XwTG6fhuHWvMMwQ9X+GfanUWWB/nct9
KHu929EK1BTpLUD5gxXE8KbJypPfyubEnXrOr54w6Uswn0zeri+CMhjJ6Jgz7Emtsh+yTygLzhW5
mx+55wYaDYDwxcBZgfNRCv9tENHekuM6U3a/z4PVDUFLQdJV2AWHWcUYPwoOOgteFa+2oaWThCA+
z9J31m+m3GVDjA+jzRFbexPID3CfRw1+o9iBC8Qz86F/ymK4psg6j01fA7js9ARNR8SLgpQvHlkr
U4FTaccunXJ8WDAU44UdCR3dmndI0YjUA/59GS/w8/nZH7aQbAU5dCqAZDfYHsyhD2D4533upEb2
85Qb4lhueg83ipYrIVmfM3RR1sJsPJG22uUvcAsNBw0fNeka9YeaAJr1IoozweuLEbvFz1e+c40+
9YehwT4Q0h1OLx369IE2qkOTxHrKiRHCzNT37xR6yrXYBKCsEu/YMcdVkYjrN3hXlb/7AaKtHUyi
5KpWjAkqsEXud+6JX+yRVgjW/rDvjdmQ8UIOZcfbB1Oo7xQfK/RkdrsxS/bcDLVdX14Z47WSnkhU
FNbx8p0AFFv/OrLwXajlzYkdBc148i6pxKavcdBlyAmxiQJhYMFh2cNZmY3pQYB0FMSoNfrzZeIN
ya17LmCN8kuzReUikkMS5L3nKj1kpbWiVgoKQdZKr+E2DbvwIQy5Vm8YWvM83qs1W6M126ugq1Xj
szfqjGkY/Ejz4n01ZUPJY9aktqWwKzInPA4YazoA9+mbdSttkS8EMhie0PagsMCj+nYa2XvhpcZL
k52FYhnWaahCfjc7rfU0/fmzyL+6IsrFVoHyKnQENRnkJhBuIMq1nyFtPnUfMk3ZIwHVBUB8ZBvp
1ljo2JbGHi2LCMpITO2XAH4+kSTpj7P3kqZ52Ccdb2h75OQ0XsCX3/s5cHTMDUDlsLIVyUFHNgO/
LQemS8Lw8zEGLFLHxxIt85MuAGe2JxRJCYT7TwoeblA1+K9MZsp7ELromtqMej11EbWB0laQIIzP
8P5Jro2FIKUoeQxawqE2azqUOnJXL96h7kq0tklvvJotwU6kxUXnilG7tZrzwmfE9tXE/Dxb6q1U
KjRLgurjUmBxLkiJs55Pywm+7TDKLa/ABqH8wMpLl1cr8D7a7YlRztuteW+dfzpDMG6b99mF/p8f
UQ4+od0bVoHms1fRFyybDt1emUoCoOnCel2LtAY0KOMmJz4xB37yxIqxJxilgkpLu12sJIUDOivX
CqESaNEllVMSKWBKAZvxEACEh6ep/EC2BuxC47yoDwXadVJ2Gjen463GO/xiivwO+BS86rKdRpiK
vEUvp5jeI1mKb+i/KXXk8b0ko3nMnI/NwMhLh4IZ1+4BJ21+aYygrjCdOSq9j4uhTBfCzsBekw33
nhmlLVkKaFm1jLeRH9orNLJsmvjswc2tTddvSxDfYNAOfqutaRVb/73eibA3U6YMK9FtpUv+B1SB
z4ke7kp6DfYzA/uD8tIT4WOjAERqTQxdI8qxSsChBzAmUf3CuYgKicfALFrvIYhMvs0atY3t/wHf
BqJLqTwwpkWCgKmwaN0K+XRPGHzOgNSzqA6lAj5veLSd86hwfikareA+azYgavCIW7vZY6WrNsbN
EdTjN8ah+BI9YoEGzdy5BkwA+UsLfeBFZ4cZmW77bKQFbl2rvb4hhhGUCZM6/wtCpsYgZioKMzcP
I+HVA/zXdDD4Xsi7m3vizQdYnnVtDijPa/dM5NGN0IbM2Ls1JnywpuNVhdV5vvuuzcKqv0p2Gqn1
GPR6uFlFy1IPdl36tdsCO/hlhwvC2ZjuXYjvJ2WYA0gEcpaN2ycOGgkvV/8XbsEI0lblIp0hmQbb
C/+OPKhII5ykKUb2Q+IQ6TqdcYJMm/eFOyPH/LEz529IZ2tFBFkpubxpmOSd43Zuf2Uw6HnMuM6k
I/b350hRul6hWieXi7tsKvb80QNkg+7DPzl38xXvNYG6oqxhe/4MSwE1v+1nqAyq9X81xCxzcJvh
sKj2dSXgf5vT9y2CXErE8J1ADPAfkf9sXrg9WSUqc5n5jeWz0JQgHMqSVpXdaEeWywRhwOMoGfeP
gxPnLiWAIkhFLB+AVHXI62ZmhqF/toKdUBOhECvlL0x5pYfjXZT0nWier7SxSFRE1e9vL+s+pCxV
Q7+xmbkEbJz8ztxxNBU7TEKSYg165AbMiR+Tqk0BNxfGhkAG1lLn9LJGzwUJr9DVFopiZoCbtP0d
x40IeYrIbfrTPnzSO53o8tLvEpYpvFCESADIiPqdPIseM9SfK+nMx82OhcBYd6vT/09g9kDDm3a0
4lJUDy0H+74K7bUHQgRYolBPXMgjWXFLF0J0mb6tJ7KcXCZofziCJetIR0mDP0cRdYIPlw/4GtCA
VcnYyBfnOJ7J6mCQjtO79YIAz6AdKr2J8E7LLJgr41cHKuRdz/MGwkkHt52tKwdpPWe6ADg+/Kyb
1soHIrk+I0qcyE1G6j5k5KYqNmqgQ1x/MG8/1TY23JrXGbR8cLuIIV+hcDAGdJBiEy2sxJnygi37
ugc9+apNH0itqLrh2IxwSVNHS0PiBJlk//CYH8saeLTy1rgCJU+f1i7mZkwt1K/kzm20ltMvQFba
rlBYFJJg/uDzXNUuPHQi5Hzvbys2axXG2aIkjM7ZYNcCwvglGpBlh6i1utFm3xHPItuOjbrxf+vk
hRUjJ0RWz8CZSheBRTjIWjsCewBOJmB3t3Yzlr+eFRy6jCllitk2cIZk7Hrgp1In4g/BCEiBuw0I
UShKBUiKN8kmoLZY3GTRIIgw3ABvCV2EMIVesVEsXqqg+YPnYd0VrEGc4HlGn7d+0Nh22eR5muOM
nxky75J25ELvStiNpSB7x+xr7/14nIT8Cvbzk3gPMxyEtFAx+IRml6brTLsIVNui2DTPQBH6VPRE
9ggM9Q8Pd/ygFcEwWYUwARF1p47z++QnEDJa+VK0M7u17B/8ht8Wgq+mH+q7ITOP4MZ6zahsvUKJ
KwBjIzgXiU1O/+sa/7t/V4tkqGFJrH+qs/LWQt30Cgz9Mo5uW5aMIqvJ8MIBvbIWT0CNevuGA3A3
mFjzhT3EYhFHIxO8udnggf7aRb80V6Sj3eN9aZ/yhCKtNsyxfLTDSE6z/kpseSMZNHzRL3EReJdq
drtBG/Lcb3j+7npPQqXaeCewcRaef0LL7ccJguQlHEEZfnpAZ9a45BxvoPMxXDT9fwQbrgllGxZD
RRHHwtqfVauDoWhzFxPTHhFgswMH8Gng/O99f+99vYOiCJAQFNHcf2RDm0q26sKztSoHMgEnKtWW
fNSBSLcuGrS9G/La4wdBNuS+bFyhhG4qTzWCYE9lXjahH20C1lGrTYJt9cTsWvBjQMxVfNeAfX/t
Wiuy81dw1Vtrf+2N1Z9U5RSuSN9m4NipX2NLCVomeb2HjqEyznnkczWfB01egya2xKFh1n/OUEFU
yvyB9SFIzOR+9POxZlD+5utwBmi60HMwTOjX+LVmHFwK48YW6XPRq3efcWFvsLZtRCwvmaHHzZw7
jlHl6c1OGgHYKg6G0OvQLcUqVi+gDaIqHacrRc8FZHVSg+ApR+941LOGIgHCxEh7WPQeLf0rcOX9
BdLQCtpsXzEdS2OLurkccDd4T58afA0dB1H/LLwxBiHXvbZu5JG3EVMaKZVc7oE+aqhwX+gFlYeX
ILLiuEU7mc1+sM854xX7tSBx0IiLx51KZoCwJJ/I6lnuqN9PPDhDIaeEpgut36Uk4NDoa0H5yeE4
pWl/9RicQCXXnhlcN+yZS//ztXxSgSW+312oTsM0uzYAcfAa+aP5T/LrF/Qtzim2C1YyB8yH7ix5
CCPKQoxVnKg2ekR4TUEBPjm4/cRH+Z/IoE8FYWRuDKDqyUaQQh0VVwqMhEpkfJO4tHfz+YqagSce
jO6nMYGgRsiknUp1dIkVdHGjPU+tttcG1t5bEt3/OwRYGluVX9Vxo1NKm3U9cy+SD+BwpBA0KNce
NHNi0MyyaKsvZi5AomJYVNBOJlhtH3/BzI3+G1Y+koSIILbbElwLjzIMIejMfwOxHzch2XuAeEYF
Taq8bu1CTrbJcDqQfVnmCD4XtD1V0zqGY3/yqRH93L7Cj74naj4bZvrIpy2fCqemiCOKrgWZVd+a
hvQs3dvhn+OugexBq+151aqoau++Qza+EihSVAoDV5001TABU0KTQ7s6XF9TYa22iUuCuGNgT6G9
Dzcg8FZZ/eXTtLgXyPRajbQFnR2q8bIOzqDZOBudsw778mJx1bIj95aR99sTZYASF16RTNBY2+Am
nS7loH+3YtZAZw3vvWHH4EqrT2/AafbWuNt6DFMnHNdoMPwipM02N4Vd8Wt+CuZfWiLNZ4PfVHX+
ePr+NkYIp0bwg79Mtc0aOaTPmrMscYOaY9maU49WEHawTZBHJkak3tE+h4a1fDKglCcmbvytFgrv
T06PocFCcrfkTdDLIuZRPQSj8e9JqPjG8mDXK6jhV/ZEiAXjZt9r4jARPi7VPZ1FvrLQI5NRlKPG
fO41VLeRftAG/cwnmWaHZkOmG4UT7X6j9POUIjEFdi4Ck545SWR8CCbnbvGLb5bMzOrCRmDUQyRg
ZsmGKwojxzFL4NiJXaLTN/Z1ehVgV6LmxH9eaL4OyGjK63hYmXZDbL3FBdFf8SPNeKPQVt8X1S31
PGt4lMeNfwkL7KiuftYY+dO88sF9jkG7SvzuQaUzTpp7q7XvmdXDRmkIrtGDT+7Se80vamJYONhP
U5G2okuovyq+2zFcQk0Ig9lfmiW6tsawBFxV+C1aQ9Pjc+ANSQ+/3/db9fHTs3sjDMqtltdLcAB2
yi8tFMy11eTzhBEj2W3oINAjDbBdHEIzLHTWVSid4N7U1Y6/pFbmC+FcYXWt0UwzRfNObc2WGpY9
ZoVrRTV56N2Y7+ctqYpJiF8ve4n9Gl4ir57LE6Cl9BBvrC4pynhCi7w4Tgn0OPZHVbVZNNNPlj3x
gxamly0FjGUZKuovfV2hy2720QHUzniU2mFblZdUp5/OEASiE90r8peocjq/Z/Pc1wi1y/bf4KMH
UzIOU60PStfOrEi50seCW4aeOgJO6cyeUDhLyeWJkgODsGCGOHGlfcs8Ceql5hWwVYYS4iNuzdBA
6MsIIb/nP83uytYKHa19jtExzuHj0EZxRA7ROgD+tCHfchGxskWJNzzUKcb8C2o2bs+kVQ9wSM8H
qofJkd1CJDSe3vPMX4I2gBHB1OFKfmp2k6Eyu+bWJumLtWF2TFKfjV+2GynkXU5Cj6fpCHdPa8iL
Xmz0Dr1KTd3QX+xY6R4APnr7zbp//Hsi3MBEGntMwaO/UHvE/AbQBDFYD/ykLQFqk8FQs3/mh2ab
bwnB8wFyzlp721hw3QytA3USa41TvgzkPkmiUGFtbWi9EasD0cf8MyNqSx3bv/voXnL0IZwXASYt
nmZmZpS95vgoJeEcJ9WWf5T52oDcSOmXo1DubUhYPy4P2SA4zO56CTolwXYczWCZ1RFyBLH1IaBg
hTZl092dL58x9k8QffTK89coWHLL28xU7gsL6YyWkfxmQ7ezxmOKbGYDIDsUwg2WMQ75IRYfyEqw
b3NwpV0uATI1emYwr4x5lX/lWheqEyHxodKNqojpqCbCb/G7hmAEEJ1R4IqU4jiMGiP3tbyvEaPc
wgSNYi8gEGvFfkTWB+7Nh2TEBK86SNT3y/oLQ6pIjLcU19x7GfT1FPiH5e76tCK7qN4JijPaYThC
KbiFucio7sZr76JjtJjItKLhbUV85CqpCPjwaRHpzdxb1Ek723dGSX/c8yCdfLDaSe+5R4MTvPP/
NTeA0QQq7EOPUbrmFATqSmvRtxDOSgQhsc0Kp0gHJ7NzIQ9oFlExyFNtjh1xqtowHDaZwa0EHAcE
EBJ1Yze47+5e2iL6M0uvHKYtV+842xS2xbUyD7Mpj9zu/sorHO9Zk5Xr3xuQzQnk1fn5HZnGUKkE
mPlFnSDpmDWXD0Z9xzt0D6s2nXR3Il2PBuwQwD7Tm+2VX0VHTt6KlGts949JwEqRUqm21fj43Oag
XV+XRIBmUIG7iWU8/aWieKuXaTvFNjH1uhN9OglhDi8YIoU766ASC65s6shY/WJNgpFqdHz77Ebv
5LQfTptZV1LSgrPxclArJWYJD6D/SGx6IdHk/8/WtdBLrPYg7ma6ff8AyXO4CLL0BOwsUgAjwAxA
YPvdAHQOP6nakl/ymm3ZbSZ5YVfBdO9yu25Vo2lSuU1P9IxCtXLr+G9lRz7muAc1mkQF1DOaqXWR
CtaUvBBC0u3nu5Vm5U/iqnT4XxdLViy6W99QgYUs3i1Uczzq06zq7lOAKoAGWkWbczmhO3VXOz34
DCImhClxH1zIMsCYO8yNe4qN8GcIHnudycYxcF8PK0vhCUiXG+yP7dicpgsCOW8mG2ncWovBS/sm
XebP+YPbAXeLp3dAlWuiYKsuEvr4QMwqUNpP0a2PWc3T0HrgUO5WAlGDP2yd8osIRdxJkgBp8AfQ
bpKmbq/9lJzpHerZFXN2iS34lbIw0nKK8Ma4Ps95LNpdUQjc7iNmQ8cy+mlmVfB1ZU9kCaGZNRES
CMCOcpech7ac19FGrY++DRVJFe6qMwLC/3C7lgD1bsU1LJz7xybxOaZbG6591G8Ev9b3s4y6fP/c
2OkuMk56hmuU3UOQsqh1ufy/AOfxVi6J8lMJpuQQsIi4nWb7mHLL6kW/B9bOD6vZ5rEpKE7+Mvyk
vl+B2dFCQLFzEa68FTvczGZqx7zwWS3hp2LwrXFVlCOW0FnY5+HcScH+3aZ7XVXiA1BOy8/0k5Ch
dFgBEmcL7zTR/6Pdx8v1fgx1DZRo0B6uumzwPm1y5Xoi0sUajeXD4urEAAanOegQHWCcFgNSbEmu
36RUbouTiCFQHRGfCXFTYwr3CQJbKMXzjWcWOXSeVwBTYar+YfwHEfqKeQo1nmm1yBU3qDTnxEe8
MWPf2Sa+JHu+sPbDgXrrr6cw6294weYeamurCu7z7OmpxcdKypr19pLzUfJrrIQ6Q2G7u7X13LFf
SiZYJ5J1+rkJCVUtTFyTYKslsxH9VRRikMIv0rqEjx17rLZ7n246roHcZMkRr6riVBf/yVezQe+A
W6e5zdyOZA4ALCaUUlqvz3xqyB3XPOMXi/fArJ3YFOLe21hFxvrU26p9U5rUJsw5z6/ZIJUNtbbT
2a7Z7URPiwiMcveoyCy/Rt4r1Qw3cRaEn4rXlnqk0wxtKXbuYRpX8b7qhNZrYNw7mGSiShA1ko3/
9q8zQXCXXKWNH2dJGtniZCdYTiG/Ttoo72kNKjScUVgmhdq3v5INlh1tVD9Mm+A6s9DqOcGQlteY
X1D/bHxDpxQKHwk8u8oox8AkGRjstuWQLslmo0iH81Kcb6rrFA4a4yXXm0wFK3ELID8y4Yi3R6b1
g3LbfHP2x2cZLDLj9N5yihCXNFpmebGIG/qE8joaDksvzot8BtZdbs0YTqQPc5/iuA1Nn69/JuAq
F3TuQmPZTY/ntsHfWvwxLCEA2DTf84yABNHQNwgInUEmYrcqe1GfwuTXRoqefP7xcN/josikE9E8
FelLIiAjCjBjK9aDwlJL0yN6cCSOCW/VGLTbvjGfY1ZrZoqtU9khen5MQaDjo0nObjNc/HkR4ITQ
AEf19LsDwKVusTtFoE93nubGIIQzfqtye779r6ueCjUpksrtUEHzBkoGT2LjouKzuSPanS56kJ11
rjVlA2r6X/6lvUaRGeXty7r6wlQUk1/NV4nSfmFisYGKdhxDBtGqtYEGuoyLKcYktPsJ4qh/zJjC
15qcWbwE8eJac8X+uQJNKre5WE48nVuUTe9SkMi8M3vTLZAP/0fiHNZtJj/JToHmWPfZszOaipRH
5y+CTCiNBCL4hjqy39E9D9dt0zQ0vz39rcfsa3QMdmTnlX3PFz9GNhzrKDAD6ldVjaI/U1xW72zf
s56zOw+eyBWFdiI9Uj6Pp4Dz9xXL4odHQZ/rKU9h5X4Sp9kBxqTZJs9a6+HeqblUPieSzSCWeZq1
qy86nW6nR8HlCehU/Q9FtBKG4XV/zF6d90/tt8goTYNPzhpZ0cUPKGT9taMwvH6PxrXhfYmO+ldm
Pmqr5sApnmYsIvZMRBfwQavK4gxPmx0CGfog5chGwAL22lNKvG5mc8Ef0YnvBWN6iT4VuzOqR8Wj
pElzeNPtoQ7SRpP+qPc0qdIv9xV1BOblkXtK+fl5G+k/azBgxnLiD1SpgDGf0jdF26cv2pB6ZWtx
X+4l1wWuw1YByZD9FBS4qiR2y7wKeqWMNNivdAtHO489/gY/6CTIkvNgxtzYoEqjDtjFW4dO1STo
xOK+BHm+JRijPR38iV/Q4oWOV/HT3dd+OFgB1U0WwEV1lySxS9IsZMwawZ491DQk2ndQb5ywRGkQ
pHqD4/c4J70lbLc8qRqJ/tckXdqT3LqnS46IwQWIJyvn0pETmYUH4U0FhksaSvS33o90AOR0HDHy
Kn8CvVVqhpghOsJYdkuv8/DVXj2QVn2zIxnjdzc5I9N3pkvCE6URc/yB7KiMJOqwi0TVvMxYxA4K
Wj6TJJyNCVFG/yQaXrmo6Xe8eZA4jcZrk89QNSWJas/OQKKYwQYGSfKjKoooJ6DeIXbDqR8al8Le
UcUr4Cv4tT2aFY/gKvksYeAIhXImdONsvde4mA5om5/vOA7/4gKafKpjsbdjA26fT9RQqfEHl4uP
eeFUs9Czme5XjHjnNtgnka5puJ2YQB3jk9gXehnAJrnHUr0DsaMNiaC6o0/uRLYAXKpxv+7Gb8eo
FYaYNZruuAVJSBnmyrgrUni/ASfxdkZJe1JVckgkpVMm+mVsclktx8PjxnqhwhEZ5UZ0DlGg52g3
hEwl2tpZKYlMjGZDPNluAG5+vHO4vu6JUR03TdcQ5ACiajaZjiBPkwFb8br/QJO1AkS9W/HIm7qW
2PmVFB/48nNGzDwsixjI1WacsP4tZrGjjbKyuHfU/nSN1Ir0msvUrYGhvfJVq8YjtFgDPdrxOpQl
tjtml0/r+Y4Jk8QFjjvphF/3LbHzQSj1nVN5zOhAUReZRUJ3BrfA8VaaE0+0riSqeonDs6uoVBYI
c/tbrzJVbBcj8KmOh7xcAMGBIvS9i2bFo1t5n+vfiNUFVEY3WSZ5lJ/h3ltyapqeLNY7/wBeWtSh
9O28XVz+RSCyAYce/bpL1CxVplUiAdWM5TazEQQqfb7O1tKhOBBF+KYdZSPqb2LxuW1Q2zt8Hvmc
feW2BAY7IGHSmN2NRpZc/MChPm5V1OTJHQW1xYxQQQSSA2zueQtK3WqO2J21QCLlqvGYeBUgsTFC
/XQ0c5/Kc3gBV5lMbEtuwdf8x77Nffsr9tHrH7R1xI7/nvrfPABYcqqwTPceIIpKKGMWW3mM/Fvs
U1mcp1gEAK5h41nQbcTLPyL/mlxn5Bm5VPJxEi1pGjI5tSUR/b3+3qdgQShhJnin84/735lmqzaT
SBRSo6g4FiiOn8eFDeTe+Hvi9oIcQGBgOsiVpdeWoSqQe2y+sVFwOjKVtPa9R7fzwvXjnk2Sx0+6
PzbsSl3hGoWEnSPRyhBN5jO4gt29L4xlT23HOgai6v1HOh/VT3MsNPfAtl16euH4MXEE4h9yI0wN
XBfdDdsALW7f2z3/yHQ6IJ0tq1AVfe/arXAJJ4KBR2Y2mMdUn4KBZBQujbQmpi1xJB3jZjvCTheS
v6OIdeLokdnuHx3GXKLfhNr2F8IYsXeFMM/E3hmIU34VgRpOhCV5bsXjPRxamXgrU1SKoEd8Cfs6
rFP/h/1sAJYv4B288XhXQmNE+QVpsPChu7mxJMGCMGk0sbtu8NDEtpQIhHoPDGOUkpzNBeXy51il
ODxnmCGlPZdo2eNnLpKl98hgS6zsXhdPV3UA6gL0ubLQxjm1uszeLADPJ52+lN8arp/Mb7KERqnF
2ZJ+FR2i7b7lmkPuorhhvqZ0HyhRfbYi5k3ZVC5PdwBb+r/klNlwWmEm+Zq7BEWg9hMh40I9zggK
zwUwyzd7ZBLxcDJxVWWMstfUwUYFWMAE1fkCqbp32P73OPx4qLPMg3qrxeBkYBEwM5ysf+OL8fcn
WX54aq555RDUjoujzC8uwrVOZHS0GhwIME02kPZUUASmS3+L2ZciBKMiTGrx4HNRR3Bx5OdMPYYh
vQSP0k4Vcmgyu/bIuDKYwkjhNVRWbiRxgWt8aGwa8M11ayOvd2CoevQA6Ufvkp4IRNV4kSI/bmcN
AVu0y1HCngXHUsOw12X9T8hh0xre8d+mWHGy03xHO8tLTeQmurSjnD+n3SOwYvgoBXAJZKzoyxgC
r/uCHWvz7jAxEgYzTLev0tsmB5RE/HkWVyb7p4RmMw3ldvZku3Ki1OF0q+8YWYN3g+X6aFAW/ntp
FmTBNiDwEWgLuR/vR22XYS20ruU4akhsxDbV6S61X8UysOfgb+Nj8EBNlnR6k6Yy9nKVcGPI+XlE
Np01uG5MzeUGJ38fdRTTLYo4l9+W4/2EDRpwexGYIPpglVHm7/cwKINpM/ZMSZfcC5ASxVz6YKD9
QabjHXWJb868bALuUE5r82Y+W2LHDadokzCG7qazgu3owwa6qZ5ve1BwpumLYIzdhaN/p/2YFkXA
+bv+w0VcaYjwJF5CSx/oVd7DexEiGLpuNHQpCzqYAyv4wKWWRATXXnyY32D653lB/y2J9QubeI3+
eXA1jsOFk9PjKFmUo7Ie9Wn5YovHWFgpv4YOD6/YcgCs06TKMl7sVSUirljF53W0qk4R+cASEH26
oG8r+eYny2bFG4fl7SwumSMdlFppLsk7oDKyDkNnBrJ/ZOgw3ikULOQhLFOPyrYI2u7N6o3fm0Pg
jq5SipBjM/OpCz77ILFgvsL9r3gBk1SuJyVRisqCLtHKjyWdz6JsdptDigtJoeErbcckwEmgK+Lx
qPTJF07LYWuZdFQQVJzBNfVovwIBpH16PEVY6KuJBytq+gCDMVP9+2R/dzjneJ8WJylkD3AonOlw
883mxpG2oFUsmv1TkP4DQInlX2/fE6Edq/TpUUvhmJI5KQLSIGSVa6ERjsNRMQ4RoVek/AKxHXBK
YE4MaL4J/TpZBDrNH82mXVyO3vj2VSE1q0H1bevD2Lpjd58HmK89a0khtlXwJzbSJqeoXD9MrhgI
L5mwbhugSAbvAvV4eivvFrwuFk/DVVOUkbuaM3bKZHAZGIkGA2GUHXMK/kngam+lkvcVia+K9enA
IHpV/nIv0pXDnPbHc2pj3b82fltGAADPpT6+HmPUm0UF8TOdBCF8+kQsEPsvg1DgKgVt2mfcf3ym
fiGb+Kyyr69zNHoKlBtTZwk1bqlCU7Xg6JAs6cFPhu0hd6TSD2IDDrZl/uVdw4bK5sPLV+4gEUjp
b//bsJ6ccwgWCfG6YAQ/7j5M6MIvR3gzueOHhoQPe11Xci49R0Wjvramb8sIkPn2U0kwBa87m3nP
wylBY9wdWaC47vENpYulqFFYsYa26bEsBqPp+oGFaCXGN7s5dSd0sqCgSSsM5r6wibuNuh3mW/iP
nTVOwmwO62ISX6h/u0QrM8LW9dc/jvnCRN4xMeohPKIN1QX3hb/ICNYIVSF7i6VJaSLoz2qd/Vjx
eGoMSX5lVYBAdTyO8K3ewJvQ0yLVH3qhyqH4n882fA+o80caQeL0fHL4P3afx4JL9fBxDsf9fuDh
vBLc1pmsp0h6h+2MnEfBKmVaasqbWHb//yC2nWgUA2wkauOSJyCCzZRP7we5JLVBvSan3iR9Iv9i
lBah1B3XhGH02gj/fGOjTN/jb5zSf6/TLUeC5wHIh0K9xqjNOlgUBi475To8iEsMqC7IWpoCFAdC
Mvqv+Fk/lNDbVZ171nS1p68aqH7k3laLTzkkRm1xbqJSP0wio4d1iL9my8ch87FUTd7fARHggB6E
EhkxQ/a4t5cGDXYygLCFEeJJJkImoj5dp3xo3T/xD8j+nGDZ+/Wlh3eOFCZxtVO6pSjuYtJnzx3s
AyPI1vwlw/oiGq++VhAC3CsdEldSbTpSeLYHs4C1O8ZqBACGHKPP+wbry9LLF+rc/Wzbr0ISYyaC
+gpNXC1v2TLxN3e3/QpkpcfzJ51ArOcO6zhGl3FFBaJNEQCp/vWUyKzNkDXlg0jxpLxxiiHsCNlR
rEYH2aVxK5py0RsaxHBAHxU0YddPlalrf5qnJE1leLuPCadEUphEah5FOw3Q2ZX+17qa+y0901C8
R4iVCBWqnHjqfVZdcKfVY55CvYCZGxA9FPyb9VqiGiPVoy0WPF1zn2o4heZvuY0tXKpMndzgx0F3
JmvdFHpSBEwvZ5b39JklrrzpwSGFBMuiLgRY0rFR6PBMnWCUkBk0KhgCXT/3MYR4rPoA8V5uXqop
iyOWJBpwHsNsZJgP1v7gcSNMO+7EIX+IMgZyVr0t4DvCG6nhrqW1S5wywuq2fJaewVl3HlaVTvzN
P/ALEoLwN6BZV/8BtgGA6WmCic2rw4hlsAZ7NH6+wr09QgzO1hdzBuRUzeSc9uD1ZIOLhcsZCx/w
o0i/IhA9QuBv98ntZHlsNJDh06bqP+pdfNNFkYK8b1UzH1fMKQ6zTAdt4h5fBwnFEUxTTvXrNEgA
MepaLC9/W0flIVWNC/oiUHUYKQm64vYiecP0plDH10POM5FQnjuotWS2VBJ2lEVCTAiQeOuoH/4w
Z+tCWqj5ALhMKYVb+BrMEm0Hwbld/4gdWaISBe3qiXcs7njZ8cgxqJC0A2KNIIPHgzYAdbsDPkbq
oni7xY7TH23f6WRGG1KSxURnDeauK88g/QaYw3R/3HGeDF1v678QudAnd+xLDJxBjW8U3xsR/H36
Oh6MoEl7Ao9xPhdwWfwLrJ1b17Xn6NRH+7XT/hSU6rcMKoK60MlJEakwNKRHJHUDCx6sAhG7Lk/q
YzhKpZcbg9joWY+/2sMkkLbmXXyl97GLCbpxwBevrrQnw2c1rIS3OPhoz5iYYpF8FT4XbupLf4vj
2Ew8GZ0sC8x0eLOFvkZN2k78qoMhudrcEcPldC97G+4hyl+0Y1jL9fgmrvoKqIS8D1dCnUwEIcEW
/IRUhe0UWzQk25HJJ+RCpBjetpqlSqB0+p6/Hi6160pUthqovQ/1VjcyxQbbG4kp4KsxkGtfgJQU
Q2h232I2VNxTQGa9BEBB9IbJNGoZeDPq/SCrHJVZO8Bgv7FIAmUNrT5w0NUBvYPQ1S1zunUfUcpP
s8Up9VY+xLFUflgwAF8+G/Il1aIi1RNocYMz3hwwn0CmljHg3hnTsAU0u8cUGcfWJ2qtqVqZ3t2d
W8kpdb1kjNX32CyRFeGvgNGv3iDXQpJejse/6bxXe+6GhDuF9spROTGKpKzJHAWlpUxg8WOaU6xe
tRCqRb0iF7sTdmPJY+/p4Y1pVnQuAi6yz8MsOHMKzRe34eoj8TZ4TqzsWr+3SVpFU31pCNIlcx5z
z5dgvZILZe1+DF8+OXQo2zoXTJY1YATHaeF8bXjFwHVyoM/4ev8pOtaAYxit4u2cI9aCCoFL3o4G
JAptAFZ9gzGCOWUDSUa0AmLBru/fQjNxdWoLqlfU7115i0KER7pcHfnhwc9pfABEX1RSib+UAOVI
Ue033d7GJHrPfglZ8qqCI3s5FUH3yeGijcYLTNjLYQFMkqoQrO4PVnUGD1PHhaFc/gJOxxJR69T+
XK57H11bROaP1xL7eQVUD2sQzmk8i1dX2jKl0B9KCnebZkGB+ZUTrOc00A0wx1Vjr8/z9D0SlBv5
mXiU5Ts4ZICy8+3dc7koe4skvD9DrJ/vI84v1fDZudwradFxgAlg6PXNvwysedv1qiBTdnXNXJ5Y
Z+xLYS4XK7vZW7RcXEjiXaC202+63TL2v0K2w/IUccUSKYrxManzeorhhzhzW09RPtiJt9uQQTqW
LIt8+kPIYKXV//NFUaVUdJqYnYTX8scCzA59/JnMWb1WGWSKsbtUTrfh4yQTPMOwyAwfp120tv7D
sASz60p5ui4KPvwlWa/TM+gj8MZwpk31RxuStoBRu8hQBoRaXnhXSbFKHRHoQtHjJ486d3CdBzag
SoxXVkmyrTMo/vO7lVcEPfzgVtWLolRp3rTvqNZlwhHb8jsmI7+wapgpVSrj14G1/AavqSXzJEcr
7dmNxOu2dk12AOtFJISoQsxP6IKaF1lEvip4VtwRU4wELTVk0y7OdEE7bltCFhXMic7j0gz4BC5I
lZL1w1UHTlyJ7ixayD1Xp+VqT7i2fF01FNoojaWEt3deV/W0Ix1sY383tilXvXreGx9xEKZlYtKE
YMfxrYpDbEdQ4dvZCsUk/dGIaw+m+ejIdmpFPkziw34tF1GbRA3ND6sT7I48cYLwtRHjk5q72FEo
g4/Pz+wAgqIfOClB4OvJm31GxnlUREmwk18OlDvT6l/Tts5mSnSvM/Eezx/OPLBnJOhf0Z5Yr5iq
kHfl9lnqm9HjND5vfeGTl9kFe2nd6HAU6pQvODxtBYFYoBio+nYB5wHTplgPnoAt32f78wJXAHNT
o5orJH4A9C3OyXLk2PGsMgeyvXP8B1YY7WgbhsCHPdsb20Qiz4V2u62RnHrVdQXR282F+Q0XT2AB
VA3eJO+eT/3WPV9O8ha1i6WtSRicQfXUsacudFi55QThqntkWIeoLYZ1w5D7T3hqATODAIn9tzDy
IMXyqSi1kMsLl8yc0sNZJDIbUYUDiySUv6VOSdY+tgT56JycK8U3woN7DP4Fayljshx7VDadsD1W
maGkdzqEqvTA/sNdys937V4CaNBoOAELFpfbZbe0r9gKd5I+3ZN6mx9YujuRiios4iu34P/XmL2r
x+eAtVDNlc7V3K7UR1GiCNfaNqAspzl1VlXwMPF7KSFirLYp+HuW2cBEhv6aE77zc97nIEcHOQgc
htnU7qmwSJC0tU+z4gHR0B9vJuT250YvFADI2ZIhhL/NYn5TnT4/uTzL+CttE1dCIn8VRkZ6evuF
/NRsC22Jqg+8yBrRQ32SO1TYE6PN0ZweHjBPVXD2hErmV5pjtCK0hZBhJv2zIDn+Wpy9tyQQWrQu
5oKRmdaRfQCGktpvHC1OiuHRjyj4BithLSKxVdI3XAjMwpQKG70HqRJ8OpvURlkICaDap7Y6vfpG
wS9cPfq2UQ0POHkTs5EIcvdFRw0/EStF6aiN9P3jpOBvkoeT1OpgulNxDHW8AwbsrCCMy4N92GBq
kBZPawqMC31VFQuXyUSWc8Ck0TeygsHNd2Q0BG+w27b5cSkrCvLtjgZIoUE3oc75gem03Yts8CzI
STZf6nDjXCVBm01w0uJkOwllRhW45gj4DWrNk5DqSlogB++ddjKaB1/3uBTk93QwsTad0rpZG0aN
/jv0pvxcXvcibc0sXuj3QsowPQwVnkhnZZ0rTLVhe1ImIuicw8/zRqZ0R882dD6e03kfkbL416X5
bwJ22N1CC+xTHrkz3lP8nbNZvY3Tqn5Eqql4HeTHArSeIi0A4844BOdUCy7KTDGqQtCL1x/OXBgs
cfJ+2g6VlhbTISoArbXYbDQoPdNj7zdFEQMPx2xO2gWmNBlDvh8io9wEWpbF4PlEudjxoTJtfJw5
X3EUusg8wa3gwTse/9E8wZXaQ9tEFjC9XpslLD43o1iDWM9+BWcia/vQsUgpSTPyJpv/R30i9Vtd
lAnMOc+l54pQB1jIpQuaeVs99h77hgpfDHzJNYXvcmQGlhaKW1voo8U4eg0gvSXxgRtkJB16ykY1
8zYJHOXdUlcpN5Xe19zFgl4Fd9d/nTdOsPeQFY4Xo3U9zHicuxYav7Dh8SNhoc6mkpHpzfZDlqnC
UssbS4w/Yjb3mxP2tkQjayQ0rdmU6h8fJOvj5vCz1ac9fCV7POvnbUpbOu8Q+Bz8TAcIvG+31nJj
v/fyGw3lE7YitIdv9yne1J6pV4G18dmZoI0t82D1LHpaWZb9AOx58Isl/e74tH/JHLeX5D/hMC9Z
1YfLwvYO9c+CdRMxplVwQMe4yeioJuK8zGZag5J2VmX7oWiKsJTchnXqBRhDtXy6HsiOSIfDepg3
CEaKIDthOj25Sm9f8R75NlbcxTdLAkryoFj5n9TjATlA6UX5HEdbzZq6OcMpsFBkFsqaLpeMbHzl
NbGtl7SKoqxdrpOwzFa08P9Hj9Zck2kyqsAjWT5dcDoJIx02tdx0n/PyCiWkQLce9DuZqQJ6HK44
b9/BLRfPXgQ7I5NKzvqiX671LbVjtOu++wX4lFYnx4aJzYl9mrlZ+xcNKfSfnooF4oHZAe/Nj2DZ
+ROYDfpNH6vxphW9J6iV4OZFt2EKx484mBlzZQSoSIStGnqFjOKVXfU939WdUjG6aUM+rayoEqto
p7jshYvL5bya/QgMTIUGg4EYFoZRqOrtChKJKFF0v+ssntkQxEhn5i9m38jtzUeYqxtM6XugtfcZ
nNA9IOQPKB/K0z5S6UGAC6v/l/bUQKj8JYq8OjVcYROLzgFyS65loQDEPayJQldvgOttpZMhRVn9
cXRb94uzi7ykjk5rfemiX4Y1r/9LRxaoe3b4kLiXXgrNh1f6K8LddcQjYBz0es61tcWXH6B/RZ/i
YGifYdHJqVsOdbCuB7/R9/pWBf0C9cTa/Qqc2LgKzVEs9VETNMPZfm5A7EVNuLPXpKY6qWBqS5El
1utSAZQxTYssS5ZVQvB7eHhDt5dHB5mZkiNCVBl8Ke17y/enVKs+O1ZLy7js6p4ItKNgcTc5FRyW
mCtgmIFmrKo8YiNTD2MrkPSfXadoMSOTTcn/m79tw0eHMCKpsl6x2ISMfTcL2ACpLCIhjk+9YV6o
amYEyQ5itSEkdXDYERZSOBw1yQt01KjIhrliyfkxABhzHNNzpxZr/1gyswKqpnisRGTl9eNw2sl2
3pkAmuyDJisjW4l3cVsI+Ee/9Ia0yzItCQ5PTWeUT7MY4faB3YdTTmNTZTS6E37spb+guKgOzZoY
zYvN26ftBEelGvi/Kc8rcmzWZlSqK3Xr9wNTJ8b72swQB7sU/y7uXD4vXyXVR5v9A7MH1rCU1dGI
F4MusZfUcgMvfVL6+H42NhHLtr/NJPmlMuLrTASJTkFtcYwbbnx9ZMMYlNg/uU6wceIdGbjmjYui
BSnmxbUEV3zuOL/XTYpyxZxAtp6cbdeoQeUPkz3VS1ITEjwiz52kfAvLJJzkEMIAId5O4Ut5q6c0
075zh5g8zp0q30OdTpKThO6/zRho5Jy/3o84tV2lgdTINFyP9oZi48V+VbI7yKKKO8XJA+MldrUL
BPZCNdhb5EW6BMFFhUJf4KY20DcZ2zC48R8M5GLil/kMnWRLrd85g4NFHtIpfkdPaVDvx30tK1oF
tiMWX+Z6QTtg+SuI2DlJsAd8jXxKXjkicTG2sdyvs1xje3B/FrKIPDa5vhUqKoZt+PGG78fmetUm
XuIw4XZ3qzA+g0sRj4EWM92QGZCny8guYVNkeC7+YdmSOWMnP5T1xyk8HevsFHkVUqmGMCz+kBxm
BiugSgYar85h4pE+QsSLziQkC27bPyPhwG1zLyPQEqAX0yTGP2L1OmufaZBHVnFYK8QXAJdYWbxD
5bEgWewd0lizqBi01idcBgsCjBfAQrsNUcw0IwJD/R9R4R7Aft0oclcxt5C5Q6pnKZFUL4f4q8oo
hpIROrkL6453U4ik2LUZtpMA6CYAgR386yNOKVjUcla4W+/iYAehfnrxk2LOu/ulABOU/Dp7EPX9
Znq3GAnrPYkH4scX6hHERbFTxgJjrU5vQ5iNBWwESdS+307yExfhUmDpBX1BcIqSV59CU5ktEh/m
vbBzBXR5QdNp6u0I6SlWZl0qI3J+k/oSXm6VDUq4/w0gyTwSkNI+eWjaRfNgf4avRfJP6lAFY/LO
/q1mjLPop8qQK24zkNpUsoa1Ds20FsDqbr7YoDPKix475Yv3cU2i4JxlKNyiZnmad8kOPxdwsuX6
nnmXCDfdMSwHMl2XFhej0E2yqPai63qEvV1henmVaz9/RHlbxXb14+paqQiQf6u20CULEnRHYe3D
G+Ckc/oGpm0lT1a1NOIhIlFFZM+ky1BpnueJiPlVhPO4ziqo/0nQ2ip7A/X4TmLqBo7XN+TErrxD
tZ3P52hnrbwIcoPIYXD6R1dSRXv7Jatal9lFsrCfVZ6/YszDHN4Eu+bxDaxI4IoWStoN2TqBIMuR
K+s9KNbNOxkoi3BPTJHHOPmCEDIYu0JlwkNVG3pWNi35+6JP9y7MSepoKvrpTtTWrMKl0RosICjA
XXCBd1fsN21hVitoBx74W3HbkdFsEgO7xwaT2hwF1zfBB2IgPnPU4fKCQO5jX7CXJ407bKTmuCAw
A6Sbenrx/+1sI4EM2EoihTLhtZcQ443GGjKZer2myexr0bsTWykiiPJfo2S3uoDJa/v1cN7a5oVE
mp+9i7ilZUeL5PhAFkisxLZOC0TpzOwpUT/BpeFqvFvumktn6GzfQjjrdQ28Yi4uD+x4IhKf2Pfk
UyT15rttCel6xJJ0NhH46FZK4YApz6J5N6dJgEOjlUwrWPMWfFAotwCf5Ui5GrRkCjGce60Wc4b/
lYNpnSsVzuqe4oaVBT14DZ8wcvD/RjmgqgyHW4BMMSx17FK+mI3VCT6mKq0t65EfLcZTjENa0GQa
7xtKjmFtIBSShT5vSMzyakczE8rE3Z16VP569PifZCeKJwuaQGraHWrO+Au3OGsZfJxhIRRu9uxa
RSFaQDZOav9bBr6z7dEcp1InpccXk9zVxu8TON9Ycs25tHZqHGtyGBKFlm5DSbvPt1KPpguqVPKj
3JZc5BJuDMu/S6gwdXGYDuGkk527bk8NPoXJ8zzFMiYixlDYl0u3Mh1YOTOKF4Ez7SGeoMo/mvXt
dXVr25hwNFX+VFRGXKlOn3EQi/R2aecYNnna4NORNGEFtD+KFxiFNw3ZjWvBmxX4aovuuSlsW7LR
r9PasqoJSO6J5Ogczmpe6zoviDexTSHJBMdonujQgkilyVDQ/QX8iTGAFadc9W7vOKtR8NtmVp1C
gjxGzEK7kC/IMp/w5XcfdYjXqoFV3mLRf0blZ3ZDC4qVA8Jhl2WZ6Khv/9aWtD25xXKd8/3WaJxj
erwuWq5fLLvKXSDjocHft4QI+ui77t0G0oTwQkOOBngWVNV/jObNkO3Dc5snr06Bdip05NcnGz/w
/UxiGAJAjC3APcknXnocVF04oysuqIWJCr//59j+rcvjYeb1hhYm6azsnprJLnRgjzVS2yD8tppQ
EACkFhxaVQzyw5FAxIhV9qVGhCcDr2SeUXd0pxSvyI9CLnctAdC4O2A66W80xtfZwuhR39WuywXn
0DFsGJ6v73zzkmK0wjJPNkGLT8zTgeeD9jI23sfGXK4mP7EfPENGuU+QnGNlbaRJDJWR9Syq93U/
3Sq4BFIVQZ4hx7IuTxO4B2I10tSeywOR5FECKCXXOXHRD67d0LLq+YpHDFq5Wxf9mLSPki5xuV/I
WPIf04qm90SW8oXa6Q56Mbq0/e6ptKzYMPM4SpqxPC5wSBOQnrljv3XVc8osYik8DgB1dp3AcS13
AsgeIdl1SWcmrP/XOKvuKpvvbHyEJ3dWrxkbK5Z9tp6v7NTAEgpfpHpnP7O2i3DFMXQAuY+6RasA
WT0T802+sd7rbG+mgchOkK5mTWQQOqr5chz2t6hrLDMHziH/1zptZXqyAbl0NukbaxB/FCCjybtD
lYGGhj3UMANVjaPflpBxXwOfK+dNJbM55cX6TGUl/Q4ziEdJirLYzDSPoWBOU7jBL71qx5ZJ2t8B
1fpMa8vL4AvsxGC8TSxkU0B4QC7oM0ACiPgqFwM0/5ywb+uavCziKl/1i/K5gq6W60JwabKpEXsr
YNgs9F9AwtSKnnbs1P7/xgcXU0WZUpPzroQJFKAhwBlLj11gcoFKcx3VqQ0n59kB2HRRUFDcRPQx
0YuZuoSrSpePcJU7DzQ8LJsTAd8zuaJ6udknsf2tj6VoATTsF6pX9zea2KZ1NbkzfcqMRJmHU/DS
OxFn8U+TIE7yZPy1H8S6LHmf/DDZDwU63uev1ON7RCJ+MVDj+a47FI9M6j67ziBO4WTd7EeZL+Mv
Ew6eslOC5KkG2lmPF2SZs3YP0mJWUrQESmr5auhpDaZbLlYNYUWlaj/ppxq9t2DXA9I7a7Si/4cl
XcRidENsG3GiY7T65ZY3lLoCLxYKsK+RIlcu+sR3sKqfip3XmfgzcxnyoF3oXvEzRn/n5ixF9Ica
ojUTRSRcC/qA5oYAERT2EpLmvJLFfhoIpZGce88NQ/SVOCjQC3Fx77ulWQODvH7/r5pPTWxWB6fm
EliytOhHytIa7EtmFLrD6clWP6pClKk8q5/jO45g//yCEcSXVWKffRWUU4xsPiUiK0dmNnpQ4gTX
4X8lJCI4ocWAf5o/RxXa5MNETxETVz0izn/cGaf2Za+wtH8VWFHt0Hh2XDvsHQVeUg2BeDKXXFJ8
dazk7p59pDV+dCImhgePFaIklU9Rk27R4ID6hie0e2qY7sPCy2vn+OUuocH9z7pcHcDOGp26xgbc
0jKFD2DxxAKGBBUyxRIjVC7bWfdgDsSLa7XiSnTQiCYTCA3yywnn9Y3KP7lRiwVEQO836kRHu9nq
hy+aNPDPW4CsPsB2ErM7KhSJTQxOEVAP0gq/osw58wwr5lpY5zsRgC+Bq2SXwid5n5GHd30P7+Av
srFQ870DvX41llMZygKNH4wXzq31d7tWFUcct+Pqu61cggz4a3YxoH7dlOeAnlel3d/gQhlUVJas
fVTwx6IOeMSwOTyY7UrdV+FySr7UqqEh/qwVKg0P3LhDXVVuaVhYqc2QArt6VztnhOF4lx24HRZt
GmmjyXb+XPhvtiq4RmdhMuY536BDfCiAQBpYRYB1VMYaTo35ZNwfHo+Agkqqb6Y11PXEBfCRPKjb
pEXRxctG6KABE3SobR5OpewUIzGLWFEqQbUNTOTxf6ZiTWz3/fafi1JjQkOGAWJb9bmy1MI1WKsl
l/stOBfjeNgAg7u8aU9CLbSxGpZ9H4jrq2v/MTFyx3ETUuq5R14xXcmS5tF5BV8ZAdlw2+voLIva
yefGhntvaMR6qc/wZ+vuRrHhrLZvczTwB2RTbt21nx6AGTuAvs5F+iPzG+tlnDBCYK1zUMe5CwgG
n8VdDZoafRG0XSgYiVsHKDbsVstkNCtxklBR7YO5ekxGCTEu0B19Nv5lNRIjpetltJ3MWhMXx0fi
9sXuXV2LUiirSECtvHlNtayQFIgIabIMx/yFaGY6ycTQJ7hNnVFJXt/59uCRoIwV5pGnkvXwStFo
zXlZ+Q1sdAZEx/gL8TEoDaFM7q9jz4l0fzMezD2LRx7G+dSGxUjUngPLAOzxp1/XqANnV6lkEX9d
yq6LvVzPKUeZtMbhevO6QZE7FvJk/BOW7cbRGJ8iFH0YpA676BSxSO4YlU1c+mywlyCe37yPmSTw
q0pTgI231UzClQznn/USvdyViVUC3DbtOUCltX9Tuv8r46Phm2Cdio5U6u54WJOE6WkynahiPXXh
6vcLLwS2s7FLMKQ06LZC363R0KixmEwkF0YykiwqPYtiC3fCjGmtl8aia2VSwQWqO7JWKnjLHsN0
n/NJ4QWlU/xW49cW7hFxAVVIfijbaRHlsnDdIV8hOPC3PSLjR3PXny9G3eKHDmEN25crOpBzL4Ut
EbTS1878lLpBF8c7BEZw104DsL5NWKYfqCxbRfW6x6RkeXbfJrJGX7AvHq+HvVQpoWKKjqrLGpEz
gYsykH3/HLxcm6RilKqnAy2Fz5S3b0mCY+DOZkUIs762QfPVMTy+jGzTpd2+P1nfyVW4qZP0jUhQ
l5BQ1fJtWXJboeHDgFFyo1vAZVOoWJMNK0TI3zHo611T4wRO8k2M1jNt9dLki3mIfNqegWd54ZG7
bnFysEOdTXd7ksz9akL2VMtIn/+OAAK08qnybXeoarMWBT8VK6rVcimAsm8IXHQy0l9vZN1UeiQD
gpGEx+pHShsawIaQAW9t3Kf1S85GmLurhjFe3+BDOTnJuMoj1QFoH3xJg9GLH+vAwAXcEsAF6oxh
gxVezYLPe+LUichwpByWyYdpgaudDlgVhnYNoZ7XujEMxs3MzARbh1kH62HbXO1Yv6fVmXKFe5FV
JIA2Oa4cSSBtIUTqfG8WIFFacqlMAymZh7i+C0jXRec/svEM9Sc2oKWS/VqnN90KLy/0a7NCTudO
qTkWmoabEqmwbXMkt60TygOwAQ7BYt5PUjchfH8x5JPBKldNKV556WuOZHGLB28+HQpsM3r8JVoF
CCcTeDGrwMhqcdXN2dZeUqssNqw6KD6VNBTEMAV6qeJ/4gpj4T3h6aUqemEkbkYsU/rzOmXvjS4U
wMY064EEhuSAMjVwV24TdQ/MCZwjsT8PbUXbFPMhPJRUS1qjYQaEIOhFrNSUmYDpU7UDdZRxotW5
7Pno5drhR6ttMiL01IS954srnLx7V6dL02uV5gTtufrWwSFBzm/k3u51SeIkjdyAI1rTtyT1nmNn
eKCK8kcC1YON+7wLUgtrQLKkavYcXq3YLOoI9jZMQ7yOSa91JGQ3gtEyrUgmC+/7UN4PEbw2i768
yhBw3FpDqkhfLKuwNgO8VOrHwkSLL0laD3tzrUcSoXueAtMlPEFDTyMClShQdYUUdVFjxATO5F6g
d/B88d/bnUj/HSlT1UnbqWwKILvxE1pu+MlvwP8uHgGYVP3sy6t0DGDWOkyexguVReqbDx47Ycy0
AqAPs93gHQ9JJaw4pqvqK9b7bN70LIMSoUD3D1tW1euWPGhT6InG3IossDkZ9tny7fbXuG5HbU0Z
K/RmLgImUlMrOsFZ11lNzuHBlAz6NILWHuJYeRa9kf7ot9lOXwhENmzZF//COQhJD608ZkPBeZ2i
amStuJqgMjm4gY3PKLgHQ4zP0e+6gVOGMQujYOt3ByILfR4Fzr8/O9AkzFAdoAkA+w3FEZIDQatC
vg5Rbx8mob57afi+nbS/5gtOsCtHGxO8Oy6FtYrmi1SIImCHvfhOAxanS8VSSNxqoiAHnFM1rYlf
MCHlmK+LvsAcIyxHU9moT1MqDjzGJFTAVgo9NX0aCVoYs9ac2kJsVFil7hvT97QIzZUMtsp4cW+r
z1lWQd8inPGh0h2VYfJRmX3VFxHOdeTtP1FxtUTRx0dLzZLenyukdtdXD7eJ9/SSxwLKfU6YNn63
H1wUGJEyA5HDXkrVqB4jZKYUV6/yZcLQCbzX+04uj7M4/dgCsENL3Co8Ons0b+SjUGIbMGtnImx8
oLQwmT/12n40m+t+GUalNlJogZ9QqGAOl4BG9+CPVU48Dmv+Y3MmPlP8rfqcPIAIc+KObhcuBGoW
cmEMyNWMCmu2DA9F66OfepEWrlmx2ISwUjkDKkX34iXdCacTRnlq0Arb2h9t8FVOf7Efzwmep4bY
ngL151lM6NoI5dD75TUTIjUrGPGGWCqPGtDClEgVjTk2y91RsBTl1vpNUjkGM+U8+DQzCzzRRJtV
VAHQFAu6ybfxzcbfup+lpuQDqwRF/yYoQVnLXVZuroG/f6l27vCJ01ljd6R5f5xq6OfbnnVetWej
I+rd4hBU5x5+cF+r934bGMw9uMHtxhH3IS8yNCylLfWRig0JTCpC43QzUMGeskMCtIb/c8UrACoX
hrUS27jZr0H4Yz5GcVnR18aTrNWxKMDJ/JjryF20O7PGd4X7lMyUefMS2zSr8EMIoIimIeR0VwBj
PAHEegUEKrg1GweyDA4C72r02TL01ku1uX5nHFVIMPpZ4SiPggRxz/YMvgX3N3zShXLahV7oMJC5
6gcbfSd47oq0TjQCqj3nVxcfLh+6QZEK0Uj10YymDfK0oszbMRXwYjQHKAITuN3vZueG4QdVu1UU
LH7wbZRuhnGsHg6imro3vtBEEIxaVbVnPkk+ndcnGz7IDp2dxiykVY8ZUfMRtWsPY8Wz6xJiKePc
4E3Wepd85hD3/+8CrB2zKG+qw7qsgJhDXODypiZ9bT3BKsCk06aqgrbutSgS++jBAiQ9Hs1RF0gS
uKjbilg9yBYcS6j+8we+a3BwkfaHCEGpoqCQKrfVBw2H9Krtu2i+whJOKIPa5/Y4ChsbmMgVxvuo
tWWqHBHUtGBjo5vZQwqxa7cryQW08d+ZJgpNK6h6OU9PJbqU7ITQ94V5XAEk9M6eJKIkJMr9iOgn
fiqnJmOgKI/xCsvJ5/cGebxBIzrgzR3SXMmMF6MEE4fXM+RVA78X1FBsBKkMW7anQW85ql7/Ob1n
NdX8rOe04CjVS6DHCARkzfF1dScHYbKtcPwwpwIyK3AYcrO0AB8zyAua98MW9K0597X6iJJgeorB
XdujpR6J9tUzq6RpT6NmKbRB9EedcI4419opvxtmzL5dkk5sVWE5t9jWqnU1ethdl1l6cLrS6TF5
benuId631DrxXcVHTDkuz1pEXuquqdoOXLHpABOr2qnQyNDcrMWhCPu298BOBzn+Z3HxhRJ55rRS
mSTbspjfGPSEEmLiJnsWZAEtPaZWUh7Oi8GZ35qYqw8rf0kkqQbpmB6BUAqz/v+MLF7galnextvc
ZDpQm5i3EkDrVdzjdxRESutb382zQF4hZtGp5+n1x0nuW2OTIXq5mANGiQSG1HuGexx/EgGNUlZ+
h2MTTW9OMP0Pkc44z1081JizT8YlO+uKWrn8iCJb3L6UL4K+O77vDRjkIGP51sncyi0Q3ow6F4s1
vJD9G/ozXUNTo0YGlDiGW5D+3gmBmVY9d/A99a0rnwMNLHUb2ojZ5OcgAV8nNUMXbdrBuQUAmC3s
OCTHLim04b9FmbcRC0zixeyINjvLjLWi9qpNXj2OTXbHW9TNNV5MQxQDDMKuRv1HgNFsGJl3Jp40
c/m7lUKzh6hqnMbRRImzEd8BAY415oeKjHF/XPBego9hLuUzWYCsKZG24ghvnx6aglT9pC/bVhro
gqvmGGE1UvLYPm+IYAoXASVoNiehQPb7PsoPy0No8TbmWKuZC9EU9VdJcw2XqPCSxKK3Bm9hB6s1
7MjvrH7mephcZhZ9VRC205vuLpxX7y4pkYkf5pS6N4bY1Yu8tJC/O5/aPFVWfVzhCMdyOopaE3Ou
81PA1E+y5Fk1965fDz5ZIy7yF3vhZDNtOZdGZkkjdRPZBc5IS9g/oQYN0dYyzetDky0EqrHgTs+U
rGlgj8qfumQ5VeOH4zwd2f6Zkw/t8qxmLYOtJOCIVVQ4pcPfi/JI0Ft9bwXh7IqZtWfPen0rL7Lg
0L2O7G7NNrkPL6rPKVq2UPk84cRheTtTTGzEGslr3aowRmnjiPDrO222Fm6c99RHV4J62tCrfLCv
vaDvDFbTm/TI7fj8SK6WsZmsf9G9I7TbOGeuDlDAGBIQB3qsnW23kJLNFZTxgQWM9irng0bVpD9D
JktY6vOLgWYMtUPWCQ6a9D4SwsN+hNcbOD5vRXFv1P15Tgk+TGN4bJsue1BIeJDkvSdyfdbEly8W
VAfDBjnFPshs0Ploz5Voa4XloNaP1BwnObzQdrMsodbF9Zl6qsM2faxaxeDVFzBw93QLNlNIyumu
tZZlKNT+TJ7yB4rcWWuz6m+V/S4BnvlYZGWW1HpRVvKyglqH1AohlKhAbohl1oX8OwEWZYbLJSIG
l6qeX8mLhzYUKwZMlMNN1HnBF/UppMcf9IjrfIm2pApDFzZ3Jmm3GflHDCNQ9qQT8HjUwDuaZZmE
DF5h4zN4R1g7oDBizcFLaP50xGpo9FH8ngEM+mMu7bNqPqVXwEiTkrpazf7a2FZdjs58ugii6Fau
p001T3iYnWVeDJ328MNvCFWM7+yujf+zPhV8Znl2+sO8/yDUAkAyCmPrLbCCtigHULVedkKTmgfS
Bn5yfoH77AllTMqMG0LHQXU8l1OxaKLwgqpS4EH2i+1epjygvArh/8UAmm8vct4fAJIOZh3CFjth
tfTGMQCXSY2rXHH9BhgeOaurfqabXTV6NcLQ+tpOGn2Ot74mDg/YIEoTWvSOcgfdx/55ozBeRa4Y
EmI7FlQqrJC9Rjii48r5r3wAd2BOniQmeRBdwa3MHMu0vNskRplsPUHn9uXs8+H8D9JXTCfcrTZG
Ikvl7QOXlRa0XACi8iNgObV7/7wTYLlGXtipdEVIQ7vGfVIBCMbGuDn8Xx3yidy7v6v/uK0hG7dP
Q1fyqqwniiZe+G94wvjvVISIcWxu2sgCbG73Pby/mcol+Shvil7IdBFAXjDuxEWorsisQlg6jLNo
xRH3xcT5SJvznYC99pU/8S+XIyIh6YuXnx2+bLUtOEXqDYK94Eyd8gWY3Yf3FpPTsLwLgGEOP/SR
nUh2oVFDjS2sBLq9BljFjlbRlhemCqBxpGVDUTJVK7eJkLZUWk0Wuxmtge1OcjxeVWFfhShczO4m
4UlzE1fNIj/G6I7UMzWNgplBSH+oq9hFzuqMGoFvStJbHNKxuHQlTwEKbcz+4AFn17KKdSQA0/SS
Q2KZdahLvzPXaHU64PA1SBSAW+1u7OqBiTkJSmIAFbzLvIS1jboujEr7CY9VmRAQP/cbwkXl4j4s
VyAh0MyciMCwE9RbTknDY+aqPt9kOBxUeNuRAla7mdFhooOw45u8dfw8HXcz1PHQV+trdBGP6rTt
Pen++xpCumKyYreX77eaE3dOxTidX6j0u0mcpVMpQhGOQMoEDwEzDHaIqoZogNrEfP14FoExmPTE
fLe7m2EVtRqzPhkwB7baeGJ9Hr+X9MI2vFg6Uklaa4A/LZTw7nfAAY/DLKxXLYVJFCMbyPb6JZ+I
/rzdD1WKS5l/9d/pSnr6JeJzUW9ii/L0cA6nCtphQLjS0C1xINX1NdagKNl8VRpLY2WUpRTthMGn
Qr4Lm/REUtWNIkp3LrTn0Kqzxg6o6O0FK3bB+56XOhya3n1OOwuCA4TKdv4cn5pr9SEboc29UPa5
f11zW20wB7Io2VkB/hDctGpH4YUv6Plo7osI0qZkWOY4kLueWJsk118FKwKVzpxR3ji6d2Yh/BIg
8wqH6L1LPAMxRTW/fwJTquaoP5eNqkiFfMMCn9Wta5sqOxjei+xdoSsWglk7MFRf6jRxoi9yJdf7
6fbFyrrG6puaHjoJ1hX5HGhW/lUkRJb+7zSZAFfto8y5MDyTECj2c7K1gLsXYkOLhWEgo1C59pKx
3Fj+Id3En7P7BqkZU8Q4BduZDh7pQ+UAvIdc0NS5NIBvyzXe0EtnNwk5A0ehIkmjuOcBmqB+cbvj
H/Z+AdyEowbD6jtdxPgOKpGj8AOGjQcb/FQt1jZ92Nphga7mhkLSkTwnAoW4+XUKPyiqkihOTzpE
gknMAlY3zO6xJ6m0Chfzmqfut10s0qgSSgQkPGoE5OxHXFpVyX8d7o7g5jt7B1vYrtMgODFgdRRh
E2z1vRg91ZZtgGoYo95eJ2OOG+Lnk5tfLPhyuLa+zIM2aI4dGHCrNXAwqIcXoNTj6mUvM+5yvMf3
7gPwSN8rl4nlm2VmrVEk+gCxitjIQDAFeEggWY6s2OrJz16hXHs0bgQHwUqxAuqwyCzIwGtRpYJz
XTw40ATlu2GwfEjj8LFsYlfpZO9nFw+GoGgN45qNYQQ8u6ORP5Zp5yxJEa4+ilG+gJxCoWFDnh8Y
xxzRTu0VME6kuID9xXKUtj6SCHHE3Z+T3DZ5ThPUzR6dcVL/7Alo1S0GlefuLy7z5s9qLxa9gPGs
eVSqXdOo0lGJj+DS0N7gcbYJ+6DN3mMg7eJ4pvg/69RMwiahw66pe4z6tcADxi45NkxAClKMH0Je
hgKZQerDBu7WFlxWrVOegj9VgyKDYFONU8y8q5VW2r7v/qSYxdImMERVm+zrRqQP3RjwMU0r8Sc7
rK1ahto5k1l/HksPI0d3KtPs1oLSjdbaEz5jB7MvVqrTrh/EpJerz5q37uhKhCFni2bGxVa0NSh+
ZQtWUMxRyVTMz7kBkdC4uV85m/75DlRE4iDM9J32eF75HWDg4qXHd/q6zPD41Vcn8SoPoKyNPB23
eENVuH0XZD7k7t8ysQJBefCxklXy7zXQFP5i3LrhO5E2haQJ2fFFvDVkZ2ANOHQa1UX6QPSfxlBf
AVNrQgPF60mNbDs1F4O038J7hn7Cjt+5cFC8mvTDczeSw2bUErIreBkZTRLyiftOA/NQ8bIpayCj
1U6vl1c2g6WteiY+4DU9W5rAPQiFAZ5Fw3i15FSwbToOZJFwQh/u2JqnzbRHA0A0qcnZkLCSxj1r
s7TDDVUedtHQN9Lu/26ORTJ2qDXXWEpuSHXpKdQAd4IiTH+rAcqp+VfDox2XVZXnbYcwXaR7r33g
Gd466tox9Xv9EnWw52x1PClJMo2TT8/RjQSPPMqIZ+zYVUZKUrB5AiOUqbroPmYLU1vZa8OFSWOy
QVsE+yDF4U3LEpKMYOyPRWc5K/R8b7UALF4rygJbIwShvthzVse3Hhk+3wJiNU1yUYaKFuKDslRP
LsB+kA084mW7sQF5OuypRxQrwx78pOQTCEruVs/FBYaQO0QC8gkIk6mX3tHvnr6VnS2BNRZUZrJ5
vPfUWAVwIRfIFkKBvFBi6zrEeBazjOT4zkIZxjESYlJmPqtVXt745rYLdvxKsz9vxB0aXn6YRz6e
a5aMjxU911gh99VmQuQyrLIgPv9VOPKUWMa1012qjwPRInj/9wH1yqYt6Tf9G4LCxTtH9twodU9L
oXiiBLWik4fmLnIMNNXJFx4zCq6vJUGGy2WUq95Zys1VPOfGGkBslTaqDSwNyvCAkDAoYA3mum64
kuFLE1aLywnrrAzCq1t36Z0Xgg6CzvF06j4Hiwi7OefBNOY2a38LpRu1Od2F2klCtQ5d72FN93R7
rCi/QMc6Z1CK+5QbanZZvQe2VwFgGU8sF9+6nM9x3B8TxzwDu3vtYWOMv6YbfmZO6cyQtYw0T2ow
fSmypqkI/wYiToPpri+kT5Mwm+wust7dxkXXgtUWfuXXQmf4c3J1N1aIe5ociOsLcKVR3j7UG7/N
Td9SJM7gkJu3iRI+YE4W9I8oruIlmCDTw/h1shijLIf+3bdaC6BWLeG64p6wL3t8PEZaVl3H11wG
8bhaTfzpPyBRhTYJMzlHAazB8LdZVPChoJaOBu3VI75oiS6Za2wV/qW3VVIhnsstMdONObd4/4xq
TnuvTmDfAN/JwUYVB3J7hlI29zDcHc7SUxSA7kN1m/Autzx9NgrH1cXe7wtOA6oR7XMW+DrX3r/n
JGKegNrTdXBADlVM/wJg1ME4bRqo63WgUV5/xhHXJat2/HdONC/JtNIPXuuvT79LH98VQly5DoXy
2ASbqbUiwC1OmFj8G6JXNmrrN3g2S0abevrsUCx3i+jqpMxvXXqLrm887RDOffCyu5QQ/havKLoJ
KNGZmegrgNWDbPuWbdOfhsB8l6EGMUZSkXUiPDwGHBwEmA8wSAv8SJvildk/K8qTIX+wXiQeLvj2
fMcRHwHKi+ITUVI+PYdMXe2GitGz6IqZni3amD5bYAaNlVZauxmLqtnHlG0KwccOzBTdRN+5T2sq
GMALsMaRPz94EXntqbgsHmbaYtntgWjMe0LkVnU74aq+iqFjMIvKUcjXOIr2HwXl9qE8RN5z+I9s
VwzWqfbDXpf3T5HmOCg6sbQdummRSkiPjKw+CUWPWEvKsXVC/M2VN2c9UYHbIQKoT/AG4BbWjjBd
zpRnjErT+WQRJ83SaAzgPnrIH3KvIyXH+o67QojO/6f1GF++XeF1hDP10l1U2/UWubPPcKTF5qGe
fhl6Rh7USIG+Vvw0BFH/LkH77lFZhh9zSkgceGSCPmnoNPZZh/1fdnA/1X4NtjaAcP7dNdKW9PYj
p4EoDmyYImTqwFrb41poUGu/e+9Bxbz/E6uo3zLPxv61w1bHJdvSmtMZ8HFzKlULeG5jeoiq0YXh
N8b7rK17p4Zy4ZUhaY1lChslQm23jmwFauUjSIoiNqhD8gs0NceCKjrDO0aofX7w68qIrlu7R0mm
q3FsIvluiUqD2iE3x0byliANa96szxJ0k89iP1bkTw/dlD5uXjz4nV7gOxXCHS/xWNbI+3f6R11s
oaWvdBC3MbZn797vghFvq8YUwXNu+m35jqq7JBDhvBdJMAJoOYygVmX2GKrB7KXvmMMXyQdZuZrM
Zshi8VFKWaDSQWHNRI2EK9yaMGg+eWbcgptXRBzuXwlIBA0f0f4M/LoGdSRuAygFUm1s4Cqip+aS
mB1yObloaCn6lglK4OSEtsdw8EAO2HinvP6Nc9VZM4eLInjyjedk4klJPsHIjfNZNzDBReOmmGE/
2Ur6Wz9pkCFyTwXi9/G9CR6IksyT7+sf0E05qGvoQ2D/E5UoIdHWBurbYt2mJQ3E138E46AlrqRW
QdSqQa7Q49jt65K2pHXVj2sFK5shQNbn2V7Qp1hgi8USWRWy7A+FxIrTM7nMpl2Fw7kVgLzlwSI6
LCSqc9ei+fcfMIBlJDrBHHoKS4+OCy58t+aIT2IO8TANuS0AgabQ1igza4CsxArg3zGPNNdHWRCP
eaCX6mL6Pxjrcssj78jMDDQMB1ojDNUIWBPZzgHxhx4ppwqkZ/lhRKV+w1e5qSLbGkBnZYV6zXpa
/Egd9LFJwwF7+14U12EzW342/334K8DCB6Bg8rYhj0VNX0lO3QfIezT22loXcnYpcTjX1IFr1g0u
p2uaSQrXJ/z5GiC83/rc8ANxRrFH/DdIYNPt0z+m6WffYcRf89/6PcXu4o57w9aWW7Sqx76ogTIl
jR6EeYU8OK+HCfSRO3NLyhou7RUYpD8StIpWCqa+1Mct1dCa3wuoXt0M3fHe+Keu367cyZ7sIsf3
BjHRIpN0kKn0Ue5cjC0nZlxTCluImA3de/ShkbD8x8o3fl0UXI1CfLhAKE5O3sTbBDJ17Nd2bm2F
1ufueE2CoINgOuperCEwjvGZr1DaWiOxwBnozspKrXArT8sul6H3udQ3TBPLJ3zGSKfe2rnT2TDp
mrN02Br+rEQmEPp42rgGXSsFAmbzdIWXQpz93nEUvIVO7eaFhE3I9pYvVWWl3B7bi8fT662pyikY
VGm/lzJSO+fMawmgJtKT15C/k9m9YGIFh+kXz3aLIarxw1yZasdM6gH8fbuM6sdyYjpFyHTS2/Yt
KU2hqHRgAq4Zkezc37R6gFLzCyQtGlq5H2y0RjKlxs9aRu2Lot/lenSSVPB5UI1UYmMd+oXFy58N
ayIVhZ57HLzSkuHoWMaWOhFNi9n4wXLhTuy+NyBTqfbPhliAsdkFY6IiUSrisGDtodEoV+sm7j3W
Fxmko5lclozk+bpBKd3k38Bgqje/zbBOrOtfRuJagDYNevHO0IIkOjSjdIQbRq6PKfhY89BuTJgt
neB+MABhB/BbpJztWhrZ6u77Nw0x4Tl8WEuNdrSEeeLwr+p4huz3WWfXOroFpmxMV+g13sBm8BtO
cWmgiNxngRi/ekAvw2/JW3lrp9RsREofxVy7KRP9pdo+Y3kxrXr3n7RgbgfOQiIaS3QlntY8Bcgx
AHglLxoyOI6cqUgyqZdtUkRDtBetbT7bVPqfOexvgEtvmdfWJoIlr5SYgOHx9hjb/KDkzXIkNwz7
TLTY1pv14jUbSGPzf966C5rktXwaIlBq9mJD9NanaFEw20lyRgnRtCRoeKKzcHNfOSSbUIAoStEA
wZoZUASwp3xURC8PTShodSOxaB5HaJQIzrL92eh9oSGIY+zRNCCAJtL18+a59a9REiKtXsxMc+5I
OWiH+WDsJFYL1IhHZGid7l4UgGKJ0CXv2Bdyj0RqyhLSBBikI5WgUHvNGrZr090cPMeYYG54cN8A
9waDFw3LnAb7k5OpYtaSLGObRDKqwPcKhEmbUgG79sfIZpNdz8X/TYvFXgfRfc7QahaPMvsCTuwR
PHoOIt6+DOftCblEGSqHTFJ6BMmvtxxMywS3gOfIKZnCO7wsBZBRLF/hTbWav/aVqz/eIQetnod2
huZM5PxG1Yy6ZowXt8/YTGiGpq5v0YgC0jYjU7OxONEquj/7B/B4urwvb+m4v+ORXvV8WSbfs4fn
HYpMofOICV0NbfilNP00Q3E1WPyoFAV21qSk+twwQBUwqN+rcn8iwlxdwJru7D9nR6VW+yJVPNLq
IKnvihDxmU+iWmcEYr4jmwTtBlgFCdQwaqILlp3vX2sH3L1iGjTtOq1sWYVTIwK5mJi59cFfvWfa
3Ibe4bI0PnzlBlRhFbcno1qaoeqaMfWMzjOq475/0TJq1c444FejQ/fK3wOybDvlch5jOJGPRz05
IWbIvN6/gT4HMbGdqMgU+dRw6neHg6thVrYJa6nCeA1LHrO0S3mgisL0jKw3gS7MibaSJ60QJS02
sHg4hptMNaSuJiz5A+r9jFyD2I3BIDvbrdimQlubuvFF0v6bEnrD9i5rvLl6CSVuNoN2d1a9hiXS
nLU8No6w1UEFzr8NJKMWiB/dErQzjbjJjf9YU0XoPIfZtliFGNDV2ASz7unViyRugiFQ+6dPKd5D
oAMr6UxDgHTx/vxNIIGqm7CywbXa9iAb4Q8sEir7xDO57iipStHjj0ECbHHJnz8AwqrZxuQ4qw1K
VnxknGRGNtlAov26su+VTLS0hovZ85FD2qp8bMHl5QZ80oAmQLvePMY+5ZN51/CZi68Q/0SnrKNS
hIskcdZUAYc6WYFqxqEn3tmWJvXrGLoGZN/E0heg+yIdWRbfCAM94xDjMHu5UJvfDmD4ak90H5aE
8eMOV7A7Pwx9L0H32PgDFYTPZ4VT36Ei0cZCqBDIcKR6yFMFCIKsGleL1PCUJFkcfJh0DiryLf09
FX6By3i2diEsFmPnQO0sIzwsXfiMHMaHR/RVrfHBrkPKOvhNN471R3X4Zaf+9zYq1N6E8Dq98OaP
B9K+ChzA16h6Q3/AOG8Km9upHS7A/6nB3jiQuL3v8HZL6y9cDw4L5LzoHM4aAc+/hpwEphNPHeAd
2jMw5yks9bgYxC0wncsvw8fU33pdVlGjPPR//aS187SWGu2qBfTe+ini/dPeQm4cw6CVeaAz4OcC
Il2SNoSbdqOxU9gFAQZaMrKYzcl/HxzKSiwhb6uGDQ5Ql/zbOSmWAjSywCeLdvPWaWQgQ8PAkH8e
SYhgpBB+rRPfiU+n3rT4m/nUoQWqyXW6v84P4hA2RDgMIusUaXVR0h8iI5kyJVtANjt+gheAfubK
uLKjWNafzGwkNza4d+NOpFRoLlyEig4Q5Bo8Jj2bLPFSuKPOEuVRw9lNUKarJ3Bgb/YGvuj/LELu
1E3gjmP1eqUDw8vOMvdniYJMH8ma0xG6qFdlhf/QQ3QFyjhAC88l4DZp+QZ7GT47v7Smnv/6MfoY
gu1tbihJmND1zhMq42sHROhX2ih9S3Gfn1urEGiFMhFC8682P37OoS8+r3cog18UJKOXvnZWZsmZ
OCcUHpNlaBiIlVexwLSM0reetIEX6opEOYQADQ83rdRlHNEUflXD1iXL3ouFtVcnUbNJInijMC3l
1ji0gmfXAUn8E/vHcB+FpUC3qbqDgGcUNFs2C9jmctBIIbOEWiPhsZLv7ueiH3SUyIusS3OKeH9E
l6uhs0Rp0tua+JIkrIh/OBM8DHp/faKedySC6U8kLZ+gU8ttghRmRUxSXY8b3eKKPsdSIDlqAaWw
8Fekp8SzENC1SUZWQtGftyGeBZf+csZkmBuIvFFhibkCo1ZYN9gUH+56ppXd20DU8S50TPVUg8Lj
GZ5YeajMPMSvU+w+3wzC9NDbJ9fVeU6YmhCF2wjPSo2f5b0vNyA+zFTnK/BfJefA7Isv1oOcZa36
YDmkS+GoQCwatTROamFPtSUl6iZVk4Xd+bSTY6F8wCbt2M9/W7OYtO9F6J5oZbbX8642QMHAbeDU
Os23xcAbV5GeoNN+a1wi3eUcoxVYuSwLtWfiltZlUrPCPYIM79xPK4DgdByZ32IOBlowBV9U0sz2
e6OY+GGDeDm3UDxGAMz0kOh9tM60IOyeRDaPR0JVo+JvCBX/2o+m1hue4g8Olmtd+3QBGSUxumyV
mecLnyG8meYMYhEutVDGQGgmROC13UZj7h4zZoVKDp+mkHD8yGtwS0YDSjkayQrH3JCV6vdCrZPM
sqzkmdmXG393rokQwiOnRP+Q4o1hublNL3I+SfHlCRGfO+Zr5LLcfEB7CoPDT+4kQ8DfBVUfoLaj
owO0ES6uc6v/1uxmZZ7nqN509kRKR7Vo/7MtyJmY43cs0mpMOKfk9/pV2bWl1ZE0zVaXByAxu6Wr
7jZNpqV2KHF2B3joC3Mi1OtZNHpmNtNCUdwzU/nl5W4RpzTwWExNFYdzLD5l9oRsqhPH8SeqTJQG
QyZoLRCIpHW8BQwCN/YUdPUY+2mz9XhrJAMRrakftL+ml4xcMZ9JBxqoJ7maUD4yAW1mtEnZ+sLS
+CZ3skE4pJLkFccqLVWv8o3hzdI2UmvxaRe1Sf4niBL2VJ6DQSKesUDFn27Q1/qZ4HKGBXJuXIV8
8X0MDC8ZnAEYtziiIKcWgTBP84WsFYdrOK3gYDCDQON/Fai6ueu2yBEXeCSef8yMmKvh276/wtZj
RzfJN8hz2XRDpwt9S8I/I9p6w7MDVoJejF+J/qIu2M3rf9YMDqCxyInPr3I4DGiU1RSdepREADik
erOP/8kxb5C/kMh6nPsyc++6LlsrxysqSk/8GxM/6KRVGKP+5Zv1EHCOBQbo7GpqMdPa1zKm3U0H
aFJkVa4gouSA+/9UA1qdBlsY+09GZZRlwon6d+juHQnLM1ci3wLvZIpWbjCIIq6RPuZX4X7iuwDF
dutG1bBXbNavHcozfhSqH1zmE7A9YB2lnZhc1ZVvzUHllmB/QNXKXZIuTN+6Sv7ZvQLEUKfHu7wl
lW465G/hsNDAj61BUsQQr7fMNutfhfSFD2DM0lOyU/v1u8ET5fnqmPbJV2v2DGRNiQ1cu0+PU8J8
iZnDKXtKGVUpnZ5VtF2XTtnmOd/5JCMZUMiNNDz5UUmQTH53FFCUZd1RckEhCkEFHfidkoXXbU8m
F+XzAAcqQI1P8vWs1J+tC0ZK5iDXThsfJVhwAYuR60IrxAqeaF83hV5R1fz1gqYu8NURNOKJ0OFa
Y2gLue+OwvA4B5kFGTidwb4QD1Z0gLra9RW3nteozrNar75PCM7adIIrqaIWGzmTix107rTBaSph
GdYIXTxt+P4PMQn68zSn57vT/fBPtjjuox9DNSWgEwBwc7w3qHdgStigY7Uo9FSP77fopW8n7cFc
fiQl4Oa8YBnHcCcamjo8MMvgHDphWyWy3zxdcjdHOH0O+XF3ZLth/b5MWAeKncBUfCjmXnqr4/Qz
IJA8cZ0Z4p7GJ7HdbOZ7AXv1lm7JtIhaBTy4sYCjlncvvv3fQPTnZtl17nGmgmZFqjZGGxyz4CmV
3k2EvxY0soHl5PM6Io11vlcFbmwxFLvObCeS2W0XNyRqTXJcu16fQvP8EwavG5/Cyg+K5AGh8vYw
GYhrwSnqEiz5aRtcb7GPSr2msXGPiQlfdRSJM0KFLpCCOj30PFDbdET5f5bsMe/eElITWiKecr34
kz+8/YsFt2HOc034L8xnSWMp2yBDYRSpoA5aslOnwS1/onK9KdJeWlkAYgppj9UECO8rH1RbXwDk
zo0g86x26mlSQYkR+iPL+eiR9etXub9zkeF6K0MwmZFdD650JWMzltgkj9S3QvVHlvTqiTHVKW5L
qeqr6+rebgUPivkZsnFb3CwsIAs5N02Myf+fO0iuGLqMMTz9ExkDo13cGinXAd1j9Km1RHxCCx/Q
/g+9rszo8EfwQcBgb8/hHJZlp0c/4NfRSCoosbkpIUXuCR/MMFFhd1XvobY1FiBVMdiALWQylS2S
ss6HJ3mTAZzgJg45HO5CUl71lAHJJHdhzWXXmDYVm1+1xxw5twoM8vj1/twQgkryh3AeAFBNAH5m
lAuIEYgmwzeDgTx4u020Yn0aS4SlCjCBqqHYoiWyjgdF4SYlu2f7+vDhRV6Ktd/tAvcdOFBl+LbH
gXWDvTPNcwsgqPATl8Zd0RrHq2FO+qN4jxQnsSzkOFpByaM5r/aqaxcwWJ1cWKTS/dSiiE96ZU1U
vw8xEymBr//Z2+pRNPvj+eu2xH1vpDEgXMrNCtQ0uBsublASARKW9JNAwJFUwvbHMXqAM7N4vyi3
4ibiaMN6aSjRMv02g7aTbOhNZq/Grd8n+4HuQhTYk2j18fki8KCeATgHZYfYtTDW9w14sTutQUKM
q3QSLNL0mohpxayZg7SQ5Cj33pq9BMPDzOLB3YBDNTh61+iqIT43HgNb8juc126lA3U/H8Tbj1+o
gQyIyzd6C/8k8GogTfpFUSGyYfiX9U6xRKZNrxEWxo4VGSbhDbmc9EikZcrRBHvooRGYsoL3MVFr
0GbKt/ik1pBmnH4TObFiRo/JTXRRLDU1flnu0cwvAMNgec/odVWFjkY2Y7wViLDlSoeYnzQQn9x+
ikW3k2rgreKP7vZefVqgTx/ZCkAtWlH0jLeGmeniH0HSyu9La62FDbK+gmh6saUSCK+U1lHu2Qe1
RYBP4tIMi4MnsFCPGBggcBi1I/EgA+ehdBGZLChwgXYgOAxEpuoNw5k5jB8bXEgKftGCBvoKKWEt
CiLIqw5AZWu35oDbaXzf50X0oa30U+H1VuTG0ec1LXy1zbkDjespPvl75Wewa1X/7JPerQ+hw++8
IZpJlaEjLgfw4LyENRHTkU1G4Eagg9WOXwe1kOutthxaxuFq6qeuTIqbY/zB1UMFlmIobZVyQqZV
sioHTcozbZL7batIxHnQPD54zun+9iP05Wwhp/rFeP4uHIPIeYVeBYFqNq2U0xvCPG75JRnd5+Qi
TK5DS4lRnKrAn8q8PuXI9mxYu7OzePiHjGhLEb2sDZFopk9FDiCU9r49J1sUuxyRJJtstcxHk5AC
WQPqldm2mhDSSHMWivRxH7UGjBMf7RMtWXQv+PF67/hLnzF3ePaO5xBGDTT1b2G2PGUpBFVqPe88
M/wNPk2u+daV92eHSHUBFmRrhtgyKlv3NQIavF31PDGtBWGQYOnEw6V2GO6Bo227WgjB4JS2z9AB
JNNNFFrh5DBYc/ho3oaWQqpwLCsy8WSAQTnjCzDxaRzN8aRM1Etqo3ydPOE1pwlsSsPccccVsote
H2v0e6+u2NtlGkGYH1e4QNmBsPlsepDGwjUhZO1vlaRu9+b7yUCCTiZ1Cct/xsNuempZNwDLWTef
omoUW2/BtR4tRvN5GnNYf7+DidJSC44LSCtcSk3+TO/yn3f72LRVySZGtbfFuD3+hGnubx6dDRRX
McLwPdj2qmzL4okfF7ZWtRVlrl4+PCyXPLc58NFCankMzc71y/u0fqB0HGzGmGlAhHyuBfMJjnfN
ZF5o0eVRfmEEqH4fmD5undGIKuyMvyhAjgscC6b/t0QjTnAxt3ZoTs3H4wP92P9zRjInzx6rqG5y
n0ULcJ1/rP6MPDvgZYQuN6pESz36ctTiy/RzKMpzc2h4jvkoQQqCcw0WZWdbSZSI2Cc/pRBR7PvZ
pPDBbmZ4LwxCsFmZV/GbHDl4l0kdjJ1ZUyJ/uphxXg+EaFWWl041mpPwRfbkAJUJBsdH+XDOBT9U
mJ7BTR3xUM5actGtSM44EHVPR1Al0ZYa2mYZS+A+warYVGubaJ+uOUSw1gpYrUlQT7wk4lc74eZS
Vaypu1epM/pxkbeiuh2meiQYk6n0uqT7tCqGI5krUne8VKPgDUTVufT+mWZPI6wqia+mTjWrbCBS
h6U483uV/E1i0gBwsQBfOlK//MYad7/eBwwP4+No50Xwx9XS3kqj4LgzvMz6TUqh6DRKIEzB6R0D
jAgTzAr6gb124EiAsjQTHGIm1QxhwF0b+V27HrVA4QBKPI50WZzZKxUjeqPv4HeaSheYR4qfo2Sa
02+/ovOc3LXhgbke2OGdqkUW0A9tmeV3zRwNBKdL1owDixgNQpbE9BJy1M/AMTSVp76gCepoClxP
AVY+oTrIzCInVHSpmRlW9NKY828mejEv5obnMmq0D6KdkxqXrUI3EQ4/P7roqtK4ZZFDE29ULrND
sa4wFXYTMI20zeiPOKv4VV8MwWDYr7qSPvF1y7ooK6e457Xug5FTEtjxmt6zHUeztarNWS6DuJa9
87706likfvfgnM6tGCNfyJ/th6VGxOlqneD8vyuaup8++KDnR0Wnf58+ih2iXQVojlPHIIHnM6a5
JuEyV2rBMgohnhxM0h1u3wjOyQ+pY9YlS2GiPUegxehYB6cqwa5Qmov1WW7ztGPoT4nGIsaFxoee
9gJYxi6dDsfWq0vaU+Xg8X9CqGfic+3LPI6xo4FIsES2yeyVdhElR1M/Xc6v6Xrf0ISh3EdXCj+4
qlMkobodgmDZvfPzJJ6wQqWZr6gh9YrIQvRe40Ix0UmQSS7E49lGbLZ/Jy6dEn3DakdFthHmzYcm
3UDet0SwRcgHkcaV9i/C4cGnrvDXSmvxhLvH6A7l17HN71vUOBlTJ3Uo/RT+BSbkVz3OcUDxJT7P
DF/AKa/Gj5Bz2SoA/I+sT5cJEO9/uF/UQe06WQfG4+xkRc4DUzt6TXz9lYRMVwi5sqNA146n5dyH
ItL90Gl9alcLQQcY004Gummo99dFJ1JFPZBYvdO+4vX72vcbfeiyB7ZuZ1E36wCt+EbWCkvZX+Xl
cbLBjvO8YJb/uxLSVD+KQ/Orw65WXMT+NlKN2G4Bz5nvIcYGvUUw8T719KCBAWWmuDXDpF40ITZk
lAqZ9CaihBas+tdTKQDKy1tIpHwStUiy31Dc4u+J5bctHN+zcgzE4RzXK/XUqu789d+xy6AqS15x
0q0BgvbhbecI3UoWfbVm8UxY6ZqRZ4GMHSgrpOmtact2BIjwBoFqb5S/lfepvK0ngXN2Zrghntg7
aWUnGxnGt40jJ5Wfx0dVZJTVrnAx9Ixmr+7dMdOx5Pf/XaCUKyN3CJM8Uzt+WqCdDZCPvJVyR3QQ
qJp+/xjxiaJbkLAD/ZN+vOF6NtPbZY77TRlC6PJDCJWBM8qpDwyBozbmlb7HCsA0diy+Wyr0X4Rt
m6ep1VhvFoZmIQVen5+Ucf9EZqFWwUz4LDBxbZlFpHgVLrPBGE34BVUuoQt4fHOlWm7PIP6AUjPo
31QzXJ0BCA6CfI2GefoeVpdRsdsCy4H3H4s8Wbgy9ncqDvGYmKzrgLl/h8MabDxG894tqND2ljkK
00Qov7QCW7x2TLJGkV8FynV/n6gSTDvmvykCDRD5GrMpMZ4eMC4Csc4yLuOo/L5X5lfCKyB4mJ+W
6d4dfsf9O2iBktp68vUgjaxnL1dhH4nVIPVZzNqBVy2OSzxtJCqxr3VhaZvZJI7DIlCp3+hkz2Rf
VfM4qL7EqZ0OaGz3PBQ8iuG4Ic///c4/TPMW6cobGfoki/U1Of+BFRX7JzPc0VrDYxI17dFVXMGU
Fu+gfiWrkDpQ1QMnr5z7fdKH+XukODcoeAVTM5iBUpL/u1WEdHA01y7BdiAU2zL2syjsVHPvJNMJ
2XRWQ8cFcJriWPcmIR+/b00Nc9J+yyz51ZYLgag1d6R4HVVv6XBEPlUY2L+GoV0rAJADbZA9IIh7
B2pR3fK8/zhsREU8rOrvsrN+X7/3SYFcMjW0ehykz4hMA8+MmfYDlM6B0ZGzJ5wHvRWWu+fDHg67
b1dByfGUgX1jZZLOxIL4jKLMbZn8ivaSEri7eDiv7J91WcQJvUTZIvMSbml4gAcKT7sK49IX5J5+
RzXpZRWDbnhUYDj6ALk5Mal4jG4u8NPEdRHCvSm3giYxBA/WTwqnIZEcTWQR8doiPs5z+9V0omOG
YF4ppG05uCkz5TpDokNTJ7O6+lWqXcbBXR6X//poNYIT02kXLaGymQXbN3OgZGfqEjbUptMGepz2
bwjHLKYgr/gT6jNkaqmIfZloUFpAcvquRCH1mrlY6/wcDX6fZSfWlS6uwcG51vlfA3ZW/lMOSq0x
IxgavOLWi3AQ9eTFa6t79ung5k/0urrIxaV+GMzbeV3Po53sF+17/YYUtSzNLoOr7Erb2PqESuLZ
EgiStSCECVXWGYNP8Xuu1HgtIjM84x6Q5S1aYGi2oKwl9hgQe2ZMoFQXja8PikyJm5yzgA73JuEo
T0DOlvI2iJGKnuoTKMToGKKQXolFGySc95cach1jYIIzSRMzwHeTWQtNRJQFKV4IIJXEYTlUDFu/
1456n+RNPdApgng03ww2c3R5puqJREcYcBvtPSquTXK2ln/BeNDVZD9w4ZZElKHNQBxHCysphGRh
iOeUOT3ovYRwqCKq5bf0s0jL+rD6fN16BrS5LjeezGuDgv+8kICCKyS+zMUGl5Q6qPx2smdD1A7t
s7PvpH5yx+9J6LpiNrRzcSLMU0lN7JGZoxfge6sLns9KUXMIf1x7ni2vUtbIp3pszln/1qQUk8HY
LZUEwGtN5Ar21msNKo5Ki7WHKNqf6lKiHKV8EYGy8qkZyTOk5pu6yO2DTDYPsfvVwxR+BjmAfFkT
Z4/VG0PB9lj3fiD4zYB8hO0ixrTnzFlupJbsywAyjmebsifwSfYPN0eOlEg2fFIF/tfJewY+RXge
Spxuk8Tyy5hsFNS0BuOZuW3fNHMFEwk2Ckv1eKUPWww938cSCoI5nCqnVjS9/JpEpw5oP+QH2E3n
rLQZvl2mJyM3J1pjOAnIo4HTP2W39JzyFws/pAXayLGyeOOGI8zW3CfbkjhYz29+DWX4jSDIVSkk
jIzAgvpDLhC8oF46fOCxC5i3XdPD1jRlZconJv8miXHhsLz+91IowgLOFw7BY6tBEgPNjUzg1kjm
lUO4wIM/dfXCp5O30z1MvZ4W0LiW2LHgVlEw8uhsWEylX7leQ5i4TbBC4K4h37viBQ1ohz4aoBTO
QSX8tFmIvyIBeoyxEDUttpLIqhR+8EBEgxd00104HDLUJSsfqA6cE5EsduZ1bPjAXM5U1e5CFMYz
2MhH0U/VpBJGvpQ2wgu1vSmYusGjOo7TppalN1dC/C35lNvOHEjEYlMRaDVHmTQuVpoUbTbuKbaP
fyye7dVK9vERZ7ElRD2A8V2uUmMqj21+fL8s7GcYa67+hUn6vWjURhY0TBPz1ZaT1s2DpETubtbS
gNGVMctu0HPXxbN2tFyBqNTHqg1sUDed/l/TKplFJ/1kFe2xdZ3oT1MbbMk/K6rEQNXK724fK2Fp
M/OXuiRygvDoPWtdBs/d3e4dL2gLDHjMpxbr8732MPNsQ8O4mkYcxeMLJ6jasPH5gQfFeTzNxGKu
b6BYFxBLxqhBdAYG7Ttmhz/9BzYRrPONm5kK6jj+VMIG8DNb5/P3nETZS4oF8/hwxxR2ZjKG45WF
pB6YQGJ/Cr6oq6p9T27DwSF3ymqa81KX7IT7ecF94grXRikKcw1d3aYXF7txWR/ZxTJtxRTHXgyo
yx1kFLamk+UhR+r/7zMs3Q2UkZU7Njf9xIRy89ADm2nR0smgbX8tAU5iPTOvCr2tqHlH6yunjEfZ
VuafADJLMh21nhHk2anE9NLr8gnpIbqefh0lzKs+ZiXDQoVwNF5+qwUKaan2lgsbRrVlYhGZbrF7
/u+nRHuJcT2JZJ/PG8vqa4iNGHjt9Zx8Nkj0bEs8iBdZei0itaJCpfCwJ8W5PAnJmnUqT2GihBwZ
W+tio2E28RyeaqszNAFDBdzezgMtCjRDCeTeFKFU1WUTTYlEtzAJllknzdD7tKk0YZqlHBH86eg6
i+AXotoOB13pMxhC/nButmhXxaQhwJeWWzrAWIwtZg41BK7jIt+VBH+EdxbYEJju3CqPlTAvzlgD
AY/Z7STq/tMq/kM3SVPHSaWr2SC5uVEiYe+crHcbD0cH6niNV1W5oORIXonprue068HNixM0+W4h
V95oA1GiaeBubxl99SsJUWLeJfM58d8FtJ3MGwSenNNVw/V72sjEvPXJPbYp8UCn++cXHN6rO9Mq
+nQaOXS9+srgXUGshCIRJkIGuJR59R0S3fpTvEgEULrwY7UylGPrITzcY9rbGmNJ5azGTTlhtINS
WcZtmppQS8gEuu47kdCTKIpXEeYuq94crYgKzpHYdNXVf2l+fEC2GZsdf1OwDQjIP2yTBxyZHgeg
ZLP81N7MoATxsDRO7iRfVR6VT/Bkki66OYpvBSam2EshfLvdEsIhb4ATtZKUEIl4dz02WS95ibSn
1XpfTeOw2CuC/Iat8q+TYMn0k7BY4W3Cqutv1gvcSDx2P+QLYYuUits5HMkqbWWinKdo61ld0AZu
mi5UN0sc70OfWlR9a5D/v5JoQHRLKOWHGkd8WXHQrSoTw+WmVXqR9a60yIGy5biy28dzldrxftPx
OE55szD0AZIjFNcEdhJo0kAnii1OX94AIDXKZdxdy8rv611FCfH0jLVfRT4zTalM+AXxwe0qZA92
UAmAXTjlo/pzGh7DD7PvxgBd3P60zg3Tcf+KpHVwIaCij6dgwaGkgik2MSUpl1kjldbMUI7ew87v
vwUE9TtIa43/n6No8VOitp3pL91HqFfRqf6LcpWxjMx0Mzfdp3wuC/r7NdQyu0zFMYMy3uF3h5X5
i5oGBJyqwUlO2osQYxGq/g40kOAopXatDkJ28ztmcQyML2oQDwvXhl+Ci1374MP/kNl151OrHvmM
DQ4lO2zYv6tMmWrBwD4serqtjeDmKqmWKcJFAI7Gj0W8hBCBkSkYR4ABm1yIJ9/hZY6ylshUMaUe
3tax065KX8DKlMkLF+DrIMi16jN5rTVejUFglaLn3sxaB4TK2yv+rGIE4hcyWcwb/Jjk933EzvqK
GGo5bLH2GnppHBvS0geeL1Ct6y8ap1ySpgELkdkybHuH5NtaRZPjnekndT0zgHMXDuA8ojOEfF9K
k92J2RFdVuC7Yc6D/EI8xu1dg0Jqby980HJtt5WTDGebUNYg59n6luRFaHDFIzjMoeJVQQTLwgJk
R/tPZ5oDfB/ZwrO7pPaMRE3HowgDVwJWUs1HxLPMRp+yoh5sMNdsG/WpgNsLZBU0khDo80ooSwi6
gyd+DZJqSoDlUUI/iKBggAufLZQjGomvydsYbsAKBK7uYVIa2An8nyY76yoETzLUB91MuuG36vBM
3AjeoV+QydFpzAVDTUDv94HhdGUQvYCpKHjfm7mJwmCPGipHmbNWSYX31jfmvoCc4EtXlCEX+Qhe
JjhN/QQRQx38CUe6Qq5W2u1MnnsNcr8DRyQTgAipy+gDO43SSyNPNMTAA719CXzHOLUhhPG6End4
/9YObk8xBjD/7JOlgp5Q2S3pXwsgOBAODh2sSn+SZI5j5LuPyWg+L5D4fUUmb/hpFskO7Bt7PQ1o
NcT7zfMP8l+EYe3z+slldMrwLTkzdvhFejB7QY62UdoXIXk0+FIgEcTLu1i9gpVx8TQNNKimddFe
qcPOVtidIGKYNsnJREIFrBA54cND5ySh3Aa7s9YtyqgOFng1NAU0sBd4ZopT/z++P9vVfRi9YHFk
KqupsTxBa/c2rQuKuMPUBfMRo4ioV6Q2QpURwOEiG2a/TAlP0lLoN5MnIQ3+ZV7w4962IUS4IoE6
JLNXM+/1TQueraFYP0EHNjrshGWXERTxY6A+LRnHbqSTSkeekprb5+g/xwhDJwf/O28+WyY9cmic
TQtbWR6nurUA9AacGQksrVgUz4xG0PYurQA+KPISs9Ixo8aMRvc8oCg5rxocv5i5oU04neYBncGx
jc+sZZ18bAftiTmJuN7tui0crEbTzNeuvhg6eE265IPfqIvqBbqgiWw+mQRN1OVY37oliAzBl3Wk
hescKvRvsE4OMypGZms7V/5LqLH1szzRL/fEI5ZY9aO37sb6oeNea2tD3zNfAbKkU7kd0IULhglG
B+Gr4tDG/SR6baX1fiRBR4nUMtTJSBWMo4HLjCUuglpuqWITsMUczFHMJw89zzY0no0QAsQoUD+u
mvtjp4uCZk9rZJaaJuSAtzDRZCe+MxTU126DwztsH3YpFnA5wCk21gUoyBt4Mm6o0HHJO/3n7uF8
4YG36CiRX4XIIlTc6jdZXTn6Rf/RyuGc3dLM6tQnfxKA6TeWBZkXo2coX1A+r9jW0TItzmxS3y2C
xphFbvZyZ4u7b8YKyKWItXFE/S7S0/c5mXbKlhA/Cfu/3YT6drrFlpD6lEDfN6tQvEn+tEjgN0Ly
Np1K4nxtS7SWvJG2x8ZYXdkSgVTL00/Hq/Yd3g1DYAkU3bkkEEKSEnuArsK9BGpF1y2Cl6/m8i8t
MwDzqG3o+1NexNHHMX8VvcZcjtzlgLkm4KzJTE79IEP1iZWz1DZ3YOoQa5wqePpuM2m3/RU9noMz
XlzSaE+DN0QkDDJvyHkXZwx6vVxDy9amM3uX1Nnrk0C7fHNCctXrG/RWGnrh07mSTdHmzB6MB2T/
K2kQT1IPh1M4ab8aTeav2np7RTqNdOE/15p5XPtOA6zmGlAVDfXpiiAt7G4iQnuj7Oh65cu3Uk2g
OT9IeIyPDwwq2E30C1j8AmezpfRnyzQfvU5PjyO2LuaK2FRic80pIcfqzGI3Jc2hVZdykVZyTUpy
ZGLlu6kiC+GN++2w6YWT35aCNQ0d0hgvUUZGdYhCd1QUyWAadfCMYS+/vjA1LeVfIBFBrWDwGyyS
msBsO5QOmaQphmVhdHUILTnaIvac6IWGOex6EwwCqgaUZBnsftuiSTf+2H1KATc94OfLFzwmi5LL
iIu+kyrrVJAGGmZbkM843Xkyjsxkm9Fy3dCvbmvBTesH4+p+aLKZVHa3s5g7YbZAX0GqKGUaXUbm
qqnb7f5OxeltD+7RuV41QeLp+CeTQQi8AI3B8a33QXaMPOjZSOlZWiNZ5CwnJOi292wcOzcl+LGh
PzFHN+y+l6/1BQ6DcYUgAt+Z/oVDhu07eBY++f3Phb77iiVDKjZtm9+L8yQaW/EWZdfBqaiI7+MS
N5lbKbtfQVFqw8HbWolHJYN3Rk9zHhgCFUEeKr4qtUMcCsu0wTXaAUOfMKE9Y2al6IEitSh/AmeK
38e9B2BoAYWytaRtQddHb/v2kaWWM4lCat47XRdUrJCZnQ5oK1E+Nbqw5enry9uAbH7aeAFDrBbZ
TdST1/yiP+XHiRzaCphP1qZ9usGQ+l2sHuj9kEcT4XIW6HaBNp+dF/aNTNOzmdDkdg6I7C3v/sKH
zVizXryRCYN3KzJIz0lIcAr3hvKo6bQ/U82wjMYL64QIBuqkuCfJLk19+zh5rdaCMA2YdyxU3zpC
3N4S7VhqiwT+Jg9i5BPn/w7XyZgRppZ6Um+yZDwQo1MtwFcgsdKwXFKYGMlPJxFvrRKUvDpsBPrL
w0t4yyOIfUUNII4KOeoQwe5vlGbeUrEEp9gDaQU5uDeRHBtdor45HWLucpYEQruCFHJerqjnlMWR
McCyzrJVOwSx/KILzOy3TnT7DuNqU7Mj+ly8MVJw8lx24P5YfK6VtrWae9vMaaSnCpBUtpAwvG4p
s1PevN4qIp2a6Mrry3IXUtyh8uuNWOqCbPLRZC4UqXwIItK4hkCRjBTF3SBDVWf5MXhgxamubton
bqqbqF0QYZy+GOE4OhIUs3KT8NMpbN9vwWpHKmxiar8iC90668i1scLkv3Y0aUv40sFqbGilc2oK
Hjrc2RBOfwviffk2Dtu0G0l6syQ4wa/UE24UT9FJiLpZWUIs2E3N2cYw1G/Qn5IWw1UygZxlsbAK
9T19tCA8jStWuTgzGteJOSczO5j70wQkJ4Rfl69zTMOT7y+rkm6Wz+Fr7OgzkagPUY56xHPY8isS
+Mxs3/txfVBqeoYSJLZegJLH8hHCh/0WGnsEK4NGtAUv0fb6Sm7Lnc3yJdl37B4kLMqZTIT+sl3V
OWrxJb8gBUe4YV7oOx08UayFKHXBEtT3Gn2hITgBuitYM35j698BhSJzJmt22+3SrWvZs91wdl15
ZWRjtt72C1WQRYOx5ZwLFOS7X4qmYjT9eCn9Md5XqyN9qE6+4M9ztLtGsMz8brGY9c+bTaAjjqdH
f9eOfqDTmrzTr6alRt45BnjFRkkwnLTteQqClgVm86fhCY/02HiPNgoxsFMGhZJkegsGzTS+fost
A1hgeptvvmhh9bHQ1bCmvV6RuBIQZQ1qAARCmvMIuRld370myiYVGq8ya9nPrVqXsje+EDMmtRvL
SVYfnmtJkZBQdaWv2rwdoPqGpeeFamTIhaS+pMvL1QLn5h8kJgvT5l1610A8rNQVLlce3djks9nm
kp5njEhG58Yn5/NHqGVuO9d9T/wuMOKUGr6sWgJi/sIJ6J2WBqk9iCC3o7yPkdOOBMl+nwtyqdpW
4Tf7HeaQ/2TKm+I5iqoAsTE0G2cbKLPrh457cC4BFfPgpip9Rnay8Cj/gmlOraMvArRP2TxY3eSy
yIEFzI6VKyHAoXzYUOgIAdRie749ROdmo8eMMTEi030JKEE/tJNf7gnCzjKxikVgoS1fPsidYBoz
qIbeJ/ab0z95pHLGc+r/nKpoKdzzubDvhU14ZwDcRl1ioVjwifAbYBkHR+Z86ipcLvvqojDDa/F6
RtVdT0VCfksEqgT8f55R4Hc0Ngc2RmxQ/rvDa29yfqb0l1kwtfK2/p4kt/2ASVKMZK9mdheQy3nE
vRJW1z7PtsWYsPOZ57Axz3akmgRPoNV7xrmBbW23a7lCxGc7q7BiRKsCFuVhcgmuIngw1ZcKHgFD
t3s8QuKipLItKqiqf4m8ZMWLy4X4l6UipZ+EoMdHf+KgpaZKTd7TxwLQ/F7WMDHdk3oO4DqGXqvX
/OMM5SzedWdMNcvs8sOWSrJuTYLGWC8yhsBEfINL4XEdntLG7I9oYSdUClMlH+qhNRVLoXoQQVzi
TmE4P5LPQjPISdnglNyQXxhufYVo9X2oVSFi8HaOeAHckD/omNQ3vYNcMj887VaGmWgS6PazCBwd
kaO2aGte9IIHUL0GwTeQ+qRJQd1E6nXxBmTRangPRQQB5LTboLIpG58Iy3eYsXvzlGCBZfX0yirs
xsmo1IcwzsALVkczwcryPArI2yfJE+tsPD3xtrjq/J4ZAi9aFrEYAN1eP/smdYCqtkl8qyEJ6LwD
kt/PNSkaIe/TO4U+BSXxKGES8PJCrduwsb2cHWKUEEqNrCTlo/Zm8AtYT3D2YU4qpzXufyYOt0c0
vBa7AkTiq4wSdItUJfkXHz6KgYKQmw8r13NetLWPBqeJWGRC39EuMFxUOuUlAV9NSN0q+sTqEa6J
5EmGfD40MxS/72Obi9KCyubVrP+wZ6ZQst8GxxCQKV2sPC1GwiwIFv8uBhh0iGPJWx/uaeGQrupJ
L4ZNaa4XqFMsJ1PiG/ezGoKMloYxFWWBhMjb6XOVxaDT0or/ZuKlj+49WVP/KYU12FRkL7ox9c+C
SpnUsKv/ec1Py8gY9CMRszYEjUb+i9hzR/yfg88UcubXubz3UgXDbfi2Nfl+KbT8GhQm+f09LZSa
0Kk1mitY37CM9aIIzQZxaBcTNcgiZCRGbO/A0bZxJUhBt3G7M/l+i3uy1/VV3v8Ok23k5In544M0
3limvCvMCJOp421NZlT3a2aQVNgqmfqAP8/YtEXml8OsGj3RZQHYjhNoDI9gBV5uKqVia3zdfym4
hxkhZqOTIlVysj+Tz+4FD60Wvr5P8UMpD1DnQpVTe7ZQmGfzCYz30+b5rDy2hq31PlrufvxfamqO
5hlHTDIeqMadTqkj5FmjkeqstFaqpt2VuWpeWfmUdE4WoCGX6zwjtUZpcgTrJUnMhWd5H6rbhpzG
y4dD3CEiKwO2rzkbOu1lAh+SJ8L20GDdZ0MlSIsYyXGKDL5XFbNUqsJtqpvFTGiNZr5IwWqBGdjg
4CB1Fqu7NopA860d2pbVwjqpLnWarHhSavJahAHmFOexrA5bIzwtvlJ361X7sq5c3ZFIizwGAIUv
1h6QUjgNxlO3/UZ/Eaeyqd5tDooGXU+UNf+ctaNjn33ldnS5qxWt4RA+BDZvx5t6uMIlWwdtqSUi
3fHnNMUrxtjiu8/wNnSnR3bJkTI/2TaytG1F4guB8LVxYt5EuKtkEZlTokZbRAlibCr3gCSbJxcw
dvraqjMW5Thd2wHUh1uGvrZNHElUm5AWdqzaxop2DsrLymyPFrJgbxfcJJXLmNbvc6MG8F6y/sCo
z6srMASOb1Ne+FyuU2mPUwnrbfB2jI2MRuzZfw8Ro4wCmLbsAnWun+k2NGGHIE8r+NHiwOENvNMq
U3NtUu7HPlQPD25uodMV2+vFGiG5DnNnd2kyvO5qsGF1wt8wycyJF47LiTLmerV2IilxTAqAsWk0
FNuoUnZjrVxuVEg1cMQchOQfzJ2hY/jHJPzopLEicrQxxiGXRNQSR1i/cYbx582FqdpBRw7tD+dv
hOT//X90Pa6b0vktsloCGPbHF/Rb5lpWQoJKmtCh82tdp7Y9GqHTaHACABkCFgko4uT5z3n6tji5
4HhZwByuJ+KtbSxDJwo8dUeF2Q9y5JzNH9U6IqFPR1ltLKPgAFHoocNMTPNkQvvHFH6rkwQYJ20u
U5Oqu8aQmEnN9j7trxoEX7iKw1MS7Zkl1GhcqaGs6YGtHQcWGkec3dRVK170valRACEQ5dNNFCJR
Bvl7mEGc9zGWfui6/ZxOPqKKYv2+Z3XW5IDMxZcDdSLLvaejJ1SERKRjQmTcAJeWXHPeOsRBoi6V
hsbQrgPAwaTd5PUuJjbMw+UAZtfNNGniPAAGuWxxFzXp/1oqJR+HQ1a6hEoc5+dVq/5Ldvelylxy
4t4iOMlLaaHMHqq0tNrR52tfjVMqTnl+W/Pi2rLKAfl82MJW56+R7v5lfpXGjmMXbh2dLnu7pZul
FV2qHOWefGD7cCJM5XKgFZkulgdOg/E2ADBEH4ddGwVXhSNoNjGSDu9a1e5Bqn0HcMwcPQSYPz/E
ejyIwR+8xl/r39HT+zJ3PMJc4hNkpyQXEyvnOvp7xjFZF7WP1fF/w+XDnCCvaY19vP/x63EDhs0b
vmnqRVW8k6BKKfZ59oLhQIxigW1pQttKlmHV9WQuuD06kZZiRZBEBF5xhcoaFanAA+a+3XoRhGUM
m4+7JkMhaGZokA9GmODgYxTqsD8wBr1lg98mMX5JC+N5Xk/Il2hpyIoZY/ucJRo0lrpTcx9AV8D/
j7nU4FLmO1EW4aGOpTHuH0aQYydheg5S/0nTe5jGStDcVYzHPrQqIwzmwdBKJSfmvTg9OkipZ/ye
J7Qhs166oH9SfAZOsDnOowQhxJYs2gEbmyeB5R0jpCK1OWcdlfgVjcZTKECLt6J+bT911Ok/0Fno
tRogkK18NRyQ4cdBNDdkjoiC4IsqFZZ/cZgkgjmdFXPGhe7VusxzGrxPltXHsRSQkLN+ebng4Cwt
KovfOORLxuS/nsl5a8dNwblal6KCWLn1+ZAcPENV96W8N0ELrKnQCWf0RbdlGYJpf490QJXdMsaY
Y4v+qKxnVLwewDsaO6WzUQlnL5/9VHU2eKK2QQv6SiNm7qhPfF/8ruXTC9oXPZIIvXZOuT9Zrn7O
HfL+F5yoh1FEkgUbXZ2nnR0Rq+4F77UuMrxCN3G7sRkQ/qFS3XVLrNOIuwxd9B+C4/qkvoFNMiuS
6UGBSfFgVgji9xJlPNzJmPfm6Z7Lu0oR72mwOztWaunedsjL4n1UuAZv4ghoAurfxdWkFuwF8Fja
r1PEzMRZODdhQg6vyaS2PN5b7YmMqSDhuR0Fk2+2hcSwaE+HJ/3gBl6nAUnV3v9iAFvnJNsp1HY0
t1U+gmtoMwCq6eifX0Q3gsmp/J0p0UdFquFZ7KRiJrgrdGcdpenQyTdYqQVQJK2N1paCE0DweEV3
63yJMpKSpcfU6EQXjrd6ev9DRK+SIPKm2QM77jeG4lTbMirz4tqhRWlYs3tdaix5dr+u3nNew31l
kemsySlvibG/5sJNHhABflr6YTYWBvOZitY5sWz6YlGUcS67Ea8lYLFIXk7kYr5zmboFCUF1SgUr
+wGgkcQgxvR9/Q2+up07CWmuPnhf/3Y0g/JCE4qw0C9QwOPTHVhdDsUNX9gbUcNT/RaX4dugMqgl
waFjMQmxoavdFtj1x6rRzBLvrizrSctfa1FU5qZdnX8yPHvOTonZN5bFSbTdlh3HJ8NAUioGe294
I23Q7esF7jKvQEYBm7/VVkphVlaMjG3ZtNxTWpHDLJR5FRqdvOOOe/5m57cNbRCURZvPzOeWJUB+
qIAyAONmyqYh8CpVxcjAeg08Fz/B6sT7fS6M31zffdTdZoHNeevQqaFqYd5ZLqr/9UcDSePG5bZo
4/iQdlDcvyxwKKoRsx6BCAqpQy8UL3hb09wZmWWw4xRttisrqdi7yUa+ISDhluiFWIvhqebd9m+P
lTWLfVCqFn5zrjpGIsa38Umm8bW3dIHXs81djbYQwrsQNH3pG6DkXAvhXjvoNOyBHkazK2BUi32U
j2yJo+Pdu+UpIhWp+VWnnm58bu+0esWwPv2pK3EX66Nv9qsOCWp5NyFYu9qkh6TtIS9gJU3WdZCC
k6itLbr4INbaoYgQt1Ew/+8iaqCpbscLUPbLlUWcqo+6gxCKkbZNDbSVIz1tu5pTmJ64RE0guQZK
8fmhfmITUyi3P+Tg2pqv2Rxy5vjIj/ckeJ88n5iC0HcogiMC0i2i3Q42xtKDCMrzecKr8quZI5dr
7kX8EYMmSMxh1vEy93hCXK5guKPOncdzBwLSJfESIsigay/RmiZgGUwAC3hy+K6iSFQaJicro1sz
hL9pzNtdF6Pupafiy7tMN74UU3m1C1mSkybx0I2YxXjMgguHQpT9y9onENzaeaLNgOzjDsM/4Qzl
hekisP6VfFCUmmWYMkdhiIVh8ej2kBTY7U8/Ged51I2VhjNvVrgVRSfAnwrSykspUcR0eaCfjuGE
q0HmLUrFukw+pJYg6rq7IqkzO6ZWLxFpksaLZ2Q3b2l4wKRA6bRXxra3G6Mbl6f2gTUVTLzB7W+W
HEYgA5rKKVpU0R3kkaS8ZYtCpdDSemaN6wFDgCRAXciFaynjx1SGVLfi6Wh4HtJQHKBFJODOhCfk
bPyaVzUm0aBdPVC+R5ODYHGMJOf0F7zY4nUw9zKYvsUA34KzW2y+woJ71lMRuRzf2E5i6V/4/viu
agQAYC5tHKqaOoBEYCVTGXG+IsgP+poXKgFBgYxoLsPvKYloVLFdCB9eBZNPCA3QNaWpOuI49Efr
DHxyD6z4c/iR0Jo2CKbheIkUAVI/P0gZRcD4NiL7rzLX/6Zi8LOIqb4gkjCrNTKrxYJMk3/uXZql
ihPQ2cTDBgvX3534sLuZzkoXdyOJC6pHHifKrSpiC8vQ/q3RyhMHBeRLjTiIv6PZC/WOv9o1L6pR
RNv8n+cdrqwNNRZ0eKc2r2K3Tj/LVPQmo8dxT7tKZLTN8rMUgftS0mHSy7V8dhON2nyYyfEf+dJk
pzMayqf2qaml+kCrQGpzEc94eWNaspWX5urv4TnS4/lB2AlhHOjgOf1z4t3RRJX0zYfIU9HMb9EZ
AU97r8m+OBBSJgikwoPwaXIDznXaTexlHu+cWJPHYa7AOWOqr6pPYSZSYOFfZfUyk3vWpaV/Feyn
FPKb+xyVAD8JVuUZBXkjAPo/MWP1oEYIFsqNZ3Zasx3E49vXiNFkumtpexoKGlDnIvpIJS5Ciddl
a4pAV6CWHYiqfokN8qHSV8oU60RU85Lv5iboB/YM17bUqTYItnSnOJVRvSxpioKswHqdZE1gnB8t
B4JChBDUSQ79tIbdkWBP1vdxxfoljWGL1kMjw43zxZTCrE8Zn1AAZEkpeQtYAZwdVE2FPVnXZwqC
OaHhC4VSqmY7gFWQBI/ODKutedbqsqViAr/HzaMyFZIqMKFNzPP2m+ZivcqwngUjsjQUe3BsfcVa
jjHeB2vZZJccy4MRHy3op8C6AWet5Zjw9ld6nsymEARsR3bJ+Y/HQL+wBuQnl5NYLYHb8dZDmV02
rW59TKuDskZXVnz9nIrC3z2VxAOxL8MdWy2ViBv66uCUoaBNVQsdM0OygylsWQJ7lweWIHAEDPbq
aqfP0/Dw+iBunaOw3QjMSIoQb2T1ROzU7ZJ7yGjmu+wgSF3kO6xjqu2BAmCQzxHtnt2s6LRwU6dQ
2eRmxPI56THYWY+3WcE0e1q4K0VuAVewrGCGpF1b4T8vKo0RlZyUA7LkDT6+DS7MspGKMuhusmaC
L7i7PJwJruTN8cp9jxJzv0kwYjssZk+lZgdu3nUCTVX/koLphhvcP3B5Ztg4getBWnErp7bG/TYR
dPOfvGESNFR+Ful7wDzvJvS1KhipJq8ts7sY0rvlN2F+fatBwdLzbdqyxkIpbyBY4T6p7mVnbm+L
b11HDiLd21L1FwYRk+JiR9sf+HrykRKc5NCms452ObsBORJAu+nMnh5gmOo9ARbaU/x3HBouVJK9
1ilcnYcMV1Ul/HvIW0vO0t0HOUHnCj/eRjCLrmgQ0CBBwuZwFtptA4dK2MMDCh7dFevVxgSDMYkV
oXJp5ka3h5eDJje8FEjvleqwgUg9P1YySj4E58mwhr8Kieol6wFT2Yqqyj5OPssm0o8nox6apkhe
7FVvSrQPVw2Xf7nns64W51NAQIOFiAEhVxvva3L5K4UNbOua4Z5H4oWMw9cEf0uVocOundVdmKTC
bZksWrcxgayjz8bkomwUdHrjfIyd/ha20EYIsPU+G7UUQ2XZWxlhqJHZcbOT4brzOD5aQJuEyFFp
n89tuhKLTkbTwDwY4ZXhna55ZN86a9C3+vUty4nHdoR3l6QeF+N5/tadYHsnnd9beyYQQYh4oq5T
CG9n8IZqErx1D4uC8c46qi1WW0DQaCfheVulnGHWbSK+biPeDFbdhSK1kP0mGRI5TOwtmEEWsZx1
SXn9o+op9/bB92BRm2KNS6xMFcvSZI94pgXGQKb0h05/zSdQLzS3Bn/R7SPHE9SUCQsteIK5JwID
YZABFP1eakyfJCw6WeoaV2HMNQdo+wdwVO4s6mF38ssH+pkyPhC9wxo7XzUNS/DYYt1cIONZ1QNA
yTC2cohIBu1t8MnDpIbziDQhQUT/7yuPvfpWcKeS3jt8y9R/BahLgGp1k6Y+CNsu1T1qB4k2tcaQ
DUmUpiwsxSUeMw7VxnZnrs4k7miWhqVr2Z7myzR8Ap/Wbi/NNU/ECc/MVlB89Q1VYE7q1EoqSsWR
lT140XqGi3mo7JQ5aT/P3dpi+EymBQTGTZWEJQxJsx6TDT4dfkUJADJ/9kRkpvRjFNyE9jq2nMrI
Rr2UyRjwWWl8UwBaYqLZ2ecCFC7sR4MIqW8c04hU82SH43/L44MuJrvBbj63FIb1+U21ne3UZWBI
yBux87BAODwFIcbgXsrJc9N0epjlPDKBRwPNuu2ew8/slmNuqDRs4ER9G8FLZRtTzxpDrAoxMeGI
BOJ8gAKtFn4NQVYNYPBWf4GAZlI4Sn1Uu8asU1rcbVgNGdV3Bvb5OXPiy35CSlGodL9g+/OLXXqM
U3MK3g2d7moepAp3P69y3IzlV1UGqxH93xLZTqIbQbPhTF3YhyaJ4McVcGvQ5aTzha2cLvxRqajB
lOkDHRslel+LNbWK3hDRHvUYGedy6yNw3FX1WFqDucEvryDN2eRqNOqAlbkOfhww1B3+qb4sUYBx
pkjmL8JrATIOYe6ko7WNuRiPWZHicAQVNF8obsVfB0at04paJ7ct2vvYb5ARirmFQfwY4rVG1bRL
Fs7YDRYsS2DYkTsfx8+XEaFvb5D9lXVhCD5ArdCqH/67/uSCBKng7L3ccvfuuRiEP3HnFZDLxgVU
juyYjnOSLB9C+dy3wFoL8HGMGONHHDoRlTSxCXe34ot+MwT/PYg5RJ7nRStyVlfWCqbq1Ku6pF+L
T2Es+3bY6Z/bPavb2eH2PY1vobe26rfnJRtbx2x4HC2x8F60hJex5sV/hsbr+QJRUdrf9CXOT28O
tNuMEuyet/sFciyB+ci9J0XqJO8Xw4jhQEhV+wS78s02F9jL+4ZxzE+7+lsPM04bSQUZptwYR3Hb
ZkxUGdToyt/CfP2wBsZJyXQg/mBJViGndl095bBf1W1av/WgrGZoUOjCkwi4fgJelUxXHVMAgDHx
ayFg8fzkDpeaUSMT4nxMUioaOHmzzDe5B0f4Dv1rJgHoP2Bcvnyxf+NG/mlQzOm9vP1MwsVNLoU+
Qt8+XvQL7L6Rg71XsjHwWzLx0fadrARdc3XdHgaUjmOvSk4IJXXkor04weHSxgEDl7HGnyYnWN5l
qFf1NLx4Ui34TFUsQJV26yi6tYRHBB/9cjR4yb3Blozxj6ulokqqfKVYZq5oxo9TApBAKbHOL9Va
T3Se02kFBsYlgdhiftNO0/lJJRkPuG8AX8dN7T1H8znk6pKBCnndTH5tzkx0VL7EZjL1jwpANKF9
vuo+e2Cf8RmIGwQJxa1Jna7ECIN+bjc4tKIZDmpOk0gKofwEJcmsijwiw5+VZqbhiZZvf3rg316j
JsfbR6tFA9F2vOx3nJ1Oo4q1DuNQD0BmaoZCQZi5OGeyqLqvMQUZ4z8mcPijPbRmbRzhU/OPDy4W
t3kmmFC67AmcbG/Oxa/Sxk4Oyvqs/3V1CwQKHFfbv8GN2LhFpveyY3qlKu/ws5kJi5LVq7wnvFMN
hyOZL4AT62mF+Cn+FrKBHAPjuAvQfsyVDiyBxQgMyZRVv9uW5DEozqZBMmylOkOjblLBKFnYkpv8
qvh8RKB1mdGa6Yvzx/6cfGfNwEdbraLedSrVEUxrpW8/KJKqPgXpGiQduDZDsTm5rbb6BPixjoY4
PxsGfG1WEHapoW8JZ+DuHssdophuCVJI38h2zeYf3NLLwmIAyZWk7TvCHvMTOLhNPoR2twS/bfAb
pDiEpr+feAT9uqIKRj+syB+72GAO3l6aWCvfbFxlgC1GgKBRCfaXfApd2Gz7wVwag2rszLQKKS1T
lFc4qw/UwvNBoNZdqA+18U8tulsZtl1nmmuoJSI4v4Y9wJ+CsoEKL1LBBw76nZMRWCxda7zjqMFK
SbnNZmjYMrM+djyhC2gVuyN2n/DeurjE+AE4DD0ZC1pYLtseqpaaEjOfGe5BnfE2VMI8Y3mco/Cj
lblzWQBC5qJSQidEiTX4YFBMwRdiSpcrLii+FlrDToy91X9L3P01QeAWLbyRgNxHMw7nh6BktO/5
+6jGNmhK/pYdV3fa2D6cKgoypw8z+tbjbqoGhEtbH3E2S/c1fdyiOYk5iqHj6HFJZUukA7tnCyaY
gqO+2+Intmb1a/xfPPl1Q7iJhxM3YL+V9laXwy5+6OG7EBFE8FnULqNYBnqICP8QFteFi7kSkCAK
LYgpFC1SiixarQHLiCHzzWodKUxejxXf7vQxaY6WJYad8hh02chVWUA3xo5M+4vMK0GGZl6J3Y/4
SPxEi7KXzpTPyRAdK+TaYLxVVBKHi5kVkawQTWJmrZaBUr8oCMYg4HQpnTu43i/Ld0JRjkSORTAv
37vJEjth635R6wjrQUz2RrRVL9yBzgYf75Q0jVP2yyFrnpV1R6hNfDCau065Fl/cDzv9hBFYtnAo
Vr2qXME/5y5nOo7EfbJQBJVnKdLYYa87OktWT7vB6azVz/FF2P6EewQKRNfbSdakRA/bq9oW+Zua
WVbZybM9GecDwMcCZjQ5fcx8gewoykqu4iMpCsSgW0utgW9WLjMZGTAfiPjT4r9+pta+Ln4r4BuY
Lq9X7VdcoeQTcpw5cLpRMsJzvC5F4D0kz3KO6FAVs+b5mB3x+sqyhAa2FBZoD/ivYNHXI8OrgBOx
4E+BaARxVJylrylHemIsTILWiYR4OQ9IqpOkCbf5xPzpdyZt7Oz5R474Y5YbfchC1MqgKpLdn5X2
Klac5i1SQ3eHf1kiF2k7ZXxWjUpL4agIgcCukyktpUHoy4u4aOLHuc4jBfBr8uSTQyTjKSAOyqi5
cpTjDWZUMQBVwfZ5RyUdejtxkTnHf5//v4CzqMlBwghpB6yzSgnNI83vwwMcaEU5byOqng70mwAQ
FhB/D97F8Sg3I231yaKUhbHA3w07aBD7mcK0WyBuRpwkvc2pnpbuFIVpvqguPu+fX+6XcFEdqIFe
6h8IKN1asSwoSgxKcl7m1NarkV9Og28RgTwezYqR8n8UTHPYoERJ18YqN/9WFUS8NacEb00Sc1hU
OdjlgUAq3cGoOcUkbgHK4S+r1ZzbuP0vuUUzrphLkJRB5zLXMzA56ogwMWZID96B1gbKJ+kroPQH
d340bOs4fVCdRhe6wF+6pgjdKiqcVlnnDDaleDdZ9/PsOt5hTLbcrouCaK7j2F+N77miLZ6QIWuc
PZo0GB2xBZ2nzZtsZ9ujOGzFrOtV67VdUNOEmxAPqmBVwfIGepET42lIIjux5xiaWioe4QuuvK2y
9aGUF/3N4E0WLc9OoHpqtT+RIkoE0va0eelNQqtMmzJPF23W2y9P7iPhmfQOTo9275bX21SVr3ii
TL4L5NfIqj87qDUWIsujtuwCv9zeAmypXQVte83fQAKtKRhtng3I8Bv3dDPqRe42Mmt52FPk4xdI
h55WI22UhFKP8UuKK2Zh8Wi0G73A0eEKVLrBin35yxOBBVLgb9qVSOSSi7QKp8fngelUkkw+/FJG
3IS3cZvZHXSZHvqLpHua6+vB4A9ybWpiogIlGfh8OiV5s5xeKSLKNkZGkg38JJskZjl8u/TWurgc
CAoPpn5cgaTw1P4byuy1orNpcBIZIiwxGclf1BhxB8/fRv6DBzsSh6IgjE4aSDj+9MJJIeTSBo6F
wNCghNONqfAXaxO9GvRYoZbHrl4nV3v3PgUuYE0mmwRM4eOnkzKEs/OMHoDVTyjfKHK+En91Pbrv
xLHlYmV67bQDRgCbpGFrz+aI+6Tf7nX6z+69+/q+C5mUopzjTHRlXwuNdxgq8nG5/7G10IO1Slrv
Hf1Cs6PPRdMSAL/HEVKq3QaYixbYq8H07q5SHqCc6PUg5LyRgPUv96yd6OIcWgcMJLUqmtNePmBx
mC+SN/yeB1q94pJKNNfF3ClPZL6YTK5VcQX/KyKAdlH1jxv6EStbzfMZyN+J1ko6hPoDlJl58ASK
0AIhYWs4mQE5nt43gGJDmhqaxUSm3x4Kyerl+4i74QUmZ9uhR9aGPVggwCUrkoT19XLcI0+wU0sU
TLEO6zxKsNA4QVnnZGH7Rb/K5xJQ4uuvAmesnauTkKSP8lFy+PFiVVJwNXbFGXxbpBFsc69UMpF9
gjvqmZiIC0ybSS9Rw/v/i76xp9aA/ZQ8bSY74dNZq4KtPs1DHwRPgTgRPxlSRvZnvSM8C6u50TuJ
tmRlB0WQxPjCB9TMUsQqIvu4LuM2PbDmp76fDC2gzcn46wLO0x4dHcno7w1K8EDHk0LRTKn2qf0e
CmQjmIIrwr8B+XEgvsZYx8xSrtKvSMMvyu6zbCHJGHg/MiPv6mkS9cuR/28ANfJBns84U5UwqIvv
s6cc7jQuhJ8wQ6J2bcZv9lt5zd402CoMqibiLK89W+0sblQ/AM0U3amChATGNnbPvze5bxNzqCB2
Egxjw3gzh8wCK8jKkAAm28HSyZ+WJTL2wJMQulq+oA8b2g1SCi3m09TLaqL8EHuJ9Lm/Dqqqahwy
QOa+KeME/if391VHj6BNCHSKjw0eCgRfvACb/1m6NhxMwAthZOTRc4gK12tg2F+7rs+xPBXaf/AC
0anprf+Vyu5X1vEBHgk0nUr00x+OUX4UBZ3s+KxLxEOyGQtOyyaih34DIgNYAJOfn9EG7GSkGnC1
DMvI7yLW+5vt5Dqf072jhpn3TkYMjlkcVdPk2QOzUXItRa9AWaJQll0kLHeg6FD6Ehd7G8cOYjFb
9Yf3+/pYarqLzLmVzC2Yg233UhqbgZ3ClHtnWK1znJocF3G/Xveg8fDQulanP9kaW0SZYkbFdgeI
AXwC9FtLONrbntzb+/xJJ/9JDDihMOg8hMQUVlRQAe64KAHLz5r05kYDqKHQ5MvKsg9acytLqTzU
I7DcNICbgrecqxvpC93/wrUfeDjDr+ak1E4QC7T8RcngT0fX++ffLsPPv2xoO8b6AJ69RToQsXh2
7XcziRLLg7ZaPpw1YeBuP5uOL9qs4uLkI12YMZAVd617EXErFMmDFeF9xN6SnVfuIk7uvbN5Fkim
ltQLhTHr5yiOfOw5ZcdCDe6OrX9fVLiKIBBF3iDesDQWzbYNkKvEDHOguTJr+cDpqWOJIIptetmi
xnifPdVtLrYiw9OyQSFQnSKE/4+8oIrOVVRd+UkUc2wVXSRMFVMexj5/bvEHHS0NQ0bYQ+8Bor7g
HJg2VylFhhOlvAvUd8bteGwWdHE3TBZZY4fKtm0zrLkxR00S7Rqh3+TgRi1Y4VygsWGzMO2peUHq
l83TRNJmn+eOgeROmQ4sI6BzfkkX2D1ICEM2asjPpu6iesdjyzXfFcUin3HnWujTI7oniqcrCrn/
GRtcsJWDgkAWrGx+EJQwruCcUBki8FEjZv1JvnkYn/xZJAO4YqLack7mlzcCWEAAA+z8F0sA4A1K
rqExLngryqTpwajvBTlQvODi3Z5eL+IO48wjSy11IUIAwxjAXITnACWVbyW87W/swSgLk3/wex9D
NbFmoBXnfdW+XLuP+B2S5o4P6B9p6Tj38dyQWwsHGPi2YvxfmPsGqUAfeJA+DzXfyj2RyuwY0pr7
QOoCzDsJEOhD/uiTATKJlmOKjNgUJZUKQFOB/8I7r/rpURrbeczI0/XkraSrMYtPLI6dkpErWi4M
w7FTMKR6kxSB5rvytaTiAACd+leWMv2ZarVEDCf+UnB/yJAKgQ+ru30CdsrfHpf1lYH3K8DFfdbz
cF4XmH2TgL+5Tmb66atEebhDy9Gk8yq2pA8a4vgaYU3yocLWsB1rWw7b0/4aT8IfJWt2LdUnwwTT
idvvV26aJfvdKLCityVIfEvP2TSylXtpZBY4UEvWxLRpW8Pci9cjxNv3brqX4sN3JQDmwlPbIa8c
WqMYcblYXH9RQK5Y9hJWsdpdq/Ebczb+NbMVZ9akkN3Mzkrr4bwnnCoRwtgkmqQOOzCeeTP2GDO2
LkT84M+dK+SormG1DGziloDtsQv2iQ4Hn6lQoDngC1Rx4I9vpwh7xpmssR9UG1UiUR3ZO5PcI7FO
g6FGy539lgjx2Arx/PDTHBf/wGATRlk05LO8tpUXAFkN4iAcrDaF692yU5pkMCAzoQ4e6kNhIaro
+QEFvmtiQap7H/jhHyuji6Ewx/xe9DOLMEZlF0AL/AkvxcZMHi6eMJh8bfYftD8VwnSNIh3M3a1o
frD6vQVcRVkCSk3PzMuNUGi8yF8vjNUHR1r8rvFRLStl5fjJjIcfMCC2JVEr2b465SL9zyQOuSns
F1/D2hbBs5bVhXIaWG+OLwuNuZEpNmq0paLLdodLMhbHmv4MNycYaKwo2YaZmMkOT40kkvLNhlew
R8dkueWKBQxWfZhQKyied+0KuyX9qNeLPi26JVPh+rLRwGhvnun5FwyCKWZEsR0USEtM+XjKKn5g
7/3djRrJHjAoJISB8eCSR0djLHouLtoFrYN1bRIfHI3EA/qznaCuaSdovRotweJRdO8nOWEb+0Fp
3O0SoAub5EF48hSBxJYsXW9s55Wu+fzOEt0ttcll7eL+uiaQVcw4/mHeZXNmZq/0oREwpvVRnlPp
ugj+SKRIwoKK1vZrZPbMBP4lfyDCo3IgVut36W/ArrSbzrj5bY49E5rogSL8eWi4SuefreC/U/1O
Huo0y6hJUmfll8sc/Z/vxOXjn9j4/g9VIKIurN+W3VzDC5BBjULtMdsq9A/Jkrqi9cecbBUAu7HO
iDsl2C4HfbV9Gp2iqyDuUh3u+e6bcb/Rk06QcvsKlmWyZWgpPTBFsjr2RtDOKWrYUdtL/meawPBr
i6uLyeUQ2o+Mtzu+0qWir7ZDDST8o+or5S9UuupX4maawrpDkUZHONoMu9NWO1PIzVQqUOU9YsNA
mXwfl7pjTU3x8iKefoIVWA7PHtRFRJCm7hLCAtIaVQ8zOuc4okb76HmJUzF+GIhUYFHvUbT6QWYX
1MBMbX5kHg50L8MT4c/ruAhenRTJ/Ecrn/Z/s4j5aivrWb6trBILdZdQAEXV3x3pwQ7ncyRrAPNZ
0Kw5H/R1KMg/8WblSZU8Quia1ge67spMKf/DlItXXHuUki4XmeKfwJaZidUdWvSWIQFbpetOd3tg
ylcqCRc0wgOT386me7KUV48I3cII1UKcQdrqkMogd7gRySbKd6xeLSvgp8qLYrTqO1+505Z2GWKu
ikQ0ptmohmOvBcGfCZudHn+f9fd6pnsOkY42Y6S5JtCj+gJVSxa8a5shJVLo1hZVolJ78yKew0di
mOCQWBFqzSpvrKx7jxB+rXUveaauyRD0Dwdw5om+qmbA4ciKXct3famhqHSQkXGrOFQDHqFOJqz2
/VXznGdB58IetGfFi/KE7EoZsBzvWQaLbMT6tDB3/SIcHTorNwUVLW7IB5YLx9hlpPXapeGsXUu7
YyHgzMp4eURHMpz43uIvDWLHRrow5GRWolgaVt/HDreNvBrgGGwEIqLxOs5PuqhOGh28F51Zjirg
ia4kGCiDJVgXRVDFUXk+B+biqd3ALMnjuQn4jaj9IymrQAoRe8JZUCZsEDHKR0tv586oS6RPdZmf
6m0qMeWbtRAETU5zbf+MUxUFtv+ei0ri5NlSiz7Bj95M/hRWdBu8LCrPhN8dOrViUWTgMMTnTPUG
A892RPvKlddbalXkT+vC74Lx5yZc46k6DE3OLPhIXeJtMjyM/zwmKHrmiHuVA6IQ3/jQN5fe+hj/
S1WNOKqkMpQkJ+KB+l52rSNEo2sZ8C5Mu6spQvYRbaLSr7Z2OqDgXZZkW8G5Paw3ukf4pnHF2c+x
89AH4NrNgK+WUtGTB9be1FGJ50GFLuEOxsS4NmRKuc3welKvvMPDh0JM28sfyVZy+/GuTMdWC4ZY
6N/OAKBO8tyvnmGIbPDiTaRJhjfrSoxkYCXqb5m0W5fUQ4dd1MxhWPpzeZ2WZtZaAydyhTqqE/MP
g5Ci3oarHjxQvuuOwNRMR9JIB09MG7mjwVwLqWaiy4qHzAt7GmISJ0ks0qip8fW1xCN34+4LzM/y
honRZwo/xMg+lbFwJkt/kOosvcq4EFeKcI/l+PFxrpNbyKgGzadmqUFa3PkRxs8xueHnpPZ91T7w
AYpqu99zoAhVwfPW7SbV0oFvGwwkC21jZNKvGzZmpUyA9mCzgKbhQG/qPc3sSL2REDkEY7lsESlE
gK95WZpwLOLm3XGgdVJKfPBHGEdr/fKd6ZlSZMQPfQ6xCQ8lfBeuF9NlrKD0nrdI+T3fDKZWHKGP
eyrfaSWkq0p/tBE3MWget2Vo7uUwgQcDqsGVGYVM+Si8VXs+p/aqKkB9o+IlLEld/eSN1hnDQx+Y
QCfFqzPu+5JjcFIGYYIbyzJyGj0/LGH+qgKEoJ3gpoBToYiCaPOcG/ka1DQtCgjJ/WspgYHiKt4v
ZHG2O4LfTna4vr2m4+T4fOinP2jvm0Rp3ZOF0WYiFfpLo1bWj0es+bgQa9m6WU1nrKoYnghRGk5A
Zt1bboliNrva7u3xVXzvNKAYGngyAt9gab235tPca2c7VK26NG3IOUQhhK5GB+NuU8R1TFRQnFgJ
zW6wND0IC0x8GXDIhr7RCqzoP6s/3rNcEccvh1wFZBwuAGr/qht7HSMcyPI7hR7f2bFRBl/FTMmB
GvEryQ5hsRv9hVqTK7zxTKT82ipsGHeZB2QH5a9uSJyvFA1G/x8VjgXSkSA3VqawueugNu/nf2ie
HczLwk6fFi9Em+E8xJ9dKFaa/PsN0ZKdEPi6AJlS+ZbZuGWUlMj8nsOZs2c9fZd2VDYx5Ad3NbVo
M7QNwjObQ72wK68BA7+dFXMHnJVI8eoAxOgLJ/T7QLRwqAuipoUIEfOPykLf48MGp9YV3BwObx8v
bO3Fx5B/sRK+dXyMQjsB8FwJPL2Lje2E8y45AQmksFYAizNqyOPHYtGEVLtTQTaWIqTHNcpHirMc
oLOz8mvJBANXHQipw+Ax38xkGkgwD/ojLI2b175euZ0iXV3kVp/YM7932wI/FKTRvj6uRZNggoCH
IP2Y7fFYlWNnO0QfdPbXOP+gmwJCcjCzfTlT7WsvBDAzEJEiULC8ftWq4oCUwL3CC4n5ByD6Xx17
59eFU78hSG2u2X/9iejghehQE4+I3nSXB//VnaGJT5dYtGdz++mdzG7/7ULP24Eg+vpxxFMR4TRk
m7YBz/O5aaAuGtbqCLhbrllHg/qBc211CH1dC2W5AXrouWgYEJyCg97rU6F4ZNp21P8/hewYHJkW
mS8PuHp6rYHcH0yjUzkLqQOJIFmri0HKXFYBBld7gU+cWAgWqGtfwYGftdsoFudssN4C3spexwfr
NtxbM3+Oz64aDX0n+E2K5qc/oRsW3c6vSha/eDzDsBUN3amDP8rUc1d4OJMLFEoidTDLEflTx+8n
XKyjxztfQY0padhLG4uCOQMoGnBSwaCcZiti/q2MukJoZtbxWE/jAhVmRJehOUau3arCXxR8nITZ
UhRmYc+jWnxnzMKlrn7V1jrUByhfSAUdStIMAicUi2Gj6zaEXr7Ytgy3BVfbp0ppklkaUP/Rviba
Svs4rRj35LnzeccFnNnnoA6mU/bFHDeQH3OTc7F9IfvtleYNhBwXvo4t9/30+lkU2z+Sxk3Ty+sL
vNoKMYEVIqIcpS5DnIQkJcd9c0DnvtBMUIiEEPz4tqBJFcUo+Z5Hwc+Kqr12yDRnNrjG/OHDb44r
SSw8WsijZ7mS/XGbYL5IjGOHp9wFhoaPljeSHrKmmm12ANeZOSs4CIoAUXTPgppVmwVT6PvL0mEw
04WA99CX4wYNmFSWiaS9WtbRKZAvvCd2UzOVg5Kd6wTyLFaQt9WXopdeYBO7N1hHia9sR7cB/P2w
j59YuUkRWn2Sf59lku7j/FeWClV9jrhjlkXfWUlEoA1W2mWFHI+FOQ5Hydws9gUBRTck65WLiYSR
5+Gk4ZxeBxN7QcemG/mJHcohnbU0QJPgvPb/hTIlfAk4HtGuWd+g7qEi7b2iWbz4J8oqth+elV/T
mRaQpoBqY2vhgAPn8S3TEvBoUw9WHKZ9zSaZKZD9Y8+K9fYA6I77fBU8od3IQAIcAwX24iOMQ+sj
MXjR54Aot8jsICh+T7W97gOvyAXSISSTcmsyzdjPyDIKOawoQna4Vm9SiqpVk06jDlFMr+ZqpHEx
lV+Wkg/6rrpLfo2dgi/W1c9BjROs163OGb5UkfVCrGKpYJnr4ARxnLNncEw5XRAjYasqSWXUwUOE
SJ85lmPj+ir44mLlXaU81xugPiuUgZ+atXd3nVojAH5aRlNPr/USvVvIVoXyVPyYjQRxWxV2hHZ3
49XKsXHt6P5/adDnjt6lRChFzKwbx+15isZxrlfn7NmaErSygZZLnYaWZaToJszKIntJfz5F+da0
IQ2NyeLuZOB3LRaIqxB/sLpmJ6LldS9CE8L6RwoKYHJmNCvTA+KRV7Owdx/XRHYHZU2lMSVqVkBW
+HhIjkZnFU0c+i5VXGubBAhCG1oeU4zanmuITpyWDUSDIJBXMWb0ExH+EWHYjUZHtdqLOgvjlX5k
0jeM9jrTJeljjjN/odv4Jw1OKpwlCh5AP+MnHKs4b18SoMiRaih0KAHwb85+mfE35cROpMdDntAi
31zVEt1Hw9MG3Ckm6vBL/1eTdz1Bl036O/3s2Kue3uyKPMDAIbF9C/zMrbDmvNF+rK9EDryX0517
d3TUkPu05nIe5fqtekS/IQUVyI3mP9JUwxK5KbihWL6bKBwW6/LqQTek8D7WyhQybWAZK1H5qcp7
VsLB1bkfvzVXQjP5noy7pzTzSWtKGoJeK2Oz5LqRbDpJ9LQReBwBWZ/HezOmSW/+WnYflvAzLqG1
QU17WVffhB4PDXh67byBNqBx6+y2IVprUO6FqaNhh5K63T/NkCRgEde1b1PT8CVQOZ0I23Zg4du0
d4Qi7t/rqhIGRze6eJZd/ZRUO9VUwXIba3HDGbq4p31H2CI7JnsIe8q3ybHQeTG9EdTW/MDUl32B
9RgSUJiCJDAHuQH5TdQkRRhjmlW3SZCsJKG+vxCHUdS0npEggrpzX3tgpD5N0RrMVSmhGn1WDVxb
d4Of+o+Xd4IMQnEypw1q0TYhtU5f1jObK1PEITEakBbtqfY24wSsBKYHZ7IHB1kl9B7vmIVpaVH+
HR071vpMuT3Ovo2JB25MOg4zR+6NGEFJyF0oHn3fYir1j4TmkxsyQbBOW42i/VQMsA6Ch2e6vLXw
VcXg7uusA7Sl3CGL1uhKG0jvzkMtYxoFA6fXf9Di8fVT5LvLMOhf6pvDRPvUxAjaoRPoNaC+xZfo
MY38zr9otZ6V91iLWrgBCg5HeWz7v5JIJDJplPLsJVplv4aB1v2J7CShFqF1Z0djRf/ZHpHwRruy
/4FT/k9dePKAbX1MKd+Jkfebl2vHPipSF3TkgXpulygj9LDslMR7bxrPA8th/48jYcpnVFsmB79z
hbY7wHvBNURhHcx8zKDynUDojSn5b40hfV170KB1ii616Q4l1b7eZuLLs31nE35ELsUpSdZc6H/v
k8YBXcSsHDi3WbvfUs5u/2w697jG4sz6bl9c/dIr9bOYBAC0YAw5qQ7h3xZ8vy98qj2KRFg257YX
l2J5lrvJYctrlFONFwdYG1QLeWkoJUaQIwTLnlvKodF2hz2zX5JiBjQwN39KfgWnKYGaC9hArgew
3ioMnbT2YH0tlqGl6XnTbFxUZ3DA5ZfwlK2x5mhDY3LOiINCeB+ZISvfuf5Xv1dfW1wEhe/Z/bmV
KmfTObV9oT8GUcEWTNqqAnroMMnEMJCBUYVfiHdWeohdk1tjuLd1TpgJuqREHtFAqxqJDA+XdHyW
LoAcy6Agf6GhCQp4UWWQzd7JIDrA/BLXXC2iih3cypoCFZs/zExxqM3h/PF/KJ6shRW7OXlqIfTt
iMWST6FK2u1yPXa9NsDUBm4YsJnvAZz7xhd7RE3ZGSFn1XjxfaF70ydtn3Rada7apS4BeyjWzcUQ
yZhqHF2oPNtyf7BbX+opHdJEWAzC0obR2wIToryTtyg+a3gN3mgLrvA5HkvezIy7wOg3sCHMOk0H
R8PlLPH3DWB2+Ld/fi/KUZy8/gs+5reAbyzE8OfbGDozhwzi4kDnBeChQT+l6/czS7Ly4+f92MeA
x2+o1SKP/t6bL7p0ErrPF0aQzPXX4h9hRlE12GB2Hh0MRmvdW6lhZRuD/6MMLYoYxHCxjc3f2cOY
ypTuqJIBvsKLxz73mhMWQPeW5zJGpSjyDwGoH1x8gLNhRRM/hLu96Q8wwoQ7Yj/e1lQtu8wL5MuD
BaiAy9pg3qmXqomugcEgpEh6j3HTyvQbgpsE8q7gsVuKdJfXh5D7meja8MYSifm53tMBQ+AWC9zg
eKDjwhT56zYm58y2L5vr0nLOivPcNwtnnZgZ7uOi9JYcPuGMYyFvvejYSBnI2DgusEkGXNSM0/cx
MFN4ZchvM8pSyAXDLrefeU8EheuL/5575NGbbzHf/b2uXdExCiq5NptRR/Vf5sBTdHGPiNbwdHYL
eHetHnye6PQBNtO0tQY9Qhk9wrWo5Qz3rKEFWoWqCdZEU56Tcl4vzNPvVM2pZvDq3gPvsqHyVaBn
WKDKVBvDy/Rjr1AcmiyBykW/kcrQGNjzfGDQgpLt9bIitkXoDHKDbpffGClDVKzmiF61un44WzB2
ljofagNC6EcPNtYSRuF10VCaZxHUdz3u5S9Z6aYDQYZKqXGvt7KGFzvivjFaI5WRV+tmXKXr5viI
tiJ0J5lndlNiEok1yT2njHDk9yQ4+mN2rj2btD1ibqZXpUhZ7TaJOqk3ADefxjfMQkJEWPVFVayA
FvEu1QudUs0vzkOFBhuaocGHLXKztRt8+eQQ7QnGdco93s4JtPY4ZsxmyRasaXsYgc4FFfIVO3a8
a1/cGY0okKQBbvs5j01ideO3gfrop4q6Splz3pPojxFTyEBC8D45dsupdPwrmvU0dP85ZkA9A+o9
83YKd40tUYJDy02AbjVf0MaQY+czlPMMtXvr8Mn2jjoH+bSH18PJFtW2YzsejTSqIwlqFQGLZccp
lPFvGCf0ENynDmbnONeqsW2d+2W30/Z/LoByqxPlOa02MH/4sPh7YOp7D7YWB1uX8tXpsqSDUNm+
jnIn3Nvjj/nrUSFb6RyryNY7MFJ2Rfse4wY8B8ciCyX2XaprHajSjaDFyQqDsSTrdtE61mLTil8/
gR4O8NwNmzsor2XMk1FLLdmvNX4j0LYnhbIPdZUrUQJQx5f2O+G5TcFbJBRHO4WZlKQp89BWwnWK
lQ2m0QBobOemJ2FypRubsDfcq6xrL39JY5WWqn1bIWsPXwBu2R2w7fx1QPb/dpaARSSqNcLyVJ29
2mCIt4vqdPBE8H8F4KqfwSWDeLBQnNms2dl/GeLJTfly7vtk9GZ4lnP51a58VBTRcGtED6KkYu9o
4w5FrDhXkbmJKIrOp7DhKnfPfrSi0B7Kx7R0oVEQAdunQP29XTw8nXCS1153/EG2+PkXyHTFBl7g
4LYHXYMfDuKOHprj64JgNo3RErJkkeODD+qLd+gY00E95er2ufid0flL0kkKfj8K35JwTC/D6ocl
2tx9YlbekjAHBRG0WgDZq8xxbhfQcfx/6qtEXrH4LhN4MTW/AxuipvBD8fWewR+B2RfHMNDSy0pi
VuYxxOQa252vMdcABTzRGFqh2sqGnLDoYurIMr86FdIZ8wqUpg7w2UG9DY3oXBKApBOteDjr4cAu
E8XVxxmp7tz8hb0Pd69KGjXQw7I5E58GFUJBgrY8QOL96MVlKZErT9JU3z4JcZroRFOqezFZz6bs
0BwpRXKhJ3plVueEFP9fNpkaKQhwIIQR6XyX+SbWUXJUctvWnQy4wQGrVt2NAEBcg06D7JoAA4eI
Gj+A5OIzGa+IhWBaWUULuNpYwqLGLOHNExNO3jHC4eEqz83rCt+1c+3RJ9oNbhW0aaPng2xNqiQI
3LnO7oCnFpPKSJbh/j66CM4NcLs3OHgAzggZJ3V9N4sYjx0YCImohwmM9YD+btRcrEDQLbfKaJuW
7u7rUp2fiZZMXBSNmOvpBE27GPZjhechNpAyCu/kdPsERtPBy49rdBH8eBvs0Cn+6has9rWF+CaV
c06R4VDOoUlGS70rBHFhcysLDEx0SDlD3Lzn3MWcpZCIFYEv0htYPoQgHL5sGemg3BJhLOs0d5mn
v+e+noeImKHFjJpeBvGpfP3wdbFXNRZMBldCRwbGW6XsMlu7C7d0pBgRAL83YL/IjHRzhp6Sk6+F
VMlBvvN4JmbHwlFYcO+w5pqP/Vua5OGfBdTJBR0lNRTzs55PfnVwWg/ylse9SCYIuPKshN4FSEuc
wOf+oZzm5HOw/SaVS1TN/TZH1OUjiEyNa/bZfkYJCX90bWve+ipmnvVjFj5/Zj4wTA+RZVRiIdCW
Uq/plVamlbVNg4AqvryZLt/wo6yFZUqjmOFY3J++ARFfz4NQdZC/E3ofbu8SfmxmMKGrGM8DApmK
pWWb42AUXioJ1hMaZIF6kDZRDP5s7IDBulvnZfzZYnvRBp+6YQyZk6ATL3hVr0LwFbIwJVbb4P5j
TjTAy8foZxSGulv6H0C41/pj7stRRhwgTajF1muGkGhFIrfHXEiC+IGzf2p9fkGZUYpiIPoe3rmR
By8rWDyQryL3eRu5+9cVdYRyyyUc4SpF11tojPWa3Lm0f7cLVZ+uCU2XM807nSqE/6d6vGKNNzbO
GcTNOeKYB79Y4z4Suw6BJN/litixzgy9saij6vZJIqwz/dZ90zAFkS+MXPh5NkDJsNRvLIMuudeR
PKg4EGFqtYxfJ5MZG11cuXV3wTRZWSZ1o8aWKQVI2YUiI7bOdvRoNTPXGXWyAcfx4hZKt+WaMyMz
NvDbiim7v6t4NG8JDK+HBSxcBUOD0KV2KAwwWgE/m3vOfxTYo3AFUtc3vR5qAKGS9jKE9splgEDr
WDyuGJe082sr4gHHOuYRGDyATN7x3aqdzOeyNwO5fyU4ExcgT5sg7YLaFgRkFrJM3KTwXBKsJg7e
LmwVK1E6rAZK7YQ64X+pw+FI9iV4tt10ou1MwILRp1LPolIC8P4rpPGagWi34TIMVQ5lksMs9Rvz
N9YOaegYW8qJZ1X4GgM4t19tMWWk8aUK/gou0c8/tsSympIRAcbYzIGyw+WzjAWppl6Gfo1vvovn
9AH5QAtbF0H+PgXBpTdjlOLLvawm5ea0otiRq2RLCtJZigqW4H75XyHbabdia4pic6sRUewDOcL7
wmTbVYcFgG5HoSdqLzNtP+ueny09UpIvU/eNitYyurFNcyELj3rELHx4LUUF+mtcVGbOX1QWRr6X
Pyt1XlmRMQ4eiYQh2RW3x5XKAPHO1DFj+KVLIdHXG4HJ4GdSjCkURKQD2z9ZFsKk+/RJP4RIaXzu
y2sP7ubNq/hohU/XeNfb8LEA1Ur+3WI10Ox3pwFpAppvvSRVvgq05HGWJnSxEfh+bvZHkSz8/SGY
lMhzor8qNj3S+c+w4u17wbSWqRf/s+oy0lKkT7R9Hi71GWNiMHGOevZI7xszkSmvqeCNQSBxmN7S
uUHt7ngzxBELa3od8kpRgnGmr91hb359VIX1OnytkSrDmSGqjsz4oWavLdlon6Ir6EDpdKrnLgw9
wieFEblxuy+fz2rljYZpa9Tfnj2H0nh9Sssegx5JtB3CC6WRB3KS4qtJSpNe3tfe0Q9c9Xmn+2tf
7VxQTQ+in+xi4cPZX48hbbypPYOox3Nt3XQhAhDoYM/C6Dl+BUkbqd1UcXebeIO82JAsf9jO3L/i
gk4bgcQRWiLBNlOL7oqOZaoEkvUeCMeMGPPTgYKu/pe3X/zoTztnrt4EVsLSqbgRNu7kKKgl/bK+
JEmYJx/ZDVr4MiAJIysmOJITTrY0DErcsxj8kXbLZO7eIYoQrMNiS37orxPA7eBGE2runRo1c00J
ifndyjTLys3lEPbDSuDommgmEuQt5rJvnOrMzJrzML22g2zWZEOjG97FLJKZ/8NF7oC2Lz/KPuAq
8qocqQBlMwl2YaqIvqvUbVNhLLX8Ss8PB2kH/mEVHfeFh7tI7+aeRti1Zz6ixi3EDfZSxnNuWkGC
a4ur6Q2NC86jwl18rdzuSjmu1uClN4s72rOsKJqzYsOlQnYU5dyf8qUisfv5dK7w5haKSJ4MPfie
GPFlKcAf5SDP5CRLOXLqwTMj9KnnCErO2HhyVjAMaqDp2Zp8UU1NcmYfC10IlTmjaWG9sLzLjTMS
FojZxtao5ZvQ0cqAtYkagrru0omIaKnzs2UpawMzCn4kAikg8Evkyvyr1B5BG8HiEAR5th1sA98e
8DxlkK6D8c6+A6iC2RBTe7smaNO1HoXT11bh0IjQGDjv30wZAuSQaoTrym9I4JgLVNw6tlPpeUa2
iqVVrpBa6If4oaCDGAh24ri51dR8UVHyhj+dQKhCB7n+9zkjUBXEBUfVSqMlwV+z8AhwWTiC1ytE
m/j1YorR5csvNiHUjzOtP/6iI8t+eUEPbXWYgKk45rnGyUYE/P4mgubZe7tqXxaqDDh5e6QVSF+/
SQRaLSdcwb7OxXzxvvOXSmcGt7r7SL1RD9cypRknSFUInNUoqoLqQz0cJLpyCfmNa/oCBvNmGnsG
cHplKH4yxYWsQ226EdhXelM4P6IIjCwJQS5qYyVsyW2OOsXf5xhS5y2olx+ePKKAuEoOjNq88wk/
AW1pttuPj7vYgRjW2fIHMtxdrumZRLMrTZT5Q1z3fSmdTFFIQUmMBXNU8Ybe3TCSg+/FUTX0uruC
RemTCqtKXW2vc6yxUxYNfX/27XCH1ZcO4vyJC/wEi85bpPt5IiGf1VnEncVMQ5sGSCSZU+IPBkt7
abSutQZ/ieC0XtDliV/M5N+dqCxwtnU2ql7hMgYIrgpWCzxBRbNHi6DebsQfqv/sog8fe8fvC+5B
3/gm7NIkdGuXDcJsczFHVPVU8P7iohD13n6n55buOqvuph3WDoUmvO8H1lnbzUw0VXT4E8w6msBq
U7KEDH5je12LRIPe+Or1i8FFpxArLl+YPZjG8l62xmnquKo5qP7htofUJvlUTT5ZmdwEMwFYTWGn
0zHGOGCiRkIWT6QRkHLAGxgs06ksm3lqotBYQaQdOaAtWZxg0hh46uTnBViebUC19i06zxUsxdli
a2Ifp2FKYKB8GYvxXczWuABYck7xAO0vqVDnojIocwcMkJWI8l5vxjeDfnLRJk1WvG6n5f7i1/zI
X3tU9q2jCV6bdoJkaptpDgWLggez207+t/6MioTKFa86VWxM6mLH7cADG5kPhGbi3QSxyspYVpXi
LnvuFqKdQzHFIzp0xBQxxTD6YxPm+m5aIGyGt2K8+AT7e0MKmYfh+amQj1+wKZ/Xng71nHr5Tk/m
WyqPnc97wVsW8jCua58p02UePRyGGIgyDaDpa9WCLP+hvnzYLpcXPMQzsLnG8HcLuuEDxCB9D9Gh
6Hpq4Ht85DIlHub5cdcCJrCeEzPNUh4rbFSJYYUT86ZlKfiUyCE9MWov1Q3eEchosTd+zzTKmKz5
DOzDido8BAmdYTq/au7dbCUzQuVyA1A1ejisulDR8yFN1Q/40xXVatjSeu/JYRPLu3x3pfMLSAp3
/C62OIGfm9C0bGPIdQFh4JUFwUVWYR6/RrkpENLQmEWbC03PJjvCQjR0oT7iJiRQ173Sfh5PZ7TZ
fJwmY45IUT3e3fGdF1FEKSB3uw1KhhHQeYl0ljpyG+SqSJQe+rAoFWodMELIj7voiUGBFIGqKybf
D0ij0zq8TOspTu/3zUxMBB7j0UqMqkTShRinNeBMebTKV7i+vSddWPWSmW0lwtzrtP1wMp68y9sN
jHy3E6DvajrNDrjKi8RKgExvaCyqDdmjKniGKTe5YcjfbkrnbTWkP2+Tq5iIAjCPBd/8xWG2p+1Y
CV+g+9s7V3Vc/yqZhNBlksLwPH2iSMqn0c8ErksVleVqRBY1oRshqQWfA2AWBoPQ5uXzUp2XzBZO
2OlEGUO7wPGt453BJuboXKXD+gD6C8AHzSY+8zmHzF24xRBaoAWUe/zfZYFSrorFZwHEwv7/f+v2
+M28ipYVrRCIvDsE18aK6kxb++4Zsr+j+EJYSMwk1VdPeQ32vn5btbyczJSIqc1o0P3D22O/iLh6
eiPAT0u1sc7Yw1xLK7ENnnRQaUu1i8JFv4fVu9NTYvTNuKg3VIBfhIY2T8mebXfvcagqHjaIP/5x
UlzYPrIEtvcWLdUrGahe48DPc4pLCpLgvAzfx5muVmwSMC2JeWHw4+JjHpmPEXZ70Uegp23ngpEO
2tQAyQYce+kpTffw/jsuWOxGcPNfqUIFThSy9GhJL2ZqvKZMeO3huIfM2sepu5VGQH4T0lioXVl2
xQuS+0N//seUJdrc1spcS86mU+Mgs/58JgmG5UtjiDcfV+RnbbIe3RTU0Gt3AjeeM/WhFSqQEjHT
Qb6YUrMNo+5lUHS1SypcTWj1721f8u35+GjMoRdBIeut5IV9j24IhkPnoX+g8eM8X/yt+MT4VUBK
sqGb9Y1lYmTviezz5KZeFpf1K/C6vIBDQhK6TjLhos7VIjTxpwxoxuc/U5fGuYaslX+o+hdWMQTt
4inT3tpNX4AoNtDU2yY3cU8E2Z5Gu24/BJbCQIP4wNtZqT7JsFmu/MOFTxJ0GubkF4pV65u3r5R8
K2dObIeOnhZbic6m607wZbAUR3RI0P87N/qdlr8N1hxqxnh/wG3lxZt4nzydRaV1l5ZCxpoHiRCM
UWBsh4JvTdcTvP+guMq0l8DgzwheakCsABDCKU3uNSOhuCnIWjC1A3yUiEihIHPZRXfGIi1UQRQr
Z9BpbQaau5zMpP0ol+lLEFbZA8wVSzAj71vGAq5HrxYHTBS59FcNQSQ3/8Ir9z1DfZsiPRSvcI4w
KB7x6CfRXtKDOZOUc1/olcFmkchgx7r9E41SR8veRDxqHrUI/kzjtJzXZKYi8+iVSDlM/2mCCceR
cagnLDbyc3I3ZlbJq7od0etfFirqLGPwpuPaMXPl1LRCMNR5MKYrEIdRZMC2z/KTp5owVeSblHXP
shbDHdg3yWqrvKKtT4Gqb2eRcwLfGQPEgesEHLgaOVp5X8LTXdiVSz75BeZGUjPorsprvsFE+2Yw
fHXsi9Ykiroicb7KOkTozQPSeMpCf5rSH1afbLnlYhCuM+obvp8F/T9zHrlZ9v1hLCjzsUFNm8UH
Vm7yO1s0gNCz9a42fFGQpUBRk54k+UQrMc+SgpF5cKFUPM7XyfOqqBlYV3nk6WlZcnYvdJ1ZXQzB
viKRYh4pLz6Kwin21Fdol+LKnsygbGsmNuGgGMeXDf1vMOo4KEzJQ6D1WZTWphFB9HtYecVOmHbj
bETFR3P3IPzUzAKkGOoq8weKUQKO0DKGTe1oY8PHibXBn9wPPKoxAuELTXgkn4RY1qxxppdx7407
T/IJSPek45unNI33xEwIorqSr+gbo/YDVBnIdEhdbhNd3GevUvryykiLtSuORy2COC8OGRdKTY4t
67vfRfHyq6HimoSqugCVISjbcaW46k8zv3w8PoD3hIw1L24uzKUMyxJVNgt5RzyTszkMwW0WAswG
Z3UT54YOlD0m0OyK0qHwyIN/JxUXLoYxo2SmFx6sKIXm7T7IbI9aoIfzOAt7vRikQUb/prcXl8GF
NgPM0sTIRSmRLQUk/vs6XNs+gpn/9yO3K9tiyWltkGXhd4xK//ijMSL9Mz0GZo6f9u4Qg4uZYGZW
tz3W08HbgH3+AdvFBLDnq2HbXrOnsapva8DtzvQNKF7M3eoSB/hQJTk90kwJWbjMtJtQz9CM9IbB
nOj7vvZo6a139gXHtacQb1QNGxwW6Pd2PCN93b1gFojg9SqXlVnV7N1/EYgBPALmbJDBTtNS1iEa
ZG/ccpGGrCNDZfwjLavl0SOxa09yCombD/3Jgpn7VYeJvEtSV4XOytsKiRNeDq4K9x+cGi83UqVQ
VI2E2q5rUeDvaoLIh1P8bn6QtqH+HWRJvnQRccQVaHdk6qMPBCnpedcybkqw227qmyZNavxlylMS
TQuV97wk0QCQPFeuPXae7ATekb/x6TJmPP34cyGnNpP+Qcm7Ke/94KIO2KZJQD95GQUks8sbFOj5
4Q3FUA/PDL50G8atdhJoPfTbwEjwlFyemHwC4x4lOxQ8wJeFGaOkkLCoepQesam4ihRt11m7eiTE
kzIKiHQ0WlZdrFeFzF9obDO7LfsCEy/m777TW57lvi+4Xan65WG2PKz+kCzqCO9R0qNPjxYHSx0z
EmPWHCDXvfmadCwYZlDPsNuf7RDTfzepFZ4zsuxRSJE3gni5l1qO/uWh6hfwg5UJI/iWIqMIPkKg
MWLDrha9rxv2f2RVGnjJq1NhxFU6+xj0loU1eOADQRI58Qn2xJkNsXwfUAUB/77aRAD9Y8Gcp3kz
6M7HvjzpSAKoR0/vLOWZ0Unjwziwhk6GjMTyXXD1TAsnDdjPojdyJbDMOxek/x7v17PboeiQDUQ2
aqCDoFSlV2hu8hBFddiREoJppt6CpFwlI5pwpP6wRA9KxwfOy6TyvXiGS0kZ7ctdVJKA4C1/GT1e
c3mmE5Zf1n63vni/ju0S3kcZX/PM7TI5vUFOaLiH8nmufsG01pg61SNXEGp7ntbXwNFzE++tHeml
GScEw2/u8YlyqYO4kCULzRGP98JnhKYbTmBhSA+X8j9NKHFDjw0SNaiokrn19BDy0X1lJ3tBPGBI
nurcsuuJS1aGKcGzY7bGGN1Dd7djU7z4Cv9Kx0HNxfaJmHNJCvMx+EL9i6ZUPjE+4B6bMM5cXwsg
m5LOletNv6Ff7HShNbZ70YoxYsSx611KK6J0bLzTrJyT/hJ2w+bR/7bbRnj80PWJl6XBwEr1PDw8
Eo1kDfJjUAZPKFRLnbzkam78/iRlcDgMAShWUvKg8lSLk4R603gYatp1skaztIdCz4XhKrUA+XoP
rmvrqmRukQb33u7AlVPXDVCxHrxfBmc9L+G07x46swlhH1tt9gk+GepJrZjaI2Qx/21uRWQIKXe+
Ks8NHaqA2BkLdk0uOTlgcwvb7/wEOdveZ0DeFbmzRVSPrw2lGfEMiMT5IaCSJmAEsggvNNoGSwti
MYjfDvaF1p/wpkvqKxFsoYT7xILl+ahx+mBynCZnvV3UiA8FneXdevAGiWCz+HJEUfjbhm6i0+yw
5aGdZFCtWdCsbuX6EOZK7abWMYop15ME5wpXjifCrEuFvP8pNiQaQAywGugmIHAIV8WPGhO0U1Hd
Tmkc/n15J8k6GRyZdBGDkfsFvT1qLfYjrnIjZfMf5cT6xNauz9Yzkh8LmakrsccKLgUwoilVx5zP
Rzq1sOQk/N3erbVJleQ49qqdL5ld3ibQrY0B83mvvcfV4yNqQdFU+2aXKcH2ChtYkKy06bg+5XO3
bl0yEMsTUXlazzPg0RDINrDZP3QmqmX+zscCkIkS/2uGo0RQ6alo84o1VrU4EaMwZHFg/dTcmusa
LUOkw4/jF20f/sB+JzvhSqx5XeyYFRGUw/IVq5Y8NOD+F1k9sPWUCNOblTEeAZqw1ITFOL8FX4BU
gHwxBe3uGe4QX2NP4G7MEHI3vlHOkqsjCb77seVyeUn/R1SsTpoW09nJil6fgxIRdOh0zg/WQmS6
LeP9yOIQUZrLUQ1dpaIgAC3yrP+lFd+b4mnY4DvIJp+7l6qRzYKGPF5tmvcuNwqUu9xHUUc6A+SP
qqVKvlEtg3NfnyXgw2LBi7XcXg0aMqKsazVmmF7KI/vo1fvdmoa2NxbgKxmNmJrJ3SsO/Ol80CEO
H7+ej5rnXqUN6JTF/khuW2KDAKq+Cev4wKCbXx/+3Gf0ZHJ8S2N31Ej9sH2i0iXPZvFwqIqZV++7
K979cKGZkl1tc7pvMlOWAhk8LWHsClTqT5wBXRU5nX0mtwDMc3RmZZsCr/kJFEvfGH6MTPtABoc4
MWNuJZ6/Jn6l9ux0Z0MW+5DgIU5m591CJJfvgkMAKUxthM4lpOHPyyS2AQfpWqNDRyZa4O4rkWFi
ovqqI23DCZDTzkcVUiqSWxGufYWAzQ9HHRcdUc70k1nKbx4KENTM3T+ch/EQ8eP+zluwVV8pyRGy
BjeXaN7slwSRaRmfIo+mUAPs/DFOKqlbJ7O5Q602e1Kp+ewcDcOOdlIHlG7L1Oe3L5VHxALVXClZ
AM6Tw1J+LJg/UCrfTxy5HvD5o8AQtK9XJBNlT6J2/Z/8Yx8MfqUr7nEMNiGr0DDvxf328Nk2UJRD
F/9tTOTIgGrIy12THe3mUZxaDJ7eDJ8r5+WinAaNkCEYPxdbkcqoxLyCvS01JfGSUf3mSU1L7L2G
yGi0G2l2heCfkwNqwp5j5D1gDc4chVobaijb/xYdfv4R2CSqwJ8B73PkDng7g0OWfJcYHS5skESA
o2E8Xq9WuBHLSr4Ussmm4A0+tEEo0IlBSacsZco6QgWeA+9eytDVej8b3xwGqnTtADtTlBkkqgE3
SdZlLYLURo6ajrribjim3Nha5Vv0hmxrLieEKsdxeyfkyi2g6sXiyoazGhZCcs5U/WBbeNOVzigR
hVUrGCARvCmeNrVpGHr9rJeM7G4yN62yOIKXF/T9q/DXpBNPFq2wgfMOEn6aRcBBk90UNIu57/EK
9y/GLUCwodB2OODaYe76xFm8cIhiZTDOP5wM6e/FBamE4N79ipL+0zeElgagfbbaDNMOp0/jnN/m
WtwKJ8KV1kgHY9xGuJznaPj+5plzWCbB1uxBZ6iR/ruNOyf6Fa9+D72aypICZlbn5JTs1yzLTQk/
KHQLJv/Qxj0IAhe/y/eEdtI4vj7xpB22DJ25DJ6CtANoweriJyT0MBwZKv5GFoLYY17WME3mDyj7
fe7M5MdDp/a2VANxUXGwWSrdv+HyPnCnUF4EcV9RI6DF1W++gN9+FSV/2c6yudiOWXU8ZPnxOWnP
+TFgW9dVWrKZm20m48/zvfKH+xBilJvTgHEByw4p2x8/w5pMeqHAJgIQT7L0wRHAyByQlsSMMWEH
m9Gkag1nYbsCA6pqyIKxL86/8do73iamMJPVVBNNElGteNIdbuzJOii+Jhz1vwI1J/Sza9fQyru3
Er6izZPgmX82nuA4btwx/rhl9Men4wh2efIXTBI/5ve9GlB6yfHI6nQlCZsMHCausJVepAa7I5A4
Q1vhZAuh7GAQobUhOcH8Xxc8DCmr0G5968Etpy/CtEFZ6YgrDvrFGMA1gjik/84hU9XlKQBrsRdG
AZh04aSqipOedp3gyNX7iGMdfRQPSAVdpfrwce+8OuHMKDYHvU0AxHL5oDhnx0tjtZkC89BfNmzo
c9VR9Yd99ENb6oFWGJjMeJAAKRtUAht0YdsCPsrvbn7TxL/dl47AGr1/0Pg0C0aGBoG4704RK2mf
3GsaRElVAEnb8VpYTbN0fTynYmgbwU8pnu6JTRUAGZvNNTI6KAlCXJ9QWsh2RgL1tqpjFLmKJOYz
u1sqLmiVRrN4/1gy7HcX1l2vvZEU639EfsLYXuO9OaYmuN1lFPTVJjhary3chLHiBuhD+6Dc2O5i
Xnj716At2CRjvetHNLF/sBo/PpEzeK8MMiqjmvQiCEMoCaxBTYetZ+lg8KGZKQZVj/xmeYiUGtUf
qkBB78wy/5wA+XBUy7fYVRxz9bw0kfJAXsOJs5tkFduF29jZ+OirPGZgN0O0qRHZEtP96Gmj5VrY
iyhuIdvyplKFmPNTSOUqf9xQwEC4+jKhA3XlvgzIHxF5CSvT9M1GhZbKoz0/ioyjwZpriJwdvbzS
cbAWumNYuLKo6p+1VSbwe3bl0p8jp9WOlDqgleuZC/dDs4VYH//nbkPnsjW7lh2WyKRBE0H1YbjV
P4qBHDC9z/a624YTyuvuj78H1UwW1byNGYhoF95JPbZRkfeywj/JpFA+Ke/UBf18FyaTapVykx+l
pwY0eNwW2ZeUQjCsUxPfcr/36zKSLXlw5GM0NTm9VmaDtGwUSZ88DwLizfFz3NOoIgBLnMZXsW87
6EF8yX0k4hfe5D4VVQRTz87KVGiX+fMI6zvn6kV6KsotzA07kjK5On4CByzLnd4YrAnthGB+i4U6
kCQUdMbI9ugancm/GE/ke4q5/6TZxnwbZWIIS7FHIQbrjIedDImP+gtY2V+3sF61JJVHAJrxDDGK
8Jwmt+jRDAj1gP0w7Zzo8MMd27JhwX+dv6l3SEcucLCoewUyDEY0SVFnYFpK4LH1nY4CtpB327Rv
u0pMG6kUfxb6M6UFgs3NtM8v6SOIinXad8MyJGuZfDgAaRAjpcS5dmfggACMo5BMqIULb1TAyDrY
t6Lo0mUJOQR9Tn/A6ggHNlg2xJcwh1tANqFugSWmEXdBIKo5YVok9bsRq5kdZ9mEpdiKilsvaHro
3KTL4VN8qTJwHRnBIoxIX+VKvOtKrx4CIhx1r45a263HKiWAyl6/i1hCbAwK/lB4y2h1UrcQQt5b
Aidp8sqrS16puG3qOXlSvytLldJevGjzN4SSWjTAD6y6F3h8ppuYoORnaxdqgDCWumumUm/lkvC8
YcQAltnIastvCVnIJgKMivz6SGQNC9WEHJm0j3umNoaNOdJnDFBi6txXlUXbJVYn8gPQ3zjQntcc
04HaDZ8yXqw4xcG/IGtZZJSN8vy3prhX+nGPFd4MDqcOvMqYrKfCRlxTQerfY+APvF0/V1F8mobf
UAWlVL8VYy4jL8ANL9dX3dII9reEnacv44NnDBFKlqXHr/ChP+XTHs9aPChEEmlEDbazMvcqxT+O
f2yteuP28HrXEKTe804etqvVYCZNKBN95tKzPPK1BU0JGQB6xbufbmdCcALNy8NiiFYX0/t4xwNV
+93tVSzEaRdzdtqqnUupydmvv79m8QmBgQWp4YAz3D3PzWjombvuGX5FT+LwtQNrPt2FJXQ0o4dj
ZxK5RHcpCX0Ls77HUeTD1a2JuRaT+PIi3BXeLh4s+oQ4+HPDPzc2ZD8N9lJgNlAFpO0UPC2bJS8m
MFPVRNg9qN9OhUCLSAfNfXwd7ME979Vxwwh6xvV5u6wI7t3Tqsrivfgg+27KfJ1KdMJs5WlM2L+j
QN+3Lu30MyMd8u7zReK0Si2uy9cGnti1GO2TTd8nmnPRl22s4J/QMMwLyNZhWdOU0no9QPZFGwXw
yXSduXUud8JjnUEzCcrsrDzgIZp44V3UUS+IKvsjiyWTHVKN+WUpKPn6DudQRugoMt4IpvW/kg0b
v7YY62kcicKlrandJFtEpAHqM2Oq4lygPc5JicubG2a30Is1Q+N/CHocWihprCdIkD8xbFXxx9Jq
nQoARBieVBjWm5gfN4KWyez+9r4IiZLeN1HhoiSNWNMr2sxH6jTRkBEQd8BMMkWU3EwS65a2lT7E
7sp0FxcT1cAy6ZrxP/ZhjtnaefPawD8knpqHIgr9jTunoDKA9V/u9ZQiniP4kvTtmS6dwnmb8GXh
tCYXLWTV7OHqokWRs33WYYgSHaudGuq7KdxDKogczIghs3kLVIvDnxmVBonfHtRlzPTUlVW+abIU
bPboOdHVeIcewcqDcxBKhYh7QMGHNSqJUnnf1A5lZUSSAmy1n8b/+cWYQ5vaNZKDfG763/8ul0bP
Z63VaSBtPu1r0J0l7WsNt2KvRl9iF+Z2y7jnR5NQNkJbefLoKKkoSgNPX5RSZ+wTU/sVrdPu5/S7
1FNg0scSs039ARZTZOZfw1+FbZmyXn470oC2ScUEBsZ6ZR3R6JglnwikfeNmkJUELzZDlod3YX+8
6jmhBIoGyNFf5UanV2kPCMSCoo6beaY9jkWZ0MWl9yFN5TVmbyw141gv02LxhfSvrdXbNVG+nLTY
9mYohN7BtBpg4dsfmhEHEtClnPfpN8vIMsb380cMIUmbuZLWw81ErI4QKGkYyNncQ5fWs2iF2gr4
IAUlIw04gAe+FSbvcaRYzcyQNwyR8GhVwtonmx2Ko2yjjLO1Q8n4rgIuDsFlQ+uSVt5WCTkV8TN1
ZLzEnyek8FtXzTw6uVd9J9MdKi90OdHM+4MID0n+SfxGcIlMOH9cD+ALviEx/xPfo6Dl7zcu0Rfi
a8w1qNyJhJW0EqCPa14PHF/3cI27Y5hFgkMj33KGSUJV6S5iV6Pri4vO00D88v8Z3UU6FeGVa9GU
CucBp7t29JK7QyNM4uFequtgzXZrwTZm8wHv5XkTVti50GHJPx7dP39qIwz2UQ8AvtK/tSg+D0wj
dh5uHqt6VyytUoSF6253l+rEB1L9+QLb2uPzhdsUcIRjC3miwzr47zAkLHxNE42YauAwL/hy8D7z
5Gc3bcYGsA3vF98mymlOPwPpw5TVqykn/5Bz2jBJFciNYp7/0GC8Y0fLwYUrdM1CysDwstsR3cCe
ENYf2N9pZ+hCnoypLCmCfmwxrjLY6RKKbSjUJZEz0bVAcWex3KKqOMOG/VOczCRHomM48xXYaLj7
Kx2Yzr4fGdyaBFY+i+1zZYlfoTdIxbcYImimYDqiDNQaffQPsI2g3mS13tYbK0qZp3s6DLeHMsAU
2p4ZjX0oTB+gQ7uOZQjYRB3TG7tcx1LEPSPC2S1DPZ1nHnqXpQhOnBQmzu3Qw7GnTS4Qfx0ZvALH
drKlKw9HQ4yQKrMfOi0uIysB21KIGGWpPUPXT/pL1OlGEtTh0X3D6pRicviVTPzh/h0q93tqw8eC
9eqZqUqfcv7bJ+iFMQ/ej1NvM469IWfihniK6AWJS0e1vEDhQhlq606oa7Qp3dCxrS0FjeloKWT9
hv9FlY7SowLrbGMC1sxvZZCJ7S9J7BmLINKOjAyYiP3lrXThCMcdEKn+Ge2pPiq+T0wTmFBVkela
ERCamkv3M4d98EqKnVk9qChJ8qjYJkwonNrFuT8zsaGS6glFW+4FzbeCrBl3BaWLaz9hJ+UbS09w
iqJaSaYf7gyt51fCS6AcEvEiYTjFT1qa7i6WO8r1Hy+5xi4R4AkGW0DSuJtQUGjAG5UKiV3XxqVn
wnK708vVpRcPxfpVI5O7edAaApwz6wfUdLiD+mJ2WBPVhnPh+M30bgEfYoJ98BFszbLSly8l8TbB
VQI+AjWhj5SqlJl2ORquZJSx4/u70d9/d+J2RXuKwdf7pJIiql1dBBQOml8h+D99wnJrjCVEgQuk
clADPf0mszWLypcFoerjCeD7AS3yuFgzvfsao4EoFn72CuQNM9PhLvwDQ3QQ2ws8/KUMurK/S7a3
wopWzuUZhgE4QAsKUk+AsmYCa7NflImLSJ4da/ZKCJ0ankvPyDd8xxyo13ShmqUywoaNPwF2ykK5
aZHXKQPIZ919sPPuWtQ+Me0g8zuenx1XXn/Eq9wQPNv3fa4SkX/zV292SemFG0bwzTrqUk0rSAqV
atctKuDBfz1ka3TJ2vFd8I6M2q/tTYNngpa21MCD1kIslxqmILKhSMzKhy7YJQ5xk4OEpMldRXQ6
HMiO3x2R0TAqVQnbvIcncXnQ1tLl97YsRuUtrLP3+7fTeRswj5lXXifj1F1lFwgbzBo62p0awoKl
bmKJe9bM/uO55sjI/aAUv6lDO7xMv+5PFDosHJXGRxJnoxmgmxiwl9oTMU6VRgv5lqnPgYUHHely
hRI+r+UbnUaNGK1I+dLzWncM4u83EbgfUGaWcvuYxc4AB4kxw5QES8/gcmVZ0KI9HwxnOgt9wdSy
M6x9tgN9wzg7Pnb5v9yNAcQI0e8yVkL8gTM9KS/1mTyuYPhe+y+qq+XV0p0fKWWhUasbJUoaQ1rx
2XrYQ0t505HqQCm2DMOVUCLLK9k+FjN1bmwqTTEYwjIR+Emk4ivasz0dYRIYJ0zuGqdfz5qV7ZLu
AVT+7DFFoL/jcTJ1KTY63QpAf9JX2XkORyeU0EIMdM3QMQcJD6gcLJ7Ph2WQzg77pMV4k0YnhSyj
U+MSZ5fReINtUEDiKqEXzsUAiam/qbesdxNgJF5qvm08O6HfLdETu8FRsJID3uEQZH47QGgaIvj4
xGvvzYFrBNE72XElI5lKExDg9Ddaa6nYbk3BrIgvz64IMV/jFZMNz6C8dBkPsv8bjS8n+M3YIWuw
RjysExjNf56sxmJ5XhKA0pl0jh28Uay3dMKRDJuVWCCyStNz1JgYT88jsL5Oszt1lu0V1Kf2lqcC
jAkxDqPNqGyj52bdU615R+sII6c+AY0Oupz7AmZJfcZLExhx7LekvcLgdqmH0Vr/rYvD1W2lnHnw
6TJPet+wKeL/XZ5om+T2I6n/4ZGrwTTcz6dlCDWLsSE9J1q9MPE8Vc7LQ60cN/LHBhbtsofXNBhU
5zgAsf4JdWCgqREWfUx2Up3Cdw2IKCKuMbdT741Z/K96DGtfyHRTue0UbrPgpU4ogF8KBjB7svsQ
dsYuJOulIWLnB7GnLvcOkuzBiP9edCqnK/UY4o5xxCtOMYrX3XBWD9eXipy1xikG/9MwYTn8KNzT
4EIF5Ht7QoYvKYpahYOl4gEoNhPbc/YCf1GPb0rtxYnrV+A4w2Dox2fhFxzASVrKBbRYcUy2p4yd
dwJs6Ddd58N3eQ+ifGgMbv84xd1CJDxPBtXvltGPh2zRCMMvZukQmWB827gpubTA1WjjcVgq28RK
MUkNSjorCm9ngGpQUJXY0dLPtjI8paNiKt0qVhbTLRym/+KCa32lPQvaeN7aTWktrvIRIaoAi6AU
O83eQGfddRyINGJIiDPIyrWJBOuuGYDDD+wmExDDrGmsVFSVb8l5HMpVnNXtsHwygxLtSjZmKDD2
5Y3pTqtylwAiTBtgLe3HdRKlpHGOOGYYoWrqyLRbXEeyUTQEZLQx8pj4iAoJ4uKRWlLZI/5q3jn7
azgRKfY/lRGQGxeX3SY3RGFde5UA7J6l0Su3lhWFu3+YtECRc6m2mOpWmjphqKQhDqM59p4mkpvM
AYq/m/168U9ssVdgMx2oIw/T7k4bkzpSRykPCnFhsl2PZvg1fUkJ+bOJv9sJxBFeqx1d2EBEaNBA
Cznc01VmADlvTMf40Uuh/MVKdRqm6CE6MecZ0zWUq10T2GICcxqUbuKblTG2RzsM91KIz9j1Fc8y
9mRTPtXdlr0PiNLtEpUupkkvu2dFuerZyi70SQ9aDlh9EWZ36drE2GYpfH2016cCteTxB/DD9J87
GxcAERgclQPU0SjOk0udIu0Xi9FC1bcP2FSYB/aumGOVB8ApiH1/cRjOvHk6+w4ZFKwi6Wj6S3If
ImWME9LKpirS1Vhuj/J4K0w/ZPgK26iZhsPgt0Mz8FJ14shPnUznCdWdLF8+l3RT5caL8ph6Jq7+
whiaYeO9RwDZPi0w7P8XZ3sxAk29VaZXH6f+AEolryMPXFJxDiDYXDnDSY4QScAzLkDf6ggLpkUH
8tCPmbEVIAWYYsz4esqXvsds5hbiG4yU6f63KTzlBf5EQhuDHZjGALXm32WbtfTiv7+hLXKOEL6s
fzJsEgHLkWUedBaPT7883A/lVwcicjyieAsijKxJHkZxpk+cYFIwqrD8s6SF+LvBjoGzV8JHPC2u
XIIl7V3ZfHL8JGRa6kihb7CuDuamCYcf4SGbFBq95yr5MDZgxP8jGASfe40G3Q3p0HWRNR+qb4+6
khdtZzeyO/V+dT27fb2G5nyd57xuUrLktJEZGlz8YhSBSTdcTVFA6CZAjjgq4QuyVTWMK/PL3U03
K8ImtXuKiqpI5l1iRyXnR0zqfb99dcEd7cuC3bLYRY7HU7KJZuTeoLnel7CkoJ+/ACaxLoUj0EvW
CRIMn53c5pGUlo97Fp2TqcaRbMojSf77ItgEeVlQB89yGguXBbWDPkdoFapRyBxm7BxXA00si2Sn
sF2t8kg3IzzdK+yKnIwDm0azeXi16KRvVEu73YSfV0VNuEkexV3CH7tg/YihQq26edkg3+9Jw0SE
RKurSqvEMR3WNRIEeLrNh/RzlsK5UBhGYIUuF0ZI3fOY6yE0fojv99WH1PIHCQx+CktFOibbww6u
bZTbRrgFHi7Ek1RY98XNbXsXyGgAXWo56au4H/LIlDMHspeq6tgYu1TMM+N76bdNW/rKNxF80aFo
U8ztdvoh6eqKvR0q9CRCYt/Jpn5fTrTcQNwi1TSqsHMy0NVcPTiX/hp2AlVQu2PPqz41JvgBoq7H
s4erFoEIfOAY5q1u15Gu6wU0hRvzltYASej1mfcJsKhG7Mfh1tt/67WhYNJBISjRz6tSWQT87FUk
mJBdgRzvNiU2aOg9awFXzypceJMeQvO2AXZ8VIEqJeb9sW6tRW1KF4/nWGNuaF0yUDR1GiXRDYS8
VrfxdDuXJA1/St/np6o8H/CTcX0NylcqJwMHx/A4joOdCQBBDyZkU7IPV2cLkapTjnRlZtvZOLUA
d5YqVKjuBtUbEPKuM2Z5H/FAwTqSAA+7yZgx5IFCeeHWL7wm7nDHvPSWgPKVo+ntNTH984ab7qfN
ujWeZB1FeQhw7kX/Cpb6TYRvbGRNSf9EhkdOPiWKfI3P68pXeQQFHiT0+BLiwEp5jJvoa9PSqnC5
ehYY3dH/u1zgblaue2NzS5Dn8TW0rSo+ue8frVw80ETBVFbpsUPuGOWxsXMj8iz/qNUNyLiIF4WL
W4iO5JUNMqPxYCfx7sBHsCyOevR2h/FZYvL7G2vtZVtYOlXMCsVb9iL6x1XvmEvRb2w7Dw+/KVqP
VYQi7RuW40LsnULmrT5WnAbZ/v9b4wMvru3AFknp23Lbs3WV0qxGdplHcicquBXbwvIQWYOY1cur
dRW7qT5gTojKfRp+dQ9lvHrNRrz4I40+ZSKydYEsCTAonPaKS53mNV/f+iq7rEJdxKOg2rkBmdht
fxXZ99Gvu52SFU5qH/ii3HIVP1okXvbkXoAG9XRZ6GClknErrX7jWDglgdOKHjO+bP0261NURLoM
DKSllSZe40To/Wvusbq0Gbe5V/Dy3CuFLLErCk+nzjWnrG5Cw1CV9E4G5+sI5Dcb9WC8K6EiVlm5
AOLf/fGRi+6EAGekBvIEdqHsZUX/2ARBYEupUeqEWqNqAltxD1qN90StLAoiLk6smTGjnHJA0Nqj
/Hh69eH9a+DchFHtUfqDIG9jnqTBi0rUq0pxHVErWOM9/yDvVJLlDKENI980TtKaayvg7ZJ5mW/X
yw7Us7k2kioc4dJRq957WEOCYJOJocTfPsqE8zb3p6MjaECE0toQRlLpZ8hKgMw0NDHiRFSWokPK
/REcwGQgWV5hp0755hgt63kgnM3rDQ/9faYQs0XnwCphJhy2AuA48nqNguxS7ESl9+x8+vJCb8ai
OSrWYgFTtJKAfulMnn8lVfFsVOWTy0Nan4BLdcHk6oHkseZtY3/SamRnWdQ84+rNHyNlQqNL50/D
u9wv/uMUm9fpwbgQr+wVn1juxtARikqtzreWtLUT4cEgxHCFwE0dbVu7lwfwxLWVEl3VCNQR9XMW
Ud4DHdyJS664l76zLeIgAVGrla0YXcM6BQrYniIwCcyGDuEi9QSjgTOaCHnk3BlS1/fimkHC8pqk
5EVDDn4a5khUcpJ9EZm10YSuyUj2XvoArRVKW5niKndafRzYu/VPFcXsgFi6SlfB9x1UnKh6Dxjr
wIYo9q7qoMneJLGZhw1fsWpzpVThIMAOk7keGMi8VwFO9NL5a6OY9p3dbCw4/8+b5TLAQCzCUllW
3Va+OQdypIZwUf999bHuCVOMnk4bxvkg8O8uvD96bA/7R4U+6UQTollDwgst5ABQcjBPNT8atu0d
zle2Ap7XcLpAO0NR4VFKRAf+PBlJrwZmcxX3TP8ALyno8jTJWh2B5voZ+WzCrOHlom8GXZ3VCEXP
7ZRa3crGKlO4Df5e7RxE33PGdYhnemHbxs8s2xZCfZCplgWTYIKJj8UXM03saG+Yzi+5ZqiPZW9C
TU3vc65bgj5Xf7jCxPl0Wq9tWlO1+xa7PdCp4PupMYBy9iVe/DEUw5yHwB2BmOBsDXpN4sCeo+td
eUfO4vcuSZrj+zNBHeIFZ8LBIy0CJAK6kc3xmUl/kXOTOPgmV+KtObtro0ATbtI55LY6weZbVkG0
t4aPHSR0XsCKiQdvVG5UTCrZw/DBvYRdQJZwLrRf5q9FO/GgGiP86bXZO5J0EyRrlT6c3l3Ly9T+
n0c0LjfLJxyfxFRItBp8mVPVaqaAX129pCuxe1Gi+OowKOVlQwCbB3Hv0J3Xk/yx88tTBGRQabTa
J2rv65/jTido5B/pVLr4QPG8XSWK4VKLA/4OG0Lj98KUhxYxi4Nil56zPhTcqUvZbY9safWpoFH/
VtgKj6l7IEpUZvwiT7vM8k13RU8jlStnn1jXwrIgdQuzaBtPOAoUuhBU2MpLOKY8Xy5bvUA5COqm
pnEDPYGldZHyUoPhluQJraxnY22fMqy9KJLUU7slcG6tqKS8wjkVssO1wcyetGVmJEyFYOIEo3cD
b9UYd5pxsOUeK/lsmMwqzELAcfWVuBTUR/Ylms0OQ1PMWGbIDpGLR5VNu/nqhwjM8+Ljce+4cmNS
DAS1qv6JJ6T609sRmQ6xErD+kaBglZlbfe/k7ZjlIx+LOxFr6TVND3ykJ44EILAcw4WYLtCdvCAl
eCEVwYUKiAsqvPIpsNjIalgdURbpb6hrnV7GlPvgGBMnjkWSTAyzHq6qWvu3iNll9fLBQuKbbeKN
D/DdyC4XLkBihsl/QTss6Gn6zhC8SBPHITYZGKnOc4JbnElgF3ZY72E8iOhUsAqOCZHbcJh8Rpw7
SHSgPTqBSyO7Tjdwm1j7BA5x8lH8yoCnntN6VC8P9hRkcWjgoD6dCMc/QbEEVaicj5+XIsPbXBIz
y5lrofw9XT1DquBelTFfwpfpl4hayqbsHKyzvCOpE4lhA0RWcGns2pFTZVcsM0fN25BBJQAwvi8A
lnlgYwZ9mTFwOJG4DlNVvSWFIQMaxTvH6Jb3dLNzk5Df+a9OC60DZ87FGlRS6KBn9biMHkXPdUiF
m0DNkVc6EoDwWF1bfBtiPjchpKPGDvCXPSjBOqv6kMmXbO+aDw+Aw74I/4X+B2v449MGFjNklT4k
2K/VrMwLEvUjaBl6BfNlPkZkQqaN/Jt4AGP0ISMfH658TmQk4KlD7sJFYBGZVBzXqb5Def1vHzpd
MFSkyX6nbmLB3DCktjUGHoNhJA8/zJrexxjrxCnYObh9A0iyrQ8UBqozv1NRxLmK4mAKEbOQEYdW
L89KkeRjzFcjSSbF5PNoFySJqphKnND6DydHBPKFTc3YBGYwvjA1GRqWhmbsbKImVGdsHfEokCcT
Qr0UATeSmB+3q1h+e6wH1pi5dyd0kRUc6fjG4ag1AjyiulJu1xV9lRKaR8Y7oGCiXkFVQVrIXTgq
ca+1rASQsUzPwE9OOTSFqI9jOfjmxhu1MbRqlxi9SDozyHV19GqKBtgTi/Hw+fQJQiJ2g0t5r7UD
Qu2iEAcLbG9HGoYmMaP20uKyzd8XEjfoQJIo4Luws3HSxn20KlVaNUWc0tEuMvkVFUjOA09Ymj6H
r0w0H1UtmRzYlkfg4ljtcEM2fSdhJSimwiLEAaSTGrV620Px05qhRVXOpdNB2VJ7tUb9RkQZui26
g9UoxPdQUNnmPzeXJ4412XccHYte+VSU6Dv++ulNrrm71+lT7g13VBhCpmljMJbDS1Gt05iZDCFZ
c76qBbMljLlU8PD103KU4BF0Ntu2dqEImV+GYaRUP4Old9p3aaeTPTGM5sMV7z9dUuexhJVZKNMP
vsyOrm0iN66dXuqCeasApwbZQK1dEEpmatTdAWvPJK0GZ9nqdAc7geMghzp8MYdUsRZImzj8vV/K
g6ibqISRujs3oDq/Fkt36DoQIJjrJkpUZiKQ30DkCZ4s0rCT+/MCg5os0PtOsbFsYxiZkIwsMRTD
1LdxqlWzBlmoeZFnolbUrmnbTVQAEys4uBJM7bjhj/sgtMXSTW0THrq83mf5z9krG6TyGLx9lSer
dPG3+eKcTUXXQZZsPGkKWoYGci6f/4NGsglP5CAqHC6UBk1KvVfiE7fDoXNcv7Q6VOigy4gU/ei7
TbFK19Z6uTNAbhoq97eSJutTr79yZJzudblGpOLkULwiIJD4suMJ7u7rdeVCYWBiNBZXdZyUFCn4
MSaCTr0dyq5AdoKNbA5H59gFTDKD9p3Z/zPkcDnWPnE7opv+53LtS3vcBSY8RBFSCLsIO7F7iBIL
fbl6SWKsmWEQWsl3Vp2HJEuMb9zGoCCZ7fyrc8RTmsIU2jP11uvGWap5+c80ubR5So2gc69IFFGk
On6PJ0b3O7qS5SM4D9M/n6p15j5Cj0+GkTNswmnYd6tQMpDDdWDsMVT7VjtyaB78Zj7WrbtSLFU6
iUYSP+URLwscySOi+9cPTCsuCiHOynQyPCjtKnVvYTkkp1zeamc+ZnkskD4uBKe3McAlXWF2nKNt
x6cQ+jHN/yUKRneqyK6yTIdtOrZwe6/viXb7MwMoQw1ieyvb/CDBie4UXWEt59b66Jqi4UVMx0yQ
/sp6z408nOomg8eI8Wc3omoNSQ6LnP/FzNNblsDv/4O1HK0jirqAa4lHSSBz5bW9T02CAaakb7hb
SUy0Z9UUS9khBSPatDfaoFVgaRuS/pQEMqNfOXg6u/lW/e0ytDgR2DzrzS31c5oWVO/OdA6jeNoT
UPBG3doY7gOkulbch5FHE9cwH2iGti3H3d7TKdcA6kGtJXIY4zwfNHgNrrOxATtqDp9jQPIFBcAv
P0lF/OYQbGEZiEBOSLHEdiwam1ond++BqRTgVEpw+M/hzPkH2s8WJ5RABr4xrQQbPERF3wl0mC4u
6bXoMOthJkwkNs2QXRJLZc8wfbWNw9+CNNTbhcRArO6DJJgsaewjRvh+6j5YDPMMFqG4LZ4sdngQ
nfE0s6a0jfu+kU5MUlH9ehDQ3l3phuRd4nPGm1RM8N7eCUOCpW3NkBASB9zX+7A7QWqhmYjniinO
g2mEsn2uuBtfUyFFx4SJ0KMdEytdGDCxUI/4He+YTf6bad8Vg7AK8UkaautYVfbVRwcLYzsX9H/B
GV2c/7FlLIwXRxSK1XaOAjUOeBcUUizaucKqqCXDaVZnlq7wqKF3XA2BtnDvo++jUF8KthiwUWou
DEZDdJnlQY+u13mMVkBLCHN5DaVsEz0FvOYEhY5H/4Dz7AM/ZwE6s75TohgQqo/FbbMBsxE5bVd0
80OwFQygV+Ls5fs8Tk+fWvg3TPqs4857R28QDzB0tNKFQyxGziAIuh0WHCnYtQYXuN8t+BUGcj+J
KDNMBmo5jG3hA7I7v1UNicPazXxQ15Z5kNtT0sSbtMEd//Wc2WU3+7bDvZUr36+Ecb/uUY+mQmV2
FSl6qFjJooWoB3ZJQbWO2m10vBFji1wAsdJUsFuVXexa7+J4HCRPFkLT68o3CMa+zg0IC7kooGHH
FGxUdoOyPhmSifVV4eXtWoGWagSDq4CXdxyuerXadOxRpCx4YX35PhTT9f2Tz2bswP03UqRhPv36
wopNtrvVaImZrK35qaz89ZDf4RiZ2kLeVind74a//XEeHm08/Nh8A/UrcrnXKpXqlyvOn5lClNNG
LjgitCRIWZ0t24uKwJdOpWivBR5EHglv5tih5m8tNKbfwiHwS3/rh3DEUhyMqC7PUUuL8PSG4EKF
q4wxpxSJV3kln3O6O/ZHoMitAywxFZxcM6HocrqcOWjrab2ydZYJd0deqFnf2jZBdHgcxLqtQ+sm
3YSzz00J8IHwgEl969FcGc6UffpiGgb3qXgeytBduvZ5mTIOoQTzZFp2xiRzyBAc5yq2zsTUtGSu
opKQBka5/vDGxyYqY+AykX+IeZENI9tNYXImaCVwpcYHA7cTaz4AOmYFS/GA3u889MJM1dkCiTfm
PQ5ajZOTME9MRrhD/+KHHLt32BVgtKNK2EbXkwPEwXNxZcOR6LBNBlHIRfP3egYSk4qtBas0uaMo
HEEWkoOqthH+WT0k+XIIMse3kD82B/sNeW+f19r25069jQha36Hzktfla92mF6aOe8wQ2j6XKFCT
VRK0vszY0+R+B2ZnFeCqp5QfEX4pTQYYITzHoi1B+Hwokf3SI8h6BrgAeXevUngmn+30/x1oyf6m
DkB13RdUpWR0/W7yleLIDxgAu5YHVFnfKGJ4o5odQcc/le7SAYVfK0AW/hzawPfYi1w1vUUK8pb6
DuyPq//ffvJqd8ocX96TuFUxpOwMYbkZlZxmolBNhmHKv8vYgMU/PzUHbkQ51QSrCGxG6cfW3wg8
grjRK0u3N2TGT6vP76zDuCKQTg+SQJgJ87Irsrfs+2PSIUoWEL8CeC7iNfDSxRvEZVKTYLa4OJuZ
3iWybVPjcLExYndnC01xaLmuVh+3CEZaa4MSm3AdnQ32uyYYQyog2OGo3S0UmHY7KpqPaOsZXN2T
gx1JnSb+xmUAFeo4vcI6OMQ0dwMDHfXP+vfTphNvZfM0RYDKGYozonqEcnMZI08zJnAFU5zcWf0V
n9spnqyU8OXada9BhjdTj1Fiwbyec3Y46IjE9Y/tE8FgJna8/eJnOZ1ktCW1LJ/bkpOyLn0Xs8Ya
OuVvFTiVleR4QEhL1gizBa/r8xQ1vQc5hzAwsGtVwrw+NnD5/fRAEEV+LXdFwec576FGjtvK6hSb
vgtW+AQl2PoieMzDmrzm9V62XLxNGOR/yKDqMNAPM3ZMpO6OJLygNi3XMyDYUmwKRHYUOyeRg1GS
rO9RPd3riqjoPRAc1aTtaX91bvDv03aQW/BEthnZtWiaELwK9YUFvBWXX6S1Zby8py/xZQphaNwq
m5UgnQfS8VP/4pk1LSe6tfzced0hSqVX3lOtSRKTmWr4BaayKxA8oelJEMAEHOk46SZyLRNxm8XR
xAJZmSO892HCiqFJiJ5sgR5xYT/nipOB2TU9jARciZXHrutei6P1sj51SNGHCT2AGQ5b0cnIchlO
+F74ahjlBN3l5WX4N1YqiT96WfFx7rnmHQgeCWGUkOZqa49N4/7ioILEuaAvRJXfOmskSkEzp7t0
1kMgW4OJ4rb0sSyLpvt4hsVM5H3FZFcV6yXmjJPLgmvM9ag/3r5vSMOOP1Jj6Ky6OqSfJGOVSZSA
z5KeTy3QAr98kVVB99Oxy9GiyyNsDO1zRkczd6m5halGa5H7LNp5JhiE/3IuLn8NndY+JeOCw/+L
S590V0vDwDHG3eT7UDDwLS0T04ZDh02+ltDD7hLgc96O9BmkefzJvAFAOIdO3kfX8JvpmZxM+JdU
jILM+MQMFmX1P04M+Y5pALthCIrAeYEIdyIfMXm5jGHkqGaHFh9Xs+g3c7Y3x/eeFtyc/CcWDTl1
YwL5+JF/wYNAB9uLFlqkd4+4+R/ietAlfOIknXrv35Q/Fr/RvyO29bu56YJDXnlpKxVllr8oej0M
+SxqDS75R1T835OkGevEL3IwCmFBHtmbOZznjL6jFYrWREyiEE0WuyaNk+PLGOtrN/NxfGjombPX
hE48fME1+cEbjTpak0ZCdPh5zZd5fOpvNl39F89Vk7+L7j3BZ2OFIx+JRG5+UsEGu8IIYoSkJpvc
WM1lCQdeCfyWZR81Py5LqkiaximCBUQ0gKlrjlJOyUnGjra7CDcmcW4Nav+TdXMbcUxNcKN86GnA
AXFvFYWA9xdzalyMCWcLeq+GcWvrUL0gviyg0o4rcVq/R27s/ucoLRdMxOuOgpRhRqUp6R+pyKS4
fUj9KorAf67JhwaAHWenOcjExvU21Y/dIfFw5TCY3N/WqAVKbmQ4cS1xaHUguaNLeybY3RCSYkLx
c4VhWYWRnXex16v6gQ+1x7bl0wkUIBfYt97FS3SlNAwuRy0gSWi2dbZ2+PpOwzBZWlHlEKRmNCaf
U+EuO6tmnb+JRROPbFu+LZyWeufpj1lmOgfdf7DFrkUqnfvQrf0H4hdgxAVXypUqGJlH8VwGmAmS
9xhnJrn79StcDd1pqA7LwlHUbtE1ah8bJ6Y0qr68uy75jg9bV09Ss9zItlxVQZ47osHe6885OGIl
A8bcJitMXn74j1qOUnvsfbojTTJa68xb55IqLFRrpV+Xsglc3othFjn4veauaebfd03RuPjhv7UW
hn6jdA1jrOgRQAKTR6frXKWvaPeXu+JNz9v+KW3G/XIio51fQHhuo0TC6S+17hRzw7ar1Rj3jaGy
EpQclfNNmQMZ/5dr20qcF3ulgPPrXL17ABVgY3/78SApheJDO+as9TXtcKv1vMhMtfcQZyf0/Xcm
pqvhVZUDJns9gOPxHxfgL3p+sKOjY5j++TMaAx/N5qhl8MFjYwjyK6PiEEEZKMr9++Go8+KOLhKq
yrXBfDvcovo6uK+T5//ILVaRjZxTGKsy8XS+zp4GmPXD+bhrhD4x2wpxEG+tt+ugErM7VgZHuUt+
fxaHoB6BD4RTF+9c7ttirajAzG0qd5BL9XoMt41wbaRmPedzpkpgIbe1xboUHhZ1POL1cf9EiHVU
S3fao8ZMDP6zD7aZGt66KSfV8N7GDCfQjTTJtOR+RZzQfSs8WWvCewkqJ0OxvBj5Ykm6zgY8cno+
01sXmk7KQfZ+l+9WZrJfiljBM4klT5ChwvTKbzCMBElo8HRLX4I/w9CnmaHgXHQv7wr5YMXxBKMN
HSVvRAonIYJ3vj6RpHZx6egymljhUOjIuuaCUe5t9iyAFKEj5RbIHfXJXbZ1g6HST0asxjPLuozk
J3iU0DltGr33hmOwRc0YSc5w1rGhmVq+W+baEZnXSMykBPNbw5SSKkxEXde3oNuAIkdo1+DOi4EW
BtPiUC+s38hgQORQRKMsqvobJ7LWQj1x/YxugFx56WVd5vEYBOsmVOeW7QljmzuinU5qP3YR2XUn
/5oEK55HEdxLHBloPzqoWjNdCSvFLzL6DWxjuJsbP//TTCjd96+YvnsLTvLoxxQI6wKiWY15WY5v
JJtocyx2dC+FX+QT4kVIF8Zy1g88IYq9gaSeWsOdxwiaLvCZgcFwwACT1ZRHLpSKoDsJZH1z+2XV
u/2fqljolC3EQKdOyoBI7IThNXZw2YIzDK9bQKjxDFZ4UY3ExSSId2SQKLtw+u05eUVxUDluT9gB
b43bvFp5QFBrfOaVRg4bB0l9ABv674YjE/fD9QpDySncMmN3Cd4bX40FIC3HKRamcrZq1k00K5WL
YioX5dih5JEhRpNjWFuckYLoqtMuLo1DJXER1+R9n/rZ/BWFGMP4uXtrq/GRamIRrCLye9xk+31/
KJspywCkBRBt8rb9BcDuRVBCwy+MyVY4PgzYz6mGOMMuk0bE7oVvXljhXhMgph25iFAe68jQ35cw
AhKnYMVBlqsUbzFvua/uxLIKOyCV94hhDIpVBuqqyfZ8NTtEmlTKxVhuwV9/Evwd4CIpF4FQpFAM
Tst8QDDqH9BHsq9BeNyJAiRZRuR6SSxswu9+siayEqGZE7LspIF21unAMaJpffOvA3/Ma2Drb2ee
YUfyW5YqQV8gmQx9EhxpxmiO+TH/8C2hXzzDuh0MBZaa8Z1nHRyX31YfFUenm1PTfv8B9cRx1TNi
+lRcd7x+KYpuRvBH4Mjj3htgjWEgMV0NuKhMVwg6RqDtF/5KMG8kQhespPsqtLePFjGdygydx9pJ
do4rEYqoIhKdc+HkZO3lc3/SpNkO9UWapJF0icm/LE0cVsBBZgihBE31cXJ1WUpvzWKjTpUctn52
JmaIk2EYZaQzwd8Z8S6LtptdFqSCmLfVAQUOV74J9iQgegUh8ll7pCU5YQeYEnHmRCkRiuElNFe5
ZNXvO+9VuWnSD0MSPDuSkSBtS/hocJaiN0K1xFv4a3NkMqLTEA2RBDF9g6ZpPwytOGMJgT5t3UpC
K/9G6b+9Zk/zoC+DHSaQ7Qz3bdPGAc7bvJZXnSJQsy/r0kUnQYTKImcBuD/aYxpbAcRuEiyA2ZhV
ZmkNvFt+9uZA46q+Llr13hMVXDUMF5IKDlnsW4BkpqfDVq4QX5Nk2PtTKugQaN4NdpC2EIlCBlAo
vTNVYEgxUfFfzOGkLaxLA8BAqvmShSJ61rOGqH9+TiB455uFydGMK4VCWAAEewdgaQMPnIUhTSGZ
wU4WUVmJJi//Nl5BmmfrYkOpDUTm9tVkM9yLUDh0Fmin7uMIIGUq0zxriVXt2eNrbHTH4HxNOjw5
VxLyAD2Ad9XiElYNC/MqImHGpwfx7IKNAtMmSZGger6NWw2Js1vbfaOA4yHmS9A+rHZZhEMvbQLV
IhrmmJxFrYEFezaVnt4c3A7I2t3zn1LXx3l6VZhHErjYyLDkAbFF4SJ1IGlNVXyLEpHBYHCO2X5E
4n8gBn2SwU/+3luKPYbHiAVH73Q32WZMMN0rckD5XKzf4yW6glrB9/Jh44/6aZMttn2VFcgziq11
1aFRvDu8cG++Oy7FMjVXjK6TEBXf+uBmHCZ9AH/uvYMMQBZsTt6BDtmXvjjjxck8ljjZE95y1XcP
Ba3OnV9Dd0Kn9GAeQlk5bMm1kAorQmFWY2o5ciNxN7YOl9saQzkTa59aqOMwXvMnKCUq3A/aaXYt
5u82ADwk1o/M0fQelWCrpvd2iDpw+3Cu7A8bN1IUqXX4LH19R+/OHhbv04cCbcvjov3Bclj6OM+S
LygjvfKnPoOOdCPh/JQPfVRtBqGra1Io2xORvCsntmZuh3+Yy89aiSRmkGbUAtwFjGEmGLe10agV
M5e0ccKYL/su08ggYR1NawxnpsrXaZxt3v7o7Sun0DafTmuE7kvhoVG9WN8ehjwBQSliD944HwqI
6Fn0NJlCV1CodefrxyZsNzdl7SKMw6QkVB4WX+bXjIpGgMzE21Cjz58UqHms18rbJ+Dh1PBkAelr
OHQ/mUwe+RtRNZvhBGXwNlqEUrPPuGf+FnVnmUotQNcm0YdQ/RoQzgokcdqOL47UQBOwGAprkun8
89g9F59w2H3n80Dpt4lXQ7lBFg7Mvm9XO8Q43UHrRNQW3f5NXoRlgopPDyEKWMtnsU6ryzBDYqBo
8mWmYb6gHcJuHfUP7vAewhBeyrCjzXJbtbpRi3S7ipnTetWm+2QJf154HtZqZiQ1fcj7Ye49jXEx
m2QJDYy/tZsgMT/NYDmtPvTd8+SqdsEghs+Vxz+78T1ZLEfGwon9z7ItiF/QAhX21jqiMvYB80iy
wXKHx5DvCHwLfSetQEFzQFD3+nlRcWH28CC+rRp4/YbJtVIjGorRQbmkhDFY8YgRZSMioKmjvxP/
kKX9LpCFaeYFYdpBREE46KrtQHa49teP4Ikhn+POGslkGNTmNjUvOlqSzRGJMo8eD5mSAT9PxksQ
NZemknanqlgRPoJkJBXuxtba4pO/cbYZST+fsHZ6zROqBrimq0Ll5nIaFOvZUB2JISocZu4SHZYh
XTAx3BIZbcd6fpodVQulbPj3koqTiwIzeHOkP++08gPzzx0Et20hnbB9eS8pyBAJOn3hv2vHVDmy
FOGyH3DZd20NQnjJ8tRQp5k+n3abLd1lyN1gA5nHImZ7ZkCRoelPjnhzaRUYrW2niRl2bT5qdzGC
nF6cgDFMIKMUqKfSut+Vvh/NSqh7SD2qmG/JQ0QYmm6IH5iHYJOX6zM4V34vGL14xLmWtKyrSrpj
aY/wyki07q+arBKTIvrHUL7ncxRGofy6b+QvFSnhjPez/8Ins920ePP8SUFWiyH0y14Wspfh1xZC
pBVb6NSCRcJMH9f9pP9bPsmoUnzIEoXF/zLRCkv3XM2sTJ8712LQuPnvPGMPyBpSewZevYpcOczM
4PkFCJSjGD2keWr4x04A2bCUObO30WR5gdAAGpK0Jr8GV/YPIgBRuNrO+67z2lIdKQ7w/PhRphld
Jtnd5oLNclUu/kLWKbjlK2EgnO4Tmc+ClRHmQj2yCQlezr9X+YEaD8nP34eaglxjaoh4UMfKnVTL
Ztn9N7YNvF8v5ZZr1wegsLMuLu7FEJdyo6jWqb5Z8104sqQVEHlMiSL1B7PmMi3d6rhDSM5d1p4s
MTRKCKwAX1C/60g6Ih4VGbaWPI5UMXkWg+/f4DCnMdRHDTSUwtSHJHVnPV6FymcYwaxAj4EHr0PL
KD2bLoEDf2bGqglvX9PDyxqf608t8MP4R68vQKdxll4FiOPfd1S1EcuSWo4JM+vFmm/I+b4/hgi/
KfGiA5wOdRaAaWrPztx1KniYbYyAsuh43DkWxhnA2/c8GmVLbMwQm16Y5XydRyI6e3NyJZfiDx5o
RN7byL32o/HCaWXNDtl8h/74JQBKk44Xynt4zlVwoePrtG93CXgoGwbo8bDU4MB3kXlQUILoTshf
HWmqEWDxfPpKlyjFea8SkmzCfolAUVw0ZCwjcbimbMFWH8UXjuuy52hBLf7bg3Kl3tu/JzDUJA2e
rrFRBt/KH0kp1VkWP2n47l/izTvG9/4q50QbauRAkrQdPWjRSNJERZpnSE4tPe5KXhu3sdqj/MBl
4lG45ELNbnEaJn0WF/LXxSuax6QFAywhnUPO1GFpxCh/QjaJoSF93pdMV/mYStpdK18aN/z81ILV
kDx7kPTzAvKpHkeALa/SblPLoZL4KNPF3Cz2nPVcIFHlk2c182bbBc9gMwW5EYmoOq88nLWLUW99
zs+iXKwdz3qRhQuUGYfkogqtBuNMXQcKX4dkR7LfpAYj7Mx0ld9KuFGdFevQIZ6G5imVXaEVJ9jV
au/RP10aO/tDG01lCGy2VciCsOfU8VA2qHeDhreMrDGDpf6x7iN+8eNPKJwRbQv+cfd/iZiCkFL/
rFMXra6q8pr8yLpNs+dQm0F9D8YYEmQ9/U1EGSrwAth6Czae+Y3g97n7HW/5GhbL9QdLBykjfNkV
FJZKs9A6hCqK3bHX3yhm8jqGAQcR5FVePj+5qfnjIf896/AgiFW+S4VdinPS8IAVAu8DEzp0dTrn
GWUrFavg0PQ9u9t02TI1KSH8eyI9ztnt1Jl+2iueDZIwqDnx+urwRlcr5VSpbSr+Dpg+azy07KaI
e9O6JXGzU2pOdM+LPjWtJbDpt9to9rUy196PdZ+CvB76mKlMQLuVNW7M34tluJWYzlyTwLWzTfsf
KhLhLvDcd4C61JqrpuWysjXLm8MkGYUHe/wgdMPGAabwFiQrGw1n/m7mGXubd1P/7vca0GVDHKqM
shG4FHRXcSVIs6ckIfzxrZohhAs2uxMen2J3/4NrD/wqT3WY/znYXkenTdI4MrOlMCpRUhMJU6C8
gTTYv2JWGssrBDH5SwuVPsbG8F60ZYeKRxt61e4CRtgQrsk25ZMXFnJzwEQQgaI8bzGBL/17aoCM
PpBoV6s4djtm9dxOMhYIjlBsKMo0v1ZNbmySy2FRMszS2OYlBwzE0h5SqjquBbSxzZjXk1WlM3Bg
88nGKKtOQ0opabhHa3bac97cowrQsVsi+XqvAG1f/lhnHtEmDizKNkhKtW9Cp0LmCiiKZiN/bNHO
/TPmbxIuP3wpG3aWz59TxjtMfdXU2RwIfJNIT1pJ7xuEFeXrJQH1A0VR4wRH1B3VnBbPbTJssApK
M1jbedgVm7RPcTEngirKTIQ9nH2he+iaqWcBnUd9rBqIfkhwKZGKQfQyEYBD+VtahCste3XN6iPr
vc2X5ejhoFfsW66TNBgV505ZOqzjzNrHWyfUc5lrcxf3XtGm0LXrgPXo79Cd9V/8kdbNRw+nYJL/
skBe0aS6Athg+5cw3ljui2tG++7YvTPSVMtCgSVh2AZqhlUvyB7T6cNenOTVYrEKRz3qTimwgqvs
iJJBZccLtsaV1nf0T0ScDDqui3jmxx+5JHp/8z3F15Gnc/SFi7d/Qsh6bqA2fHTsjRGlS9ETe3ek
FQdKsGY2/s0xEuGeBi3hjUki996p4c/MdUVgJ8DKyL8zxXD3P5oXLDCEnicgZyvr8d3ljnOS+TJj
XXlp/qo4tnBoXg/0hNduZE8ivCHlA7hx8ndiWVpNFEnwy2YdoH+31B5R5fe4xVwy+E2uI6LaFXp+
3RTFXnmO86tqZ8kLqVzcmgq40AYS/CmwiQSa8Q0ZMOSLGgE6t9HBAbJown8n6Gwe2uvYyEBYjjbd
8CVtQ5PGNzYiBwEhrQSl94YSRlBtH6ErPxbjQeWLfPUFuaiUu9q0yp3WUIfXgiBKbiI79lEAyYW7
3rxp3BZYTM821mG+KU3qPtC+FSemnw2gRMeWWFVpWz1tFwlyB9wpGeQkPlbIo2+++2NbCf31TflG
RMuL9NFEaWgfsuJ6McrjxRZ5DhLD+1CUMYNnIzxguShkv8ftHOiOVppyKAzdly0jzIX4eteBEOyu
lZFbRoLPyHDA46dKCnx1yLBuesBDwD2+YrPwbK7Ckhm2m134RLI8+XuaoSSRdJGRkpcASwaZukyx
kZ8RzRb4rQyKBZMB02gAKhXt1zgujDQ6MxsM5Uf6J7O/E5+g8DiytpHjqfUc9GHNQzLem2dCjqoh
x6mVOIjY1lO9eXrj09rdJg49vnQm3clu27p3zEpSZS3P1BIE4eKn4xjrU6PdM/utUYsJs7dNm8xH
fDH/YyO+lj88WkhHdS83OVnvs10AMrJYEwJHHCd+IIdGx3SbwKtmO4j/1jYV5oEvHKYL7n/8A78S
wCN0aklgZs7fLaqUXxNCgmRuQFKSfbsqNfDOiLvpww3jiQw5EFVjMs2bhIusPj1o0fdncPzvn+/u
eDk8yKTk2tRcF1TPA1qPXgwLm7RB6f97YEndLM9R6FtXy8jhsEtAvN08O3ugtf02011HT7vfIC99
th0Ey00Gg/iCboF5LC6rAWJgsBYgKRCDZA/gvYIC68feD42YXpUwdrd+adrUfv3r2TLe1JGnnlEq
3va8dOjMTQDdAyLG7ZjwKDPoACEPGbzx7p4yJlb4lCbMKykn2vDyWoygBjizY6L6La488Tb6Iil6
OIuBf+c96Qi4sa4pQS1v4OMR+IQqchgAa8Gj9WhCLCtHN01NEgPsIfNwhqJMduWRFaL3SDpblLVw
J1vRYzVySKeOLRhb3Z99SHXqf0aWwng4x8mMK6QcqBHCckRpikoZmvCeyHREWJutvnXj0fBCIcvm
F0VUHmYjSTCb1BAhMejXrLOoH0xuVIWtwazT+aRmYUq74PFRpBD0DA0MAowlXLxsq4w7AZLTTeKD
WzJ2IaTv31HdW2WvEgF6bMAorup8Ter5ad8svu5LS2fR3EbECobPcFDY74430LC+cDbnWEn4qEtc
e/47DInGzLFQBSoHQU9iyOBfprAblckNCNKttIQ/M0+PoT4Je+skaUBBltaQuYT+wdCsILlv0rNz
YdiUeHy6LllU0z+c92bR6L9n53UPUxumRgynQh+GC1lAvHqOwi9A7F+UiUby70H1MX5U/yfj5BFu
n97GHvHYFhm/mjb0nBQcY6OZB4Tnpm36sRFQ6rVRV0ZHZOVEbbMSnepXed3LoSA9Vs96N0evf2hz
3hVG9XPoGn+1EOojMICoUw2cR2nP+2bcyZHGTAvOdlthdsQRK22ciT/Qsm0Bv4DcOZgQvMMQeFhv
zGXWXFC+n2byT1973KPHZGSyM7t9Bqah+ybamIluZ74GDqdwjNYJStfnCe/C+W61cjmNvxicp+7I
mP637LCk/3WxpMWdJ6Ej5V9Nl9Bk75na0exLLahQz2i3aaIzrcXohxe6g8EkqjAdzQx/iLYyEDGN
aaiZb3YVmsy+1/VKYssN3Rw3+h/0fmrcnK98EvpcKaQS9rkXTRb8iX1GlXJhhJAhKMNVPk+5OfDV
BqZR4AXBXh1/S2LsAp5fC4vvee123Z0UDO/zzrHzguqgpmdBKzJYTRtCPRqOI91k/QnYzFRnzQka
JmDPWvl8zh4cTABVAgX8Ou5TAvV+dQ9+p1R5Dj5+cbWhcAKHaeLRIbvlBg7Y1TlXPmhQo8qDMXbi
jmLd6ONICo1CY6hyNODXUCXsE9DTyBy/4B0ouyNkkzYD4H/E2YsviV3N912TU2H2RGXA9uL+uNkE
rCy5VWUGHtfS3tip7bsIlWOmBL0TqZOBnidxxZ6c4goaFzDhRnM09itmwaV4th3FI86gBIsSD1tk
w4aiPOxKH3yn3GP9f2VuybWXqTtKradWP6uddTN3g/jtAEOVZuU+X+DtJJ1/xk8UdCfo/12VRnGy
3Ln8lTYdQ6DQ8DChXgvZEpC3OHPxt+FoaDoQy+fWAxufbRtzGuiYAz5T+EBP5yv4qCEM9mvqzUgF
dVctJNwExyj+GkJCqgBDEwY43X3BVfj21x0hD7uyaEUcG4yFmFL+7Qqu+aDYhwUWpvaUw+D/335C
cHqPRBaZxylCqQjwaCnOsc43YH7LSI4ilum5jmoGToVCU7DvStos7GfQFSk35WPpFcRup33hJoSc
UbBQw9PV6UYmviX48kiP5TiPB+1KIzHddqWzGOVjuhhfg0dAEVjlhAOglkbnqxDFbJRjPNhETArV
t771GGVwjsqdVxAS2WL6yqGdJFf8hjk7X+ytooRPxshqhpAw/mRyL2zhbsx0Ymo7m75/Syt8zF4b
0GzFEYytO5kE3EyAB9Dzj8iIEeq7KdVQRJGabe13DJN4b1rXW166MVbeK5TL+kunTZX6l5d/QwXt
c/GQpi8TeW4C8Ysuu4FdMHk6c8A8XGulgPZp6OTYO86BmAPQXZ/ZO91U2zAZ9xAkdsNb1qw+ataC
1/o7AXNWuXssUqekvTrrZ2FBiBIr2avPMJ6BpqWG3bYMtDbeWc9Sxsk2UIa5MnSJGGmhMQyvs0B+
2D+uqQzY8SCiBOKkl/VANGJgk6ogR+GgMdNlFIL6QyRdEqGnAEdomENBY7Y3Sm2sUO6FtqHr9I/7
SimXa3eF9JjuZ7l6j0DtqgcsP1JbOYeCVfhjbbbaZ9CVagqN07waSefxTQJedWSVjI4Yzfiy0jlT
Zqj+9zOTuIk+hPbxU9XbqBmAJmJ3i/LBVkDy9ajOIJDp4Ka/N+PxNIlpwsuhkSEmlmP2xc/8Va06
/tGKO35MHYmU2NDBwSqiaxHnjxvj/6dpxtUrUZGnyh581LHAAFQ0HSlDqrra62j4vY2E2owcqhL7
IDL4TfwiVoyFpX4diOjP/3FrxkU4m7Nxvzai1GEtpUoITd20jdI2Eel9c14O0JVrHyKmmceBgwhq
s6q6Qx0q1y5SgpI91Xqg5k2oNoZqziIioQDVdsn9S8HPGqByyKEFp7EjY+gc/VcXRWADcrEN7GGj
byZwtyDKTcftAnbYTbhJtuAExPQhs9KvAdw96usSLGGpX90k6has6PIIGwGjVwsGhCVyFEHVJo5k
XI/I2/2Rtosd79E8PhufxWWNJJv5JiM35OemDHS56Ugfp9SeU7hsi6s38bEfEha5lFiYDmnVKqIZ
1rfRi8DJn7DPuN+eJo62Vn9jXzSQCkTTuSKupEVXLzkpXYFeb4i3qMHW+ntRA6z3bgRsSRl5QdIz
9ukPI28vvqebeESzU31aAPKPjdFFQ2n7VOIYQIG9/eMRdxk7fqD3DXRSxh6w4Bo8DQWWpzUZVD6d
lDiBONQkvpvkSH01kQ45uJdFygEzNCU06wL8xTvwMrPfFeX01Ziqh1F3DaaJO3tev1aayP5X9VHm
YqDaXXUbrx3pB5YEGQg44A/0gXZJ9sKeWhNd8azpaKiK9J5dC30PANo+oiOaGqMAfuP1VJsI8khG
apEvy7EbMqGsnEkCzBg/DOnC6eFCuZvJ3zmhyt8Ppp8Wr3oZd71OnonIC849EtB9eIcoL/xVXIt9
YjbYANcMqc0aCwLoDBbdvQt+Rl/tEzbD3u/SRykaVuvn4ejjvIDRZO5AKY2Uui2ZtU0Swz1uiX7C
Co3Up1PEByG6L+4roU0rbo9M7UmSb61RfUHsTBVRrw+Wii9lbnxoH1yfiC+u488lxImiEFKYNzG+
3gA3JE7/4pydYQN8N7ujQboaXZudgqDwmffitEX4j/3t9BseBgeiyIbbb7kMT0cVlr6lbVOYHRk/
W3ZiBfB3cFXniixZKv0v4pKIWk7RTDWy3ous88+APQ6Y3vu1oWy/NAqjV5DhMq+0M9y2IzmFICCs
88Ha34TQfxdhD3BluqgYunGxVG7FgkyQqAIPEGgUI27NudZ7kiwteR1a6mQpWRdsdtJ74vTV34Mn
BAEh8NVaKGQtoeqoA8YPt95afi44/aN7GCNncKBAf/MN5lXqxaFT8Uu7xqP7SX02fXlB/dgHuZma
jJQw9ZLtpu+5ifxSo7UgiDc9W20bdT/+P7A63f3tbOOykkoJlY334DsC8r/m6lRWQ9pgvtJqXVLO
o0Se3Z163IfbF6p0XxTdox6U2JL2r+MR5KTJz2QXhOfknvT25VCDU956T/ztID4mUFotwy+8sNY9
sWSS72bH87OD9dWU0AAQYTx0DaBmt4+C5Cy0v0zfmpWDthKWtZeENe2yDqeMqMnHVjLB3qEgr5i6
sytkk9OouqBYFALWoXAen7nsadkAZ94rhsq3MTJ397965jCIgvwmp6pgUvkUHOX+O9mMu8zos5M0
vIZjDIhYmJ1poreWGh8JwnKdRvwoPiwNcfRpGG39cS7EGk2ptgf3Ex6jMHnL5uhKdItB4JwzaMNO
rypxKiHEhZMiEH+Oz3+uwjTh0NSBnT9IY+IFpqjqdHSO77IQ1TdfhtYIVpzws9QfzOKqLLzoM3GG
pQtNz5GQD0NIpa04SANFuyREj/4gpM6Qd3eilN/MZFGJ3szHbNpQW6dn2Fn0+0sfJmh6b+HmbOWp
wr6OA1w7VNsv25zIgKvnIsu8CLZsDfj0lcPPIZ2Y8AU5OjVT5x980p41H+FeDpeFJ5AqiVhDKcXc
4y7m8w0klvitxZKzfHqXxCUYdXUtQ5jS1KRF09ndr3NTdlIknjnmnH5wTkWBmuem3i1hhUH48E0f
2Vd7QVgls6a9Kohab4H56mKwdyuGAOzjQwOlZkQqwgYRU1p1aofhKaxFbo0UP86uA66aLF7cQ3Fb
mOJYJMGWxXZk+MCsMrEd9gf3Xv7VW/a1kwrUaPXEw29ebnP9IJLvXNTpIlEVJw/T1ZC+stS4HndA
/yfP3uidmqAjVaEwzw+pRDaHp0EQj+y0mIf7ub0ReBbVES0PtWkAWrSy7zimnz2okK1V1OWLttf+
apPLNobofnx9Pe5TrWYxxOl9r1uZfx0Uxr0PFdPmgF2Ey3xpNUV9HPCtUA2uG7zjWZ9hzNs8pfg7
pbn/o971QPTjggvoXimddN1pbXj9tVIXZy08Yt3S3OQj9wxVELDKFFUysv0XQ6bDiAchqhu0irbR
xin5skCg48ITmHlRMtYYIPzBvlGHJm7O93Z5rY0C+XNeuZvlM7P6JL/O9xyOpPALhPe5fJC3PwZU
fc4n2Yj6xCm4ZQvdrwoOjPvQRkgOAJQkBfyQqfw/zTo13bCGLaI7c6EC9V4Kt6fRd7ZDfIsJnGmw
6a6y62OVsjAu4GeV3ttwaof7jGJ/iBo5e+yIoWgevlWOlHPb1hNG80KGe/79RfBFciQ8BpBrtWqb
AWR6iYNpVrMQaGDFGzg0N4+/bghgJ6iISRQfuNC3GbhchbR/FL7Qrenr/E+E83X0dP2mF9CFNn1O
EmRlBNIdHP35t/JW4iBLY1iPe0vUyZXFNzm+zHwcRset5nOsRjwN8qaBrySzB4TYBhh+YKGQ8IFg
cikcNGzw67XPLRquW8g0tp0/e8JF8b2tV+6DeLINzOjyE6WJhBDmz7t2CZD24+aIFD65qdDkkf5g
iQjqcTf2injpbu7NiKUTsDs8hT9NM8LLrHg/dkekPJy7GP1QPcsnprxmNCroT8N0lLvwJcOiIV6m
CPxc6MXF8SK7Q7+R6dPV3VTQ1vcavTWAg6Jq4e3/p6PEsTjCon9SRWCLsd+exTfk9BjrYf+cSiMD
qcyzudFOHD5eOaqdJptOvYoyaEaNnWDOnQAuGDxRkuJLPIJMo1JZQwYDpTCsK7WprCK1XHH9hzyL
vG8TKG2UTYiAGG9a/S3ybEe2FUgrRusngJ6YLTZjo58y5E8r4+WwDXNmhMwndYooKfWPUJR31M7N
/cpmKqkseGImGAZiJIIoaL7GCYuSxHPYUIydXPzjo3hMEhz7cJq/v457sf9yF772AqXBeNj+U5jb
LvCPifCAsgq7coppmqzQN9Z5XNKj7MqDZ1D/UFVF+x/IgV45jFTsNKi6fMZWhmsu3s9BoqqonlMj
aswR9R6rdFetZ2UsRiSye0p8qK6z+8/9KeoMyH4Aj3E4b2JJIKLasrKMkJ+ZUy+bJxOu6bJ9KTvH
Gt2lOqdG1wsO2NvEoO3idNErkgzm7to2I4x9lt7wEqWlrNt+uN3igXfd9SKmnpFvgRqIkZbBSbQW
6OOzW/d30JOPISBcQeVdM05RKUHuwnx99+tCNKoEjuWOFhM1kxmBLcYmFQS9tS99VofSaPES7OZW
YYWkoTPyBQjxjbswhorLUUEzq78qBWFM6ticczGFL39O11olTRoEgIrHjc94R8A2i8z0EUptk/Zj
xWnUadEr/nirUOzwQOPI2RYAY8fLgqf0xiP33R7HyAH9KsePLcqEy+4axUO/vWyCKg0frxn4+t0p
WTtKhEmK/A0hJhT8kOAIN9xYA9+wGvKIz4RpR5ubZkuckENjxM2wLUZ5m+/4Rxn786l9uOvT3FcL
q5qphZWZG1ZlRhl0QlOQ58SEWpfED5Jzc+/Rgzgr+RofgXubK4FHCXv9HoY4qrASy2AVGI2J9MgK
ZWWzGrE3rXEaVXFqqmM4hXQnEFyW6FvD8iFb8CzzU8zyTeqyrooaZX+LnecKQU3b+GvzMwR9ud1h
gBm4D+KoqiHabqEsXDMjiapRL1dg0yrjjDC8+coBYR3Uxy/P8Rt4XhSVPITKkmDtOAZgbcouCAXj
ihFuaaJuTDCG4DYiKq8m/qzT3yPhFoSVascYyij7hkc0STCg3EmwgR9r/q1LwQM7iMdNGZAhTFpK
NmsGGtWRUF+BaHerHOrhagR3358SWRd8qB+5lQ/+ZflshpLK26d4xEBJw4i2jfW/lfgiDgbrDiFL
yt+GsUD6xUiy/HEFC7YOfmmpRdEaKhxr9bXdJReFP8cREnnjvQquG8nSv33T3bZcF8hOAon9vs6E
yDyIpD9ijrygNtTavFsCrYcSk1sxayq1ncwRIFCqLVlsHGX96/Qckh6/d1z723JQfRfFGSkZG3uD
DABu3sRRiv5g7MQt6sW8Bu1kD0DEudb5cTlh5vQ6ZkEEMIuVmyG77/LdC4T1xi0VWad6YCeR8mDw
CQ++ITU+JdJorghwRkSAo63Dzotjx8lyIvtCYBUrSu8TMSnn7gzMa6cDSXAGt6jVgCLQ58gD5OJ4
1N5dQr2Bdsunodx+HQB/WbKsIvZKj91PMhEFd0V5YGJaObHqVHMe3ce9CIzm5wbQM8dpnAwbcaff
chz7x/fq3i6h2YxPkNbFxKE1diREIVbSHbymp/SVZyg7AzizlcdsrfY6vB8QErvmovFOkvmkHf5U
aAWXVM/xM6WJG7g1TiLxAeff3lbv8TAXqeh78y1V0b9++qtOBouRKKK+8GCBP2a3D3pT46LVhbdM
EwUJTlSZZoB/nZKCCeQ+cOvkUB3HrGcsl+VilEuAArmaw4pDvsO71QuTXJURWlruNsyvUV3aocSK
LGTrOPuO7HOMuLYVnQ8X0/3hHPbLphTrYDvrn2eluTtxiaNPIH/s5q5bL2VGz+6UBc7YYHqZ1le6
e3R4D39q502NWYyYi1nE+4GsgzKzOSH07Ocb1TY2/RisxGucb+HLNGh03YtwOj0+Ao0Lovhw9TIH
qakaLU+OiAMHNgXMmsVMCc+FZfN9VvHUUvamxtZOxPoIVfVdtpVmE0bpFizViH0s7FQIU5CQ6Hyb
n5eHQsgDpuhxlT9LIWlmDlywpWtu9yzRlj70FJP6ehaO4W040VsoXyStzn1pfdg9wwIYFGvNF9kZ
EfrHGnwS3LYniFxKpzkc923cdv01+CY2IyHVA7epWfoU/8vwmPeRclBnrWLVDJmmCBrw0vPFGs1v
t4jyhLJXKV5awJ3A2jmmF/9wXCx45TsSF+0HHPP5RU3xzKCkuccnhyosBVsOH+o+In+WA8W88p1r
ymu1iIC5KBKph1L2TwBN/D/nZzuqBe+yk2BZULoCpGeqrIz1MQXPfwigaAUlz8PXVwbxV9vPuNVr
y/hsfmRepXjhK8vHsXzV4Xp3ER3p6gYf9UeOflybE5RQnKlaScs91oQ8ym31A2IoLGsh6isNLE0O
l1eZ8ZQydYG/gBcXZJtZjcOGikotSxPRd/+rKLHjKAX/yY5+K9RsietFSH2iJ6yCoTT6o3eVsN3e
SA6MEPvWMTywPeSF/i/cGqS9nHYat1krABMZY4F/IsgoqAH44zdaGvPh3yWgY3lox7AvAXmYgX1+
rum7hTatZOUDUZgsT+H9F4caObgAhL7dEliogxna3+VxXYseKpwQKfARTr5d/BpoAIXoVHXajo9J
IUKpZ+k+Wh4CJzxDF6Py7aKSNotF91GkfbEcNGAEYXdZcl4Ra65GE3R3XcvtmYb5CSJuRiBIq7TI
lJx6gySDZLDziYruZvfylln/tYruMQjLGRZ0CyFhbfZQ/H2Cx1mhuL3YkKD0Qr6Z2D4Hj333y5lj
jpXDtvrvZARKFrC5EZxC5nj+XF/MWZZ1gb6NjphsDooM9pT+tUB9W7n302ILLgalVEfOv7acYfCx
a9JCI6b/yXRJKBN/kPsTuDRK+mjUWnb2h3xAYyLUsSaGI9suAdoFPm7FAVP/DalNUSXf543APk87
ZspDM3XY8JkMDHYS4E9+CBDcd1aNGF2+aZTWtivr69qqo6gdOjRzInAtwB9/BWRE+2VvbRw/7MCb
cnz9IuzeHiXIlTTjvrHEBQDwe4i229bQc17wOTU++aRvKwBn8oKA+u9ys7OTDljNS8PZFvxaOjF2
t4+FvRuaYG09wIII87X6wg5DQ/bsXKT1RecJlPytkceLPlOaHFJVXrT5kwM8WRrAwTumxDyLx82Z
lTP1Ya2Qf28DRkItPimoOUf2Ypku8vHdoLl/f5/l79qVYT3FOE9yeE8++/ILWmS3DwrtVYNGflYk
8msZbJIA5Rkoymf3tRQxUBvUGRMg7IoElx9zXD1/rDByDeR7wpchfFvw9NTXSxSoBFp5W7E7XaUv
ql0uhCjUL4L0rfquYFmnuRIoIZsMl9gk34AiNw7lhmak9cylrpgp3iF9XGB2nMb/BoJcFKbbsj/2
qIx2DPgxZYJIuSltgS+Iya3b37rX7lf+RDnZPYBNeRM5te9TEH5BakZpoyKVNu8NvIf/Tc6a+tt6
oXztxnmC9umdOYCVb5kesYDfv9W8nkagAe1KHZMejIGBzjFNGf+nJrB/qd2nxVFM6Rst8/0O4dG/
3pa8IsNgga5lrjbDFoPahmyBtxQzq2Q0WN/sbnme/eZD/+fWq8C4d9n2JBn5apUJQPE3DlxCeLFN
UlhuFV9jN7I5SDpb57xqDYdT1xtVWEAQjTckssq1ybRovJ7e8D66TwlhL78xWTUlu8mpwTR4HRfb
1/04FdL3OHbDLY6D1vMFzs5F1vZGpqLQvIBgUbO+fTrkS1T0CyBj6T+mWrVerXvzkQ5+unL/m90Q
yQwxa0EIX/9PAAE496rpLgG1Btph9/DP0vve76AMOuZbc8UvKkmTwbF7nt+5o/Pq6j9RfFo4t19I
I6/fdtxyzUkkwJ+dye5jfAbhDJo+4HbwELBHtqjQYBkgaV2UtOoy22z/pMM0F1fig3gyPpPeYrFB
hXpoXaqmOxWrBRhGR4hhCSlcnk9CeN4uTm4iNCXjYVGMcmuEj+lceNytcmMnVdN3Zb3RCOEUWqVV
x4+Obl3Dd+cAFsO5cUH6L+9O545JZPeGAISDc/td1S1FJqu10L7E5MyxLvjJhctwbZp5Zv0j+vS7
oaeuaJljb3i9z/w3ulF6eG8uHYqDMB/I4CKqjm3cvVFVUgA13PD/GAU365zazWJa91ZdaLjQsWQG
YxY4MlV8Yt2qBvBIB9JDUbjY81lTjkKUNX0kadrZFmir0hxYFzgnRIn357fmHZ88tFdeD3L/JGut
hFULxtNPhkGtGfUHOSuxWqZysxGWP0lNUn0U7ByVK3vX1ctKhj7dFi2Ot9xsYEaOApubMbLXKcDD
n73/1BKO01Un95sZYoyT8YvZze4DwDpuOTWE8uuM0FLPfHkDgy4d5IdJ+Phx0VGhHgEglD0kYL7t
3Q2tCKaXEIpQ6yEh2mwmP36sZe82CBeolkF3dxJSUcfFmQ4ulVEyQHh25QVV9TsKbJcatju8WEvL
g9G5nMCgC9TRSkefP1xbf2ssK4hWtchqjKHclAO3eSXSzb7yChQasSkCMLpD8/nXK9JbZ18KyNGd
drDWMQSE8MotyDUUOlJH9Ai3Tvp/YkrVS/dH8n18OE+u9REsqIu1fUOKurYyFbBIo/3cUWoal0YN
jICW1Ynzd3wspVPDHHjGs3tXQgd/Sd5keOICqlBgBGpdfYuTv72GM7uqhgbdMFg9hQXmG1s2aIar
kdr5jEIO2UsyxFNq3N8cm62ksv0jRu/fUplvFRGcIoPzZ0jjnl1tA2jwfvxOiViyI9yID5wnThi2
HZNkeGSl995HY0W0Ulb5l3Uxi8AZVd18p/q0Y+vmmS599ThgxcbJhox9lphZKi7iiRzjiIhqrQr4
mlDw8NAYzi6uocK2IfXDAQ4DEEUdGj1WmwuVSwIYly+InJEcjloHLHc23a2rusJ1ir8HjSfXMnN/
h6juRo7rFl1165A46y1a1+jcqzrLkCCf7IRdkWBp6H/aRyl20+WfdeFFB4hhIxY1cJGsub5UA5xc
wJX356cC1WWxaWCx1GSrznTwbnX5K5hmEkDcWlMoyNyF69PD1WgoA9rZx4VXl3YxRzJq8xE0GW/A
dXfFhrVfMQLk66JyAv8SIfYuKj8eH6/Y+VV/BGexWPFet8pFmC6uu5gvbjcRPaUSL4HcnU6eOTAc
hyd5wHilirFZjS4qzAzoWBqo5PPYvWIGGSAougkC0aJCWztbPcII+MUbzvbXAl1a9HNtVl9xR4k5
LCGrlykGPV0FMyYM1KFXlGEgnh9hIX5xOvXb6T0MMc7r1IL4UvGkyjAHjUpdz6QZkvv7RwKlJxB8
IWW6WgKw4QXix9wZRq8oPIkGwony3FsZQtRe+Zhbmcnp+tT+/wT7ViPt+bqrepSg2hsArqiR3Z1e
Ehjd7vyvXCp8ZiKP5tOFsU2WNZ7dPLUJioEDpZTRw6+XgdqjjNtUX/J6ZTs48hcMY7bRrpHhareT
NsAn4KuQh2IcWV+/SSmNFCDVKANu6h3HdSw3Mwg6tlniqcl+zVViMLheMFpj7XAg01hn6Jn1HU27
yfpRm0uIAL+5xkvgnTBqsPsBxOGBzwWbP8uxPO5hdhihn7l5r1/kg6UFwRMHWeXab3gEwuSrvdUy
90eTrEUiC3XMsEjodfR9iCL7s5yGXg/JNz6nIDw5UB1/309yCvmLRijKcxTOUSE5r38XQRYHOTRs
yk2cIZmtaeQEHQ0xlUQSODmuPNRwZ7aPrntFJA/jzd5zXSxheITooT0jPQNDJxPgDhpB0DIEQB8D
LwaaJIGNDg6qxixjkSzGWnCNGLi8gVZZsAq3/Re+wOhyGUFfeqjtKUSXmIyGtlOFQK+m0NJn5WBp
1gR/dT5GT4Ut2FJBMhV5fJYRwBQn2OtH19y1ubnRlmIg8wpIssIhjJRzfFS9AMo/HxHNpJRt3cJp
l3RtDMR2iuPYwiqmI3KF70bPiOK/b//0PQbvrhw58z7LEWQph1KmTfhT5qv88nIFKu5qYLQL6VUa
axIUn+NOALrcYeswBmR4SrXRcFpvZn3z2B3qhd8nqnkTY+EJYp/zijoyDip8cko81RkYYSft/XCe
9aPUnrrnCcE9F5dwMM7xvelpmr+sGj3r4EbRvNN+qdl+KwAhz90E73nToNosArU3WxRjzeQHbIGg
T9zY6SFWR5grFP/TJ/EH1N/drK2edO1tt7ouwpFrAHJ3ynUmrOq2HuQNlycF4VcmU7yukXsiI6pg
aW+sVIH2zDJIEdgCY0f56c4yA7zKUQL4O9BWzpS3HxjLO4B06WTZffShRyQ45nAOUK7vXDJNxJPF
qYjwCmOwfBKvoX/rtHAi/TbWs+gOLQaLeJr6nDWOMqixVl7c+WMMh3/nfXSKrBB9YR9Ap+/eXLjo
tO2dSAXUN0I2oBYflAxX3Vx0kV8ilgMRjgyQfwjuJsXjGlSsna3geK9KDEnz3QvFTUOWyvVA+XBT
7k/Doj6efXvOWZW3G3Hoim0Guc7fXh84m+QQiKBPTtWT4j9EJmAOnanqOCM9e5SMForR71wmYOCZ
s69HoRK5pvr40DmD4M1LInyUjHAfxgdA4Y/LDvFaZ3uI+p1SJuEhaQHd2A9eSnJ7mJmWPVtx8d5v
TOzIYmUwJPfx/emKoTDyYgVxbmkIxI9B0IC9e0DMjz041QUE0P/HVeiN1QdmFrUkG4B6KfRmjUju
xUQ1kL+y4/EAnN/CCcM5wdVqFYAgBgokujobMDjDfNXe2g/N1u5GztCni3mkgKeCEdtJkNC0BEe+
4GcArFeLmOX/XgdGOKc14LiP0xnhJPb2eM7ZpgTbEzFFOKQlBgURysG42qiUhGPxsiRB4thSfPC9
40ofGy0FJqSOqc+/O7ImJLk72LAbY6Utm4aONN9+R3vL+zP2nyO2OM9Nzdgl4zVqIYx9AXPEW231
bC66c8pxZPFfeEqdafOItBb+oDD0RgzUkURQ0QDhgz8nFSFitdIw6GZrAKPk5X8n5+hiADrw0TaA
2aGvGsqw0cVicy8l8jGcPPtAt+a3p5HEgLcOOFzhfGNXGZyq3OeMrDqpZ5KLzd588Wssx216E9+9
KbmNwwU8GWEEJgEVnR/AUCcabZwck+fVdFusXo6uETCDO+rOGC2DJoJAS6jIPYtRgMtymVZo89zZ
EQPqvlkgCt+orjj3YMY2cvP6X/HAkUrr2bafqWhl+hMRFI901jSV8zJsooCE1cfNnZLBmGkXyjXP
3M26sF0x0e/LgLe0pWAVwliNDKH7VYdsgwmnTQEc1bC4Gq+6Z80mIZIek4zfaZ0lgBqxvUCk+m5z
QJsvLlOcTFtQI6uEduqbVlFJcvUdcgfm3OqESeB1HIYPEqx1CRhuLVgC52W2Kw6yzSwi6lePNkbT
w/QTOdyrYnzAd58X+oRK7isuoWqrKYOMaaYGmHR0r6ah6AzRm/zRjeDK/JNYcq89ckTfwH+ouX+0
jccgXZLxfCgkBfu9eTmkKqmu+kkZOAL1fr8j5R/Jzt94UV6hbsOGIJT0z3llImoD6MMJV7r9i7+u
Fj98R++GCOFJGnNPb1n7l+WmtUGNiQLiKud+nhl6R2fLBe1pke/CQM/KGMr558+IBdOCVa4cEudU
DVVrqS45eXdGZp8fBGmJqgs0yx90o2mK4yDFhc3S98WfGQVeg2nKc9+1Db/U2gM2aqP5cZNfXtv2
8hofw3dlMS8AY4SompdS307DnK57IPnphcmXwPvmG+6aDdyYrdyBDg1ZjUIpCMhnxyTDDCGY4e6i
Ay/L+nlkLTPWG5cGjtn2yJLkEsczbFbPTGmpgQHSpfDOYwo3LYDlFC2pco+fXnIf0lO+NZbP8ZLX
FRBqmrux69qlcujmDqz2hC6grbK2qYtX+p/ttWXAysCfK34Q9D4MbbxuS/MoPnMnKDIyIuvsAYoO
TLSrA/HLWjTjTs6DGJIvrwU3tfkCBewxkbZwBzC2v3gDle60tWEMRsokWuwRlxGa9a0XptkPpziC
aCgsWFnRFHvdPILsQmq3tyhhle87e2IfrpeStFcxUSGneBW+864bMyWN04blQ1BRv358X2/ZQy+W
mfUgmBz2SsywGYWwXvtlGXDRP6x8KGzyqcTEmUiPbA6tEEJEPy2dognTatkvGqArsmT+sSLnTBxp
T0XbEGOHlauRP/srXvg9jeCGVLdcbW05+uQXLrbDkymowFdnR1wrbXHw1IdEd2DsGSqCGLfp1+ZS
jXY+Q5VmJjhmL9uR1K9uIfQePTSRHxrf2DD1Z94ArnhmXlM+UVrenS3ZfCMzwtP6+xEswgc23OL4
FMLL5NkoachKE5J95Kb2lu1isbeCA9Xye0VysS1Tc1sr4swENbEsp9XQdl+RGdcDc28dNBaijRp1
EEAUVcTH2uiNR5Se5pZSTdWalSUpD6reX6JqZZ22JEaBL9m9N01KkrI0O1LhpFim/ZUS6Hc9Kw+7
6yZLHtT04FdR+mP5x9rVJwHqtSG4lAyQO0OY8jYxSrQchfd0jILjhtsdf3dnBYPH8a7lo3GWratO
qzxtvhXTIbLctl8ohrVuxdzqiHriCt7OTQaKhgIP2JZqQcb4fGMGNNA/dAqfquPkOB69klAhFqFF
b8zq7WFFK5DS+pp591JDPMCQ/DXpeSqLyc41Pb0YEVbGqJSCcjhinI6nZFlDJjr34vpU9e/VSg4o
yploPIDc/NBE73bThoxnZb6rDS8m7NoGgc7HpmhRur7ncJzt3E12kUx8CrnuK6xD7GRMumZkKQRA
/MZV7/lLgRTizX3ieUG6y73XafsKby59ok+mKlMOxjWcKbui/CxEaF10RjwcjLA3ZdoORiNvK+Um
Wk2UHku35tP3h89hUTGgqrUjes180g8MNOEhwcz4Ztg+E/lmXZEIZyF3yCpw5nqH2u4Vr1+pVCtO
V3o66yJ/fX88N4QEt8LrqRQm1gGRpZPWkmUD6d4/OOUdH5DzHxc5celJSPZZx0Z8GvkiR+4RNR+d
pyCLGfj5acKFzVNbXBMuaCamr0ypKJxa6YL+qh1YZoSx59Um557dlotHjQ8+Zj0cMDDBuk36D5Kg
5l5EOXhNXPJzkM9b7/+UNdPB2V0spngpNlOnx3fMpWtWBTqiLs27mo/UAxnsfEHHGReYrPh+OyWk
7//r/9mnExJFNwsLekicIC9JS48aNWHbO74RWjWoWi9ks4+VMcMyAMGYs2cT4K932H1naMMkchcd
bAPyOfSLzTRiY3Qap0dAQHsZwe7aimRSG0v+o+HqccfC0WROVU0YwWnopCz2aZf6JOmhBPqYpwzx
EvlYXkHCg0apqsPJoLhRrKAX+xsVBtslYIVeMFVKhVv+iNhhEdmDjKdTpG3HtTjdpNGOvsI6DBsU
qbZSxE7IQrJvudi/G4lT1PwYhG87quyTull33/N87OsOyXD4TxkJ9Yn9BZlPCIa5suZ3EKeuo2uJ
fH2bs2Tu+QGiSb734mSAsC2Xou26BE0fI49hv9R0ruCiuf9/RQifAggjre0mYrQfEuIrytmqZ5qT
eUoOssreFw+aTNWmh1it6ExIlGn6n7SDNBb9zoEY3ojc/h4fU2M4lNyhGV2o7IP3YAzSZ1FbPOpW
o7fcyD4TY0YmtdIWNET2MAxs+dS4h1RJDHS6rR7I9BxrnAn8cy2+Wk64/4e1Tms9brWoenv7enkj
VHjecn6bWy5EfttZ3GE9KcpgW0Yur3sJxy6QHSs57aRE2cLa/N2m8YgsXyNCHJk9O3tV3aZDsMqr
qUO/Ktqm/qeZi4jnCdFJyKK9sHtz9oZQpjuqv02nfWrH/iZ1VEB0XBt24naLDP8cLQUo5Ruydase
g0kJX6HRUhd/vRQPkD1lOuSLc/HlCTV14qGG0fb/8Fc5APowWs3bROCtwg9cVEj6dqOWkuvx+S1Z
cl8BvW5g3FTI3HdJZbSIKMszDjLlXVcxSCuLImOA1mynw+3ZF3H0wJCOrpuUWPAaGEB1NfCo1ViU
o1oTrOHcP1M7dDl/4gdyLIYfjdgRzF0LSRKXc6RC18n0Oja1jg5NwsEQQ/oBDwDG9suQyPZXsSim
NZtY0GRFhQq5Rvcom6v3NFhqX5xRSptWQs3u/J+S4+pNDn6pxvhr698FLz4/JYEawf7OCZjp6/oI
ekh9jRCHP5fWX0V9NQXpdv3GoYW+vWNHQu0mJqAEzS8FHg1Z9gmI3HymBr1z99T07y3LkX+4kVQI
NitdyDZO0EB2gm+99TMSEc/cA/6GxCwJiPjtwIoytoHLD0LrJOC/mfRHd0pr0GOK4t3S94qDJcja
dsHbS4VYHTcVIk76u6X6RXyt2sGt+Sp9KdW2HzY4hRgFmVhyEroLjgnAI1KF/pQzRh1ZcNowkcnp
kWgnpQOY6EuAZLmMoEPoDnDwDUKwWaJVvNKnXdg5X95fEiWCSny9LbP+S5JETtYvILIM3/SOQ7ai
ujePN+SNgUK61cy/yLHp87JgfEVNwuY8aXah/InxrsD3cQmGIjvFGikI+0Eq+A4FnUyGCNe7yRX2
nt7zTmJBw/BMS+RGSZTL1PgaojGj3kqYrbzcMzzOhszE/5h/OOIkBg0IiQHKT1nJXClTs6p7EB7y
uJdWFVseiGR9ipADqiZ9u0riPBaRELdYpGrTqlnoa0Z9IxIPCZAseDhCUSbgNHwouM6+ymicUiOM
58+XMm35O7Qpq72k04XS1vj6loJo5b2XUsbqZ2DhG53YmhtV83flUe2avjbqWWDkKMiJ2lYlhAXk
Jix+b6bJ6RB3md/7xuGLYx9XIeL6CcoHg154ccVxIM56/WAo8H8yDznIVCDQrG8RnHEtGPusPVel
5rxEub3U5N5gAplnfjyHwFbznmG6axxciSbx1g+WAI5A4/1eieAKdQTt57Ansv6Z/3ZiWXQhLjOE
BlI5jXERmg2CgJnqhGPbR3zdz3j5RcbNrD7AkCve6SDH9dgeh/5h4ml8H+fp01AfSRfeckCnmZIY
Su6WAhii2lQ5JocUIBCBGsEkh2QtNRIL9RQaFCjJEIA8cDR+I59XXi2epgLIy9htQTsyb+oLjLpI
UtOLX8mlnBZ9lObQrwxGrGeqq9h/h/YnyiKB6bNdzbooIkOTsmdpKmB+7bR8pPxrl54FJ7S7DWwN
ARDTJReKob06vSQTQ8tWUC+GcSdSLaESEs4BKuLvVrvikKncjmxUtu+vXlvWm8Ig0Jgqatl4Engg
R7wCgqlDxqX4zVuOW5VKbOVS5qFce5AF17zxETZHk19aMUCaCAbi9kIaTTpd+CsgBiZPXpOxpK+U
SfaAaSt/IIQk2Fjcpj78bFGQA5V2d5eEGEdiv7XIjqwEIFk/a63kQmjF91CBIlFyCpO/dl1RJp4A
fGJE71fCMKT22JMaggcr1MkBto2haHfIzhMW8wRon5mM3bYZgGJVeDqZgGAtewPh4+i7wGAVnyXb
VTvkVVB3um1C+Q7DSTjSkvrUzy5rK8dIvCo/8uyWegR5BFqGcHtilfVi3ObChqKu8SIZCClVZ6Mr
k3rv+RdeeDqke8ZkDVAODcAIls3wtg/jGyJmHzF4PgWyG0DSH+g65UMGcwemxSWtO1ChK73Pa+8r
Oa2qQDc1OqwwuVydC2WFDRke0f0YmX22aS9U7KETP0EGF13xnxbv5ZZ/PqiwCItMDMrdajklUybn
bf96ZUj3kQRhnX9PWcxpUuzQOB3ca2eIA2++lvkLbk23Jg1M1KIn3AE7Mbsy7YMFALI08lXTzEeT
+FeGDAGoRrc0VMfGBfmK0YuT+YRHYZbcZsuHL+CQvlN7zD+oqugYN/6POoRAM8KRVZuZ9auESmUw
ed6mjimbXJR56zPs+ePnM1tcx0kLrJ12wwpfchkBI5MFkPqXny+jp01Zk2bbXaJICSnxPqW6YyHK
rZQuE7K+M08pWhQbwARoni/a0L3aDdeFdlY1qHFkg/AbLRuUqdxWbS+rt7LETW52Qc6mH+U0oRjk
a12CqCgtziFd+dnYPVlMXlJZp4P6XPzckg6soTJQ5i41Y4itrMOsA/l3iHlJAfonXy6ttiYfDZV/
xv9HBLij5JHkGq95l5tJu26nB6raoYMeHVxlfKBI+9BhS60rVDHWlOB9xs5ZC+6Ii/gCzvmo+Wlu
ZNbbxXmHfg914gEYMvSuDof52CCHGlAmVuhB5rzTog/WEkr4o8ZMAbw8ZVXiC7PG0bnBfrIaSp1L
XTpNxCro7ZjxAR5ZKVDcX/JIwS52OZM98yiqAtbDV1bFYHdjjPxcysWs1bdEU5mHQkHFZzE7e/h+
RLlO92KUHoH7/U7t/ZMV21YCLXUs6h0N0Oc93Zl6qWMqwRJG/5sWY4ApYGE/IigrDTcC0QKEAc4U
RV/rO0tvopCgceLBPwwxOh+Krqt1UluHDDfp1tZGMqwtWLb9RIw2w/PYu/4TIlJbjWJrjAUR3n6t
D7VSZeGkYU6BYQnb3gl0dLDuNE1ASZuLxa6ybo6UHlT45T/dIKtI9HquTHr+tEWjHzgIff439QS+
tGXMAePsakPYhfaW+FzWnPptS7EEUf0c8QxNxYNAyjd34pcHpaBEJgfYFnxBmZxZon6nIoSH1NkJ
/Zrs1LffuMQRfoE5da2BvhE2hoTW+iwhHcPI6Jw5bWtVEnvP3iSoZSYD00dKzHBiTmu+K5EImZgR
es5EaRYJyk94e+ijczyrHKckcOWdsY7otSsHg7B7ooezI/gVYQUC3WtvOplhBLQ6a0b/cw9dt49K
AuKgI0z9CM9fqibcTy2d4Ch8YV79CLGzWaSaKe1aS9NUEdw3dD3aiVBlBNIztP/1dbqr2QVdGM73
V8hMCHjfZfNjOh6ftCbZONCC89JaegBDZQrK1Fi3lelO/8L5qLX/tHDkd9yBUej07Vn5YwjLPToI
cRBbgp6PZH7rON/Cf4HDqIgGHqjQzJ6o0oGOicuWYzuvJsuLcM79vU5DE/2ENFAkjh+3pn1HJC5B
SWcP3/7S/NocXK/T0F0dTWGFpz28VzB12xVzM7kYrvk4zmkFoh+l+KP6rRBzJCBIvhu1xxHoFRrN
1Jjxcp6CMl3v8FGPVqXCPraFOOYmID/juyvZvFOkXEP/BqZVCb/s/xa2APmdAZVaUS0pS51mryq7
1XMiqSGHtXLQkAzYkh15mpUiJef6skeOBtrwBTvHJfMY90CGH89rSrkKve92VOgOaN3H+JikddR4
Mp+gGq8F3VXQJGBkx4mv1iIr4ouAXJCadHa+zEKsjdt2GoBAZk5AYzIglW7wC9g83fyQKWPmwJtF
yfE6/l0a5BMYwQ8YIR7NKL21VxrvN5QKCOdvac64ynkkD9ARz/qqFGeD165TpfAX9uNLCMbMI5RV
4k5rCZbqHIIN5bp481ljOp1JHjSHf4zXs/GHO7MgRTPiQ6zSy1jqlpHoD0PIsXxGYDDdm50JsC8Y
VvdH1M/7vNhpIjhkvAm1kUdlQoQ6Hju6kRGhaWRKZB5p8FOL2gCoax2tCuixTNNEhc+/rTD5qLrE
IxeeYjhMHhYOhhupo87q/gDszvBtaZaxeRA0BTN1XvHjKUoddX//saHMPcILAhdTvRoht22CBb4N
7SZDbxu1R+ug1XWOkonW1SoONpwUdJn5UWaUzMgSEpmTLi+E4Go7jkQfw30b2jxBw2ct/tIh/a3H
Z6dnUK6KMQ32aethQC4fUyX3hp0Y4vbRvgkJ3Nq8zuFarI3Sex6qwLkJgR9Qzonbo7H7KJdf/8Ad
enUOXvvLV4eVKHYOoh2c3NL5K8bGTFb3d6KBK8nqvAQCPBNt7icVQd60JcP0MGZpAyJ9ZQU/Ypy2
5rqKA6+LXykCSx3LHSyLvZJu3UWKLVAOLhAl1BUFz7GoOdha8p1/2yXsLSvjXIn5cXgyZzebkL4b
YldYrz+J2s+hpuQ8faPQwZYWZ4wtdn7nKSLUJG+a0Ms4P+sfzXV9V9nAlv24tlHE3UydjMD6wZDF
W/dvRVwgGVcolKtBNrM404xUSJSwPOHE4ZWaOdXBixCpIZ1eJ1QaOpZTM04vJbUXzYUCs3vIHc8f
gG0ytjvTwRCMoCu3IOnUsgdRpVGFa2gpdGMR/Tz0xAu+HLj20HXc9+VHPAd9YwJCmC/Q+ea3cs8b
OwdXG8L8lKc7riG3ujWLE9LRv2HUZ71Lnp2AjFeKlM1GN03+BeSMutkaseEhOx7zwhaf3+exMb2G
DwDF99l209lY0WMJf9/9QUhre6FAcF/a3445KTfotI0sz34Kg6JVlm01UQxHPz6wh8RYwF0f3/tJ
gPfY9zUzN++TDEfRLUEdXybME4gvesB+rjICC7dLaFPSjMlktDmpdTn/u/8dpET7VyCU8tp5bjqZ
1sAp3apcFmGFKd7D6Pc9jS8JSsquDbnhQLmwdgM/+Ucq8ETsWac9EVZGH0kCZrEiXAALtNcLi01v
O1WQfyBRIlugVLbikoPsyWvoemRm76vBuWjG3CFrIyKaprYmlsMSTRWF3Bt+jvlhBUnUOwuB2elb
kbMm9oRj1N3JRjm9zChNiwCbz5gzFhbV5BzS9Vcs4SMaQtF52wYDqa8UScPVCFBhnEo64DHM07aZ
vbQ2vQC6y5GMAVuRp+xl4yJdx7mAQSXg6CSSl/fV87iV7mxtCtnqopLbqRY5AxumOPe5e6zaU+Tn
WqkyprnWlH8VBpLSKdSV5meB7YT+x3Jaxp/jvmK3RyM0wk5fHNLeAqiN5GyGxvjRYmAKc6L8Q2V1
HT1VvIE1p0NfaNxXYUosrA8uLwBEWUPq0Di6ZFOAKAekK4uTCSZm3/KWxMATKRaTKP50UMsrhLhZ
Gttvb4+z7EJDG3RgvIfUSJHHdtwJkdBg7KEhhb9xe4QrO0+opLRAFz3m4qNk5/2UOs0lmEIi0Gud
T7JrZNhAIIcMcb+OAMSr7tj2fiAyPf9gnx6yx7Gmvmei3ZAgzR0J8dlg2qOet0kBv8jvY+O88tsR
l0k8m+eyjA5x7FElx7No2o7n9qczUm1pvvVImQuvQxMaozelL8lGXe5xDzNlv/z7IRGO/0MfRuzf
1DMj9HLY+QcC+YVjurmcJmEYBTGlwzNy0ChAkrEPAcQK2jaTDg0hMcZT0dlygVSZvoiYQb5ESV+v
rIVKmU5dRO2ZReHLww4+sfCJMAiUFzG8AuBBm2nE/lnK8wPAcy9gJ0oFbBWWSAHg5zndWjPdzoew
pWe9d9+lK+84wEoJaLArp5nBy0GG7JG7ohXzOgI/fuyci45KHkk/UwlLNgZvShFGqpNYTnPOmayK
ZVg47mGIM9FDBAuRjPLd2VI/rCoDRxnwqjQmyj2PmB7TU9ZYlE6LAJlI+vULJj0JbakYKZy3nOmL
qMqHT8dQIQAk5gKtuWOS4t5R4w1C9ThCNaRGU6qvV7o32DfxlVHtT0dwcxkiuo32g2Ya9QTvzZS/
GxRT1MLz2Dpr2BQ/pXlHYjrH5K53X/DhQNKzouOzZXJry4X55Pl2PPUsAAC9UOXn/NLP54txYVRd
JueZ9MzA9EuYgJUM11+iuaSjJhpK4D0kH624ePvI8yTb0IF+lGh1Dqv6/hL8PjGpDY+GOz9QzQ66
nHIeXAWUNDPftKVPzvKHGgwiOIfkNiRi9E+jEOppVW/YvlqyZ4NbCPzPtNjYJkvuaPlQ/KxcBKYH
s1favsus3m/xP6Z8MUhjARG+qYVAkrNaX7p5hmwz7yoKHPdBVWbfldziHjQa6kuQkyveN2SwZ8Ui
57JZBEkp5R1RyCAmeSA1d8zBlXhDBVNt9xUlXl3Wku9anRvck+rJILYPUP+GXXI9ckABMylEsa4O
WZPD1Uk7Z8Vo1XY0LA59sBZ8pdWXRLBBgUh1EdiKEWS2tvK0gOBQvhLtcvO9GDQbTFp45ea8RrgI
r9fd2ePyK5eTKnW2l2Sh8zvbN7zZ6o7qKGfJOQUieZPzI01A1Jy+PdlTYuaZoM5ERVCSEsQzrd4z
sp4oEohE+aHJGUNi0JBNw0MPYqABItLLFZx/95+FBD4gY6BPJJbL53y9wh3oRpnPI3f2p71/eLTy
Zh4LxyibGWIp3hNC00PfLNozBh0ftB3xgeoDMzxwy0DlG4Q1FfKwBBYvl4omxdxTMNjjAAuPHK63
imE2iWVXCv2sIZ5XmJBIyYGLdA4HNqEUZSvsuDGs8HFXSa5rQ1f43t82a6U2WXmfiIEfGJ7W0DHs
vqJc/+unNlbKd0I7kcZruJgKGpZsGoyTvRvx8BU18UrFFJQ+NdJNfP9GrSa50CplClUZ+jQEGw9q
c8ytn2Z0ikoBrXfuSk/b3J5es9WG2hnivnJS0q7eTicRGOYHV6MTfgsnpMPRB19yG0rvxvQY8nzv
blR+kLEFszn10PMpQnnSeSQAkfI2XWNiA2akfrVcmyaetzPegMen4hsTmFoDQgjPGcvC984IFT+u
5/kD/oo+kuOaEPlVEQkHPLor311VbH55pKGKXWzPbRJmW1un/jXph6l0MZiPdx+1Ck7joyNJqqAR
3nJbIMrONWSZbeZJmYVkxF0JuFP8e2I60qEN+AtRIawiTrRY6JCcwIGOLXMNbPZSWBSzScwYKuiH
jOF75DODiQlMMazoUi3LkaHPtQVBJIwyRQS2kSXdHYcNlRUX/YrFst+AtU+/KZ/rm51q9Rus5Giz
2x67xU/R6ybehgFxMS4gllkBYBBxS4JVbLqP8BOKCfqxUEe+j89nDHYNgvUXLZSDA6Ji8o24hYjo
zwB9QxnAL6DlaBSLwllzuLg9WfpoUs0T12I1W7t5Iop63jIAWLPN5izepJO5dwq+4gyPuX6MVKsL
baOZpl0VPuz8gvg2YVLSXBnNmlD4Lx2sy2xP5Kde3lpmtvcmNcivFsKRhfIBx7xG5TCai9Ny0fNm
khWIGw7A+2APZMWFLq4q7n7XuTMxCX7veCKsrYon6HABQZvqU8mT8MD0jMN1/0uiaZHESuAyOKLA
F/y4DbUwj1GyVRagOJ7xb+kBtLEqjARsLmKaOuM+Gc9ooQBO7WUhTR72g8VQZosTgZWHtL1VP888
GzGHwdn1t2u9OuZf2ANWlowD5Lplh3HnENkKqIe0dDt4w3j2873sneW7fwsjrJs6q9ZeoIXamqQt
N/qwBbwl65QOthw4V4ZOcI6nSeDYWbSCE6cGbnJuqY+CiXHNbbtb8bxVWFB2uQjn8O1THencrSFA
wXshKvG5eHP9PMMTP9KS8N7IA5D4wazjvwLXQYh/wJtnQAQDqt/fjtGyS+dPim26+xAQBVwkMudG
eNc3IPygrSy7zN5SkpwomZl6fhi62P/6aQ71JmgZGPKOT4ntXF9vfWmbPiOSYRWgjsCeR2CdQJR+
FTykJVMEggKts06gIbPB2+4Qe81uQJ7vmfMzCfzStvJggXBE6oFyDI9Zp16SCpf2FVZgKeem6ZLC
Dod9FdnyrmaMa4nbZC1NaJzR8i1SSvoYXOE5DXfHM913ACekKeIMr1FQxZCMxGQnFEzKugAraKud
6RrZqAW2ixF6qdWZKIq5LeEyvXfMMh9PEdE9smSFmnSFZgbuTXjgg/jJvWYk/zsuVUpJNzVrveeP
3pNIJhkdu+yh04Kra3nZSLL+1umSFpvKwqOeGdO20u7fnpnIuP4h09WsaFIFyfw1+ASlhZmafloK
aTc0rOh5Ur/zsoZvmvyhZQBvbWJN7Yl9PERvYMcSkWLlgletJAXWjthf/OKE/ZSp6YEOxQVEFWsQ
Y8JonH8MDF1A3j2N1IafRPQOZnV7KqJCkahbvdYPVimMq0eQvUiTKOwpPC8pQMinIbuIMNYn3Yw6
CMlgOyL9bLZdx59EUpgheiqaMriJjjwt0QSk0fdDQNtSlA+pn3inwb0LPrgAB3mMO59WFnqmH9J1
8U9Up8hNbLzQtzUpyPSusVkNUQ8iGGxZEKsAQNicApfhbOSRL4TZrDXvNzPV1dU9DBA5K1mvMS7f
8TNQKLX8nUUt+UD/y/L2o9zqhUjJTFltf8hjuv/d9S2Z69zYYYwrlFTaM6JLs4dREcmf7fVrZJOz
njV8lZoT5X4knDDkDqaI6KO2ZXBHfOwoPsWkxG7Zdnm4y98zW4OP41IVwaFLYIuBixgupta6lpVi
RWlcmyc3xBHg7H9lAU9lyhIG8LxVAaxzm4HkT7IuLpm0CiTqseCFceeMQApeKT/T4Zslmdmwa/eb
TFFvOU3LkiwKderJ/kAfq/8TXO1DZzRbgqCX6aztz16dY+SWWcwSSiFI1ksVkOG/a3bVqTVVJJyL
Qg24kY7JCGboi6avQeHr3O4hO9OVEtnchrLcFPr9iIzu7pxMLSHOAeMI/jcfJRhCdePPzGwm5PFX
jC4EqEaoLaYrJRi9y8bvkn2SxzrY7xwcya6s6dMId/7icJbSWcD+fbf6kvhF64abI6uBejGHm1sF
dHxGHU6RAtwnxSgT9VW77HzALKKpb3Aqh4RrZjY92GW/rf4uEx7DnKUOAm3TSW4+otBqafkeVFsx
sBJtlrfB6HsCJpGg+HUPPjtQc1Cf8/ONncEziT77axFqvBDtbMoGfvFv5pOpuuxpNbtIdE4JeFtf
QJtMIr719p1b70wAohwCbY58YHBhX3nXrqZSaNUPliY3eQxDs24PM3HoSE94m2WI9Y1j38O+ld5M
tT2EsBj4fF/jafKapaenTbuxYwOvKOPbD6+pjn3rRgFkP+YXCfsWqTyhoBfGa3LsPyJdpMiUfhVQ
PgF8LdA+sM26MM9vvVKSzBGROIVEvzbexxMeq24ZVKvlcQQHjLtoBRNcXdWLtwNR6l8n4e9u7PQq
RqveA0j5nFj4EuWmU+XMoao3tLs2WQ68KtMlM4GjVz4EZciDBcIOo16Pj501vj8B1yQuNGLg+JaX
1t6Rbrbn8VdtC9l4PdMleYaIcWJ/LTeR/oO2SNFsI3qxU5QTycVf5TBSlXuziKDz0WF3yE1MXaME
bsn+qdLFk5XqHAwbsmv5AgSuqaCWMU2kD4BOGOj0tXNCO3Is8c8S/B1wbeS6dNSPrbBvWHlpksL2
+Z3AOKKHwtGdU06lSuottpEPdilkSGcNJv3xVGWJzvgjwNRO1MRCPFvGzIJVa1/3qlrrB53zlmnv
Ob/BlCU4OOVEiq2jfLCdSZS+bLjq+/BRxHNTdMOY9AzE7fCRXV4+7/NtsSDf9Fsxzv3h4QGua5e9
/KsB+9yWbDv9Wi1jiaba4b+jRW2thFwVj0p8nmEuCehmCQzwRqnnstJMlruwOimwjKjLeJGGZePZ
c3CSs2ZKK93bOrVQ0LyQiOEuDfgeTj9c7ipikZTfqzoBEzUUV/8YUnGoQYmQsEJpRfvVaen2JgY3
Fn9LTwc0RtH+s61kd2+0IUhgXCYxHZJ17jPSRVkxN6NUcBkaB8H2CmH0/9QM00rc6MPVQ5LE3PUj
5uxdWvuF8uOjN+oDJ1awScouqfSQYJG1C6Kl1Yz1hsrAvBL/J0qDOOUlUGDF9rMkJ1VRITsBD0+h
n2wccD0Vw5D7L1PvzUjXz0osBCuuDPRQnaHGkZJ1q+IaZuPOLpg0sa2/GCqcqXK6Pbxjl9NxLb1x
zD4D7xyAUHxwSya35nobxd62felFMeUvRfvN/4474M9wUrPM4wuxDT8VHBzwzyEEi4kK8FZsvcE1
Ss4r6659iieXjy+x1VVBiPhU1l3FbOAGgls9cB0dXLpnr6acGqI8JsNqAKYI2qBbC/FAdq0YMeXp
hnsPqYHKx49EQn62V369WyCDSgxrX7QyLbhsbTYg8j0wzudZ0qLxp8lOivZxto2Pd/DUQiJrL1S3
d4vB8XZkD2XDtqZIsx0JyXqR55RWEWpcGpYEqmPIJ+vM4eKgPKxSWh8a5Vui0Vaqv9OsDTA2SbAm
ya1iDROUfKwvBuyr35I0JoJloaMaa5rA3/hvw9yChfiP8xXYtjMLP6gTr3wE72QQ8yEnn1Ub5QHY
rW29oZb62r3AmmbG/YBMPdFTsl4VJxHzitkoCHwcsdp2Lduyfb7jl59cqSSzaIjFeedgoX4YVkzo
i6sEPEeu1DGTFw2FaCePxixYnHPDvSsoPE675Zj6G/pDj0F/HbeN2h9JknKBo6Blb0uOCkOgX+vf
TC5jVvYLrx4Q4V4TT2Exj9QrI6cJ/D7+C2A/aN/mxZVDYJno9diqhLLnf5FpOrhcAiUuNrCmM68R
1DVH3Q+FA7bHzGlI8HpwnKOJp31zHbGMeD0vsp5n3FXlxtCOzZ7AIMRpjiKhsBW+N4NJoXFIFPmO
wKwi0DjMp64hb4TfHhTRkY+QA7O9En3c6EDAy70F/EO3sKmnjHgTTAOdtvjpC3QfdOGZrTa8evcd
G5oCcNZbmxeaZshY+vetHfkZvuyxBzrpQbXTdsxrni8BIl8ysHLdv2848iEOCSZ8oR+pIxuzrQO7
36BlKVJ96qIE6BfmdO3VGNwSBQKxzhlDsLbzsXx01ZuSGZ3ekQoyoyt7O1WGPIF7V+sEk2u+42lg
uoiv25Vq07uh9kefX4E1vqtdVUmpteXQF7dWWCgXb2dYNQQr99b3cmmhzc/HlScG7G1SXd9HQGHy
5morE4/GF9ZfH7QUnURJrG5ErGlGKarYYPbCdgdiB8rQWheuevrJmzbl2ZpjqQU4KDEuCMCfHOCO
VcBb7+TrnUzNNTEv0ZA6SY+NKR3Wk3FNPNtLQ3K9+83jNA/ugSbS4WuHSK35mAOQmxoYG2o06H+n
ozQ4jDkbvZoTE/9soulm8oPosR+FTnVXfBUl4f5dc+jQoXfX4z01FIR9QaUXEeEwbkyQ9q35qtIv
p4eqoFB99pZp4EkUfRChqSUU58ksobCW4HWMUlbQEVtvGPlxoTFUPjCQO31oGHDoPSu8J+/YSvLI
SNTIH6UjHmHQz4R4AbgGy+MGCG3KJJ05NwICw5cNCnmn0VgsKKTujLvb0Cdr2be446KCRO7i6z6b
53RwIrBSsp90V0JVkiYwwVUsc3WY603JN4uBtjMgFa4QDN8cWBwsoDj6IxmzjtrsdUsFWcCPJnol
vhB4Aoh/QqW+cNGTh7GSFC+n+kx71ZKFZN2DleLJzmDmYDM4xf8Zop5vjOLtQZzYt2RIi2EwZ7d9
2ugTBOvr/jHyGaoPj2yYccGxbMGC0qgdOt9RjDl54RDPC8Fi863SCRFkri43K5cGG/9TI4vsFWhE
ULA5TPttjM6oSUGYn54SV4HdPrTr+VYVV0zeveztpY67JXrPAAjT0oVNUe7P1WH/Ya+FTF8/1bG/
bgH/e6A+O53MHmB8ODrzQ50q+QOakHd7CUTRgbTG9EohrxEJij/iuBoF9LqD9+ficCpX6Ei0nyxc
UgIJ1AH5meANKbdFY0KEvowbKeGJ9kNUj4jmZv8ocJmpLzWe7ToA/4qHPzui3dppOYHnGIOTHjMe
QMLZBYTYzKLfNCCX/pOiqGtKXBMty/3XtB3in7bHrW7x0UGG5XPf8Za/Q6sjwthrt3t8y7oHYqKg
GhsrNhnhEGCY+QJxybE/gd7F6W583hntIkApPhu4ocGELsJAcYenE+D/9I6QVV1ugOeFcITE/2S0
YT8kzKOTbEAiMcn+gr53N/mlODxHpMQTvK63cJcCR/g0WbIEyQyLLF50KeCBduO94vRzWVEIVeKd
pVj+ZcUNG9T5DmBm3K4mw/EHqibA6pRGUeJuBk0WsWHuhO6+/6chb2dkEAM793WYPotmG1xqN8Rh
rjAqdtEoV2zX8Slm/kaqIQxq3nqMrWJrASTG1PO5+NHNBoMPcDuFIhyBcLOGR3Ud7szvirMZhwU0
x3Gvl8h4hakEGb+jNLJPZTedmMa9Fc7IiVZBB3/maefir2XplkViko7Jp0ZLiHIzzsHU847wPUIu
AJRSK5Ou+2JhkOnw/oktolxTXh8Bx5Fsr8NvFdrzF8SWvJi/SIO/0iWPLTbr/1HusCjYt3EeY0IQ
M4PG4BnOYtliM3CDE/H1g5D4cjwEKKwmw5lWKnRTVzeFuUeJNcBm3XvZjD03Q585dFF6JTWAffpp
XqyqcdKF8tcizj2aiB5497jMYJddv/u5lmMV80461KCdbuNRCcOMtGZdLkmjFjAhmIv9bwxrJNWL
snGNyCf7AqQFMnmWniGy8vvLgyUjsRglUWESDyyfXvjBjVIKJ92H7FFo7J4d33qXlxQ0+nlRqhOk
39zZtByTypLTkZfdfEz13eCVq2g9kB+sowxzd9LLuPZoa03nht6ODaOHBck9CcZ8miKsjb8DWBtc
ePw1iGgUMOymmi2tox7et1clnANVBrT4bCDgb0F+eF/V241JFqV4O7E0VRdWadXDFl0aiE/DdLhD
OZje6xpsrApo93VTc6AfxjKoY2kayNlyhucPefKZsqm7lAbhj1NEh3UEh/RJSmAw3CGST8l8uQhE
aRW3g336IQmdAwlJphtuY+KpPziQf5dO75UYHlP4VFNo+pX9azGP8/Xxkx/fpGn3TXlsSz1nMIWk
Kl9Kpdjr3ZGOpn5xa6JOvfy0cj1zXNJjIUz8miQ+M1Vx1qmJAL6wqPh5Rfsj08PU9yqsUAVnfN9e
wKI84np55ZzMQu1Y6TKHetcTFUknjvV1/Pet1Q2qhY0UWfD6YnNcUY6NZosKlOmXPZAFtYihuX5B
jDSmbng9BR6YF3V+7Vv54ki6XENyVdUAQ5svFgSUFk3J1nirirp9vVnx8PVlnNv9WIGX3WG61UCk
qiDK2r/1gvJ8490XuEAsNkH4v/dyAomtd+Hb4mm76oC6JI6ic1CWBZrUfAkyLoneAs7KWT6qaJnd
dw9REm/wAEQWs1qVunS0GzagXvPM5+kQU9lrhCjjFbgjBSxu3bwYqWtfN5y2LAdu5yIyPurcdn4p
MSUmuNRHiOaE88idIVextYhjxrE1mnlDXm7oYwHA7jNEhpcahi5KDlPY5rQ9xZVCNLjlFDab8Dmy
sNV/wTOJ23RpGDacmVXSOMMUzEx09+X7iqKtPORJpAxyYE+t9olMSPmFa/IkmW767ZZixY66A+BA
J7yoJ7ixw7w61jUIT5e8K4YKLrfurOzNDr6mSg7jkw5OCxiqZGoZ0v1aG801d5B+AF5jm/4wzN48
HSpHvK2BklLkQjob/hOI+oHvKhmmUU6Rm26/E0YSJH+B13pggHIK9wy1V5QLXd6fpf6MEaqVpliY
u1zBD3bsntaf5/mLfr0qYKxfeoIT2s5RSG3o5A2GhuTCxwTV8vM+rU7rG12okP4R3FI1dTKj/4Pf
ckZzLp8JhYuIlXN3VFIs1rpPXKW9Qr+GtPgO7AN2XEUhFzB4UyNpp1V0YyfTKRtSqNJaoh6I3M0d
3nHMA6qPc3SexGYw3Y/VFDxzFdvLyzr3MCRzr2lv/xBenNE47OrfrgI+WjbossHWvjj1JtmIq5HZ
Hg07e+LlRA3nnht/kfFb3VQISbwPHES0q6pvP3xzEUW1tPEQbCLtJ486NYCrRxERNj8MvNVspOlX
vYOciMnlF0tS01wnp1m268a9CFxevLPXdwEMKP3WRWJSsJqTigOPnit2nZ1ar0IFAekqKA2JLra2
M474hAX9Pjm0Vcy0EV3LJkMQHYp06y1uACyyArx9p0AaAUVVBinqzt+s58XVeq9QUYrWspHTzfZG
Hn3Zm8b4l6EQP8EwQl8I9rS3SpE/nhFw177mllZAT3ufy+20LI9OGG2VCFX7uEXpln5x2NyP5x4E
wv6YWVjGpx8OmEpoR0vwGm5RAtWcLOsxcGoD0F7d8QYrBn4lFNMWVEJ7qljzC84BcYBCKGwBsL7V
Rnw96oGLKfa0Nbq1g0rzZrngoedK7pwLAh/dg1cj+KruKh9LpiIjIi8s2HSwPUNyGnVLIQFK7C2t
bhR7xlAnITAnw2AHWnbeAJRzoEwwy8fLNmqXJ5gqmDz8pNYrbEOedOOzYJfIHLinrd2U9mqM+GnT
QletnV7ZxWYl4Mg5GnkhQgXExqTV4qVpVZmkWZ4V/z4fHecxuBfYCPDaJOEAtlsxmYcKtn1kpwkW
7VUEtFDiytptR941nnXk+zV9KzJxgIJ7hAM8FU1pM28BY0FwgdbHECZxRJDjl7x/c/Hg6/YzeyFE
zUEQ+zPhP0sZqXysgZGVAhn50RMIqQvabGywIpVnbXU/mAPSm0sMlSjAcVJYtImDBFWh0P/5OooE
fsf0JH2iyxCTI1wQ8MfyP393OZhF1bDH7vU0Q+6jaKVBQDBxPCVygMZLfgJzB3+ZVeoBB6YJsEsx
rrbo03XwXzXxcAu8VyPVEH1M6vQCEWNHn01P5HhadVw5QYmcBRNqkDQ/hspwE277VxdB/ns4KYJF
FGXk2kGJs1ZevY9tS8KRzvQblB7F0H8SirAaDdGi3rf9Fy8gvrR/78ljSNCOg4jIZVzBpga+gBap
2i1eqffI9K+EUCO70PNDZonGSjkHTyBsLcgVZRrLs1x5p66vrfCnQURwD6fCaO8BzQPdkwKS6Jvy
rQHVhebgOthZoxTu4U64Z/tEDdOQ3069zMvYxiYbERNMUJEZ//eKo7OuKJQGo+Xw5pK+aE4Brtxm
bYNTr+e1/uO/glK+Fd1YCFIM6ATutFsTG61A8tsf6VSWszQ8rb5LlJDjowE48v2ecbhMcSVZzm9G
rU+zx7elIWn4Rw5HLV2whS4js5DpLii5m9yfnJ98lCCmowxDppsyvn6ZRWc0G9wK0Xaoh2JkODBM
dDVHQoBIcHgiXJfpgMf0bsgXqlkPPYexleAwPQI15jp2+8SFuK39erMjAIm5Ue5xvieu5gp46Sea
PsyRQ9rKqv3ZJml2GlCwr2wtSe4MVpgKSXKF/aOLz57SsYgfTvswuUJwyUNgoadiWCH5ljqPFNFV
KB/e4Od0t4mT8hCaWOrXqZHF+HO+E4bVcYGMLS4fK4cdS6yZ2+KaNFveQhR9yltSvSzmljUbCcBK
zSmfPH1k8iQda8k0q8OkRfOaB+a4+PQo5ZaknXFE/ZVhA56bAKh8vRnc7BUfBlkpM+S+tl67tICV
QGzXs6579uaIQNTT7T/owu53w6/6JHPahiENOLkI+aCAG27OcPcvX+Cm2hPsB17lJiIm4iDwteRI
yuKuGVoe49JppnRM1jfH9bicPhLLRaXeZ6SJoeR2jDpzGm6djiA6xj9lm8Um1K15HYeMWpC0jmXV
g+kQeT7j9qd6E6sdUQ2p6vKD1GW6KWGOkSMZkzuiAuwN4qNR00thF0EIfouONCT+BV9pU1746vYK
oMXKwxDt/xqTNfc/v+jFZi4upyhPQiri8Pr3y2hwWkR4REnDR/ITBaC3Mocm9Ny8YIRmism+xFh5
N9e61LV9lnaDEZNmTovdaJOU3ItTW+Kp1SYSkVrtT9FccRoqmRQg7Sw3KkNSXvhswNKy7738yo4W
UB2/kNTUiKAo0zrd9G5aBPzFoqo20U/ofq/9IDspfAZpW2forSioheIXhygoY8ZIVyxSF9VagyYo
rXV0ClGKAEQcEhUrLd4BUwkh6jB9Abx+IvkKhH3uUL5vN0/T0kb0wCIz5VURqNFhHhlVj7yWAnDZ
KE7jZFbTIsE9Z5KgwKhmq4FXPDyparFbcoPa0r3v1HwP/q6cPjjS05MPfFlA4YtPz48r/3ANHNsf
S5f5EZz0CqdLXdl7Eq+VK8HUABfbrzydnkJ/JfFt3EgoxOTG/2xxebX8ClyNYWj1PmRfNgSQDBvU
+1kx2GzrnYDBg6QkEnk3BEo9wiS9agKOwXTTy4jiZ3q/1Kiff/cXE9C6eKzxk024VHjHMTO3e2GC
9xgTxpxBNO/y3VslbuexNPU0RqHNA74+wa7VP+biY58izi4aYLp3yu1X7YXn0UnfXMyua8ggXKbz
ZVLjWFroddp1iG9pNb/k8nrARN3JSWAZZRzyVgHjVDne1S7WyOx1w2T+KXdA4zNn8d5NBPjbN5CJ
T0DPBlwCfACwsYeAtFSvV3B2oUaSXoAwWAuYaIBFapGxz7WnBOewMJfL24Aa1b3lnrecfcVoTvlP
S7G0ujeeSoalEeSKjQi/KokTwEVvy0nD/teIwiMg3ZBxQsLUlt5+gjmjsCllCMjzXWBlqUTK4Lwt
UsWci5Aj9AStH6Uc86JW94pMp06GEcYPChCWlzOGBvKMAPNV8ETtsdiGL9UDJgwIJoPsMsM6LCfn
ce8tdt+s3gISz8XoLD7Nl9QWUy9opZPqFZmkVSM1hncx2Kt15eiw4qhkaRW0VuMjHOcUsAQszuzB
Qwd8oWehC/w+Mlmwo9ljr/7hQSsabt34qyoPdvR11Q5tpoCmGnWjB4236B0KNueUZ9dKdgJsrQ+j
eHoAvp+A25ikJ58UcOD6rj7YMdbgzoFhthCKD2kWdV9/pNswJu2RDbnyaY2aMw9/q4kDyNgwoncw
JWwYsOr10M3O3bP5cwHhOdUIgqAliG4lq0Qr/t5e5V3NPZEOEXAnpf2qH8MuUTaHS4jK7GIWdvjv
WnfZuTKTp3QMYkQX0WZl6Rjz6wSNP9ZWp22NkvNsrJngrykDO2la/iK4l72VEHVZrJwGLFbubgl7
DwqMNpXkynBf/zVZgD6At55A+PMeqSoUpOAcFb9ElFmWFPJIm0BqQyae7S8CGLHtD4K+IzKV5XpX
2Id+x7IhqyZgRRtv0eZrr9ujxKf3GrcfN1gYvv2MVEwVKxcDySQkt1L/s3rwEX6UJJrX4JrHuhjj
WzuviKIOaHtEDZYWWvSvsZC6Mi9sookxpvVaDpFyvTN3tsEmf5ndb5siaDrQdnk4djOEPnX2lZ+T
MqwnkRoA9OuwDNsQuuoUn3FqpAzdN6KnxZ3D/4QYEt0tMDm4ew7uRi14pYL0CPQEECMgXek46ycN
tYuz0+St5OIM6wfCuNI0dIH/UEqfxkrDzRpZCYLcl/IuBCtIAIRynv6v9KxZ/PTTUptu+BK98jzR
UBZsoq9Jd+noXc1+VYrFjmarO7puvo7ZJDyCdn/vS2ESykMxP6L8sFv6WJtAUKlRBdBAn7LbvNJm
Q9ivPt4sbtNXO8Y5Juse3N9Td3GWJO52J17Wov9CW3MBI8EpefYytF2yejpxs/qppzY7bhhTTlKg
W+osDDmHgQoKBWepeVn8ZSflGdidmQp/I8ipk92tNQCQq50SrYc+ejpuvcnoeNwbMaFSIafhm0wC
sY54YexZhkm+eqFJghJlkh9XvRZLjVBweCyBK3XqmivhCHihhUZvEQIhpiP042dxMEfQL6hie22d
Ke5uiREmsAfLeBh+dppC425D7P9F/frIZf/Gqp5h6CUppOXZyxlP97/dns4NgnVYkLnfv79r2hxv
yEbJ7etNnI7/3jcVsJ4JDvNVn0oZC5NVf0cm0zrLBJ+VHfWT+Db/UsuBiOmuWk82OJqBF2k9m0Gc
6Bd0vlcyRE/EFWvskaXusRHXI6DtZ4fiUPfRIV14c+D0ru/gCC0tph7y8yuV7cbamk+MaHeWCGjU
DxXjlhNlCLZ47Rmlaezy4Z0g2VTMTGkVjjyVaR6Oly392Jmiz3CP0oXjVDTBzSxYwWq1flaHM6t3
KPFl5LMQJPG/+gle4Sz2dswnMOEtgTxSzC0vKAFDkVuZd/zJwTroCnZcgYDzcA7lAchm69l7RDao
g94tqaU7ios8Yr9xvxkxRBS6jEcXfbfmrACDQWsTeHo72POxlsecFVUlzviMJDKxE/pcMd4M6y7p
saw+BLKHlB9yEzXaiOFRkeVXgniRwkT0o/Dprdz6B1aLMHPlcTK6Ky+nhC3Hfq3a4hv6bt8+A6YW
/+S1PYMxSez+eDcMmI9FjyPwc2uACwWIi4M13TNa4xD9Fu/El13zorYIacwLYlp9suMpNTuzx9If
naH03/XqzaPnX+OT456j5bmLvk7GGso+SiAw5nk5B+KbC7j5YYuEM17f+z8QjRHlAzz38dOnJqts
gZBwGeKNp4Y6tBwfROuzG55OT4T4VIK+IVN7fBA1rXrWoUsduS0hM7OcMXJfadKGboU9EbAf3O+f
nu5M+mEMqnpXADcVEpipr7oXIU2dbmZ+CpwzSaljVPD4F8egFQvshXd3BoPnPyzU2VmMO7uvJ/2P
+irY5Z8guHxxmqzRCTi2ZCavqJDK5xkHxt5JeHVoN3DLgVDTgu2Nv2n2YOK6MKvYkWQsIofu3XA1
L2xRVBABiJ54F2pUmO21cvbNcgn6IfPop97r84CvnuhJBQosD+4c3aLO7MyyANIOPdsJTag1aNL2
MlQgrZKD4Yx1a6juO5oNxkQ0Y0jCGtUOKbPnLQvOu2SpMbvXpVMKVl5pUW552x3bem/fAsZWMZwA
P+pEIcgWLad1aQ6yrlKHpylfmnXlEuiNV/7kcVlXLMYfYx7IjH7pvnduz11HpZ1Q//vnP65XGUAk
Baicv7Q/+yQqTN3nb4dzaBEbj2LomoSKwpgfrrZMdUY9Hp/HF1zd76ooHBKfIGMp+m41mGHJak7f
9DWq8Phtti9y3RVecpAAAR58xOSrZDbNtC7YTQWJLXqUwJPwuh4SXAqhSjCFPbpOcQ/OJ8Oo+Lhx
yfbkXsfZ9p0PkmKbhlkU2pHBTnJUHseT4PX5C1cPa9jTCDpsPcDk96gsFNYFYxhF7un6HrBi53H2
PyQERTticqiNddf1gO5Lo2uCclqT6n9yY7U6rawFqHZd+DUn9M/YEVaWiUbEXJoHgx8I/+sJ4ElT
FHmil/9pyGWoAxzQU3ReVFEl/4Su8BA25WbWZSpW8V6+2pqI+SDDClHABNRdLoTHiIKcqmbpZIkX
p+xkEF5JwTeRYLEMKMT4svESNYRZ24n2Ou4YB6sfbQhIdeyKJVcIAamarpEtsnXKdzXvmptF4Bvw
ClnqYQGGNQlt9l1OaJUvtXGrmKGdxcWaAjNu5Rx+qLzX04dochXIUCIz0FRLSgxkYzTmqSXJKODT
cmmU2XMIbSaG6Q06VgjKonGSIi9PwF5VIIM4Bz+i+As3vrj0YYrhkcyhGJnKWwWOZTwZMQheY79T
ZSlUGwl3sWq+OK9VvZBGgRTuvaJEV0RQkcsdl+g0BK72Eheeiz1GEBC05uE7U+B17s1hd90hK2xG
BcROJTVI3lJ00DBdsbRfFxwpP9MxVFxBCSb+HmOJubWYEL5Qn+S/Lxz5BdFqJWQq3nTNxhJxGvVU
uJuMly66nFCBwXF+JR1XF0hC5SMb7YkFyeSd5J1SdscnaVTQqyYMrQYBg5Zodp83Wt3RZkC2ubxi
FL7ipGOHckCoc0MF1kng8OnQ+sUh99PkG8DMX/54xCQ442HA92oh2ud79JEyzkhkA1LbOq5eWPn8
ImujUOaqfA7kGm4Nd5CiaPkj/e4Z4m+oKeQIAZHPEXR6cZN/EVJVw1AJwsDsIuVLBbMZFtVwsprH
GYQKs0eonBSndtdNsv1rTKpnlbHS4FU91hAIsAr26vhKXVJ77qPvHY0r+wvU55jkkWyCBeNUqlHR
9i1vqhmy8EuHaKACKvyfDXR9jx0XTuGjll11a9g4DopanI6I1G+P36Q6eLZ4YZ1b1wxTSEIDut4U
GYu8YNzOKbW09zCgVDcsnwxFjo4+RiljPnGTwmxFIEHwgc3vwHqIqBh8IbFLc4XQ86kILmi1yPxa
gzAaK/e9tyqokBJXEgEiOGNwFPM29lZIiXkZJXG2+QmKbgW527PLutZO4Nxd5uYbYBmFPT2ttnLq
ajIecmj/PF7IUr5kedz8gBhZX7bK3YofaaLhYc0sCcjsZiApfrUfDZ3R+caOC5lZJsxFDDpvFCDj
is2W0aKbkh+8ngyPhCOQREWgZYVvVOKzktTnGX/u3D3S754xKNGm4c4fXFrBSkS11kWqX0JL8TCO
ep0M81GU9QG+biLLZr4NmMKJdAsCdoOYF/6yw/vaTa893A/VvfO1A4sDAJi8PjfMA5rrImMUEKwb
uzQpNrbHNxk2LJzdVW2fpsXi45j+uhfyJ2qgRGs8V5WCaYBimvjfm5VbbfPbww+83DSX+3P5Bt7Z
oIvpioB6Cu4kxZ2jQwEWWC4u0nw/9h3UqXBP3wTOKV448+revYO8loEJPBi9385FTtr69kxqUgjt
Yoj0Ll/AoYnHWOCzMDxXwRcAI/v7uxC2DWp2a+3pT0//rKw8zoHLGEcp7x/nCyyDoXG8+j5PiiP8
g9XqfyVWBq7fvssQ+Z12MRwnpgPoGT9x5O4MWKTCgM6GVOWZ3NdwEAOPt/gu5fslfKCB1mklATnZ
vgFjcbOw8KeQ4Oy3EEJ4ONtWqE4snharu8tS/lG4OdwDUKSAcWqVU3Jsi2iSTRpx3IxnLr3+452G
DeRfOIcZn+vc/DovW+pXV1F5i/EZK2qgoMGI58uWe826mWwY8RfQrog2OUaAEeBTSZ7DJdb5/flj
Qdl7TqgPFGwu2ZZ5M+ARdSsFw18VoGLx0ezY/TtplnD9ron3hsCK0rzmwVzPVaReKJ5JJJKmkn8z
50YTzHtzp9SKG8DkxTDSNw2e/sr/Gdb6eEP8bg4HFWXc+G7h+Ak+MwXVK51ZTbqFT7c/sTLpK9nH
4ZwOQxT0x/z7biJVxZqREuKAD44UJ0G5jtWbYDmivtrGMODcruhozs2CLYv9+XFi3ud7dAswjjDI
D4/qTIGrW99jxT5t/3VQW3Dsf3gf4ABBAMZO1MMh8jvk9821mc+brGydl3YRXxJ7XQj6dYhes1mO
gtQOaAdYuUjOh4wJsu8f1KZmYUguHTPDpyRMknhfAUXPtCMKyJHWnac4B4VOQ+eSPu7hqGedKug5
+34i2CoPpP5zvv1p7qGlV5OR79wXZZh4IX86OpraG8KPimJZEufSlWpi/vDUECpg7gTRbyKyCsZz
T+mi0u3I+bDpg/1kBpkM3WJdNXHE/D2o/rZucxkFb5e0nTqzaH0MYYZ1uLHoqRYfc3mYrbjv0vQ4
2nG8k2Y27hhamsM0RTITDJS23zFWkxcj4tAXUvbxqGgpnVkRuZyru0j4lvjPuUz8RKpM8uHKraDF
SDb/oNcFjIUtMpBrFV/taegjma/N741aere4E2i7kWigwe0Eac4q4RUOAZDTkfOyVCPb2HsnHP4S
+TKgeu/fM4em+khx3l+igQDIcrqedwrIqdcwX8tqZBxoDvWwp4zf3i2aGLXWcn9z8+MqtyuzoufN
3n/IPEcmWVEaukCyVRnWaojluj3gJ+NVM/QZ2+gmQtenlsuFFUWqTgEWW/9Or5mHrd9VyLBU8lKQ
ICVDSnczce0z4tyoVLjwmwje30eAhM9GWeArlS1PO+Q9dhcSllml0YTl+xA5nIocTh549ls0OjR2
/5oX/MeJVtBuWtUzcZJEV2EuyO+u+CtGLdOK2QzQQtsHuIvA8SmVVeONUCIYj/02AXenP1+I6g2T
hkEg7TW9AaS5BwJ+BiF7+qPrQg1YEObfK4K02Ghs3Jg3MTfSdv3UGGdqJCpRvEwipdwHkG9Tu/Xo
8HJ1Eu3+TN8IBO0uYnpgk/WWT0jua0HR3B4dK9cW4MTxRkRwstlSfz4INAikV/IktRmIWeORmRcj
m14qH4/9D4mx3kQkR+9Yj60o9D54/T6WjZ6Fjc531OFJPJ3bP8JgsFvO/aXipC3Wb4ant7F0u7Tu
0Ykj5bQ2/QbhBuuGXa9Ers3iwhOenmEfpcqSqmkYXx1oZoTqZbbLIK+dgRmJuBQpJgYu+bhGuKnD
hzlsR1PBHGbx5Ogk5It3aULNAsW4gmjpgzBEGyDoN4hWaO9kuJPRxoG7l69GJe4jYmB5FJwIhK0+
uhoa6zWMv/0RuEGpsEoYzUdspoyKJQ++QYJrXE1ThQPGn3nKcB6qAC64xyHD+Oj3Djj+EpaNQhdx
sqQWRajYe+MLCiaSPvJEHiI2EYjosbxs5O6ODgAn14ghhzaky5Fxg1il6piVOUGYhmnRtvgowAgM
OVYpVooQrGaRKduYhSvLzBRMBkkxMzc7e6Y0EpdiF2VIlxHpvAJ8kraRr+ApgQQAg4hzLSOSxxEt
bUVnNFTmZAQHBFRTDLmzUggYtobB3DvQ0kjfJoPoHxWdTYPpdEY9vajcbDlhtYkumRtCCjog1Qax
wMZlcNJbxWZ/HnZUq/xUJ2yYK81LVRftf7S1e0704tWHbL0CYGVEWPFoR87S9OPIWlHVdRWe/rRO
1ZY4UWZIY9OtHkAsqhK5wBlpCWTXJ8z/UOSh1sWP/2jJhHHv5BH9UQ/zqe4x/jTrgLLIA9aqIHV7
o9L+0ZrIBNnwruIGB642s25zNXIN8/E55/GzPONOvmB577PaQWv/HSM3hmVgvju8fiH7QiNqHdIl
OjITY26V3SnUSTbV/52iBdEvjdbs7Xkd3dAgRgBkJhswazbA+eXd3NzOKmSivn9cj+xHwuxg7yw/
Jx8RR8u3h+wGFXxPWWmyaAL1332Sh7T1cUfwjelqNz7I+1RmokUVoKo4i891IBGKZzzWiTAleyyV
W0icqG6StkbnWghwfBv3x5Phcc6WDbQlVQUfJasNod3ME8IjjV179d2acI40Nztsmo5/gqYkPMIn
FPM8HkMX3x0vPLx1+jLXN3kcuJuk/WNO4pWEUTHIeSftDMP9sjyM6cfD1O+aXlKEkxdxwaSkr7W9
uINxQ0HRguvy3JyEVvl1CkGVwR75vUzEmFK699CYqGWzFf9K3DFahpFLpw8I+a18lRN3IYAXtcYJ
LRWd/c0JJWWuqjAGSj975iIONaK9ckkMUJ8Lg51cEQOy6LGlX7gNpQXx+nek1nmC9mE+7HA0ci5P
jLPElqbubqz9/+IuQZZvftUjtDecM7O7OIpHgrLc29ndRq5n271rxW7JNWbcNQx+Z3NwbrnEBLg8
qO29nPzInEbQTFDSAM9oJ/KFlTziSaKJwc0FkKkg/wK1MJT0Ny4/DPYVI7M5pso8/fXCZ9cRM1BO
WJoT1HWTmtByZblVyr9CEcv97R+4ytU789BlXuU+HSyiTIgU90bYACDcSj/KzxmrrLvhwS4f/JIK
4kiQWAxd6lCVmsZe4MXmYhdFv34wHc43Qb/VYpJ5pJwF67NWGsgspyuUDU5nqcbQN93i5EpQCKhX
n9H6ARgHg6U7RedJpSTKgmj6gLhimhKPLnHYQ10PFQAnX2FHFOuS3OXOsK+U5oZ+BfLU2aKpepPg
cFf0TWo0PrgktNx5JcSjShXwGfbGH6PVqXhDdFxrcWeUo26YKmorXytfQz1NOqEo7CLfSHIiILa0
YANhwkYSI0mYG34Sqz7Psdmm3nPYi13VoxyulRFVI3crMvZLW+8WwBlGrfWKAEolrgV5xXqP4g6z
0jyoMTlXw/ciwNmjQY0dAUp7vlphfYAeACCIUPfYlqiz4k6ubymPyO94NvkuEDEOxr69NfeBAcSy
RiLLgUBrL/VcCgbAE20weVbXOszoScSte/ow4P9rNopXc5mvvAsNoOK2AzfW0VJ5SShQnbJUfGif
4Og4sUUXdknuT4o5IayhlOOgaLfD5//IjMUzERNCnJiurSkdB+KLjCjabgKYPm4+M/2sKMiPpTxf
8HuVV3izMVOoyqCTwUl78Wqvm7Vy91twOb2ZKyGrBwZ6rY72BGA903FqdiiDgTxKixFOuh4jnvJV
w+7QZDxU9JnD6UA9xfoqgHE7Cd4dYa+8ZSw4mJAVc+SQSYF0bSEh27ZAjI8prseIBLidRVSCnRJu
foXzIi3q/71DRvvbc4kFBnBLhHJSsYv5w0tYBDvs7jklMAs82luvXGuV81JR1NjuDMt5Ot2gbpO9
yCdPrVS031GnyrSDgpNaljDXGTqZBSS1Pemcflmk7z/uzlooNTdibTMvVywCR4pjG6gctK6lGIvW
Pzxicb1xSPv69EWiKvyfl0wEmsky8M9L+YhpMiS9b0mEVlxIfFYJ+qo3WeB+6Y8/K3SwJmyf+uTG
fcbt4qwaXil7XA1txEhnHlyZ+tcvBrKatr9iSSTQJPlZqOuRJ+n+O7Izod6cNBEzBR9WXywzT7CA
Alu6tjk7P02MFVK4F0UHcU4IkJAXyKnmJ4UhqxgISi060kVlbO7GVVQkTM8tlJ2hVGnL/pvbKCYA
TgsDvDFZ14P8/n1FE1x5Hi16gTWNyDUCxbZpG9ovvY/hd+j+UgR8/edC3+kaKCWTUSpWOsQrn4KA
/hOJ6vb/m238g1pr8hqegLvKXuVmVIg6slTG4APSS0MBPiCtU/w3iYjjQNHhlxu5jeVJ+hmoIEMp
FdliXTGMKK6ocy53OhQT/Ho5fDo/Jsef57DF+ECDjTjx5wi0XBUHmzg6xUoNDozkQsIzn4M1nxpL
gbOuaOsMTgn29lDKkTOYdT/lcda1FgoPKa4dHPIz6x/uItOeHixQiAua7M8xu5kE4074RUESuW+n
v/L0TK6R6nh97vnPqbW58402yig/bwhiLDQFJNntvMttFs8q6fRGbALcrFyLkSeYZHBdMaMgDqfb
BNdYQXhYDfdhI8DlVqrgYpk5Rg0U8B1nOuvgUY2wqnQNr3ytwdMtc3UwAEFdt9sGh6CcfvXjy8Jp
97ChDvA6aQik2WXwscwvQV7SLwDnUrZQYpL6quajVOXbGY5aMQAzMZeeOpbkmcLCtvJ9/udhxsnE
BAQdq2i8CvDcuYuy9AaxXh3c6fjFsmRIOUiQuX0Y350mJzWawusPZUNM07jJAn5Fp8KQAUKOb2RL
8nXCMSHmgstNxPX6eSV6HbIXlqGrTSSgjtqY4IT7+OepgOf7P1izttEZLuys06mIak80C301QOGq
LxsmTAM+pJPqPIbHnsz+VTlmZ5u5qg5Gx4ZO2R1BBToscnNTBdEK1rIJ4JVZK3BHrdpvPJRcVb2Q
g5MuWcEnIaoq8YsCQCBgbmkBaPZJAB8FZUyMdp46PHq4do71FOOix1Kf+s9v7xyZYNgCu2tPjxTj
jo7/Q1QGY+nSnuWLGo5MbVIKsRfCaaF6gmzh99CPyuBi88XYQ5QpxWc33nxIm+HsJA8Tu9eye4nI
opZBcSGX/olw6V9K/BqMFUNPYf43kJ00sk3dr4USSZACbSjuqDLH/VB6eZi9wn65SOLY7ciGmqfb
Zg4ETt/jOr533Ik1aBpK+TpMlFvUykHafadpXK8FTJE5YYBAUXDCfxYQ9KnFh26t+Z2eZQXP+f3z
aFdNROs/xvgcXZkWyZCXfu5QO+zbYlfLLgivnULZVHN4pooOtmtlDCIW6u6/6trWaFyv72ozd7Lh
m4yBbpUgmgWItanE9cmzcAUuIjO/AshUU+hFEQENEa5A/QGy7dXYUzEBt/Pkweax6mtEraSvBmkj
iE+HqFoQq1FNj2+3BEYdk4/IYUfjBiX+upB9Tw8UT+Lvstq+yQQ2wvqxQpfC4stn19AQ2Y4EFD6c
LGc9kUG9ukrl992fXQHj19RyjC4GHxNABuh4SzJ7qDi7FT5rGRxa2134ouzwWMSfysgEc3xNhtyy
n+R1MNGafZjTostwYxrABJfL+XsueUMNzmWFSwPl8sjJwrBg74EHUGmFvssfzNGIS3ge/u7I2Klm
qTCltih88tDHL030qge/F+KiBDTHXjWbi04SRSm9tK/MP0WgvQaHJGhdDaRV+EKepjllz8HQT38G
NBJORlO4PjvmhOd7bpNLxXOydGs0ZNru53v7kTYBzxNCA2b/SxnwfBJj/lTDBP47MS0W6PqAx5GD
tyYXP4aPdypynhdXr/K83RA4EqO7Cuye0mlLRk9a2xm+utHVezqxbq8t9128XrMYJLPO6AAmn2Z0
9hOC+7xZSTnAqbtg6mg5c1tirTHUkD8lrNayccknkON1kJ0yjPAxrpnukLHqKunaU3Yu2/t4Obpp
dF+/ht+x6Xcbnmz4orQp4v8sG5rNlHTFZ0atwaqJgdyslRCmZWOsn7sSEGdgyRw46Y0wbWL1ou+G
X9Pnildl1aQI8Oin5GDCfWiIP7BBGiZ4+l6bxNvBhV0sYWy1uX8Wqaiiuoh7syR+8ysFdDBgt+uv
zpzbO2ZATRPPMPtjOoHMuLmBvz5o2MrZ/7d9fp6EW/ZJ+rZWIYwU6GCekaCZk/fP53I4gGIdTezM
ywflpN4KQyCLWrmy6vGzsVSwmSD3+c/GUrkjun6qtkZGu/f8LVUeDWQT2hnFx6AtLtBz0WfVZHj4
+CyRoTpLqsleRTVupSimn4rvhASFe4PxXzyYvWcndGKdGtWqv+RmcKj3Fm1+1mSl72rzGVgD8JER
CXZX8L7Cem2+QyZfd+GkGtNfD5dZPNC70Co+TJjr5PMbqyswGsbH3C/wEF2lpdW9YTAz//YpOKjS
i0PsUQfn0kXjrX+2EkMOvEPkr5QsRxhLKE3GwWHADn2NB5K6/bUlMtezE3gRuIIv0FcZhtTZlpAB
zTU5g2Z3y3jCv5zqFfMq+jYEXm0vWyxgeWDbrPyphjtpm3QotLOSvwVTT0NevZQ+UapIkgY3mgcO
Ipl4uiFgFqcVRJMLIMfYbJmhCsVdP7t5qWxZOr4JpQW7meW93fNIshMdksGBGoNK3QsCY9cVWy8g
eHF9uVToQ4jd5RE3Qx34DVV+DjRu8t/wKJRNYDYiRyZIgel2Ve1i7SSupC1EIT6i/yvIY5ljp+GW
8up8wNlIzqnPxHiMXCZw6SIlw+yr+AvrMw2CJyWhy8UOG7fVOsHPlEvY8bscJcpkPutMU4KgTRBi
TGPZRk/41bDpn5adsX6e1e+du7zXLdPfeN00mxmqYW3HoJ/wtNvBqGyHdEuB3evb4UcX515HTVbK
AFsIrfOzTHX9M537f1SfXENf/1Yg+cXDa5RWNTo1NpEQv/vxA7rprYMETKTLLJpdF7GnRLx09BJ0
AwM5kVGC/AxRGAK2KCuPy7Q7PRwWVdZLi4eY21g0E4sYm073qnPnu98ApA72nEHr/Pf6QR60QxkK
+i/dmAiG2nwW4Jr4n7o3bIsDx/7TB0fW7Xvqn/DgfM5yfwCaQwLqZezG8NPriS7uwDJ1CVX70m1N
jgE2YSiiaVZ+zsxl4nv5+qJMbaq7Z6CgnBbFK0O+1CYSP0r1W+cz7O89rXtZppSAMoTGbLjvKSn+
zU75d2+L4gRgZ7Ojx2qZUo94mCLdaW9VD399DSL+gS2oLgqacYWVJHwCAdwN97FmFiirMkcX0ZgX
NBc5LpUnIrg8Y7A/T/OK+pZIgAh3DEZVhixdlOVAL6EYXVVep6XE11cQqsHKhg8HQRgeviXq0aun
KC9RaoLhPdlZmZSVH8OzlZFiNEQYuevmHLew5qiwpZzKjcUVC+0Tgmev1z0L6ZIgLDutj4H38isM
YOczOW1a8D3yu/jwz9Hzp3kMkNbUo8tA5xXRwcbPLjq4L5Y/GPYILZhfE5uaNKgnk0rLDLIZolQx
0kMhLtgRfGt6XcF0jwa4vVfUwGmueLTvTovX5nRq2KzeuwJNau6omSj8edfN0rKw8iQa1oAuTIKE
/ZaNZm2ecwEet+UhKt9FkV9xmwSAqde9oZD/aNcqJfIDt9vUZ36sjX8kIiB/F2j7lc6kAVUrzaVS
yPZOdITu3X39qgDbZF6BCQ10zb2pqDnkQ+4YzGKlTwnN7KPfcOqYNxKBaMR21UqJuwrmOGEKDq6t
U0uuohBELY/Lr3qGc12dPj1kEh/tWptzoRJLDVljUhya2PqPVHn4xxHKApUl8ZVZPPZsadyn8b8p
ae9v5QDDCNyQ94BEKPQNUV2BxGqcDFZdGlyjOEOUfGUBiYK+91m4ASyRPgXYDqW4b2qupAjgIbn4
tUv+Yw3W1SDnxHnKhOMWyouUdvRfbSepwBEZ6krf3DuJv3MiqMwr2YVk4inkojOY5ATLl4E9sYcr
VJOnu6OWsKmUW+6uV706xJSJmZNLuT2FICIN/ekKJKSwRtyz9duzD17DozIbinwHabGUXYK4NZZy
nbckjgvmonOQha3aNMWgqssAvfNxGXYGjhZ0spxke8sPO1Opf5ShYwEq+0WLqnNg/NQItxHCIXNx
mRZfwXNIxaJZio8wFM8/wZuez9bYfSbaON9bssYZCgw2/mJQlOlAuccJYyHa7EvWmsLKA1J8i5pU
pDZSGxQSI7avzbgWQ7jrcyyCxXMDI1Pov82b5YBmHRqPcC2N07Rp/7cxvWyKH8ZzMOqwP9wf/E0F
ej6Xwg10Tuif47HvMN8JPO6LnT4+1skuS2xXn33U43ybQXwNkpjfF6fzriXUy6l9az+4fgiMQvDN
ApDmAjBqW/p2mnMaGYmCB8tSDQmr+bVT2dZmpZWNSqnQY9HynVst5DhrRVycTafajNltvQMEKB0k
f2Jv/Vc7cw5JoGLOPIP9vsQy+Q4z2QRnMf9hVYRHWeV9VqQn2bcYf9tfNyE5VHjcaWoPJJ7pv8F4
86pt4heTzSv21RZ48zQGrKnRin7I47kBHmxQuq+Ml1B/jiWCmO4DIMpU5Z3p35qewaUbkp+7GvNU
mRP1rWi9xRqOkyD/dJxxoEFdYOF7vEv3TQ1Aa4auaegkFq0o0tYXaU0rPGRe/Fj0bARZH+Xpi1WG
23n4xfxXZuX+gTuQI+oQynf2zWx59zwmaugLmwDhrjMqGN3MINWMbYyX3yXyn04G7Z49G7xqXGRS
gQ+UfC/ck/05ESGbwZhDlpaW0ZCgRuHLw0LoFcFFClxNvjZFp52jTbeyHG4FLF1autOGuY9qFa2y
v+rNcZMgIV78eW41PFOhkgIfgqKVoHVaqA1W6I618Bj5bVZ0pCMRaRAxgqfojYtM/fgkTk0ZDuLL
DcSiyp2bpyOWQxlfKb7dFaIsRjnPWTZVR7mmXJtv7v45lmizvxKFwz00SIUrC1MegYUJEyJAH5qo
GDjm2ErmYvOTsLmXXF7H8VyLYmNZ3n4vNo7Dz6fctIMR00iDvF7BX4CnOZ4QMD/hGIi4SEXBo+KP
oUuWscCDOCSgCEv1MEC+JD31SRP6EP6/br4zXkB8KG/gRUXFgOXEkmkqolYHcDH5gzwb/8Gxik9l
EOqCOBsQcyArViOBVimzyxv5NXtpSG2xXHhwYz5f2uQLDG7r4GWMCHJW45PWWAQFM/rvbvH5WTab
cy96CN/j5zw9ArLei+LEIlr/X4BgNda5PzRlO7857iVii8QR0M7eUBWo1R6NfWmYKSePYGLqHw1y
amkG8ZhU/h7VaFvKC/x4prgVXpJrwoVVu1yD+n4UHaV6R+NeI31B5IhTWSh893K4ddZ0J76FHmBE
BI/aJFtLzRQjSkLIB+MM7xXDGayac+tB8a9t88Mbm2j8INy7Thjqm0FOFN79fLXcItr8J+L/NgpB
V+lqmsZRBY/pjH/QnhIOuzR+l5TG3LvN2I5seFKnn+GYTp/lZ+U91vkDlhMtGCWS2fd9BZ6BHYY8
H2Rhq1SIITuDy4SMnJ4GxVkga5ZXJrns2WMtPobdKprJZnGIBLGGAtfoawtyM9EPoY0E9ai/+Kwd
Y5N6nFTZO3EjY4tULeBhO1CM+PCqFW3T4PbTVnOCWKETDMnMi5OepXKakDT/C38ZzQ+nXnRZacbv
z0x2vmTQ0ouC3PZdnMlAWTm3dzx8OBborbQLSlw8IVer63idBG+NlHST6GbQYWN9p4AZAC6lmb7/
sX1YAfan4dZ+zIDVFQ8e4iWNlx6PdsiMuC7fnpdpRXULiDDDNxe7JUByKlzpnblPs4m7coqrRYbu
jQDz1OeyWKlUSICm9TpVBe6U9t1hy1ZkgxWF5amSNyJsz7s59uNfyiGxcZoilwf9QNtw1dvDuchA
kPwwY7CeaswDoevI0PgGfz/zR7R8vcx1et8kQR+OKEXiv9X2zKmQ9pqmbg0jCxXZI0dg0N2TFYC8
PrQjCorS9nJU8JtIJzAlxKQ7F5iAc/1uV2Jz16P6AOE1xfghxNxw1Y1wY/yurhD9nvfE1EcWv/xb
0aOd1M2Q0Z/wisKmhf6q4z1+llRY/lyjGzooSsdJP/UHdolgiEcnFPjeU/byB1x0LnjU6Rid6An4
s/6Mofpm2L6WivXV48anIack3bwT3v/vKbwowURL9efv5dK4P93NvfbZoZtfYyFTv3/gqt3COR9G
QyFz+T5VIv46uqIBZh3txdy0ms2cXmotW0hpv7XPk/9LI6sApbLjbhkRWSE2NDrzXA5f3qS7f863
3/jeSmiGFKhHWHFMXiWOnMr8qsYPzqDLLeUOpauB/tU6wk8TLARrms0sUa4r1POkZyjfq5VfBTAZ
c/1kOGpya/m6Iv6WHbo0XD2H7jLBvoB+0KGS9Jtjw6QSK8ji1IvosZEYaL0HgLxfoOYX4OMzaV2V
uupPZwey2XEqrO8/SmesntdDrHvTQ0yzOsve5tQZhLPueZJ/HjfNLLY8Pq0BTgWwWxVD3y2bPLjM
9/yYf6EWPc4nPsKfTQEczuzYq1r7iJ9H2ownXTi1VFYp5XYRidSnytpGBYaGArqz1Lc1Sopt98XI
OHlXm4FEU2sNoI3x0NJ5CnBEjHy7+0GerI8WXTXyBxOUT0X+hP1iBuPkNT4Bo5pyD9O0ScSbsVq3
0azHd5l8OlunrhTWrtURboEUYDIabbdqk6UastX9ZdJgb1tUmEdz5s4my/PGvF0x9no9tkaDSEp3
7qB+FpH9AEc1blZuY07Io05yYrMEvthwILqFlc8UjK1n4QbFToOLmdS1rBtDWsiDuUno9NZtNkRd
cd1PVw+ldE6A3G1xDthS0F0fbgN7e7w4kvqXUzwLoWFjCm69SB1eiOXnCOF9jL9PJ1AKrm4OB+5J
0njeuTeZwA2f0+zSKq8EWTVPrwW3ZUu94kKHeqRb00aOJ6y0hkvtN1w1pLv9lp1/mO4I65bBVDxr
it7dEMmQk6PcFEFbQXn4g+qVvwOg4yLu5lsiGAt2r1fjZTLTufoQwL7nYt4OvEtLYbeUglSOzaQL
dwG0uV4Y/jWq5zigTIiOFt8bGr5NecIbPBNzTqvOPdtft7p2RyeUoSrgEy7sa0ndgRZJJKGSX0qq
zU7RvLOUxuCs2pDSNGIWaUfG8aXwhNkR56YJ1ktp92VJI5r1M3iYgCYwfWrQjFIJ7s6CUwDZ+H5m
Vka+Al9CkfoJFm2miGznCRjcNXjj/p2xThZcJ14Am9kUH3OZ89L6m/iRdDGSvp7z36urSM0t/zxW
CHaYYDlTjFO6rTWQYlSZjoMqrqkZHBHx7/SjGGIibC/o6iVqkaSs1/8o+yntrdSP3bXHhOVQk3ux
mE5OGcWW7UYDdUObXq438duwtvE1p7gtbUQUlfFr9UPxBWxohzbMPiqe0++CU3jeV0Hc/11gmmFB
kjDMBNrZmo8bQv5EknEyqLQMHHoKCyBqnG42d6Oq0APluTvXhGp0qMQjdq8RQRR+wlVYpZWcAErw
Ehs3jym42LgHrZmCenmoMRhtNFctytdN6SuridzYqnPPLtvqYo7fMsHRg+sa1TJiuB0tFU7qFY/o
4Mf990iF0M/RnfBOpCi+MHockgefWdw8rbU7xlhvUeLd4ZJvU0paQ8QktnTFlIxYcBRoGmpUVdnm
MniiDhYUY/Mc8uhCNSDMeRl5yQJ12t34QbybHhsj9PRM/GmSRUHAoIAq8L4717rArZF8CsRxoiHq
vRBJM5c7hjP+SKqrfaTzRRul3XNXPX3Q3HILochs9Fer8yyA+12t6/7K+XDHz6CdMqktzzDtxVv1
j5Nm02yg6SONY/7lnz51XqYki9zICY2dCDEZOZeKxogMd5ALqE/EbQ5qlcQsPC+xnd7tbvdusjMo
geFkO8KX9H7UedJgzDqLBorTrwTRTW44MPZYDjz1dVJNFmOFtxRgZ9l3ZCztqJk241AkZ5vrGceY
/Q/4eqMceO7P18kgjxKDZNB1stpvqggnKzHbT9nOtNipCjY5IHcntz7WDv8pA8TLw/+OKtSh/cOx
dKE8BP6zqzLGXdTdj/+0kdjQniTx9jHjjw+Og9RJnTy82MYwRvt0uk8eGd3yW4yzOIwgVkDSYTaE
lILrX+0+59uh0Cy6Ub/Q2i7LFFMhuqp0dOsfOVnkq5Av9RhjFwLzEnGz2stORHaIuGDkPP+r4x6o
dQVcvX91WgxaKgAVlQoI0bhl0NKQIl9aT664ZDHg12B3yRx9X5fbBQgFI2Bro5FaL/lggFfWOK3/
A4sD6i1cETxzV5GGHT18Or8x0rVfwbErXAUlHD8fxqTqTuClGQ8WGJMR3FhfJ/Y5uHklwjPyEQ1A
tfYFXIqVjYil+e+c+sLYi5n48WZ26jxPw91ieOCr35E5tJxkDkUQr4G6mxSlR6XFma3dA605E2On
2tSLXWFnvVLtWQ2Eu9D5znNsyJJgm+VdkDseWGVWKXwzUdOAO4/XPrd55Uq2P/Kutq+9sO4/AjwY
nVhTtfwpsap9QLoxWOa9tdt3baIiHWFRAeLyEWDW2//cTx3E3CNhjopxT9iMOYBzoopCzzbtZ8Da
SDBC8ZC6t07X9oB0Y/dVp1JlqaCYksOBCn8AzjDVzBPC2vz9rPKDr/gnFhWcZbR7cteYS4iEI3Ll
BCN01/CUAvwqUdRrYWYjEZo4ZeBgFjV8RaZAY8tghcRWDAeOaK19Z73sTHQ0rzpIwKbplB+3Kslz
48K1CRoiEvUcgtOIHVbscZAuwR7npWt9b3XvgaHLPg7s4dqBaFk/yksRlZ1If6gZtjqws2iISZnp
/I0aUTBQ12vm1uuF3gwKYBVllB0g8DfOK+qpVGIkJPSKNFiaLQJep8BlG6cUSL0I2W/jw2tIj5i7
molx6ovt/Foo4Cvq3MCQHEpMv8CH28BLBvW6Q4hzHRfLQXgxtMcARd+SE0/2PSoVXQEdvkWLpw1p
l+Yrr+z9PMN3ZRsePS91FZUD6wfMdqmYQ6UCJYZd6MtMzUoN4IiK79wsVBxtS4UP3VFf7XOddKu7
mPPpIP4686gyhemjCcp5RbJrtlK0U8Rl6tDZIMxLHYNNzKNVxg1uJvd8YNeEkG7+167b/MfzUd0G
ETMyLJit1ALsSAzDhsDp3x8pf6H1sCgrhh8brNZmc0jo6+N22Y5tbj+E+/jux0vC9GPh+DgleZbs
Cw+KVn/PJ6qb9TaB1J2HWFPY51hf7P+HXiO7BM1zKw6qf7tcBeC83z/9kXFTb/MrjjI5/vdaKyFC
4WvUjEZsUf6ueS4MGJvGTFt/Chr/CzaE78dEv24PsyBDW9RBROH5NWaT8p4BlqQrKi596o22A4gM
FBh9R50AFDNpm0dzmfw06K8HAWECWq3A3ubVAE/Ha6gfpqW6riSJMu8+uDl50Mah9l9SuzR52JJu
+Upm8D1Yyu1+Zynyz/3frxwUSsh0G1gY9ooOpwyHS6yH/kPJXI9Q5+U65C0ip5UkndqPs0Cqfs9j
WkdaLYSZ+2eff7yDbxHkrF4R4thgVdWjfg4xop+BejawcJgYfiutd8myXA7JRlpArgIBNIv/ZLPW
0RLyj4ifLQbXHj8nLmvjgtlslccTfGCSpmYdCfoix4BtkDxOlmE6KC64H0orVdQn8RhRu/XuM4tL
ex7nVCQBtJXPO01eQ8faFkz7QIJ7XRovYNbiWi5wI02ShCbsYg8TF40GpKV8F/7OEwWHFZYqoFI+
aUVTjGZzUbBA0Shso23eEbgkQmfP+YNvOJnQlyA96Lnmn0zWihMInKXNzpXBxOU5Il6iJgEOcgvX
4pCQ6yHqL0Ym2xRa7kB90c0flFvDkLZNXXfP2NpUkTZ3vbGbhLM171I8zoQlYOtudTUvfrTOYVqC
KTOC2qfd+jtZOOBdblLPBrNzuZx8TvypszLEdV/onkdzzHpIQu2sQbzuNmYZRpCg0hPGAWlei9hB
1Di6oIW471LJvVagd8Xd1qDrx3wc4nqLVZ0XYfHiWTbOknKRyIDFJHimt/eGd6KBozD+OKMXKjR1
2cjZP8EXncsk4wfeoOJclS8Vvgrvi+z/xSWHf4v+63UVtjBl0gJTxtRJQK9GfZLszLhPuCPRIu7c
23Ah55iWdAA90N34ZJKkWSSLZzwa1qzKpWYnC7CEl7REUhyQT2cy4we9kCS76IkIv2ZRFrvvaW7P
DsBwUColYR82VgKcWXeBZPOqMvRzI+CCa9Uz3a0U1yoXk5QEPh9aUA989b6Lu1fSJxMtFEQ06XNZ
G/Vq+U+CNYPvW6s3FL0/zKiBawYxj3K39pONLG/LmtD1X6R+USIDpbwTDatju8y1BofFJINd9DWr
GWKYquwKd41mM7Cwiq42CdL1JPgVHp+QDw0Y1cDeATRTOywsyOPyTBA5lhmMf6NomUz9/q7/zprz
oxNrcUnextMC+ZYUMDb95tkFQ9nk/pZhYDpc2EWF/imHhGzXMxt1gY4ZnJlWLt8hnHV9JTf6VWxA
oUUeMqmPMMui+tYnwBYzCOw0t0qoiQAyV6AJgHAbapVeeBoeSHF0zTN+eNciG63EcW5MxdmGVREf
vnz6601bwR1ZhaKjAphwGCUpOK83QcctpaDN7VNMr5gBTzImllrEOTWnXtgHJ6dko2QHJi+kO9R4
h6+o1dCJ4rji67WNAVWTOCS3CFFVAiP8a73YXRkfuVU0QDJMMKlh+4c12BLrjIl+zI3t4h3ipnUG
xDndbmgY5Ea9+kt3Rpuz/H8p6wP0P2iPPCQFTQ8bu+Ei7MjaZ1LVjpYOFQKFYNAN6Na4+8tXaWaU
PDcP8PJDv2Bf+lLqCZqx7N1kgq6/+6JW6Vz+e+/ZQnG8DzvbJsQToP3HjbQrUzlP2Rcqu7HqKvWf
WjOMC28374jvYkNIGk9jmrcMm0w0j1fcxQEiw+USF8WScGnpTj7t38keQxcImIKk9LrOGc1fcRJn
znBoy9MFSkoDefx2sUzkDX3iTdtSUgsXnFz9Vp09niidUJayj6VBPo1LHEMxSt61j1M7rJUyLqkI
bpMrtcTlF30N5lgIBo6YOxKRHUGALNwSepcYBxATZYIQjZAopLBL0hGh9L0iygA+Abu8yI2VQzPg
QspSlTc7mhYhTeCC769cmQLPqGdldMr5HlgToKI7T3Vf445JQ2dm8YJ8RKSgAQeXueVA9szBchIo
BzVd/kterTjY/o+mYsh8HuIzaOh8QvNzB3BGvRE1u/CpIelo7sxOijN1P2RhCtVNH62HVKD7UidI
eHI4q2ehP381FFxdSXMyTHsu8ldzwmNERw2Ht2zXFAyQNPcSZaK7ljuHoyq5FJ+FmiGRx1xXeB0a
Ce/7TP9vliF1kCD892hI9TNlcNolBAgf2cP5v1h0haXkgwBPWTST0TdVHbJzOFZgQS5V2+SoCpJm
ZIPacsUQ7rdTrdmdzN9tb4RAfRNb4ZkklMtuabCTjSdD7r7Lw0YaOabvsG9/lGkqHVaM2OSYCpDZ
NtG3X6eslOXGlM6+6fb8ufozaCm5Ba6/Sqa/gtJRzEA01PdyXEbbBBTNTWq99LNhHR5+o8jobRtS
fOr2gVSU9CNCDsq2SfAqkp1cobgX/FhgNUgB2SorlxW95+pRrutJgQcMm8WtvocXG5RCq+bpmZwm
NfVUUD7wmvQstX81Hwg1Lgt2DMyY2LVE2N2lv/69mxZQ3trftWQAZxxJj2KQ+4BgAxfx4ijdHeYB
ohsY+V+A/dTe53Pbu2972DL5Zr5ZNR9b35Wv8WJpwDXxk8XRr7mwtj1aMM+F/eI3tSZeYhZccCNf
w3a552FIOFaK3p5V9Etvd3NufNPk09cskshLp+AXxTiFlE3gFd4ISPyc9hdU6GLB0j5njvh9mpG1
Ekw0LEcVU/iiSUF8dV9s33bq0NGyCzMIG0W4nSuh/DF2yQxZPti81mURnaOJm8tkOOre2s5pCzjD
CEjihvhSRwxV0FJmC78xXHqDpKpLRtWid0z1ZyjwmoHnSVeEcvXB/tErCMKVeck6P8DMxOPUnp11
N7eyx/kkilIGbvxsIMZoY+i4aSZkEKeqLAUoZ9SKiu78n5JzQWjISX9/Yu7A0pM/G8VSIMt5ldGg
frIjdsd9dajP4OGmEoGbLQfyPhf12fBjCt3Ynw2t3z4/I4sXdxsBohJXQQGuXbrmX18YmGwLNG+m
skrFrffdmd5pCcLZBaZ6Yx6usfgQqBAjMmLYjOLy4OeeBR6QlAZR71znlLXCRM36KpGVAHv+HMXV
bWHIbgJx5uI/8sMR4L+vrjeJD88EhTc1vF66IKcYfjXgTyY6uPKZNYnQgSD9jDJ4RH2sKhmMke9w
lB9LYdWtRIHKbk8WFdtr+JCkT+kd8kmkM8ynzx7bq3hthJ5UDFsByfd8yGf8LZKlCDVfh+jaLndw
cfiiF2A2G7b+J49/p9eWJKqC8gIV7v0fOdp6cXWoZES9uyH9UdcAUEglNhwdHMWvpxk36yrRAFoM
RyX4NT744NIiUkezdT/t2eTB+13Siro4p7cFJE76Iq6pNE3Yb4WeeLPq541vlNXlpPIq7hv86czR
djtCoQ64FGjCH0FerZYk1FDL4CRmV8UJXmNZv2p6AJA93TJAdffYBwLWqUSULWzRNLLsULiOie39
sjGUiRq/2z+MLl3vTg23Txg+kNX0j36P7UakzdGqMJxkh8dQ3x6Mle6LeWQryXoGCfwLXWQp+LEC
tjjjeS822L8HVwyDUSg/DQyXHM1piUFBrRT01q2RLSeuuqvHthLDauBtF7sgP4/B7WSs6jsc/FXP
lKPX1/BJDK4IErcV6Br+86XJRmhGSoOS0Lsr42oHK47TRoOOkaT8MbsEmhZCNBRcuGfMfHVkOqOm
8C8DOQFCSwGddxb/XYhMfF5g5nKsnm096MSJYAgjvNMcrxSOAP+sGnptU3+bU+pn8jInpSn7k5tD
mbE9aH2s5tJs+j32JwAnnq6O5MQAF/Bets8vuOKLRg/fM1G4kte2eAYjMxXsbSWp3Vt0HmglRjHT
jch3xFBXoLHuGcrOM2rYtLZ451AkBOjQnN2xyx/T9CXucXBGMWxbBegzjBU1KWCX/ONjBoWkkVi5
l4G7wKtnTtBC1Nek/CloHrxRoPO9BFYG0FEG/qmofCEEjHUQci4gFz54DLlCBkQ+66lq92McvO3t
tdr6goglRGZxy7111NpiXXNBpKQzurKR/vFBhqUJdKL/BHBOnEucnUqkvKe4mHQ5VTHmT1eG6hk1
Q99GDw47QxHJ68NZWhiDsjUouECPwPbRR41IYNDjAsIY3WkNX+XleXjcKseMfPDzVDeotDpx4fH8
AcGTCWNX2shDQkJaQKzIwbX1NJm2OsyT4su1SvdMkOKX75KeqA9dgqesmYBcvliSHDXvTbOssGKf
O59kYYF1BI9rRjaxMGHvrvgSYwyE7+fgsC6Apdi/Lhg/vlufEL3Xyaveb+H7EKxLCqFEBv8/yMaU
qxXYIY+moQMwC/Kg6dzieNYyyngZtW1lvaYVgtY1Byh5JV+0at1GNrZPv1fvH0wGTPWmqNmPJc9W
A1lLU39EisPieIYuQGZ/m9kbYs+VcuLdkj6jqKsbY4JgTGU9rYzGjh/Urv6n9cNyXgGWUAkYotNI
HO9jcC9jAiztOUbBcQHPF7HFjQtArtAgtAy/qNMRuXd08eXjmjMB7e1aSYhbDMRBOjfzWHMa6BTK
SmDgKizNkZMAn6DaPV+li50MDMXLZ1IpS/nTEs/CzPxUS07b4TnoNQGNJptp8V8sqjU7vzNgpca7
b+nlxaGY3UvGm4IpkG7+FM0TuM5p/PM6bfe6pyVWmHBQLloUsP6oRMRP2gc2LpB9qo3wnINpagjU
YgX84KfFxhiDLQX4YsIBaDs8Q/c8G9k+w00HgOm4nyYPPHSIgjMZaqYZ1t6iVAbQzSipX7XWFrxM
hnlw5RgvwGTKhXTjUYJaj+ndi4B9uXah68OLbWrrBzW1CVPR9QppTXR84xx9iZl3m0Yl2JP3qcDG
RGcVz7H7S7i/z1j1TZ/28K/tNm/FQRr1gRRZuClm4JbnnC43uVH7E0mpeJiSdPVKRYthXUumdJ28
u0aM3snhwHfhp0aeP3pGSqFvR0NE9aRPGyrcgIpK3zu/vul/k3QyvnXP3yQRy/YzSP8A5NjnjYee
FUOwM5sIUXyT3lN8YGu8oDAERC4xaqm8VMNDehH7ss54uILFAlbeTxznxU0tcHDyNTl87MUrosom
FEFoSDn/8s/cNl2E2FuXhjAt4xic6fTVJZ7363KQgiKa5MUr7v4B6cERW/SkcNe+1N3qq7VeqoPw
upVbiKyMD7s/YexNsgzYm1E6X7LnTA5vderseFNz1zC3vXkwDLbQIvLnZ1Sgq+gcfgNEt9bV5Ugi
BGhVxun/1rn7jIbWo9phIM8IUv/QxSbE9wqsidTeLBF3WBLJqtgngyPPNTWSBC226posKOUav327
uJ1dDeNLIb/sxDA4H2dqzZIYCr+IGdeY8WTdkj7y3su7qejM7lJjCy9Svss1BidTCW1rTq5CrUA2
oaPyj325yxYkBXDPzE7DsfOjz/7wiXGJWscMrXJC+VNuaPqOA1flBS6kZDM2J42CC4cGFPeqqX0P
0atuXMDUezohm1XGN3BVSq38Zp3d4glHTNMirZNgPT9F4zHp4TOjWbRsNFASCbOotDlJiPVFpRIS
FQg28VZJ1Xtzu5/lZHolvyTOcrw4YLQrrV5Gz5E5J0gnLwDMst++A0hpZVrV71XdbGDDYjVY4hwX
Ri9DgT8nlswWVKLQB/02nwiyfeMC20PfUA9fm41oRX6CaubC61jG0Wygy9woxtfVuEaq885DZNV8
O3EhyOy3TLO6ajafT5WVVqzJ49IG+71kgc5NFALXYsChZij6opiwlhTCSgCEcKEwrQ9/tAcMnk8/
voesTxfb1NImDpBjsvk2XK5VmSMSHeBbhl5Sg+HjdoZ+Tl7ufWZY7fUeNxCTE91DDwucRgjkhJyB
VAIMmNPbdqegOiOf6rU5ARx0cNv3e0wUD0ZZYYt7ZNxm5ULKFvDE4m/TvpbFuGBRSiBmKvlNROTV
mw0cP7HI684hjiXoWNh1PWGoB3hJpFbR2vJRQjFDdw95KoIm2aoL9612bcxlJPY2LYerr8Ab6ykH
V3wu1a0uvaqUmXw0kCtOEXNQwoMoY/fnlwPZZUC1EzXWbfr+bBm3W0dXIWODA0Gbp8v6xqJTARG4
Y5MVBZ3Na/UyHo8vvSwFQX3ocnWKwmFCYBMjhGbJjdDAfxoODU/z9iZo14i40TF0kTwCW7r4BQuB
nq9+hDD7OjA+AL3lb8/vbqxhAFinLZYFmpEX+5TsLhYfy4clYSPcsDbMV0wG0BcT9UsDWxFtTw8f
DNtSoj085cIIZtfzCMK05CpgvGYkBM+Al+aEm8yDOlSARryU//G4dbTGU9rx/fFiBs7Puf0GjLzV
4CNdBzeWBSimORFh3qzxse2npLb8fQh/8hup4TwOxpPOqhk6epjy8wcwQ1KkANJqoxzXKore3Sfm
YnjiKjf6n3/L5O2mzGPqJrSEiY6udzxAKKI36rUgWk+8BRiBqu19ebpDQMmG8nXvcPPALMU5ggcz
9KOuu0G7kjhjlIGYGkk6JdvUTHjQwd+ixITDOPNGns+EM558GnJcy9MSPT6EPFaNUPdp29UvY2lu
ZNimFRnRE7sqwmhe3JQTIXu1Z8gljgTwqqLZ5y+5unvLoIaf+OoiY4+xkU8W1xnBAp46F3yKVXHU
swRIKQV+tk/sJVxWBHUI/zONFv6K31wEmJ6W/IeEhACCrtClEWLWYTTtDGOB9FojdxOQVqdjUXbe
5+xMGqfkyVAbKOUx0GK1AFHHDHBKo4oI9J6T3NTArmKE9UrNwyczwkwHuS5eFzp/4zAMVhF/l4g9
t4G33pT9ZquR6N3YvouZARLD6rJ4Be54FT/AXRs4ySlq8P6pY+upKelb2zQaPsutO+v7j+OJHXGU
9XegNz/fq0enSe8wWF0hKKpGiGBpoIMOEGxQJE+sFZrovQ8IkrxhxVzNXx2UP8FFPa9n+EOFY54A
93hv/4fG8fJ1sFbUTzpd5w7wWlHFMtD6WXxIAx5WryN6aRhgFY1udDvrLLfzNXZtmHG/8IPUErF0
6BBpfVp8Ikoi40HX4u1izC54XbYyNkLvkz9zks0FYe6OTnTE4VQjRM0D3BWnb35UMuSK8WtaGf7a
KfQDf36uRhbaADQhFfLUHAaPplif3NuiUQx3msfwZMwfDgo7j790W1zCNCKIoIEIXsHBQj2J1PAH
C5xdW+PKLg+N1KYJPIKy9eGxqJ2c+rY/rKlWeSPqLRnmbVOlrrd0IyFp+QFZU0yxlgZ1uuik55yw
S8zVJJwUOpQIp7ya96argqeMtKxw1AvinQp4vvY9xPl+OZWecPmYZ2oraBqeJ869LGoG7i3mLE6r
uzeDMLcdhISEq4YTsqlZRXgyovQ8Y6y2eBaj0DioeS691/IB0RU8gsN7NYQ8eaBSO0GTWxY6Exdx
xCxWIfvYXc4XLAc/W3U44bckULGv86gYoiw0g65lMHNAi0Km2DljiHBr63rOZvKscsav/drAHBBh
obYHRGKrfw0n4s2Sbz+TSmeGbavR4bW4qAKocIhh39aqViCeHj803UQNgsFzS98fHUh2YsuCEK6o
SNsRJAnRxplkHRG2zzekA+ROFO5mHJSuFVEaTCqq45iC2KS9NEkzCZJtz3yxC98SlJifLKK3hw7V
lUrMUlzCXiye/EsjF7BpX9aTbo/silvWwhjz3m3dDKGIX8IQHtkMA/bIbwhgsf2KkZKLyhwZMyhK
RF85L8SaxYDm8VusnyiyhwdcCbqQjX+VAz6FSn5KlZ2Ynhy0elg6ZU01IrGnQfRh7DbnZ4aRjdmF
kQdHr3LZXBdqSPsR/AhpPxjYh3EF+SR7buvvhPm9hZI81DfFLGxFyAnHF5tOL6QFgFN4Ptl1TL2/
uID/uCW2pXh437XWyjLkV5Ct9Yp/1YjKl/D30UVTCagAVtxIrRckKDRu1seF1pixVky0VIFP3+2Y
cQOOBvL6pjV0O1NGvKuYfoAV2zbJy6Yp+rEG2d61jQfKQw3RzdQi/ROKWhzJcRi93rH6P98KmaWp
3T6XhhLc6yV6V+QBMS/2gI+AR6EGtMdivJG376FooeZpxej+66dza7JhysocJysE2HRQD3UotRGC
FU16L9ib5/uA0NaYaSEJ7GMsFadexgHcOoCIN22RG1ZO5PkWg2nwz/FU3jWhk0rXhoNB/bbfZpMk
fJOhSqG08k/0ENTEdAOV0yuc9srCZ4obaWOAaogkpabffmdKZRByjQzKXMTeHxRYSkQ9g165l81M
CwGXALGeSFhRvZz9J+GDx3l25zbbhIIecc15NjBLY85iFaeZKIw4S89O639UuiQrHrikj8dn5nfA
3MN7rlFgnufEaCkws45aYrg0TX4aGc2ZBobDUNWzjM7K72kN0ku5fehCUhiAYG5Q2DHzVB4D7E3U
mfcy5lEv73+P7r6g3lR9VNHZe6W1+2n9uEDMNmnt4VQfKoGFrn6QVcQw8oj972gUdab5MyHbtjZ4
3kidMbMOg/Ub3cg1uN/VTNx1CZQee3cDu5prKirDdY7ie4zNY81IdF8h9c6/+BDVxUUj3V0HMH/w
Yqd0orpMPowR97Xq9drFzwH0yyXLdHmetuzGCNFebFKCfZGiCVWTVn1dIGm+NeJe94PNd9EDA7zw
i1YYfLICUyVmD34L7wkduf58zl67Z61xYd7Cf5UKf4ePmEp69CZoc324LBsZ3+kklmJ1VT5bFJu/
MR395dK+UEqklrPe+72nR8SEMn5RRKoilD/dtlZYsM2LpsBHKN80US4M/QNW9KoXbUzABJumTtSN
GushTsY1jtnTfgMgqWuc0TIofSKecbnyIrWg52HIi0PgImHM+bS2cshJXSyxHmiXpCpTm/J8v50K
TXSDJEHZafVQP6RadFfvHvpzNjO8Lxsv6EEzeI4U9ej/krhsr4GK35UYI+cHrn6ixRt/Tp6ieVxc
irG15rnVxzG26ygTrK1kQLLOXhyXTTGiqTdoxkoVtG8MgouZ/8vDslYxPzDbAZ04bR5/XXwggbGZ
8zY4qMM+HahADjfmXdKh7yb/0IB8v7oNt4NFlUQYdpojF4ui4asjM6/32Cz6QSJ/TIhXxehL7V/y
7oIBTV1qniIOgyT5L2LqUAELx1mh3jiSrGrK14oR6e6afGpRqAVsjW7qRbEF760NLBtD0dgppatR
41QzzwxMrXnUAhdnm0rEMtNo2spEU2i5AQ3blVH2usZPqcbQgW1mJ8UIj4r3NWJFfSfdSzecJKZb
TUjD0cGJ17w7NLN/133q4P6qpBtsxkQQbQIkZsOIIMxqh+qEq+Y1lUiHIv69TG4dlvagwsazKTvi
9UukMlOu8qwQhZoG/5lVGbB1nVafQkmqq+YdxIv/jdlisoGJXsKwwT9zu//ShGDDrFfvQCJKjr2p
XLp4HDexiRoyNKxVhJFrwhpepCbCDMb5qjT8nUO4wRHPMmxCXIqlQiE1Ag+/8c5yLY31AUvR31bp
k0ObbVsyVsrNxOjmB6PbRS3d10JfMl545cV/0fARHQojnrSdtqMh0V19m1LtGN9p2TdEO0CXRSZC
PHLTtft1N2vjECnoxzcxZrVaTI6XzTRvgZkg+oc5HfPV8pZizx3KimkN4gVrpo0zeQtal19QEI5Q
lrzljPMqDfR8oEe2qAjHU9oQSsrzryMDnFdog5WPamCXJkLS3EkJb+pEMuc5MPitZ6nK4SFyTKy8
9iCAAL8WexokKdm+Z0OsjhK35JzhldXJov7RPM+RaTmP5+Mi06Ay8zEMtNXA/pYx4b7mdmYmmJ4x
uc0cevSxvXoiHAoLnORDoLOKM4/u6WnClXZClyTHFaFH700XL4+NmuwZneiL0dfCLn+WXvKmJLXx
YXcdRaR28mXWx/2wJ/Pajvv0QFbdxrf9MYhQOThXraLYdZdXPIvG17S54jQuELHXDIVobqvaL/q/
R5iFsb3XOdq+8waedEsbeEE0IHMXz21hJSzROkV7MNGcfcA/bEDlHsQ55sNlm3naOtX1e8zQ1cEw
Tv5ToiBHYJe3FhPCfUB+glR6TGZ0BF1CbBP2+NDtb2jdTqV2LBOZT0oVevzx9Ej4bqu5WtITp67M
DAU8OMKr3fdl00JPGkRAb22hmqC5+qiDPMlZOdUzkeUvT1069/s3RyYnbjJgME17iihtua7WOaKd
2kzcNHEEHGF/cb1PUdpK8tkL1h3ThC9mKw/7WK3A/cNzQ+tc/kjaxb6bz3MVvKwIRjg1HoOZWnuv
NNn5T4ZNXlEO33g2OlnsZGH6qeR4YJbRqZYnwisHJyhlsjpOBFFSVXLKSYEC8apevxD5kRqFo5Oj
peLkg/SO2uCAl1tHy8j0mJPcPrdsI74BvRsVd9k0nf0JjGWacAUyENzENbNCdJKzC3mar1mPkrTv
Y+FyPQyHTKR1Pwbfk3hue/JMinyr2LdP796reffxVB/Bi/T91r/zXyvHI9y7Zz6mjRpk5pSMLhDS
08sa7iQ1R6sVkj9Xi8UzAyZ80VgyHuY+NhM+h9nCI8+61makg+ySsquZDqZtbX3ivmxw77jvYh7S
u2kK14Vk0FI0u6GNXfU97CjZo+pSewBWiXQaofk32cz7GLPFHfI5d5/5SqrPV0SLs1sGYJw50H1k
UzN8NSFItTSN8qRYAZtOT8yb3KZsUn0emdv5CGppmcZwiLNUHWvYJfcs6wXPofdxBVKa/40IJIrQ
ZKkdazv1peev5jfx//WBEtgqoUkmiluUqGREiwaONWztzQrpjv/b0mzQjGpBFN5Wsj4icz/LVvaU
AHfSIC0XqkwyqCspKYFX2z/btTFEvxCPMGz2WdWGIiQiBqfaG8K3UZ+SDI2PayLrwWmEepcxDwA+
BgNNi/EVHiKFee5cVHootYkFQJkotRkBmz9ZdjmpXFNBXIbtOf5f1tzRa2TjWYlKmd7O+/+6hzEQ
E59mQT0zxniU1lDRNwjr/jYpWady5Ah4WYwKLMKcKfLK2sgrsYskDKI6VdXRNnlY9nuwytrsI/Rp
fxG+P/Lb0OgNAyZRK1OdAq/9UPf6Q8hXgwvVFytvXvsIzeAL06MFyIaOsC5uM59djOZpsTTVNIDh
UaBqBqwTTkCdpgDnB69sXlX8uxLqxJCaMRtCAqCqAOEPWNMLpW6AP+9/jWUcbADeD4gH3UEGyser
aiyW6vuafYSkwfRAGMEM17Fz0qwCMvp7swWBmxo8PqZFUUYpGQD7xriCb9dr7zmTVAtf3nvUdLQs
O4OX+GbVNPUabFwDj/REMdRkP5lEXid2gPxJ1e/op2et59RP1LjTu82XyEWnDJAyLIeOC/ptKbX1
GPOXEsWCrXfUqHc4XXMOvAYi5R1yYN7/HpODcjITnW9LAcL8VuNvY54mCSjKQ7N/OnjrvZIZJbkM
4QJQcJ0A1pybYrwDEhvg+GkqqM3ryHjQUh9vZ58cfOJnImx75GDyvbbj+uft0ambPxs0yoqpls41
W6YdQEK9yNNJg+VKVggpuPqvSfQ9EYTdr6snnAKZpko0NmeJX3JqmS3Aeq3HngpPTo3+opHpbipm
VOAW3mex9PKf8YsSHOFVRLP51oUaM3OW6loCGMeONm9hkyXQhrUfzjZSPpM+GTPPHNU6OqsK6diz
OqsyV1j+kB5LPSlfrW3BvNTc4ctt7SJlUumqNPoCok1kCpyqV8ZhrMPEXuGuIdTf2Qf1uU079/tq
Kr9WRyKHlGfFEDqMc0FT0hVUWFGRhpNX9AurfxRWKejXrOwlKrMdunCq8gQq/g6PEMv3t/2aiiVW
E5pXvPNg/okP9EDmtFVtUe0RT3v6iAaib58dum5Jfw/IdVMlRf5rE+rzg93Pr58EfE8246KR78QC
FU173RfYCB0MvPzmR4xaI7P6T9uEMF/0PXKAPy74GtYDpl2XuOoMrJ/r66AAPHTjehpRFrMKCwz0
v8aTuMCnGp0xUmOcCijPtkX4oCr7VDl5r9qseZ9NYNqNRpPcKKm2vX+9p74rTMjaa0mei6XXKkiL
sBsBSkIdwzwz92xBnqBXUPIfZD3Q7inXCMtuTTfkqJM6dfh7gZL2w8KNxFTdWBcCYqyBzkWZkhPv
B1684z8zOnv83AVtEN6qkwfxYJbMGluv6/sOx205Aam9lSAv9aXaSDX1CmGN9hOjtp9K0zggjSAX
zdUS44K1etxUGdgXFt2SCPN3goNoiAQKfp8lQ68mv82c/Bitj9L2c0W/M2Ht90eslTdarazAgFzS
nKcVVscwz7CZFCVo4Yxi7jFrNEWt32BdlKtlBTU8Gs0CXeVXHMmw+fWcqQNqlbd9BH2tjDogDdAE
qEWakUH4iUoNY0hIOHxu6T/HK4VTOcHqunFpoKbMzjjFq1GnqJoQ6xjaD6KEIePVJ7CJqO0YYEWr
jux3/0H81Oj9xwxKcaGNCeKbOc2AdxQnJcxslNkeinj9Ge7ZLYt0rpwZJJJY4oqgdEZr2yZmfzjp
57uWLAkDVGcYXcXSKxV0kwLrJz+9hRV4jOo0r4bm+mta+csl83HTYOFJzeX/DniFB52+WsE6+pAj
MZNjVEfUPBuRuS5Kemzuf/BsVXsKMH/q8GBc/hxMs/VtopWITBZ8m6rZ0FR6zcjSUQLxytUODvhM
E1NG/1ZM08/9bcbLUrtYvXIlH0vQVEGDVxTM5MOAgOczJNUaZSS02GguLhjnKnDwbZM4vlqj+h5l
MlNmdU6w+BiDSpChuxi0Yn5XwPmrhOQytEuwQ2M3JOCkMc7PCQggeOcaloC3v+fF8ykS4Cpz4/Wa
fyeTZOUE7M6XXdsmf3tFkX1i2hvDA6NrzStomeNWog/+3qqM8QwsNA1kZKSzAmh0VbpJooc3W7x5
VmHJbf6BxCZOHGWqrp1YZHiGvTlkDWSK3xUgREG7n9rRG+KHh0Xdyx5ttqask9MZyyT5oiIpGh6O
Gv6DmS86lkHA0bmfcDwYKYV40UeyUOT8HHjU6h9/hv8LgPN1ZVSO9zegnaX4SVoyBRLaKpsY8oKr
eNtpSkR+z+4KTeenmfEO14L4Z7h8QwA/lU2ZbC4ATQoNglM95DYNLhh3ETxTZNN5LbUw02uqakn5
c+fPEAl2eAqXjQDO5I9dv76//mfYeIBDrY9S63anP5kIJDAND5FecCIguBbPy2QUMwiM/KIydETd
cf0ce5SVeoIqJw7JYyzBtYNuOsvo1jcZhrhbnPFrMifXL3aprZMHvQwZWOT7MDJQAVNt+JYDQBJr
HRJl83M8J6d9e9gFsEswGugMeex00wNG3IYtKIzTMezBRooIgvZkTDjby3zkPvxVSH0XBCDZUNmO
ry7gf2mbBHbeloGKfuQW4EtnnGUKkjDXmymZqDqrP/e7GYuyCuH/Jen5vdqPyIzGvwcIc7SltqYC
RvSs0jHzfCOi0ZCQgstR80mwDyLUxbhr5GnSpAoqde5EshiTCPan1ISroCBgzbXq4oY9ToDDBt07
WX3H/zmCINvNEuQhnO2TU1mwZOkhUD5dWSSZK/Wc0AWa2OEFb7vb0y32mhNNMvu2zUzzolDGfD14
bS0mSJua4bVoJONZDuepI8VIAcpsxWOhrj99jB9g31JmNjNbhVDp4c0tXtszoURKvA3zAx5wXzzz
uyrzDOdFWXXWIIt0tc1ejr9aj5n0XdN185jWM01g9/GxOxZu3YQYFefOBcRUBbORNyoHaADXuU1/
x5TD2TL3hoRenqQO5tJuRH1KzU7mylQLz1B0sx7uD+OqkwsCosC2xehX/f/EFY044Gw8jCQJZTUW
FHUFxwUKcUnDD9lQSsPlYgJBQMNgVCrSOgee+caPNyb1vVJaqwCKI7BZEyCXBJT2fT9+53uTnPst
i+915FkfBMYCVndHt6VwxZTjiN2UVWHHQvD9xNOjrV5IZKz62Bi749KdZElo5AiGCjOI7kSgE9gh
/6r/KLk+p/bqUEz0JMBhM9lTK0vhkE0kZIL4/NuMvQwPIJ9q5N5ttAHjGlZN+RHYXvBCYVJNjTyK
mODDYrhr/vx5hYZew+iyULn1gRifEVDjn9odeNELOR52vzWLIWq5V827T9YPaMxO4oR66guADV4h
KO92V9K4lRvArSTKH6yKkssjh6pD6S3BvSHcYYvvYs/LQ94C/jut7qEGzxQvNCYcs3+GtmjNHIBT
JsIHNMCHUOlSW66kQOOJifozUFuhMgrxrLNRmUoHCXEIzijHrYazE7A9gUS5rG9BChqYkQP12mCx
Mj0VKG3WFvompAJayVOLG7XtSq5XRK4/M7is5a/LgddwTKshGvCs7HhCnObGZZy6Vu3HP8JEkFke
1isIzi0mZCAl7zb7RoJ1W920a81sxl8JG89b3xVKSZqaODE9s24nY1lb1TAbkaNUj123qhIjVpEn
0fXH7cMPZXkp04lddN9XxgbWCdgMTZc8VIIBMkMlSpLLpBkt5o7A95v13HLHWYB8M6aH0+VODkiG
1qATlw6LJ4YVAlfsMk3FX4VE/SDqvPynwMrYuWdVGDVk8AviC15Z4kVHmwkYMB6N7gb++ABQZuRb
Sod5uvtnEdJcS72yRBuuMWcns+sFEe3dWMEaX3jk8MBom9PaWF5tDcwiaqPaF8rf/YgWharfwM5u
6EvIfzJY63q0b/EUenFsz2DtnvI4JW5qYMtiGL+b0JZyxWkAXYDMlULQ60T+2GzLMN6Os/qRv+NX
ZXwNqqHXn9n4BAZOujmcs1f5wJ5bJTy6HtvLfZevD1JoCoBuKYun9+QtVWjYThG06/qCo31XOndC
qbeV1zrRlKQFeWr23oDncWVTU/a/jOD9oMD8FOg/+ITlEWFe3B+6jWDfAFBpNSKPiO2Vh3uN8wN+
4Xi8hVEjnFx0WLv8cXvpTjhoJsZhdUruHvKJL3UonuWKtrduHUHCKwpcG+5QsEDC3qX3THa4kUm/
r7oYypUNwUKsL5+6Oc+bckWaCZcjdaf098enXLT3m8dv6dDKIOCWeEXahvxFxS3hWOlxc3kd25h9
kjRQB6IPtaam48nt07OS6rgap59clQ6fyKpBZ1kAdwY5fMBJ5HbFH7LzHJ5lPQsZtyeHFl+2LSfv
DVr0UYa5yLVqfT/k9QkmcbwpDAT89JNg/4bxmZ+JOMCsRoFmsvKm7rFWc4bpdwSgOOPvNo60WWss
pxg5V2Yzxe1FVJ09BIEtfdnoLyCvFIqsAc5r8kUy7gymrydnjL+wSpRbk0wRDwMvx2RjJypacCp0
KpGuSk6gJhtYHUw1iu6t7/XHiHwSY3Oiz+PXW1/TgiCq78KltOzMvnjA6BYjs1FqTQK/QGqX37q1
bcBUYGK04YeFYUEA613V4Qa5syvh7RSosaCUZcVNHbskVfWhbdlM4sE5yfznt19qj/xxfSRcftp8
Ex9FrvdQEN38xNLqzqw1JG/8ZudSzH7jEUAlngYtr0y9RzYXgUIHuYueAgojTC5oCjga2Hs5kYMM
Q+HWUpm3K1d0zLZDVlW0eM/MAZH4r6at+ZKkq15OwsYawo7EqFgn4QQ9ii4r2aSgcK9NuSXj7BJU
sYQXd5Q48V5tYkNRTEu9TRsACd5ap59VyQH0RG6o0E67zzn7sQMNVHwCa9Y4BNJVqR8FPBjuv0tZ
agwufttDZsfhpfdVsKD5YZ2P7rgJPB8TVkeNgQagc9eKnvaBPIGnEXyiJPGpSW5qGgtDdNKwaM8F
cVAS0K1XHGOd89r88pnvLzGdnM/5DfIUiTeecbKf5P952SJEJ3jjY4NfZ0h1FqXexGe5ebF2jaBN
kyjpcyxUH7WU25B9fSrh+INhYPTRh+5EvqjzE4ITZHDcSEVTTZEfi+kPLDygKYMWNe3oqfXwHBHu
HJQjKPRAGkVFwCeBhdEsEHXaHIEEmGFGzNO51IEdBD4bW06MXui8lNro+39XrKUNXZEVTGObvICP
nxWMvb8VlvZhb7k8Vgjn76VsVe2PPtUJje206lSIVeCv6meFPOokln2uTKo+hR1bkA1M19tdT4DE
BLxAmSImNiA/tosHsWwOYLRNmgIPjksmz2cMpq/PXqruxATc0bbqxU3A/0CTXCjr2Zziru3NKJHa
H1Vtni/hhrw+TOu3x+37iW1m4haZuUiz15iYG3UE1n4fFKgfVYUP8zE0tc/uw9PxV0bsOXX7xAvW
xuxGJomTtA++AVJNCFPXtU+rBn/HBr8GVU9KhufqoWtm+xO524J0sfzb57wLsGvOkPv+zG+Z2aSQ
8+5liG2+PNLXTjfuN7+hWHaiM9uBP+ZyHGkLlyVmpovNzJMvfWifua9bUunz3a1VzH6nYK7sU9mI
EsMii7w81ZHsTl/LeQG/gbYt/sD/kKIWIduJV5quwJ0QbDSPQVORVrPOUrJILul5DeVKd0mxau7o
u1x5KwmDBXGDB6smlOk+YHoWwACeTk4rAPobwMjbJO/T0HRw6HhJfxcSW0y17HqdIi1ZZZQo1sVy
WT2XZHd5EiLUnzNzScct3iAzbMVMjRlXEzPUvMcqVCC+Z7jJS6fHA72KbbzfW9tuhHJmoKg4Eoi0
D62kIkmmDwixnPK2oI9ZfXEV1RIZzKg9lZx1OExeHngt7N1oAmTNKweUH8Ci0QSBeE4Q+9dPk3ry
pPjzSQRktz7MjgnddPB/4EVgjUXKztvopm6QP0PXXKL+TfUoPAmHpm6Nnvyx7KGF1Iu0DG0jx8sT
b53MrJ6d0AMUKkgQDxvAO1ugEha0bWfiRz5/uks3cGDOhdRZenlnTEffIHS1pBlTCnPSMNPbvuXh
1DDMa94nMKElf3lNJ1kjzVDZaDLtdE954BJNyoSbmMnMAqBKGIlvQj/76JeZ45V3gtwamON2yBy0
XfUubYo4K1igUN9KO392a6yHm/O15907zxEZNmBBgId6NdvBNXJbPq+d7HIvx8eQ3Pwl2tT2sq+g
VESCnquBsDaGr0uyj13tF7+Ilc/JlmjIYK4F0ydj3jUIAHa1Dz4ldhIES5RaVHBpswP93w15gsr0
pgAmMg7haYA4BZ3gHgIr8wrXpDoCs3VhYmONhynisJYOjO5YnJkInChqKYDaoNs1clsGLhBkOXsZ
B0c4QSFlgXdkkDrua40O2C+00k6RSQBCQlYAIrj7yUXRJQFTGQFKki6Ce7QeIvTCGhzGd6vLmn5S
wlHMGN36wsU17lmyf31zS/zP01uwGCH7etZaY+JQc31pwQa9sW9pe9Ooi6uqQR+S1zNK8qR0yldt
FiczZ8UVQvybnXjxbt+hWj6bjtqpjOtzT23BNS/OPocXn4YbQWcrhDSP3c3FIh0f4am35PxIsXm6
Bh6CbyVZb9y7lHRlJUAom0F76Ukcwl0qCFslqLhZ2LQDUplr4TtguiTryVkNXfnwNaNVYzCF8I0X
L7XwSO0463gwNCGLOflx5YmlvpVUvKeaLXkUkBA8btT9JW/nAfQhYOiHm4qwPVbdBfgEah7gfCbi
ZIQSYJTJjVWXiDSupEErnNrr7BytpiJmqUh5mmT7h9exLZh02aklW2YOq3u+5HvjLKjJvzZxF1WW
6it1Uv0O6JMoTalp8pWYrXpTD2SxEOqVLVwKDy2zAj3B57XzcBgFtN2QdI6YYgRlmNrJapCo5Rdy
PKodVSgMjOCvDI3S4oF3tnp5dmwc2StDfxu5CoUQKOzF2M1As48sSUf0kYhzScTSlF9M2hHIEerE
P+QyeJJ4JY2kFaFF+RgzmNQ7jfP4ahK/SVI1gyehyssk4WNZFJRWc1efxSHKiI14riHas1XbAVOL
iMZeMpgKfNpjQibRp++j9NMdZrPnXpmASl8n9k4hsbzTTbmTHly1E2pAPoGgXQRYdEuMoHLzMR4r
ZdlK9LrIVcFcGwJiJhL/iZxNawu6TZnLNBTbXwjIbnoWGbzpoemAAezMaZtnxqDExx24ULmqlWP4
TDg/D75K0e+aI+EWJnI/FaS15tBATDT5lCnQhiP+tGv7enZ/SWRfxheYdIcd8z2lu/LsFuB5/Xno
ZjbuTHq495qq/9tDEq/sFe5Q22AJz6geFxyiGqVGPKAJ+q9Lbb3YKezUfXwezvQ0gPza02ubLlHa
OjXEbPrSU3egFI/DpnCPpqDEKjBiq8Rc3zbIBo/F+6EIe7s9Tt6wmbRXu8Yh+wv0EdCCR8nsvX8n
04qHUpCRhGaYcN1ULxYp0JjyQ8zLv4SDXBnLfYC0G2LyQL9GDUaNnC2ihUjPiw4TbHn81oJ1LiPm
8En+xgVaM7PGl8CXF6+1vE2IAX/Q5lnKoAmVZctWverzOKy2YExlRbMXND9B0pa6f3HNJyEbd4kY
KySVVpEQoIu7rS71XbN9R6/IXnzqDhVF2MEbpke74aMKIhOPzw911Kv+vjWzjx5szfvhTyvuLxXi
T85nwxvbSoDZbZT/hVBR8OAyS5Mu7PYsW3Kes0hQpJyAt6tG880beRf37h73jzh0WI4KAtp/jpPB
1zAyHQyerH1PBLopMr6jVzMxbDCRqqZGQIiH02CHGD2qnZL1sS4NtHdVkECfP0qe6QL4nYR/ljAx
Qaz0m6/cAOBaaKPgWAyIdm2cCal0FWD32td48w0Cwo/vw4QCbtpn6GmKF7xXJuFc/jxzKxrYLHgo
pFQ8mXA3Arkq664zCnXjTMtAwt9vyCWROKHRLH1m/ziUu3gRdJRlLTImbWTswNAnAtZSEMDFRbII
bxYYWU3DaoQH+p9ObPe0L4MYpkdrlv32/bgymZ6xPn5AY1krQ4ROGlNY2Vu44D/8GAfbvOBou75z
98Yku75Q+F33gX2Og1w47fePi3hxXKVOnHKgeoUDv1lCsyM7/W6NcKnmeru6LQPXmQpmVx3simSq
VmBcw72qqyCDGHw0EpNQNwIHWtUtk+DDiDEtVTFk9AN4ZGuoADMIdJ/EoNGhfPUuq4KXD5C9Yrpb
JkBSMFzKhKPyNx4r75O3OtWdNhh+UoyxBD6nJ+FBM9+lXkFrvNY9dBQepV20j9gEuO90jmzynRd4
ycpKoH06b21rkWaExYArQUikx4AMhvu+4G3GnH4lUrYnfXh7wqIQeuNy+RS4gslbIyQONn0o9f7t
TEJO/21BKhec0QSbOWzqYqDDsX5H7MwcBH45yWZn971RuIz8+iyKWeBWWc4v6FPBqybJLi6E2Jrg
XdbkkxrkE03NeYCioNLQYJiCuBseBguIa4Q7kdFZGPlTnbevylw1qdNQ+oiEDqmwMOUYwVydmpYy
egHpIG1W+D3eV0IuSMHgEV0J48WkRnZGnftyiNeV6b/x2kUGl1AE5dxkZNu1SBciv7so3y9whCwN
fdEcpaOGfBf9Ys4ODPx0Sp0kPxTpnmYD3/zSm/B47M+aUChQwctHAuSPpL8OyI9LZqQmKCvVFhUB
7UCdHUtWxmuSOmpQGoyy6frgyGr+h4+Yy5XsPcMQU0YfH7p8x0Ev5ph+FER2Nlf5dVyurGnA2OYl
BZ0NiQwY7g70NdFAaEbN9PYH5rTIAqwz6lEBIDcj23/hmRUhFxzvZGYD0RjvHFlNyaO4xRWb8ap2
fNDfphbkrKfRul847/JtJmaHoDdYAOVtU2bhm+F9sP5r8gL363059JF2SfnCiyIOIvfsG1vVhJux
zSPZ57cI54KYKaDHOtlrqLxVebVYA7N8ezKey4pdD5SpPon4YwMUgWGICMNIyoFBuVhToYFHHgjX
1B+H30LCjfAhl0tWtxQh1VrCfhFq4gQaU0E8LRl/7c9xJW6r8LbLSm5NUyt2Hg7T1hO7lpIG6O2R
PWHYzChzBRBxqJ3GjLz29HEp9y4LDMMH0nVPGInUGtLswXDmSl3U+Oi5o92fHATRLZzKU6rf7/Ub
JtZ7qCuYF2v7GBxbZHgYfbFc8k7WqJbBO+h+uFcQoTaRDlDNkMNSIWYHRrPCwCepEx79UWcKtNN2
meEiwlPXPV6yOPGK2uyeKXvWX5qU3++s6aEVaE7vFESTMuc9hYEz9n+VB/lPdTVjAw5Og57FI8ba
2u5JKrY2wzuMZmZxGalNcLmLRCBMTPvNxUoTmzr3WICoVgGB4jGYxH3ntjmpUniroRYYC7R9A9Xj
8134buNOZTEhwDWWuYfFSsPBXTi8Jt4DEv0Rw/+qVunuNy/rNYOrojzJYPt6NqF/9Hbhlhf5jUNq
cKLwN35uWMGP+Ucr7AQrah5wB4PMvt0KdXbKoz8adWYuirCiAJKK1V+5/aITudGgfnXScNWLNoAJ
B5hjx/qVZozpi1bpMygmtXSNwruXzFLGYLDBzg+rEPYcug4q2Z/pBET1L5gLVhhh+ciZg3lel72/
F7S2a2EvLblx3w+AYChBkKcTlGYcpNC8IINjuWG+hzDMMoVvR1SYM9c5Rbvfm77SfF+o/1XP9Wot
usjshC8RomY1L93Jk1tyi/3cb9DUDpd/GP6mHHhFim3QaSO+2YUCCoSfKKRo46UnVh/rjI++n34e
TJbsaMkpkHs9qgfgReLFT9Y/gMRVw59mdR0m5cayGY96MvLTcAzVzvDLj450YDL+drPU/5fOSzQp
8oe6/KaUVcrhyXZlReyf3xQvYBBrhaCBqThrkKnd97yrM/8t8jq5/wAwe8vE5wOsfrOuJj4c2eSl
XjTEd+gF2gZDUrFlH6Eb3lS9TJxMaiT3UwMWzddkOZlULJr20cU/8oMnZWJLtTaKWNz4lmsxK3/j
eL3FA2z4pJQ/TCkJJ/86j5GZepx0M9JjHldXvvj5CYcHTyIamec9rVQUZMre6gLJUR74qdbEFlkL
BA79zgXYwy5zcOUjpPTepFChQtux5fd3D6HQ81hgT2Eye1hg5MQKPIY/pNuzJw1vV5Waksy5HpYf
s15qtPmadPVFoGgKlldFpk6fZ7a95FNxuQO70VixUOPxzVG/1xAFcf9rmoGqRqp031N2OF1Yma1p
qYm8DknT0w1M2txj6qPx12ybX2og+p5OYuU7jeSKHPiNXR6ISXlHEKS+NdSUFRWLfu6xlZ5BTjfd
iJT6Sc72+bp8S6gZ1JCdBxpxl4DYlGm9nFGKs75IAsg03w4/ut7NQGlDVhb8QurAb1lpZFq/2jSH
sU4GLsQnm2SPfTfnRbm4Yd+gA0+4PBgei6fMNdJ/TaOa8hNXueA116DWYky6HvgmrECGKNV2ZeQg
gKuvcM/BfiltDVnXGHPIudu49itfW3Nbl1iLBzPGA56LPHZjYUXbuniW1kL+0N//1MJf/E8KhwpK
kKDI/JewWrmlYqYEbmaxw0u9t5C65lwOqT/ERPiT8kXMyQba/U/AWpa4k9Yk6u+FC0LPHAaP2Quz
N1FRvAbSVys1IXdh7ClXlsy9ay4/3ogEAlce+bc8oSk7I5+g7d6kmkdNGd33tF+Da1IltOoZV/pO
IChiTunci+Z6Q72quzBYG76CiYX/77bUYip4MPnuJXF6KNWPEXqUfvgg1XLX6c0eOjBlNrXFBMob
Rx4M5RqlQjtb7+uFZRVQ6w8CabyomkSeH7tnfOH2laCbjeA96T6nbC3za1z/9qJQ++swkWiUFJg8
MBRrM0q/EcEC5JuDa4+MrXPDvLgynbdoP1n+hVTyhF9cQfvdVhHQ5rvDv7ogHRbH7JZTc444YRvu
EfYI4IYicS5VjVf/PzWZ1KtLcFS/d7W4zOVKhSELVh2J1MtqMlEyGrlx0fQuVLuP7LqlvcNWInLN
1EOeqeHGA0FmXJpRZgI3AJGfLYhkxHs6h8go9k+zOapyt9Lmn6bY1MpFnkRJUHGfTz9MnaD30L2a
wb9QsbU/FczKGnxCxi6XSyiDnW3lDhO0kgHJBzcksilyCH4DfPWVliajbfx29LouwooycBysNeDa
Zjku2z20tQQZG0riHRm9+BS12kfrmL2QTnCSZhD1EDVBqY7W5CG8oR47/TjyBF0tKQmEwfGp9mxA
JVRPJxx6Jzrhkt7kzN+eJ22CE6lCOuTz7XKsRhVK5BgGcUYppOMwDdU41go4Xn2tUine7Kug+Jz+
TPXjGjihJbD4/JwkQ9UbDgEjS1bZffE1Deg66FLWce/MMHIG49Ygi8izmUz8C59yVZfyjg3YJCSS
RV+WAno4fPPwev43o7Ea9F1zElivecygACv8R3ScJa8UZIfiGy/o/S9SugIwAEfJ8POk7f5nD3V8
KRS4uV0CZEB9nDinj01lGPTPzf3bYmMD66IL6Un+BZiJ9BiIy6vc11z6Fn8SXGhovSHj2rlBEcEj
/S6hzPV0ZwMoOb6/sewMYTIDfj+sloAbvVvNL2QdGLesxzVxKbpt7m52Fu13g2H35GVv+g7vJN2+
aowDt6l9ZVR6uFevrMu/seGn0f3xr0cPUADQrsu2Z7ekB930zFwg0VtXwd21krmFs2y9VnBWayFY
2idQmc/f7RkYhaGjC8B7i+qNwjY2sl7XE2JlbJR84MA7FSr6dCubXA/qlGhrWN0meoKRWcslvT2w
2npgbW4dhmrCQNJaGlBccvDnDrMn+2DYMiz/71k7Vo0Pw9orMHRETHQHAIBgZG9/slGy6JSjIZUP
bh2jYk69COuUeO8LdoeWtDQePGawUMk29bweIBlpoS0/NJH6OuaV6hivJT7z+46X43/CNkH9DxDJ
GQhgRc+rZ8Hwg/bP9xE3bgrWwV1eKQk7/3JVyRNkUYeC9GPkT7oUQzq6TSYemEMip/9iNmI7mjvp
VWd7AM5ur1cOSvOkNT0/M4X4Z31oRL1oF6iMVn+Y9GU2qP1QVDPrAvnpuGlRBzloLPzIideZk2gv
JBRhwH7Z6UcHd83sBxh0SiZzGlwO+tQU+qbwST8vt4eRYtcbBwysPYQRe0lpwRl8dIJM7EPDO44L
dCkt2aFOeKALBCNZfKGa38i46qEsohHXt3yN5ON+J+aFrCwFkRgJ3w08qQo+dbjKdHv+D9IkPUlN
g5E9IRLLKHIs078R4urDi6G/jQCCwD0CZ7PSVhnLI9TJ0nxv4VcY36W4aqg+0A+b5Yg2FsWUcX4R
nB+NbFvUyRA2/zsGTdyDgkHbyYPy1I/V5pV+r8e/dGlBzT7QSVF5B8Z4skv48u3cNlLYvOpwrElF
yvspeKgc/N/H1+suWxv9Dy+GbcCniTsNbJPcKvnDm4Sv/NICJeupxkseHwff2/nv0Zq1oV61pv3I
Du2wKfPs9h/9CzZ6+HX1w9vUVdAuodMD5AHW42NxuoDCEw1UIRmif6Uy376rDWacxXUy9UA2Tkjm
j/lfHQpLama28Ke8CVxyeD5x5CE0gqxmSULNmcLOkhTMjzY6H0Kver9mkn0y2s9fX/m+tmrknvdK
gCKnipSzSStZoBFtmwBeNobsOG/zUJvOHbEDn7uVVbBbI0HMcHiPvpQt0xsVJUuUFHVeX+s2o5Rk
7Ln45fB1EgMglLGjRgj8v7ZEak1RRcMPPYwv6rztbuGEKG3WgPyBWgw+gQJdt9Cj1wt6Gi/bAxR6
6aXxBKZiNTKN+8RjVPoO0kFijfsGHr5q7KhEPhr0GrWASX0eLvOW+NTVEIAA1WeuFGQiJQYTBiAs
qD12AyI9O62cVkoDwcbn+8g7K+9fr+HQKLF/mJ8NpA0OsPon5Px7an/iPD3Pcf6kllmSDzTKF8f+
pna/KWMibgPSYuadeZ7joz32E2oGCFEjctWhEooYgmE7U/ulZY3K6t05nws98Kz1z+kAUCCISEYp
a7vZqyaEwrYnws6EWML0Rj3nwLq+7DWMdD+yct/EMOSfqRqR4wApRshlXzeetK6skDlY4jdjUgVi
HOKsxXqMPOeBLVpuylMh/0IoYlKYoGsCBKtO/tzLmc/NkU5/W0SkJmIRCSFjt71+uLhYsiMzam6J
6iXO7jGSSZd/6rvwleCyMnyLQ1iNxLW6k7XUzdT0brrbC6UnPTQ08GMvB3Oil8/y7EV/TgYPbMG4
B+0wSlj/0OTTHrukNVYRmRlSLYOm0htztNXDjeIj/f3CrZNtqgaZWMmUxdd/Rz7R0PTlGgAPN8Ib
wklys6++cLfFDNOpUa/Zcwhaab0EBqMK7mjltJwaC5GWv37gWdKjX05Plb5FoC/c6WST2K9cdUaJ
jpvOavv6g/DaEQlA6xJumjoEpEiqb0WKUduRYa5papnLR1BYS1VnRC3K2l7J2dp9SNSXtF2E5AdH
H5TmuZKQMONiubtchvTaV4r0lUhcy8lVC+4/A+qjmT/gaRBlhZ2L2bNBh1GXW88wsoQpkghGQ02o
j1Mpbm4q2ktub1Wa/matgAyEp6F0tI52LWOgtII8SNHzCfth0NCqp39BpG2H2f6rS4b+rq5VVRYM
EDulj/6XYIPubLkU1BjUkEhauQNaskludDfAWrdgDUgd1IGuNmureRQ1P7MB7/uQOZJVUuRnmNJS
W7E9L5aqmF27HDfU+EyqDviuRgc+W3Qyw9bjrtXm7lrDkrglnvHG6ytZ/TbLILTCJ7PfbkFtaiPm
jP8XFFQ4pJBuo4r2uv+YOKJksZ5sIHY1DFmPA8AOyIqer+kvX4uX17guXLj6f7DNcCxZ4PoNOcun
8gR5wYox0xqVqFsoZeOo7N4erRIpFl1tauiiumBIU7gsoZM0DPLA+OuNbN9k/9XPq3T5pBETe3p6
sKiA56pLntqGE/nql3Eieo7vHVOz2JQJ0SnsJh0ePO0fDBrKRUevpSNCt1R4t+cW8gZzVLLOLqAB
OdJR7RPSOCp7HEO/hgtRbJfL5o7zLTxzffWliVp09F26fxYUuFjVL9y17xRFZmHshEunsvbj87sm
6qPkvh3NPL71KVhZpHoVfnkVogaAtEfoUzioEfSXUl0kEqN2f6Ws8Hv5Qwqk6w8pvW9qORyVIP87
pb/UtgbiubmsYEfwMkTWScIkoc8IkbyKL0XsO1H5GalhzDL5/8l4uH+pXQ1QdzN3tCJ/rjJ9Gf6C
EnSH2dMts5GDdbIDuURD7UZwvqdRmWhzDVne4ooI9nsnhgDbIt0Df/c2CIZnOS3LRsdyo5YRg1mf
0ZKP2obm+DHWCCg/S9ytZpMh8QtbfXf9qLuSawtpxSzgZXsNRx55z6BlbTiLZT5L7PTC5y7x1Ewz
7JwFkW+eV4y68EVxQKRkUNxzf/myYoCAIlZRrZF2an0jFqOUdAEVCI6sqJhVn1gL5pvkkp79EVgF
JAB040RaJ3LVavcB0MXofsaacYkyEasBkj+NHjASqxryFCnvEmilzDs8Kuhaf6hv4SJkDdJglIzG
WE2Rg2GQGMeDwjLbcBygGRcy/lCuqSSbdHikcfnP1mB5ge80eDxjW4maMtsQtuNZgTc6AlsiAZkJ
cEDels3HEYiD7WwRFhUrba0WH6sVFzqLD45728AHdUZg5vZqV/Ehnx1VUStcqHpRURlb7ak5lEaL
ft2qN+QrpQjvcEXzVFIq2JJK4altgvhDgHSryo5qlMsAs/n/4Odf5zQXbpj+EWu7hEQBjP9y5uCt
hxsBy7mQ4uSp/BTm62LeqM8P9D3922ZisAj60/CRsF4gofTywpD+DE1cYab3S/54bVEMEdUxn35s
spaEbXBb3/wzN8kt1UODF4ysfyw5On9W8oREOMGwKLe6nQ9zX8Rnwgt3E77VtIROQCP9pdTatJC9
1zjoEVy904NdzOqXjONT2upHfsVuhyQ3EkjOaZovy4Kcg+qcSbxqjUdu5I9oqK9B776c99P5DMNf
iJLq9LQkS95jWayIUx2j6zZFiNT6fJOd2Ln8rcDIsuLccOLazzU/pZkFUFDtOs0M4OLMGDXSal7z
889QTnVJ/vEF+HuREgIvH+1TqhzllK/BjsiOCOq4FoYBHUph/WCG36Tsn5ZahO2uhJPRqri2O/lL
Si69msEytAiLYqG/sQpgnJ0PBLnuxsrEz1ZPAtIZvut3q9q2KkP8G0YDKsRDqdX/YqNm4U2SgZuS
dMPJJLk5MGIFD3H+Xes+DdiHcOgCVebzKt/nCg5spc2lI0JpNysVeOCNcpjr9u0jE7deviJizOD9
UnKSfPNzuDp+OOqPQUna/sdtE+CFt4/TQuN32YW9JXfdfy1uNwbmBrcCaGDbePz/lhrH4o5voUow
es7WYVC2cSYwXuzx+qyPXa7Ft9k7JJGO3EdheWy6ujUeCjPGcvZ7v8dZqqryZgoL0zDt8udwLjOF
JKbRMkdjsZgdJMp82sNpuWN+2g/qdf5zfXupBKJm2robjMPXlEt1l+RY2sQ2RMB9BnOC4SIjKj14
K7HvSATtcLKTanFnIPGi4BUppQnkQ2TCR+EgJsSRd4sH6aT1SRAsBEaZdkoFbxgs+/ehYh4A2UK9
oH9f46YfSneisXTk5CSmhMGoQNIl/V7XhoYxgVe2yCNoOiZIQlT9Ek7l/e39BLxp+roryXEHZxsk
P614uUbK+qwop4aqxZ02OcDDvR3p8qbZzxzH8685oZ0MgenmLrkP9uQriinwTiNo19TdHd1AyEdc
FXvsctVLgDOCl9m/dlmS3g63n9QygBybniMkNqITdfVWZXlgIVCGm1lTK/UNzNFZDlnlH8yxxI7h
LLFbnYY3kDWEjvEofXd/jrXD5hDlw4oLUAi4cPY0rEPXQDjtZuEFVyn5BLLpphJ6fokg9gNyhJWs
kUFAsW8xn2QLKv6LtuHmT+smd3Pecx90pl3mD1Xcapjl0xzUy1JD+mdEcgBbenX9FypkK9Xg8Mj3
wNIxpx45toauKqm0OybeKj9hJCi/RBQYZA/8GjkzqH2mH5HntsVv+fFe/e7Sw54++RIQMX2CkUgz
sx8rJXJ5rof16UPM0GUJmtlL0lhqBwW7U8JdooM7ssyDdVL3Bw3rNjba3o4JGIs9iwzx5mGrJ5Xw
OMyKPrDAMmsHNWyTikOUMlhbRCxzLl/ifA7imVifkHcjskjY2atpn22w+luttf7/h3zM+k51xac8
m3imI0sUcL6MT9426ojtmORcdB8kUKInww0ASBD7VdYp/fszLPawP8S9I/9/gT9edDSSJ1XMPtO1
elXfvTv9lxNJfl0H9Oj8OZuwsyjhHntaDJ/9/MIGWTKXZ5EUFuoQBKxzn8xNUPj/6rRQIb3zUIjL
Z1kcL/Ph1vyj3A6MX0VuYVBf5CzZU9PaqiTGssXILiMLhYvOTYLRePDSMpCRiITsrGFy3p3wSp2+
HxRi7X9TRkbEl+OTN0S+FV19STwYMZiphcr03O8tRCLAsx0RKzECWRTilPjLm3TERt0oohwtsz2t
7s1D8KIR4QDf2W3uXBGqFX9Sw5hf4AJIX5qcsUcDcDhqyRCBLCEZure85VUL8f8yw5meMJ0UuUkI
M3mBr5dVJF2Cb4DVB3YZ5v/+G5tPP527NsES5HEDC/7S4XKrn9yRw6daXR3uURSPR1ObVkvBI7Kf
V7kBvSrFhJkhYu0xelVs4dWJ8VAMSr8K8OxCTwklWRveOdJtXgtcmvHbdLzngtvX3rQtdtKZ9Wgz
fPsVhHrI3vWrQjsOTeNyDfMulEAbDXDAEhbLqXlBlLhR3sctirOBnkGeuvLJxAr/QB0s+k4iPzMc
6y1YKqaYX7Iq9Yo3F8sNhSp5d7F8dgwIbirHMBJgd6+m4mGijjkiL8hb8b1o3P1+RJ16kYit1j54
tHzaLvLHcIFTQmhGKWnY642PLSCXuyBauye+o+bEyMVWE+ld0MZ9aGA5nQ7O7OY8uS0BYIfvhyA0
9GTPx1kvQt+6+WBmINm9Ytx1Mr7npvQA91cJE54LpydXXV+J+t36KJ6OnnQ7Qs1r8C27/fkjFtJ5
Z6XM/cHyfxNXT9Xpj2mFUBgJW0xr5QARKPdOEOoNh8pq5bqLoM35ZDLuHN0iIOEYqb6I6SwWHwcq
UmfFuXIvaPddWqdPrKRnq097h0y4u7QmECvcwMxvpr1ZN1Z7AwUDEwmCPWcAQ3rWYfffbJRHwrbS
WLMQXHf6MZxr+6JmEvWjW2bR9UPEr2tYh5kQaJ6T8QLIUt205XbAJGe8he8yTVh3dm5TzcaYUyIm
XHKiln1TajmdYWnYQa195plbt1iYXI3pZ17/pAW1oXijksMv4tm9YwJEO0IRVBhwFKodGLxLBcRP
0Ln9llaTj3oyBYS6iXNMgin1SLAAp9+bdOdVoWsbYadFQ1hs776v9pheIEwiZ4CopQFXsxSKqh2z
9tm2EBaAowQRkFRVN7/z+YNM/2M0JQs7c9C5ql1hea9mAHlo3oDkE8xb3qC5p8jHt4Bdlt6Pyk4o
WTedrqw8qzad9/h3zNYDDQsRVj0/4MweS+ZOsu0y3wShC1xW1VwMZyFqdMFtCi0nc+CRWTOSQWe+
gMYAuWpWrXyL64nkLnD0gkrNPBf4aYRtnT9qvHLrXo3PMgRMjx4+GPWaF3noNhH99v7ii3NOb890
UxWJE31M6XS3cw1VT9eutuFdA1+R6JPUkv36HZHB3Hy9wXsy8+vzcU7EOCrbG1jurc9WNuoum9B2
n8M6qWYpHh5Ux7Ray8kqxLMu7UkTmLx8HvDmqa8QL1AYs9QnYNHqxPzMkKAZLwWATh5DkaTWs2Uc
W2fUG0fl/l3KYUSOhRnochJoc+5PEHa5uAHTyUu5x8jS+tANdhk4uwqd+gOGNQfvKsedxcxdJrQ7
hEanXhdA7QB9/vjmBPcZCDdbUgrATEaklrSbP/h7+yAcasZ4wtzOMS1D2Xg5Hb177bDkCzuqeETT
VEbpXVgbShAeMSsjmYi40RejAdgf4077t+McqeVbYxjUg24HBA0ZDnNcfCVvWfAYP5OUg5dI3z/I
slFddHULDXUZ2sPPstriGBPnYGUfNy3SLLQuHS4sTEjb135caRQ9m4Y1S0d+/ACB7CNAz/evUokk
KO11BwCrnp3Jeu7TeSTOG97SWVNxTWw2P7XaTc+owMqS8XEg54M+ljH/D4n3arU2gBiB0cJU9Pei
OReN1fNG7cQPuCF/YeHHuUYYhqB2Vz6I1IpsgzP1M0EF7FEpKOvMkzTWA1REO6IaGsOSIfuC4aWn
VVpcCZ3nr1ngtfD61FKDeaSh0fwFLrj0y/B1qZypF3zj2VTauVllye2JfqYGVMwu2MdzypSBI6FG
5uAhi0SHH3E6at7GveqMhjSocD+/EgqKL5UqbwnsimhKzt9NI0vt3cMY+AYeS6rWh1tekFhxG7po
63fRaOryZQlXpBpu8QN5JyGl8Y8twW8cmmkWjeo5NDRx4n0fBktNkfoDbyCwSygLlNSSqDti/YLF
tR1TqpvF+Acks2egxak+D+cRctQHTA+HA831Ga7ZPIQN7+qEOTihIPU6zo/nhpnpsjFuO6a4jN9+
1SLqyetnWg4SNE3UdmuQqcovUwpqkQRwcynY1B5IjTttwD7vMQCiTMXOxf9OnM2iYR3TKCx/9KbE
KB+evgkjinLP+ykSMq8uBAnp/d2zVmO7geBQvXClXCSiXCk2S7V5Z0ieOdCSdvI4oR2tQjDsAHQX
XBDTqaxd39Algw8UU8RWxsiIX2I1b92EEpuklCCrANxgEuGqex4AMTx5EypOQ7A9FqgsjXrrpsth
rxlfOnXKLAmX2I4PGW3uPDmixoS2QwIVHvpxtwwFWdjgTJy/4mBzX201LJQlkiIMJmh5GfV9rraD
Dkdc0BVIg1kl857KNseidI4mmMxG8AcKdJ6AfNiG2C7S+HASPDezlGq3RA6dEleWD/TQZY7LqUOx
XnA8E5FwknQ0lzWw1vcoBzbsd+lqPoBJXHniIv2kIliQ4FebgTaxl0+wzMmI3dpJndeJovDWOiqS
mErzmhqQjLNMVzeDlWovIfgVAt/Ks1KfVMUYWJMx/u+R3I6iM0uyC05vw325nJu6NktI1CCL953h
0GBqEDBHKpw6EDjWiQqC0d1c7Q6SeWERoRXXKcO2/FD3FgajpIBXkj+y/O+eUbMl6AUtZI4pbp4T
89qnOzso2O5zVGVI778w6z+LMKYQQlPYqdti9N2kSQZxjhpsUMcEXavqM8NHctSxBMTfj9FcOZv7
Kwr5XkSnxpdzKatwjK+0o4tPt+SBk/IFvsy1bji5LFAwtFoXuCI+UxGs8CwxE9b6nM4Pp7m86z8i
UrldFdJpY6W2Ebj2irieCpxul0lglVvOtCfS8VSe32wQVRwEyM6Mr91yv7VD0TI7Cmww8ytdGAu0
GsO261UmWKgfX8l/PVDFl10DH44DM2U9FXdaCLnNQEVdQNHYSmKgwBWI+TGTHV/ybSqSPV7lRc8g
Xx797Diwp4NafuN7MPOnkhwEiyFJLXjeeE4iTdeTqLVhkiguFD8yubuzQGqOjsopExur8oHlbrcZ
4mFTYVa/3bn9MsE9dYkYJlE5crAN31m6QybDrWz7mlTBnRJExTdd2ob65WMDE3fRFXKS68p56xdh
uUFbc7CAgPxqv+4jYG4v1NFaMAL9i6tqhQbv/Tiukjq48MEFTtH2LN1qx2Xa4uvkHb7NDwhBoHgS
XnRKOQ2XqvUD2JAjcCvF/pJuDDGeyFinri7A+1kqq9WLmJ/nU21GWXhlYwkf/+oO1vUQoXjPmxaA
cLfh+YJ7CQhhro0QDvxA2NH1GUxb/EJCiT4aoOmM6ywZhyNjTtkNmKxR7Gkf0iedcH+ytvBuf1KU
NtUExocq9ePhuxFqi+XP9tQ5bHsTD9rjDXXXd9SuxrcshvsIFUtxSsAx4c+5T9kMTVf12Ntkyza0
JlayTqVU98M3dhTCfpsKwKnLf1j+DqOW0VcEw6TruSEuMlo3F2TR04VPnvREIVUsjc7tOBQeZoo9
/N7RRDqOd+nfQz7iE6eQow3cFe5foPRX1qrYMfaKsiFdByF50ddlQWeQwBPmJFrxfoyPoPnZWfeS
avQbFR80vKEPj7Z6XOuva9o6Ah8xA15MuEMeLQZqEUOVMIgl56AkzZ3anYuJfCEl+frJy57i8e2v
NbNwGpsdt8IIXCQmVr7X4DMaGvALt7aPcLCqmifhc8JJaIGcQ11ww0j1OkCxhSufsr0Q9MJRiFO5
bCXuRTNlR1nb/6ZSQ+9StVFcLONtj+t/g7RHYBAtSbA4dLnSWf1fiMEJaKp+q/euzB9GLTs3f3uc
4vgOzLc7wlPkq3cMRX3JUPVKahW7dElL9qwUmfb1ggDipZOchnU2DPWftojuf8hZ8PJmtDIUNsHD
sckfCTkWJWwGOUtJg86jjtby5zACQvUy7uLdNpsqGRlqfIQo62IDlj2+7dkoWiFXdCvs6XVEcZXA
O/VseSYdE+qBBgilYUeYWgdWgJ6UOk1pXsDchLra6FzP87IlnfGmDGbKpzDe5xfegR4bfaxbh8Io
tnD3Whc2e8oOYWLFni/yPSwrFsyZ4lNukYd4uLGM2/ChJsoaj1IVaNcPb8PqKaMuTxIJKq+IA8Ig
T90v0XLrTPPJd3YWNjgTVMw6mZE2hIKhRlHbDvEFxhuOcwXe5Fh/tK4vo69PAZDiV3C4BbiZ49Na
2weP9/3x8T/WieRIXQA4ynkOhA2Jw6AVv/rhrjT583Z3uu0O0T7OqAGJ7odUpA8aKOztirc7Tkwp
VMNq0mwqTHbcNbs5LXen8GmCI2vrQI4cm4pLmpd5R0s74tKc3oUEN+HgBE2LcjanDR6qn0zwM5gF
UQyytwUlTKKYmVuKiFjGqU50c+UQKolCRYy1NxBWEBzw0nHmK1ImYNjOhiNGcGoTD5+KzWpHC/j6
/BYwHHdngXy1cbnosB8f1uI2YvqMAh+zEcqCJgL9Q1to0FhXjMg5awTnTgPWkNnAipW3mBIk5I+b
1yNjcU4SlaUVKi2DHkbzvjSz5a/bVqB31nZcsObMEN2XkJKCUwZyALGMEmxudUXd6m69txRnGj+O
WayPAC3uHdgK8M4SCkLwMEda8jLK3SLb/09NRrE2Kakua8M1NSeUW8NrWK4ddXOzCJbPIVhl0vAJ
pe7p9idEzuH7AR7hNbRa2BpbpkbJ4zmvfe2bH07HVj28Ka4mlZ+8AZyxmm+zBzTZmvdEAee48GcY
pLf9vHzVd00pecbKP+FXp2k9N3AnGlfQJGZAtYOdFiu5H28JSF1eUh7MFLkkTg3B8OrgbYiiM4Eg
2g1j/LwJW/jvHxWglCzljhyh1eHBByUZoe9aVqQIKNsLHcYcDAHGM0OUFuWYzvCWCRJkiWTKTKoY
a6NuYiLshc26EKKiO/dhjLDlsR/ciQ7Lb9lbwcOYV/3NCWPC7BE7u6j7rviCcQ8+ojXEkMOEkwln
IqvVjtfqcvhgSbl5+ekBEEvJ9y6jkMlZwV2XD94hN8QOomizi+yQSiAz2EK5IRTM8Edhq23WTZFt
ITIEaL2kbLX7IQakDTsXvh2JwhxIB6rcSWEBxzsnip42ZvfX8O76FSNr7SS3IdTZlgt369c8HZEH
iLwuqdCwQZ9xF2JmoB59JlJqYVsRimZi6YS0B4GrrQaM1pJfACimWVHjbiFsB7Cqm3Q2VDBlu8XK
S8yIK+sZcAM8fVSvF53j5qjAAzbGi6NQi7gbpelzYXpnYDBWnxObSeUIpghwx3lIdC9ft+Mx89b1
szcCohXNh0CVO1q/uVS2v0b5SKgFDan+fPxtMH0N0IFUeFJLlAOy3XTTO9l09OsITo4po8C8N6jT
Pu6bulNHsmzRCmYdD9NuWjkqw+5Tz6xsQW9jhWcYPfaLqJkvSAfwKF/cMeE2m+6CZGdtwECiqhX5
t9Z/V3fN24Fuh/wc9pUzze1LCX3yP0WODn5b1+wwvH5tsC703s0Si2+N69SVFAlOh+ucrpS8DIe2
ZOA2xaPLH0qQ0wqHvApCU14c1+rWkAsOVOcJvVPI48TqZfO5Mwqqv3grIfExYEpi6Co89fUFxQjr
pwzBJsefv0LqzvprrdcZa68e3TwEOLQ7zREWL2oOeNEdKsHBMKqOgMlI04fuEYLkReOEEUkVSNOQ
gVmuzh8Oy1pmEizdTQJs1N2ryrg7F2ermPRRuw3jW9mm5doLwt8hHPfhLFBarbHGcTyKV6an4iD3
cYkEPa6cAFyiC61bWbwdKgf4wki1EARhsTqG0A/x15jpaK8X7iB6f6JaGolXxK0WSXGQqD3M4hSK
yOrpcMa/vlDEUfu61JGDJZCQ77U+z95DRBLKfr8Af54gYh2uTybiCGLGBhrtd3igfS94u4DOnhMJ
SVuuVfyaTzAI8zah5XPlh/lFyO6EtVAZlsaxFn6QGJHORkuy9hujqYr+KmmXd5H0Vr36xEslANB3
Q6cJ+qu6ZXR9W2Q7iVABVx7pDWIXhewTSvgewBX62zr+6ueW2r4cnj4y0lSzW+JAN5TEK/L3nmMh
nb9y6d/FG+ovAMA90/AUd+7jOmlO+3KnALJd1Rrj72vQb2o9WAaMlCK+iY2RP1nNjSy8qsANBQ5S
5JQ05yCHfJyBdbB6On/DbqfaA+R+ypRdprjNi5KXN9dv9e7YbyLRCGHHbOHYSGdV1fHZRJHTIlEi
WLetYz7v+IJfMOJhAi1Vq400Z3JZG/9sC74id0/yWGJuuLMaMLLjkPUePHlYI0mV5JZn6A79PFbL
X+Kh1bbfDF0yE53r0NRWfbnQ0IFwdEYCLA8rY7DpVzgBaPDtzwi60CX+Yv2gIRUcxidE3vjL2DTL
5JCsI21xF6wmjzV9dc9w0bzTPqunNweqel2/6hH+CpSX/McpMXmh16/Y1QUZWNR098PWWx6b2MlY
fsdrCPeWgECbpObJcbagcvS8GSJFUFk7+m0muarm6t+MWAwspg4aXet5N8u5YGK+oLyzqqsMzums
sJl7SUtxXt2Lt1N9S2B/TL6+xbP8wYW7MmY8qYZgfkqU946CYidWNz2co/zbPldF4znKOobKRyc1
yDQ4hoZdKphKWF4/DRsU8v7BhS2IRd4P2Oh219T+XF6Z9/0hzGSu+tiSP66fAR92WnznV/YX1z91
/orXYctVqKd4JgjSlwq0l6mOVvxjWrpu1WFCqtNNH3PSSQLGUJhjBbEgH9Q9bsoorbwWnxfxaN/v
kbmwXTOHg916y+NfvqywUMjy7e0tTwz1Ks1xebQRWfAFoZOaX0NuHiov3d3KSmmhVCpuS+ghdQqp
K6KWoejd3fB1Mj/qJnDmRqre+7ip3DxZ38MHQHkygL8t0pNLuJZ9Ah4c7zn0oSHNCPjHdKYkXUIc
/rK2G/7nD6YWJ6bfmXW2BIi3luf6fS6bkP6z+KJAWb4s8qz6OGHxk7K+S4u2EWhf07CBUgX86UIO
1gLMcyLNHrFYpZsCwQISVNpDgoTd/Xe95q6YOFInJhW3a5k5RVCb4Wbnvgtw5v00fKZkgc3eDw9C
kkcAj/jKknsWJo6sF+vylGk12CYeQT4tJQK3AW3GuuRHLWNU33GGQByrvCusKl1XxLkZCokmIm7B
gAmC+utVG2iOwnrxVTWXVbpIjswSA7tWkopbkxb1CFZzPRMDNwmY/gSWFZC/bJyQyNOhUDmHMwtt
YUOZ5U2OYv117fjjT2dLH4jN0RUDZhrcgNSA+i2hp2emLut8r1JaGYThuNWaJ6eLPKK5AVskbM88
k11bvTgQtFPOvtGJiuTx2M0p08um55bsXR6AOeyJL2JvtG0W3cNwQfiMqOSQoC8/cfzCQlCPN0SQ
f3DMdht70CrQtc9uQIFloSrFlhBYdpjtCIshHQg/o9nhId3KLJC2T9x35C9kbQkksPfq21U/Fo8w
Ode/UZKjG3FqmvjM7hyVrL7wSr6wSEhuj4L1JM6mO96yYjRt3JZByjvw58/y9DMGO/n402mzT1q5
V878MI2PuXwnuw+BWj7GC+RROIMgInDCAWtas6M0YyT3WztX7uCuO8kMWogoEkrswb3caUvggnkA
SVaLrHWjvp49lpNwtTI0zvUjDbxZlIbpw9cAOIyOqYTqClOwheMS240kskA6a16v6Hbs24R34R+9
VwfxLiYdgx3FLfe5gjliaFQz3gFz3R4OdELHvd6/9HtKdPlbTe1S5gNq8Hhb8BrvQUCe6/10Kdex
9U4xdkxtrVCZgw1hGz/ytsT8E4xdUsKwkX87TaG6rSWB45v+Ff9MGisSPaDGCeKnt3rSCE6fYbTH
yPzPE19NJCiimsZF0xlP9VqyBpI49bMSVyGJEXWxqNi+SZdUk1SCBODogdNPVakmC8CvweBPp/2P
UGDqBDkng0/txOOlYy6EuhjK4HQLYn7BGd+mp+MnERcFAwTt/lfMqZRijhZXyyZSbQQDyZ9Uvl1E
uvCzgrYZGL+kljQQRYo+R7AM8FoREuUXg9COIwD1LHWQyMO7SV9m+uuQ846trKWtSVVrBrOoW+lu
cSDFwtPwNRsbvh43Hv7UObyyktIpVEk8rjtSbXP6rLgUddHGznu0UWniAbZediOC7IGLpMuOsvqM
Uet4fiChQ1JvRo/NjPRPj4ApFfdfbNgNJr3llG6ayTkZBOgMZxHfjifp61UsKynP3QSJXr06hSZW
IbS53e5h2pImBp3keZW+lvbNaqqMug/PdHPHhaVrND/0nFM7CjiwHIpEYkgOT9q7EFAMMdQ/QStF
971GtAtTV51aobNAi7gQiqEr4HJnwDLF6qHbvdpzvkI/lylPye/hZDcShfBneo//oW+ULv31oi2y
mtNTqOohw5QiVbvIXhJEtn8F1Eyx+2peW5R4o0F4A4y5Utem+CAOJtquMqbcRId5dvWwnIBOeJ/E
AVk3qc3cbjxr81IH/R/1tdrB37JlRDtNPqPVbNxmYRY7pKVokhxjM8HvqlEbwQ3Z2fXXWgT2z0ec
Je8qUGAOjBovXNIF0gWnufNNXcFNnPl6jW5dyFeQY9atHK3+B95B6hxlatAkvtpy64SB5LgnO29t
ElcF+H3xykIYK4tiyZmdh9UTZgOlWtTsBRmmrP3aOZTARRITSkgeLVDvXVMGJLZTb02IPB24HhIq
vkvr3Y7FoDvX8zWVu9hSH25OAZzao46uomsem8H46m+1sPdO+vxgaRnw6w+1vtLICijpOF6Co+Rv
Pu3BIPcu5CaCMm+DN50HIqXwaV32IDTXjXLo+3tQX64/D7LRMXBRmo9qk6eCml/TuY0ijHl2X0W8
Ku4XK70il0y0TiH2jmx18QJHAgFLWAWgbMRhAhXKwJMO8f1EmKHR6O2T7/RZpuR9PWDSK8JEP38g
kia+84F2y43J3P7d4ld/hQcNgvRYcvyST9TZvXGjhYPB679GaaHOjlhKLf0fsXPAShHWWR2bILe7
ZDefdGgkA6ith+3sncle/616ugcTFJeaBwqz+6+MxmtKy/l0H5OQneJEKZLgJDCTuvuu2vQK4tKC
nFmrhNsej4yL5ZsAmWwX19ivWhjpPtMax9YRe42gRJAhUPrKvXupJNntRSREvgWs5BCN+vf3bHaU
WEkZ6r7dtuIwTpxNAQZ0Doz4icb8VbKCeUqdY9I7cpoxOfc2ayy9KK7aio6hJou9r2eJ2ra1TTvR
8eCxWqvv0qjNkGtuJLpOxsYZr+pS+/5o9jTKT3UkL0frqAynVwiusa89ZnPPldrT62joK+LSOjP2
uV6LRpKcsgmkK0YL2swzTHoZruCeyj4ge5Ba5kD1rcO3byr+43eoBxruJTjSz1sKVQ/xqULP6FkQ
tDGRcE69DdID/imV7I5LNvyRFGUD8np32swZfRd5Z+8L4vEjlAF/fPCUztAPiltoIyon/G0RipAk
pumVqvCBKbkWvhUY7aui2Xa50gsvPfRzG/TGYz3slzXhIzSF4s9iAUXJ9w1rnYiAN6r08CNW8L3E
6lwldpwHlAM0InfKxHdDzv33UEEowAJ4LDWiN0/fUPyCsCamE9AhYOkjuxP21h/fFvE0wRca72mi
t+H6eVvxFuWrMf2humEDN1ZEzT3dPYJi1CDz1D2p39nQT1y3MhqAO7Mc10q6d1/HJdbh8enF3K4t
hq7eiTt3K65Lwdtvy4ejNqDoMc/ENIuxuBvdryJysP0n1c8hNk7boJn9a4nfrmo8sXUvSEqKT6UK
jQ5W/4yHmPMBNxx+6Fu0By3GiAN4usblNrXtYDuovu+aEcYH6BO9zJIDZeW1S0Gwf2RlTCa/Bxj5
HWdt5U7CpFItUNVNEDunObFavyOIt6c7WGwRZzPbC1Y6LGTZwSvFkKJski0EoYUAtTaFSE55ySg3
rMovdEs/JQvQj0EofL+PJcyHXncezFi5hbMiD5fYZMuOizOzpQP6wkKW0M6+e5nzmsqUa5tSkyoa
ycTtQG/y3eudG92nWOchki+rRaO79MGcoRkXXvj+Q7P+zz3K/EPmdUeCcscdfp3rsbcCiMm0e2nJ
c/yYlQ61HekD1/FAyuCFMTDYOt/lm8GFy3CsBddOqnESACC0DeNBWFU0iGmworBZ2gqq9eSFmOIU
pEUewmqH+ViQL/IiMkGyyLwL7ZL9Je72qDVHK+fhbJZDEH6YvuT6R33KVgPcF+V6DjfGZPRzpAkw
xhy0CPJfOaI5iUQ/rhh1FH+xNdUBX7q0ME5pcHzZmJ5K1pEuRkMYH05ZKUOolHI35/SCyUvNtfcT
El0BzGpBXvo39DtrS7XnQ0qHMnKDLog94YrumBRcJMopFogwecadkfwHw63nOyLRVE6ohXk0crlK
3/3As7jQViEKCNRhBSp3XyQt/7dxsWKA415RjV9CNEctdt8MgkPqTLEoEUPN6nwyv84fuu1HpB8g
FdOaUkqYVW1OK6zqrQ1lPwMq2/GTeLsiMs5EQipvO9evsPkrMjPkNQuyslwEEHrkWv33witPwagk
l5HGRiUc8PmXQemmFmYfCf4L2E20tKYfS0MKAq5BfSM8DF1+TBrb/lIVxl2Uk7+UA2tze4av8WUk
2KjWUlWTbH2UhoAYe57zrZ/IiH64ZmfHMm9W52H6uI+/Fxc0lEfwOUwWrQiwfXG9fqo/NRmOtm68
pJ2ugwhdllrPvTrqJd3s7sKOcp8Dp30O/+Esedn8DXPA1ba2hNUCz8CufXL4UKlMb6WI4uPU84ro
sbaxnY0DLRs8mC+BVDp2i5H3YumFuhlNsqLy5uoXU/emJ7nrm4cHLwrEwIldck3tQhAfiD4xypXu
qieu1KxPbIEEbA94LOzomyo+0ogPOHWOAQCt3Ke7iIqtleDSn/uSgeYuRlTL1xB39650R36ToyeS
sh3PKQqHX8gUHNbJGmnQcxAM9+SHefCiJAAFuW/OciXiBq12Px3+60inuOYGpDNiJD0rxUlEWU+Z
TToPInYRie3sRv/EIahPYDU8FPB/hRyXbG/tDB6UMnVjo11DJPQKyTXwJmp/LqwgXw8uw/DCHFdE
9SEscRU4MivMgXjDYsZjBHS9ssn0Ik/izVVAlVTAR74sXl6vDnjxz8eKvsN85+ZW57rOJIAMl22E
wWW3lN1eKUPbVQkqIcbocF2akxCyfuUd4wAtNrfVGxOh5KKurL7V8umVe93TIi37TMHQaJuNnAMx
eQdMhbL7HcHrvpfWrDlqJS3rJmBVQzcXrSu3S4s2t2579FbJI0UXGZHz7sLRaa+Kz8+eB/EdxMme
WPm932Ovwfg5Dw0J5ziMjFKPLo8ONXMNWiUrXuUNuG4vUiaPkwxdtyyz0YoTey3ULoDJR7DWUlvg
lAz4l6jMBxwwgEUGteHrhCc+hAv+70yIJQR85jI/7SRDb9l3T4ENDdRVoXFX5KBZ9sHORZqVRukl
HlyJAE12xjrcvQYy/8qirvWKkU7UM9Pt48Z9LIz1TNCMNABwyXv9692xDrP/gGz2tusJbY/X9/nS
PTgHrQxrtlcQBO9UYvS4t5tEDrHU4PuU0+8yk3swPPc6u31i1g2mNey1PgyGaOXoCcOTQ4RcU0+N
NOIvz5YG1fRV3I6sVJg92GHzPW08Jerp0LLNriZe5sB95Jg216R7EPurZHu9bhBTTCZRegjlfN++
MZH6aBQ9cCjGulIo0nRjWbwhwcHlsOvUWi7kdpqUsiPNCDLyVKmM4owbA3Lm0t4sP66srPWp51jV
8h4UUsdBnlLNGr2MtpuLzF89R1mPOawvcUPJopuD9di2Z3yu958oJAzxaYMYpGB1nPjrxrFwSYDq
GWC+I+Nabu5zLOe4k95+QoYhoJMCIJ5HzPFVMOmK2o9sGwkXIr2QLMhMfSXihSPa45Crt87eM5Zp
aU+rmp6egfVn86rbZbMKc/BbbdXVLir0k4rzvvmXd+EEInyzoQt7tO9wWVPVqXxKLOtk2ezKgTuS
LKFzmEQwB+6/ASqqbFs6y4Xn7UWwPWIL9UEotW4/NPTll/2xWZe2LUrnlihGBOtEXcleFPSYCRC4
S29/334HZyHRPwDlAXe3QB1asXgGrlhvgAcRgabf0v707DfB/ej8PDLseWX8bVnnNHzspkES1fqW
PHHZG2fKOqZbXrB/UZTHSD4h9yt66rdYTRM9fnnc44cZCzn2ZUkcvM3XkPeORj9kT3OplmG3xGC1
7eJ+4vfjhetxBhzhEqcR6PIz8fUZMsUhUOuLLObTdynqljLmzSMMcC1KkF/2Bc+bYQfXMjCwo3hF
9KBoybEDMYrG9ITVJQbtjGULPkXbk5LBvF/4yum/JBI2f2HRjZ6WX4aI+FQYVxt3L7njUemXeCTU
4DiXkIDDbR0cBl0MWLy28yWLc0f+KScWPGs9dVVLBGOeJeiWqoIDxUvVtq3pJVh3wfkXsC+wacBI
lHlqq2IlkLcut13ElCP9A2a5pD6hP33jmeN1pgkeTKkmWlCG3OXKcPlWwztSwwOiMKSdQ9/4yhQR
g4N++2wOWWV+/ahdAKE/h+r8fdyVITkWa3z7wSzO/hNTAZtuAU26xYmuSkWA8+ea9g8X8E+eXHnU
ANKOsbUNRlvCWq38MLlVa2PE8rgi0Jo+ugQZoLuWbngL4fG3d+elQNzm7e3p/0EfvOdro7FPwntb
4KpyQlyOKav4GLG9hSdprb87nmg2iCpOLckouc0yPkgMsFrmeZXogTB+UuBEb3h2vK0+NUWTMGf3
w+/j1C29KRonMTp4slkrSAYUPkf+sGz/BvI7C0kXIc2Oqse7weg+kChfh5DY7YgV3UHLPAdG+ZAO
zEB7IhHeqgBdOb1aup5sUINV41ydYVN1hJGFGnuZUwIteTFHaJuQsSNnFhoRP0V0nlJuhr+d6hOH
UTNmCU8a5WPysEilfmF7VyvDRIeIMv+soJDSGWmDPnQqdTBK6GW+wPFTrAJMJWjMcv2p2eGbdZmd
6OEonBZfUVfuejfdcXCVIkx4FAlsFFJL67kgw/QVI3blCoAm9UwvcRCYh5B4PB9f6jA7a+wmzoos
FMcP/Sh51l1HMHdmTAStBp7J7KQYdsHdHRloPzgjMfJVMeSNYWtzPwyloFQvpi4qO/OXnkSAyKny
+9YOJqce7g3A9DPIYtVR8IaGJ+dlGRb3b7L5L6zppVjVpuqpvHGVTWtxp/dXlLQ+WhqlZZII7bZB
OWTPzfViPeQjRGyd9oDD5oJK10Nf+UOrkiJCmylLdC+c1QTBGDJfiHj00QSaNacrhtj/zHLYoio4
sBRBSwm9+GeBXD8zOfhXARUF7/Bcz1uUg5J46rRpsKxDhkEhrgFBmL9h78dVALAhjFXWrpHISmzS
Hjtn4cg28/FzAR5rNLPKuhCT4Jbzpq/4jpKi9+k71+jQUZ3FqGNpUhALPxCbwPD8UgvPMN+X9aEd
hJK4ugkXB+XhC0DoB88+33HCrywCsF5Y4kw+qLMi8nyAabyjCVtXm3ZZksuWo0XsrUrbeFIl3xGJ
DMFKEVnMWxq9RXoomppbGnXK2yNWCXA0NJU8Q2zVDYgC844cX/CVDogzlKyBKyqiDYX8nkMwAuBk
X4YimOqZxcSYre0HJzsnXk1RtEWjRK7+Ogdsqy8/JMjktwxup9SgrG4hm7LZcLog8+pV6n9iC6K0
A9+j5ZZAPF29MOAjWJyCkpFu7TkDfuzQpeRnlXjAxxnVgoZ7XGq3g9ZJNFE003DToq1+T0z6u2ng
vnUilO6Oum7Odl0Uh76dGIeXPNjztnLoMMRKL4+dMvFaFT8VQLt7ONVedlz3BQvdSI8RAreEO0f/
1nEn55brh8l5eqgIP+W4MKVoTqJ4iTftH+luKgA5M9gkDDR4w29wXWcu9wakHsHRD0SIKtywmfka
1mygxCvW2jNZPOR1plqngTmvRkeDo6A9xNTqyL7etXBQL871smuDYgHPYHLeSsQs/D0UPBCkRxSE
gjToGR9sSSHj4UEp7P4o43rNYAe1HAxvU+c3ONnUVojKQWzXwTN7wwGAisf9+OweTNXVReHY+IAF
qUTCB2ptPGc5UAVY5hTwgD6J/PRkVXRWSfzzhSPD0cA94gt0Y89A0SX5d0IAtv6yKecL/nspH9K6
czxj1pZgGT9njkvImr5TdsoZ2OCGoPQbf/8dHeTUwNZpFjjm6fKO5Kq8MDsGxYR8hPwZu4mJAuXo
yVUgl3fpHrss2+YbnR/SPDkT+u6J/D9qA4pWL3cBJh5oHr1f4yTK5/muxXPytDbFyp4oifg8BQ/y
cc9LsTTgZWxtlSdQT2Jy1Vz0UjoAvFnogRbLofhOExQTB/xC8qIbguFVKlWlRdlHykRN/BQoWNja
/3kPClganODfllLv1HjiO8+VfzU3f6OvOP6s3kXr8W1I/E927oxw6vHTiCoTnBNjnai5o5S9nnB/
toaU90goyEwn4DcmzyjtLDocJXsE+g7mE5ukWEQ85OxspQ3k+6+x2R35upjY4mmZj/RZ5No5+3nC
yBRE2CkaYZjopNiA8mAl6jH4mxm92k37ncn9i2VJ7XDWBe1xkZwHtUlII4mHLmy94fevIctAVrBf
EeClsfkHgOduUp3LZzbLYK6Mztc5AhnrDYtBiX8+n5CfRMFPbVQODYIFRXJQ28LBGdvmz317fHBM
FCFUgH6LUIEPWqEyxSVsSalYzFSQlFnXSlF4Y3di8KZ9dfdWJNMbnhNwxRpQpyRnoT8QydCbKENQ
mTHfdvy3TApKPKxD1DG4+XRMNP9zIGtaL0N05VM/VoPWTvP2//VQqdxGnpjMqkKi/OiMZt/Si9RX
o9xg6cAD+ivRhcZsEng8mM8i31lYcZxuaaHTPc8aw4mU5DwUxbmRD/EpvQvw5XCHJxRtqEMZF1FU
wrT/RTMRhrOvrSYUwn9uUOyA6poD6PgGkln7fF1FvhkXsrIDWab3ZLz/rhKX2fvD1MQDeNN/jHiB
xRA6sDNiQUzZqY9URSQitqVkerVywb7TuAOrF/DwCZsSb9Y+frDUjm2cJWGEF6f5dS/FAbwAX564
kgbsASsBGdqLeDwaGsE1YOaNn4yZIqTqQZ/ogHtc2Ck0sMh0q8pCJi5cR9nrL1BM8TxVkhiKlFWQ
jH4soqJJbZHkC8IOxTUE9Vw5dXTls8iZGVJKNxW0FJ3T9ZN4XuzOv3UIozn2ypy82lhC/Sghltzd
cKbQbsEUewKYkWZ/jCoy74HpvTXpUeeCgjKwRfxgs98KzjHhyVCA6PWKm+bkAkBdSSnChL0hzoBn
fm5VCLml0364RNc1rAigZ5PBAt5ImEr+gVrObyyfz3ibs8S3BWa7Q6a+xeV/WbCclRW1eGE5FD3m
tjv0dVtMPJwS6j1hH4Ra5i9lx4WrlFYNZeF7FehZLq0JYOZtVqDgqja3DECAgoD34VVJh5D+gBlJ
ufDJ/a9SG8GRTnRwuw4zFnBjCRqbnhCVXXH5fNIgOvHTv9n3LLjJ+Q5jkmdLELPdM3dIRzX9DNyO
d/9gtWqLztjqm55k8NxUExWtTA2G1K8rBVrMh1MsngxMzsHhDKyYySbmZCX3pikKaALIOAslcbJ+
g6Gia5xzXs3OT/h0agCo1aZkpdYpL6V8jh96llXh+faY0J22flyHuzKxfdpu3pIaj9D/qL02MMwY
KSLpKc6ZETxyrYdlQXiv8oZaopsvUWdEhQHxznYJRTSTwxTuwgkI78yUYPt4Q77HWd/7+9T3XLln
To8ae1jdIw799aYRljleq6DBQtg4o1MyVseNKpQA4pAyNL6rwU/PVPY1c+EMt0DPXIc2RAYugBWS
yvlebpS68akYxwxstOFWsCQEKVG+AilytNbNQ5INyd+Q+W15Uf4PWxC/06B6EfRnvnoOLGSe+ZWO
9uI6c2hQmoLt1FQCPd8vQxraR83Wfac6+UQM6H5gQu8OgEhPLT1lZKXy+wdDxyasZ1IzQxpP4IlS
4/gSeCryEsLpa5r4ZjASETe0t5J6lRtJyfsQv2kPImQr9hW15nQyzgXXadsLY6QLwSnONSSJOCW5
KWhs3562lltwegLZiQClTQ+76+S8nALNZf220uuBcrD/0tNHTwmhNlDaZjD1hQrqNOXhnqkn4d/K
kakVmKP1TsWJH+UgipVoUiPuwT/4UMY/C4eJha9Vd6oIPfvvQpBgsX2DUjx+RdUlI6u9v1bQvJ2O
baHGxu55joBnr0HzLmPF/Bt2PTtKGKa4mUUdklLnKvDVfO5h9GVyXYsaRXdTqbZ0lyJFF4XoYg6E
9qmFDDq76OK/FR5DCme6y/hFpUFQgshQ4URjolgJCQfhZE14+O9MY2YsfabtZrxvMlrKVlOsNsQV
o8IJuZvSBTRtU/ghfFfvAsaKmzDxKyDJxuTRsSHcPYmSfbdV8eFO0ztT2v3TlCfAofwmjRTimT/6
bZnexBzdfTMNm+R4Mud3q0gwV2hiXHb6IUHG+DxSHbUIqasz/zPfYOlH+/Q3JKatFUitn+uH5q0A
smHnEqzWARC+EFyukQWkrVQ0wRGeqVfW75Dov0aHXYKjK1ITUJPwpI/NhpIsgZeHGy1l8sDhMTI/
T4n9J0NXGL8HyxBxtwz503qcFYRF4fljSizHroVEFNRpnDV/l3QIy6NtOXBgKe/+1hEKGwrTRfzk
5AN2GdynvLfWO3Al4amLaGDkLHiWLWRq/dyik1TZuFHw0wwGDet4GoeGYJ5pjNibU0L6yw0zlndw
bRzs5W1mb6hV1CoplWIGMPMHgad9ctE62zfJdq6v2uhPZSPQeJ7yBGgl9ZECbDhZkpUYySZFNVfH
lHY3pKbLAhLBR+jCAErqG6mPzCfvsbloniDHM+xhj5XTN8eNNpGNnvbOXVhlnhiEE/afzisHNdhg
2TcidffY3QAHnyMTeArKDIMOvFYtDNmaCZoklVBe56Z+MmUouG+xwbbC5UVREUdEtKGmoctZrJkP
P9ftu5w7H2is5jntxyV4kbjVHPEvat6nWpvlFs7VAeZE/133HzJadOMI9vb3ohtE5X88DBnlJQzO
hf8B7mHnggWLiIYl5mxiXtQri++20EYsEJe2fLZaHWifugjwp/8yE7+ldIdI4GahqLNPjKDGY1QN
bqw5I+7Zg8FmdarByPl046JHxSkl1KyIs8brNUgkuuS6+k3dsuy+XBOGKcCGB3KXez179qwwMedz
FXKwOkPOtxbuTFZf9MykEYMrMkhYK3jRBESWKqjqxiTO0uQrNuwZ2oT7vxkz3ntEl9mYwd1dlmlj
nTQKEDHhVJ+7wODz9O3J4WFjDm84/AFmM2xL/hKM+DPFmiuqR11OrDUuX/DaWSVOAQhdbV7eYM9G
gmHlODzrYPO6utc7NGfsW9bfPCE762EbYGXTxZl81RXaya4u90F6EgXd3tTznQPkP2Gs0BoK2/Iy
v6h1pLz//qB/WGp82D1rDPjOPDBNtlXeVgBG3bFQfn1cI10V0x4SX4zeCVEHk+naUJDVK8E2lTTq
ZpFpY8lK9/kPbDrUuAkNx7PWp37+5N2kvoC16Dkms0ktTX67B5BKzQtlI0GEpvbwziDahDyjkGu8
HHhaWZYnucWTpeUr2PUiRXah+cRz+Q0ZP1jde08b6HsZb/7Sv2lXL6DxyNo+nShxlvXqRylV8c4/
QhLOmjT8yCUNeHw1EtwRnzPf7GVpTJBry7TpKsWRajEHi+UpLpihp3DT/FdMepsf+cL43Vp+dtTw
Wk+lgrny78gfn6RCljipazgDVXWBr50FjVOp9RcbGAs6kXFiS3Yir6pTGN13CRme8wbadZy6u7XO
tj4BKFWny+mA0lb32W0qg/8bXfJQE+Y89SRUGq/NL6r6PVXOyFP8s6VtNrCjcgm7fwQq7p8oJRDG
ALawp1oiaksCZ6FMZzo0ya8RjNHv50ZDjv5M9G61qd/x61WpwZauUClulPNn4ifdgJDU1XFA7QH1
YblcVIfcuAn+GVuBzctuSeQLajIE366vzTMbaqusQl8HyVzEvWNYJAMPLUy2r6MXHubQQUrVsNgW
p7EVCifEQs2k0J15BKp0pwJwClZeIQ6y8SSZN8sqvQIh5VHmuz/09Yg/pVjoSlUULzg4HpcUSj3J
1D4q6V5waJMKHvFqAX2edEztcaLakNCoJYDG8owh1sv5tS7O0hJBRdmc8xEkQ3pteWRs1+pGTYao
3CjGtDCDlDv3/24Tc+1GQZlPcykk0ouUsHDsWQHm1596Kc0iKo6zJ9rZ+xKp7B/Eg0TSUqyIEcwL
IvM/qU1LUvQRdhjrGlkeYo0iA5pr8nL5RHW/xzgAkmiG4zmMKbSC++cXMgafP06Sbn+keFHkQl5g
cMYUYUMdzJ3+HiYfb2JeLd2xuk1SqmyQVGR63ZIHXhXxEpWgYsfmkReM0XMmPv68uIs798cFpqy5
1mT4IT3YQ3GoDryV4jwCrqSkYOfsp2bz75ZfCf7kAfsuaoaoCWiwDHdRll+PbuxPlL4BSsj7Lhxz
pKZQgIMlwAvvT5eRBjvbRNn52CM9Ix+hKEHO+O/Z6tiaCvVXXzSM7BlsDD9Sh/YnOH1Rmtedh4cq
DtMxR17xUz5xfUhbPD4f9fQasBqtplbNOvveueEnH3SsLMKdJzNGLUC8aDNiWFi9+hmSndrIOGBS
siu/ml827Qn2Jew142NXyZG5tdR/mrNSw5MOXcxUqZHGYThcu5bTGIq8JA0FsnHaC2QmaHfi/gG/
2rD8H71ygqtLBIx+MMelaJxpFPbgQ+3igWKhDUIsV/v+zR//umo4OUcYj6/GGgtEtp0UjtIVYLh5
IhCaxicmkVG6NkuN4C8F/v7Dstr54f1tqYH7LYKfcmlWpsXzp57v1XKErbt9d8hosp8a9bm6afnf
oT4dWOSq3W4Q2ZLbgWLlJnECGQ4d/AicVbd6K6eHHE7axjfhAUgXG+HLPDanTaW1YDvrtMTbV8HN
xaZ1lThFtRUZtt91ze1zLotBodkOTcZ9yh1vaW9zRy6OnVpbrwuRerO6gHng7P2yZAtiGQcV3xVt
3dFPBpf2AsvuWT0Si1LjeFtduAxwn9TbMseLWwQal1gUgmGwII3PJk97XY8qP0WO8Gl+jAOv4o/d
tNEIjHxZ3loc8ClbIbE6qs9a7BDjExF7BZabh06ShQsARw4fHt8kfLUiUJ5R0cLa9QzgPAar7f5l
C/7DrK/sQZY9kQWiz5f3CjOgSpnzYlptU5S5bFtud0qq+eHLBZaiRvf3vSuTbZp6pcd6aT/1sOxt
f8D2LSn1LeoeU2GynMnTM2HEMMqnC4opzrX3Jg0Wmc6qgYuhNrxl2X5dKZxK/PKDyqNZScTyqTv7
BobXiH7AMKiJA+YQz4n6hqxtv2Ro0MilfU/oKP18qQQydX6LuL/Ou0SxS8bcKbX6uXcX08Xf/xRO
+yRMSwOHWx/NEs0nvRt62pblRYu6Aaz/91o+B5SFoPXLVTqfhGctPWGhVB2HTjKkvfxmCYupr6Io
dY1aSCvqRpCNZCtWGHV/VSWj9g+MMXBco8YlPJ3PlxKM+Ubhmrw4PVAyOUizNeJK8S2XS+y0V/dc
nQDrGc55nQEQqbsXpdwDATSeIbLN98UhsAzxMgTNVEsezIirEVXFttFp7EhJ7Vzlsifrrs2dZWlk
0DuA7AXQYuMp2t5OeXSZvkQUiok8Rmj9S89OI5o8fan2o043MeM6HdoESp48z/VDnGBTEN1Ti1JS
/5t1tSN6SzhVf/gxhCi/ZRZ4T9KB+YY8b4M2vu9RPI6uBoj9FqKczd/g3/zfaZ7WhThLNCZCa1Hh
YEqB0YBZvXX//Yby2bJlq7muRuydh9gwirYrKgW3MTh/Xp2LlI5GhegkgybRi0SxiYm55K2o+H1y
XukD0be228FR3tv0slQ3H1ieo5t/NpH3ZrW/nB++RE/zyNQJgtuCPhVhCjXAlg+FRPvDHXNPEzaK
Vs4V/TJZP1MtFqpGtN8OE0ut//n1oEjqKCIMrsOlwTX2K82wfAGIRTcAZR/ZK5fCO8tXUrldLovd
s8Yg0/6JsUp9D6+EJKssKjb0DqSO5W+I+8jnKL7a+Ge4c3X3bgDBFVxSjDLbuQzCSF4JE1csW50g
C7M/r88txNFTkXn8QY99kbj7CPqEnOWXhR+wfTfFJxhvM+pxb8X+L+JNZg3zifIvREnpsmCG1dcg
6DJJz/d6RKeQz084aNKqRnY4ZjtXyUBEgNbnWXMEys60VQAuodqVWI8pTDOGkGrmuo1xUMt2U8vY
WE0Kxt2CLWjXd9UaYGobzlfNmFQ4cDAA225vZ95Cu9TIvQuLuZ3QKWYqYhV5VQtnjz4qPeGcsbzd
pKD+X7jjQ+b7nKNIf38VgPFJq5EpeZWikLTwT68xZlFtBadwSQXP/TpDYgRErz4vpcu7M4oZ9EiH
CLmYFCY0tcUH5cepiSa/zPHDb4sAY+bm0THGqqOvPFzubxVBnCFyLIcqe5c2LhVBlD6B/0hIFg9O
1i8/CxKvQcWVVA+knPVn7XvRUMMlv+eoDad0Y7LooY+qo7fUYdz6I+Hv7D+PVR0dwFV3Gqt1/QBB
nkVGJ35E4SQnhJVEparwrG2v+5Mfzz2LPZR4HQzAC6IwD3yHnqFHgNNcOgKi4BLJGn3JQoUa1Ikx
i691OafJFD9/sYlYhp1hHioKDv9/U67WUa9i/ZDR8fmGc5UVe1rTjHmW/Yl287RhZX+T9hcfrfBU
uJQ/CgzzJjAAvzjyxZ3KVKyJrfEq5vEayJfg1rug7QUefVyFRdTNSN6N4Ekgi6chD/ji8yPO0cpJ
ldTx7C0Em5QI6t0MdayXs3FDmHgqLnIEwJXYDujh6L0luKKiMk80QZvYlTjJ0BgAFKKXJtwSK39W
32sDDkfZX80OtqGWTA8UyReHNfAwmLPtMTp1EhX89Gh2kmXxo0WQvLjtf63cOdx24ZZDQyCrx0Yq
tLR2lwMv+pJyh/AgNWKnAkxyYTc/QCV6J6RGqw3eYAyRXR+6iyz84UIbNi0xSSGkDHNbfixtJctC
fjU8zZ9Htm+WfY9lr4HcJ2eBHQaZE3bFQdlFFTp1V5djy74QybGyvEqnaw3CJNtk2aUok3YEL0Yi
PdsWeuLyEw8+w/nFztDivewqgu0GjSdOoNncTutA73si6klim1GSsYPYoilevU3Rvx5giOnqfkOh
dkY1Wao5wbTZp4GNzRJlmjWvLtnLAhcIt/d0rVvwI7AjoagxUFQd9UqKoz0NkhV1/hPe6ih1+dWl
OJz0xo44zpNovU/R1u/yGC0+BrB02WiMEWbn7L6Xxfb6BaEAmSI8O0G8H8FqPXqbSwZTZSYp1D/L
V0B8eYvwT9iQIxGpzguhoGEYWEN9/d+d80GJtQieKCGiK9P2Zylex9XqFmPyuYRjku6NtRNZlACq
APLhKhBtoCEKxNogziV+v4cbwN8nPZjCw0nPDYm1Frxxn1lvJecwGbTL/gKIQ0hsDAVWWVkbpsdh
Kh5bUoiQuvhee0idetq8/cWMPgdDy5yCSfN0Eb8Ql3m3ytyChBmrNm/7xuQ0udYtylA5dbnitYKb
+BqdkuY2uvJRbzfGz7pj1+cGgCWUGwKRdLurbZ71nLEeajKVK0iN6DVpBGdK5GqMB5dMYc/yP8X1
1J/A8o/xVap4v30UYnOD52g0P8RKYzhCQaXsRb/SFHgUpdn+uUvhOwL8lqcx7KQATwiR+WNImYze
zVXXFoi8nzQbWHK8HR4G7q8p5yGGPwuJJAulVzn1LDl8Cshbx1Kjysc++RmDvfUBVdF6U/fEJzaz
u/sq9dv/8A4w8PMH25y5Z31ZfOsrhbsdOdrTkaF/pZcDvyOKubRT/sG6rQo2BrwLcco1ADt/7EdP
+W7Yv+AjoZx9ZBJ+hJB/HPGx4jKDOEL5qzpy3CpZFy2D3b62mLiACOopp3aFCdPlZll+OTIysx+H
ynIVRsTAXi9eoVBLGIydvqzJk5N5wkzQtzI8OQGfAKaREaaxU+hviOBPrNJPIbxt2ASVIsqMKuHo
APXZpOXcjFJaVwkbSHyYuYBKOSi4KbIhM/54gC3yQY5q1oaF48NgZT7M7EFyDOZp3w4fn+OuKzGX
p5riDFtK689kIcfqRGlFHklCsh5TUuRr1bOCg+8RVDBf1wXIKlbZ7lDQOehjCdkZ+a7ekTKyr2X/
mjnQnErjV+S6sKiEW+lE6o/SZPabd33LfulhnpUSu0z/cPbCqpJTz6geTOvsmOxejKoNlqm94DLA
9glPYBEljCQvAgs/5CYY31vmopvsEyuiDkkEM1tVX0E2UdCqah+t5gXGWeKPJll9YlkQciyeIiU4
TXTdHX8oaxWXqgR6wqGuiEqIGG+H6y4GXcIWgi2eJOj+5LD/FW/Jx6YvWILfh3KcovuFG7GyjV4/
b/Fai4OPyKoKTmfxjeaiXPjbDdV8F/8/sz3sdb15FdV0LCzKBRsmThoIQUXkYHGwxBZULIFRVx/o
6IaTSgPSRwKslaVxcWcVmwN4Jq4TxiRbDmN8zO61Q3MyUHUTBzkwc11K4K5hzisGou/VMt2LEyoE
uatw8DKTtJ5VGyAQqL5BUpdHnQsnGtoBWgtDDPucZqNNlGjdIL4jzKnLui8i4+FYbILewAh50/WH
EsyYA3iuScgZRom0Ii2Q9k7UEOBZqVdSlD5BaohSdzSPg+3qxCQuVec/NG4ulLNaFrCcG0GRvJPy
/CcF0iAcLwhVjSXdmm4rCmDCZb0iSJiU9U50auGnW8jLPb++8ot+jeKkktDCMY+Wv6ZKG4vuCmxV
FEtWr9qHgw7A3qTDvW03oaFEJKPappo4tIYXzj+5ecwlenAvlTueFjPXBYA8+Dm4RyFHWEAAMESa
RAg084OtUStysXtgbhqMeFbW84uftNT5N2ZUeAgsQ1kfPMBvUbj1u7HbSvxe7r/ThV/xP5xLRB0H
LLnwvTa+daAaYxcKGD4mhbDWxHCG+7+SF9xZ1hbkL4xVXoe5xhcnfu7le+osxwAq9LBg6QevXaPA
rVkeO4k8KHua45dGxIJERPgsSleTecDnPaY0GY6nA5aNlSGROlr+4vbnI2LzTdaq8zMB2CrOHLyI
wKKRBMvJacawGLcEQ3qKtnYSugm0qvm7SDgll/t63G94tDQefeiNJsdcYOxtIa6X+2kkJw5QozOI
+zLkrgtlJnRrPP+2kslwm876hQmbGMw30WM8jvc3xzt/43JKFHmHSr3eFbQ8yiVACltJ9z0dJaTe
T6sMNFr+ocddVtvB7/iFcYs6CwMiDV8VYekAk4Lysxqjpj8LrunXPhmfBfBZkoGPCfXL/UqSIE8k
3eEGrb3kaUxTHzs4cySqdXtH/1fEeTdgaqmJqLEdGIdX/myKZHjQ5VXofd+Iznl56jZgB59xw1vF
Xc7S9jlstpYtOnz47g3/Ppotaam15OagUsQEaRa0eN8ViT8PYOkNajNIFcJ1Xixlj3BIYqlsvZz5
ozsZfvTkEHcIo1UtOrKobVEKtfIUecI6ji5ZGg9DusMfP+GWk+z+5VhPzz9xFfRr2VbwNKjOU/sz
zQ93t/uUJ7K4f4xMGKTZTvY4NRJ2WyHNhVR+6vyEjlYXb47MYjf0zOyULIUuzE6B8cFGsa2b6sAR
RUJ8UEXXy6LJ0MRmKDwzjADCnS7ei0UtVEM9DPyUVzh8lW7oYQ+wfpwgXJGEzsp+eiKxFhtYgVc/
IRE72ayMBEB8Un7I9+W2AGC/jw2BoBRiUre+bS6jZfLjeSoS1YzA+EDYJLfiVRPhXLeCb+o3OZLa
gASg2VTCCg1JlOvZTXJA0/Q3kFJ2/3fwWhFHdjTRLnnuFKLM29IlSEwIEpn6SojmzgD3aI9BhiKW
tiseRcsKf93cET4/jaj3p1SMqG/N7Bi7Z5qW6u5ywfdk9Eu5tI2N9b0YGe13e0Hx0QVWdckiccz0
ZeVOOArH15x2wOYSymYCFYjnb9JweK/NtLC/VLDzEwAl9TalZLLCZACsFAA062QNe9eludQgkSqX
Yq+ABbzIrcp+MDfGst3wPLUdDQwkNySPjwelb1ZVeuYRSf0oe5ZAg+S9ZGq6Vrg/xu9gsQ49qvWH
KfN86zpgcgJ+XOz5qzAreiDueo/sU2dO1dzP3wBKahvBWcy1vzd1H73YrVtrdG1VZvDjK5ELNd0k
SzQ06ZFDprLYzywFVYJcxEjBcQPn4fvwmawo8DJ28Yp2wmp71KdVJklv3MzWdLH2kiCDrL0KoP1V
aFNKTbaY45OGScDFpNFX0MwB1uzzsIyTG/m6PQxI4gIDJdx11+vdl3i16Z/ohSTRh0+nbecStnhp
M6+iMq5n+MhlKtEtVbeDNowRgNk7DKHeUV4LZU433og6t1l4GTiaLgDnZUIVCzPt+rPoGh8XHvSa
Jmegw1ELw3p5zTKDi7s2m0Ce3rKopMiN9f0yblpqS0Q5/1sOw02Z1YGjSWBeMgS6clAC7sZq5G/T
BmRiNnlGQmKZV5d22IjbWoH1QLPWUWcv4PNDfNPivyFsOmZMghZMxbMhtoPUOaIEnik6plsFTx+D
G01e7JSGQLGm1/EiXtq/zIzjRQ20+/g1ZROqdhtwVAmROXUVBp2fU7d5iMMZI43QiKHlXDylOw5b
/1VQlouwRt4A3ZCeg9Lv8f85AYe0XEyoikFuSnRAK5GXgzF81X9EyXIuYIRnYjTdvB9oPnaVAJLL
3/Fp1nfXB/su+Qyxn7WuBZXotQvYGzP+G7qIp9SGJcHaOw3lmqq0or8wricj4nvUNgqOLBgKTq+/
Kgfa5Rf5Xh5W6jj0f6cp6Y2Xrdl8jxE0HF3a0jXcHdKnQ3xMyaArNRpJaXsUl3fAroujWePHti2T
Xz6/t5/RvJqwcSaLaH4loS6V1pf7LfSOFTtSvhua6+O+tc2x2HUW9sJdjTJwvNtVv5/DeUHKiUrS
ZcYFzNsG5RxWKgWxG8RZYdBevEsPEGQWPEyXw6V4hiFE5pVckMP9sf9Tra6RpCpd1xsu38y/6ooG
Wd0/w5VC2rdm6Cw6wsOChPYvFTURHD/BNn/rz5sSdDwE35coQvW0JJHSHttQ+Mgo10Ehj74I2QXM
zqxNeqWDOrfFyhTvCObnDhBrQgd1LJDuXELp7bbw/CvFZ1TXl4yR/H1AqtJ8ofrtJT3x+SU2t2gR
29nFwBJQao30lbYARGRIgs56LQLIjVkHCt6RZE5dmbNgF8o43BcUbOnEicoJvmtMANlJTW/B/q9a
sH4V870mpwPCYBSd/xecnkjeRlAGUXm3PLb8+aKJ4E4OQ7553upl8BWYnymYT0rt0xXh7R2Z5yyP
cVBSpoeMFrqcGvwbDFeuBdVI+B6FJgN4sm8R3ih5lhyD4FP9nH85PIfSnOfDxnZYNCvYKCtoUsP5
rySIq69oGXwec2d9YwLAmGFD5Xl0CMialfZzx26uvwDlm1R6oVvkcosVMPgRUPIn2aV0Cn7nuYkh
SheGCv0h09jq3FF0xCUfYHOKWR/8BNeo3IoG41CXVkLve0sl+WMxnIom2MlYJ5VfBd7zC6VxhFzT
VW3EEUsgsFYC9Mbdmprm5NKHnIFCXUYtMFvOHHWlrc/8+mrAtFMPNtGg/SDZxeig0TovvD0IRgUS
2cqGXfBnKW5VMcVhdaWDl9JoXBH55d6KjLhjmdZYwjoD8rhKoKMHG6jxzg5Yf9EZlSDzvOLOnGzQ
EzDoTSYmcw1KauYNVlUQnb1YNkQ1ln7dtyBClBQQC1NLBhRnbON9eX1AgWStF2IGIL6EuLHs3vnj
FeW88Lc14ZjTNWq0Gpj5V+Bax3FkonH8xzziUiNbWSaeL2XZIsimGo5rq7hzJ+eXR/sDFPp/1DcQ
kMsMNTSzSGOPouWPgdLUPjBmgfHC2zVagbGFb6AOGAOiXA0yP56Cwl93zXKuv/li9s5qxN8/dCdD
rkc4zl7KFUmnp27FKQtZQCcPVXIJfHtYl9ZqEKGue+k/SqIY86pe+2FIQqF633ki/bn8vWjfmWnC
wVoeb43OnLx8CKsxZg+z1cYqcaseA4IUTGIXYApLuFN0SV8MlsWsNx+fxNCiuztaqrNp5LRyJ5of
V/q5r+Pq84pIxVoFiQhYijVNSH9Gl/XgLGzqm7DITI86YQXH5MzPLBYZSYuqbln9XEmEoZ67MqZl
qV+4tKUxEEWDivRdGuYXCTVkJKB07Om3bA6ewkxpxpRvAaQKwtVT/LT2iQddPk7p/XDoQbmgBX2H
tQhW4J1zEU59ZYL5BHMKgnttib0kHyVrPgFLVK6HlqKr25iH15G3oeE3QBfItKLS8fDUa/KXPImq
+lwEIWAqIEbooUVh4AKkXG7oLjeMYjaKVdlodJGNGSgGruVNGSPyxnt+RLB/zFwuJ9MLxO7dbJbH
WDT9FgP/UzkYg4T71nWij80So297Oc128/ha0Ly2vXFyQQvjGVUhuNZlRgKQ+PaaP82hFtyBcIQ0
rH/eedUKM2eQ0iAFDCN0U4/n8oZjLu8Bqj9KmzvyUNNMLzwN6PbI80VQGCRMpl9v2VNhbUQ2fZ8f
wMvDKFhnSYCGBgWXV23FiPdA+ggfOyibS7nsvGgQfvmiEhr4UGddfswBqRTLBY0i5EqCppehvrLQ
8U8H9/+0sPRLBPqjThYtau6KQkKBOwWKPnpvFMmql2WbuzT7wB4UTTy9cIvisDwaz9LA0Lgwq+Fv
swpTBDPw7cE5KA8+/TY8mPCDbvpdcNFJodXENemzYmmLZv/ylalliPNM1ASJ9IYoImsjz/oFNTgI
tmy7m7Wz4zc82JQa2W4Pn0o8FxOp2Fy97P5IjTReByonKMPgy40/n7BMEnB0PKFHE7H6+8j4Cl6q
mYFZbWzyJo7pxIM1VywmteZiguUDzhwc3izao8K1Y41paMMMpR0JMmjGEHrM4AhRlVHCvQ+cmtoI
vfDuQoyGtBLLFhq3VNCN5+dRLMJTEOZLpiC+cjupJ0rYfQvK8Lvpe3cYduW7qiJk3CqFoUktJIrf
+/VFxTkKMsEqS45htxrmGsAPK6p2aTPUgCZ+LU0nqW1cPJU9Jkw14VPwrHkcuF2KRktllA5rB3yo
gB7pFgjEC8TcR039N1cuxvVp6ekNLNnM5YLn0D9bD0RiJ0kWNMxhYZ89ve91jd6Nj9jCngCA1VKf
o76LEU6lGlezUvGdwETKBXCo+H0WrFZXYjp4SjL8vI2whVrRIA4kMvGQP+rQ+gHRf7B0f1G2W/Ry
ils74uRQWgDrF1jrW/NmUyxPldTO24g47ZiJYT6liOFnYTfAbixpNgTxWaQMVBHLYsvBec1QTOy0
PAeMKwpAE8n+nIxnigCVdyCY48mJL8SVUXjuJzO8VuM9zdRob5A35iyINpw2n0y9Mili3MCGQ26n
vFei76SerNMIpi0UX/k5N+HdtLmzRAsJeFqZmn0cfS8UztcOb6p/cSTYGh/aR8OYf0tU+UURa4Zy
/prhOJAMstRz2ddR0Mn484dyRcGj2+3SBnOEXqAwdjeU8q7FFc8HoI8dT5VNr2Rw9xv265es9+/6
J9pf5EvYylZhtNfU9gsztNR3eg+r+UCK+ZerUf24FDsShMdPzJN2ZtySbOE6HYl707u1d//RbVIv
DWewjctIToSgCB+aaDtHD5Os01ckjSx9DRaZbALrh5lKIlkTqwei55VN06d2DOJj5diprfe/1YFQ
IHAAkChkD9/3ouc1TG6+UfD99DDu0BCkmCgm37nJAioX5SLwI22SJNVjr6IRzC2vZkXkHEr7DKa+
as9zOwUjro13xgDpka00pGkCMAUWpvd664lf2FD46Vk/kq/mXlZqoTxDN8f7CgVOC9gL7XmpyoOf
XMTyopqKSS0INHZ9qdtYc/aGJaeyxJucmrXqPo8EyRHb7cgprik2mJpLGX2+WT19wCYBO18/IDOA
FwDgQjzg1wkmpEb4JXNIznnEKpoy5TTQDLG6w36KkI0fmzi6XdqIfnCwb1hQWzxMMr2xPTinUhw/
QDjIibPT64izX/iEGZRFTLElpd6Js648uzcznbmJDFp+FY7Qj1BzEgxffjPGJzkDtowNWI4673bg
GVlvwrw/ZBj3z6InrHcNkkMPyZRAPS+PirGmagBsFll0yC50ud2JPZT1aFiBlaY7u1Nrcy2YDUcg
7xeRaCXLKuETtrZ2x45JSbEf+cQrqr2cI8eCO60fDZ8165zjj7JTf6k+DDohFhRFGs16T6bYVYOG
LScd9396VO19suWpMiqqMs4cc2TOXykgJj7xlPBD5XMKwx+5WCQWO4uzqjWhMaHYFDmTsBl4sg2R
3dfBFeuS3PiEpfGnwFlHBQoYsZgxZMEf6mvprpp+E0xYjxkjEDYuLcme8/c3VIdt3Nt9YEhXZdQJ
BKzHDXfYbS3njTXw+YucUqJWwwLjw1wZo3W6O2cqR96ND05y1hORQbZmJZ5XyrEr2dfhjFlOLtlb
XuCiyWll5HUV+azXOJTGpxxTcp6qari4cmkjaYOBBcS3NybCN6gCVqEXEpss/mLX9t1428xp4vDD
DwdaqXCAzwSiQstm6J4umGj0KA4vqPhIlhZTX3KEE352RYIpC9lGvpU6XZ2kjqVd0TzLidpaM6uY
8tP6dc9RQsjqhRX7McDUCO1nibR81XMz21YukQi1UTIAI6LlT6E6DMlCeqLa9DCrYiqPdtrqAFzN
EUtUZgUUE92lymGanBpgKGJ2gyuxevGt4ae4c7wMSm+06/JHvB6WKBk11keP2JuBZmIuy47W4BaS
Lo+mSR+DDWZh0MRDf3jb7abOrFHGB2vtgBlc/HrH8ZKhzIG61EhHOUsTjlnMk8ZpiDW1qM8+w9u9
QHRs0Idnzvq4/r6ozVGkpoS48DF4ZraIJtOumXKhhyJRle+uRb1e6GhtV6vITbvayZn2G4iEtb2r
oMW3sQK3Nm70uRtjt2K993GN56x/XW+MU6T82ZJJ2FKUBn+y7nSTeTSOqcQuHrkjPsnj/E3x5FoO
gkPq3+qy4VWyPCFnIY8bE5Fn6rG8XPVTf4A5AlcI22Ha9UvYmMh8uT8t3dDS1wYBNmbq4gUnAIY4
AFZQ9CGixUOZIi70Hl58rzhdcIxuZ504LoWMuqSeVDrkxWKoxroeuWg566rPTbn8+UErNPOYER6l
ut6rnRbd8wNYom1KDWN5TXaNaqEoS1/mKxQJclJPutdrCQWdfq99I7SLe1vyes6bhjqxLv0r7pUu
3yyIeeuyrklHtwD/z2eTHjNzH22hh/gMJ3404Ikq1iTUs7ScUEVw4wgYIVtdVwNdiFAXo1SHky7Y
TWTpZ/W4GXXheJkR7c1bcoMvxMHrk15lUkCG/qCksIOj9aqz2M6t/cXqJvbjdcOT0kG7snWWnrrv
5o2+khkybIqrqKmlrHF7/gMhKyBMrD3qHlZpe1aD73Y0CvP10q+CvclgQKW8xe+6VwRPEzKf+Dv/
GJEqztRAOXAuCHUYATRobt90dy5kVORIWajXOpzH+7GDrRUrq69tz4MOOd5DdxJAOk+KpF/SmVgk
IvbLz0C1810cJdR/8Ny0oq5ruqKzRszSerBRrExycT07ZNYHAu+bYLQSC7dO640fP6JVSo2Chm+r
ExBXEajE/COzUJpSthwfLjhpUNdIw7LZuVKhq9fGaQ0/xWbieQSQOwIzlw01DGz1MrNTXdRj+4uM
YPlNpKDCuqU/FO9U/tSFvnc6eYkJ13LFt0zZsqe9QRMlPgqzFdjX8Pi+adghY7cXqBeRv+Qh543H
4R7jjJm0iHPFKzPrKubNNtindbAipmPpzJkl+LEVRca5RAcXjRKCgoWSBlHhcJ2AxRlSBn+U8O3F
d9HrjmdAHZ89iVdGho0384uCrbzE9tvG7Mo8avupIzKtiCd4NqMOF2zRaF3bgHLqCUMWrv3SrA0z
hWO47woQ2+YfKHtT5PTcHH9XAFneYLPG7YgVve1fz2VgoAjtUN4HnI/GNauKdF4gMxkFT4YUG91x
4KTiidsi/HOFI2E8kepez3q6YlRHpdJz+OYFuoZiBkJNhaQiyhDSuA4Z2g0iAmex7FYbZDk88wqi
UaqpDYW0w+FQ2Jod4t9U3Olh7s4f/QVvvpZumC5iejqwqGtJXCht/9sAcIOVaTvNbkJk0oQMlBzn
LywUJXINgSvbr+mL32LGVXu1Shrkx1KF8i1V82zpfFVEx7miq63ONkiHc94bbeksa9HTqTuZlmy0
rEQaODAtV5x2LM/CZW7rRpH7JrlM7gQK7q0qNm9eRZ7AV+Qhl8cVMyULPZpeIqK6dWyIOAPaAyte
4Jp/0yNrOmELb4qhLWAFAakiv+EH8JUlGv5coqH4bb/gyFBQD28bsfVsq0bFE4zjU6p4DBVyWFnv
oyfegFOzjbL6SMXDvABxsOZGovOOY4j/gry636pRgMyCDWExjbQAggJmv+5AULgW9rUp3OCOeZFC
QfVOnUUhIKkPATlI/DsSo48H6/11jM4dUIwcVgNCreCWJLhPcWqMs+3VChALHqYyOdRoWYT9zd43
d8ahszq6cxzUnx7zU5W+yP5V267GwTyvXZhrkILW59TQJP1objtqWKGd3adl+aizUQnL4I/HBdSM
H+G9R90JfxakVGXafohyKeXxOXcEbDbsFWgXd2xA768aJqhdKMpiruKeZJQI20+d3Odr+Orbbreb
K5Rrn1ZQprtMFSJdzKTi1NdoSbl5FFJoak6Fe7tK92gSx+kTscBRdm6zBliAiN6wWfNAj9xpVIhI
xSdHYfFf4dXRUvx0xh/ji7KEKMYruL0nCl9T0tU08B/bz+o7hX6u1uj7OnLA0m/DKEOoMGQYMQiM
/9S2g7OD01T12zUh82HLROIQyhQrzHg394+xSd3NHA6mOioGDg+OGH+KR6Ok3bcMGedlYQL0SIPm
ynV4nQAy0qV1x7F2PD8CbnRzWfMjkcGydkDky2MvtvjsvuaS0t+oTDPostx8EnOpNWLwWpjnqNHX
T2jDZOtRLk76c+mISXaw9BQyrNNNntM7zfRYj0ABcsVwejfbFEDKmWz8qvC9uWX7wb/BCDNNW42Z
hRscrMrFtAbJbODtaKpDbH+pXQhuAbG/SMaTj7UTsiYbEwIa6aXvn0EH42/eqFrLNTDKoWP/KtdJ
0LWmwuTAwHPguO4ziEyWEdNFkrT7DrRElKuA9TbvjjkNCOL2qwEyZf/mWG9ue95ku9Gad0diFPeC
lU1o4DlAXVM1kKDdYUHUiPd37OzcDIqggU/mQ3kJmgH0+KQ8NHR4QsXi+CfRc5U75z6R8jA1S3xb
yJVVaHG8aYR8sX7+mLFaVMOprFcR/hLce6YWp67asCua7EM9Pz/q6z500qHwod+DX80Ouy9XFsZY
cEnLAqFXMjcAlG55txUJ+7lJM881ZwxjFHiQHDB00pljrhsD+5yigqDr+iVtpRZEqlho2i1WAd8N
mt1bg2jxL+8L+NbJTXlxx3Yp09PP8EgqIHCwc/DRIh6ONdVEEsSYZ2vx9sdD7NQ+muPPvNDh6ZW4
AcEfrYmCos2pj/XGJ/wlmqw102R8QxrGDPN4xvBTMGb2z0EJh+JByiEGeOL5SZkX+KR8AzyWF7Da
odwfLNzyeNMnGJ/8xgORmVpy8EbccnK5mWCRE0A2KXJ2Ene4tcBKh6XRk1/w3S7qcvORN3YNNPR3
Osw71tLz9EeXFRp7NvhV9kUIAkyjC2DdTvH2nB0ufvdw3V92Lsz1pz+KoL+zu3Avym9xKdIX966h
9xRnJtlMzvPduYtagQuvvrx1gU90fvUtBo23B6U75DDUDGH0gy6tZ4NRcMtHLzaCgOx2DszqdDuJ
M6fLiyw0WjE1Wkqt9qyGjDFTOeiKITLGPc0etbmfvsLP+th3ZU1sdR7UjKkooOMbfMB8XNlPYI6C
jOwYNDqT52izRqTQh1ayDXTI6DZ8BRJL7SdwZp6rtInp7RwTqBJkON6esDMwjQINOO6SOXEJkF2e
5k+X3gUHGynWc1qZ9m0KgOFkhzHPX9Oyi1OsFff82Ir/ZyYYbNzf63odkS5FbnRJtUcG3itHxr8G
lf1EHTyW6SADekRPFmvOOyRCrZTvniuOIX1RUchH0/xpzVL42FXKYghVzMUpmJgTJZzl6rCaUuGl
ojl0FKutbyzjad+FM0GBlMyqMAYjoVeuug+20/pOhomWpMhNeZkkHVLekQZv66mIGTDU2kVfk41q
UpztIlnHd2RzsHxkHFgdvmGNerYYtMTeczIytY6oYsSapNtRZ9MfhQe8wiv5J9TlefPvFUe7rOR7
hf61V6RMSMFX9hlxBO91QU6x/h5TrYt0CS1sEwtuk/3NluHr/9SvJ+HxqsraIz4ohIpFq1B0IzTD
GeFXsjlc590PstF5GBrP5pO0Ubat8dbECA9shiHcRowyW1sEzf4csS4kcAed4p2Xzknrd7N7L4dJ
HdfhVpt966V7wi3wr4gh/+14xbzksVlrwaWfPeRfUMeHwd8dXs1pwTlA7po5QVvf//1ZiTe37xGs
0a5MgfqAmJZIaoDtPOu6vhsYv1ph9eq/w6DNDRh+qeZDu1kJI3d406K0ZeMktj4w5qR8ATxLsjdt
urp+9trDpRMOKyhMlv1cwZsaGED2OfdRGuoqO+PQDhuAtq42pMYnO/9gPZi4aXIeKEpzELntI7+8
h+/d4UAkpWHZwWQg4ANual/HDmQWwkVkx3XikcXbgA+dGpI/fDdhb2eNGTuamczR4h/9VNPvxzCl
ScADDTIgY5VaXrpQkx5pSFiQdurARQtP0eoksuK4VTOQfMBvvP2J/awbDWLEmxczPY3u69QZ4YDH
Ej1EGWX8ZzL4nIIwmoAVN8lEqqb+uY5UwnCad3rS/vfOEtnZxeaY0vsDS9burPPt7fNmbGOZ94mI
2MpDhgQ1vkjX2FumEvd9gp5LwMS02QFbe2jIFYtUWl+a51/zL5pvF14dOM+teGQQ+yingfoalpYS
bRoFazxSIxDCBiNoyoIKsywocLU5JSK+KOwesb1zPvjccJltQUclj8ztpNXzmadhGYBS99gVxE8i
URzTD+5bZHISP7p0Xq96v/TI7X58ekL/ylqF2c5wR7So7ZEHMp9cUsvCKR7GotevPT7rKuIBdu72
Wkq6+pK0/GQ/P4mbeX7L6KphSVrdqGAieBy/Pwf7N5c96fDGj0g5J0zABcSbIO74TIujf40+dEcT
ONJM7YI8A7oHXOMDPIaLfrATMbVxO83+RBweZY52Bvx6k21cyHGKGkksKSaG8juQKL6cX1oq1eeX
WPI0akhJLPyOuxv36YXFqe5PD4JQK2l0hL9fZUnLk9zfLws9lDzi0tqNiLssKPnrrLhsHw/u1HSi
orduVA/6PWE4uI0pgeXJAboLH7pzU84BA1xpB1UKQ38pqsssp2MbiGX/UoS5ZxXtM7XWhFdsY41j
zEn9idgd8pyF9d4k/JjDh0POU/Qyus+9Y0zZKbj5G19tv/ySw8xJLMdxcmwkBaesflsSaTWLBFVB
CGlo9e/vNxksgthelsjgJT3KdLWju3w9glrAO938/afXqfHY8HCNK3p/m7y/rboZShirN53QCt36
ujrHWbGZe0SxChCiv5chYq48uV/fSy7wxddHQaTPi3rmPLBnq/8DwtujmGGT6+eiGTCeHVa+yPqu
GLIz2qQ70aXq+Hv6Y2V6suHbD/sfbUqGEWgGgTilnqrtkie9ySSMjux/DkZ+zSeNAHVhib2BLTI/
jCkyw4MZDKou35GMYvgICmzkoNNbtpjrEtEh0djiMx7j+A4Ul3nuL1qrU2nC3uoLEFgyexaw/Ah8
iApAT+r2xus4LU/3pieX/MdRSU4QYDDFhjs36NPEmZ8CIoKJN3dGhsNNTZkoIZhdKwkaJ7e2Gwq9
kYy6Ueesvq+vFKDP0YhvGKQzqAHAueSrjIZ7g8JP/iNU+p+wr0Rqe/iIaj7UduuRi22BdY1Bx3s9
+p8/ShiW8yRuEs6Zhn7+fiVrioC06k0F9Bf2xHKaDeduDaFFmk7UIfFxQY3WTE8vfDiLHEQR9GA3
6+bG33ynEaNuCTcrQ69EPaXk1OGZjO5CRUHcTPjabr8d2efPL12LvXETAQMHD7J5XtLZuPnWVNfk
ugA9FmtRX6W19IInLfJQjIJgpmFQSdCrdOVheDI3a6O6333qrGg0RRUjTdb8j37A0TaBrqrrWD2H
XRhhuO/9/tejW/x5LHySWQ6JQSP/5XT8Q+YQfUQ46k5ytgEirqicJsv/nSvM3SOIrScFKLcPmV9u
MPcWC4VVptVFz22JaIBJb6ru925okscMHD2kNmnHRabMEs9gNH0c0JkLUIH/tx/o46SS/S7OBRfp
rJJfg40o97oX/7aTUcF5XHW01EIqYBVHBXgfnxQnDA4N2bC655gjcZue18QhD0sSy7OLbxD0z27W
8SNFtSVx4KmpTvmtGcbEewDNGiWqrCiWlLVPoMAtn0N2u9zDrLd1Slmy65NM7kdzn18CEoPGMQgi
SbJsD0CmOjo1tO0+p9eDj09hiGGzsPDWhNIqs8aqWlAzvsYpgx5sciwIDlbjWmIiaAVJ+vqtASDg
b3P4UunwJBuzhXnWMUJOWZuedlFI5BY2QwuBa+YlxWa2nWdhniGdtXLoMc6heTW20mrtAZ1nySOU
NC2pG1z9Wc2GgcE6Co7ivfpU6N0PGADlCoNRe6ff74J4hSqb7TtQ88yt0UbEyAaaqnPDJd/3thY8
KVhsDCXaruP0Mk4uyO61YSAX75qwKKeehNmkxTeCSNg4FWMEsaMTF5yUgUl8zZQNMu5Xj7efuI8b
hTkhWeeTNbP4jsv+mt3U33s+Q6nN1KY8vv/bJRCSDpEtN3qtqBjcFEh4VeQYw0m8ZKoORmtYnSsh
ttH6Bz40S1ht5giCOau2OZohbVOehsveKd8gkaz0kmhFslm7B20CymRF8jUFjZX6jpuSGmw7dPzP
H08AlsXa4D1Lqjmy2fl57Wc+SmIWSEYZXm74cS3Qz3pYCrK599i/oMUrZWzNlTFJUEk+4RlEzQPO
r5flczkGespTZI5HHBqIUU42Z0ph+/Zt35ZXUmFqdD4+JYv+45cPKNlrdz9CjkWQunQPcB6wAZ78
lILxHYVWnM6MXJdRRPiAlnWbexRwaSIucVMUBN7vWBIlyUajAkOYZJVaUn49rpz9zjSO8LUDpARE
E2KAK3K/r1pyQtRuMklEj3LKJfjtNaSRNLBgNcCzAgWYLVllZkupWLfesqnjOepqxSVKqrT7JbuM
Sd95TyUusG/WLPu4uHDSgps6thMUl1Jjnm+CEb88aEgK9u9TpPhdqxkSMfFeqkGOt6nj3io6Uznd
FT4ZU+bv51ziq72VYtnGVx65fJVDw/HF2AOrcg5oJ+95ca5mALpCjo+/YXWQqvVEd1Q5KUafoech
Q9OLNejzl8lSM1AJpWcBH+sWRxu9lezEsBCz0gICXD0EXmR1Lh9q7vh1KyOu+gupq1YnoQyiFiQd
1hY0Sk23bktM8I4KQ12e723yNALQq5TZ86JjKJ0h7ZMUWudaZ42xqk9PGAfC227jJm/t+AIgQvVT
nGNmOWdEU5E/hZ1v3ks7BnGnNFIzGk2BAzsU2UBhOIpAfd5oeidb/Lfb58cI6ikQPnlTi/t4NJmv
rc98UVlkUmc6TTHbHcAJiSrdp3C0M2Qvrlfhephd+GCCROAN59ydZIGQNgtN4FhAbcENn3kqZhHp
g9WxSUnApZuvho4Jv1mPEYFQlnV2MZaKa6bnnwrgGBG38g9fJiM0WNyq1NcaKQac+YrtT1HWW+k+
2j9+4MB/s7jvVmQ0eHRqALjLQKAViz75WTrqV19I4oVSCJtVuL0l/7/jVdSUsOsH4/Zt9WrIQNAj
GIK7kUDBjY71JMOZkCxQhcFluCHJVoy4DpfftYGewhcNHJ8z5dHsM7CHkvEwU47+AzSKjj3AiE+/
8EiYGyvCaIbBazcNCTRgs9tCJtttRCF1HzK214mlLjdXYNp9co/BPjWPcjhuWjjJ288ZxiZ2m8IA
f21QgUCDVUc4fIHc+O4QrFdL6s9YU+pefFn0GXCRy5IkBtrH+1eIsWuX2Zah0az2O1tLCM6p+CZy
Z6UhMaQbXsy3CYAVNqQCvhbJYurP2MG9QRoq0P/uvm0ZdpdNwYKZn3XI5QQnmRUKYwo6YHx17xMa
DC8ZLR7U6jAAnYgYj8cgPgulA2mfVO94CFUFoyYhZCaOaXHbMS9ITcBNgzBvmjb/1V2DvZuuVpzv
JZXKlNA6Oslce1ltIVvfdPlpGrCRx3vJoWU6x1bHi+Cp/JqRdGmT3txKbiQjCAkLNmqOIqqEKv40
++Mjc4NX88m85YxmrATb4Unlyo0YgQuVxtA5mLaiawMMMKX9HHy37mOnae/pmcwzShEopygtZOZw
bl9gYq3RPGtkM3TlYr1Ugct3xAMbcAOysqh6BxRynkyFVLafHh2KF/paw+Y03WTb9hp6+rjLh7wM
YSE76L1zAHTsv0Dtzgyigl4JOp+5SdZhAKL0WUBTRh6U5zz+GCBO8YqGsXxe7wAs2nBTMt+ArOl0
YPFbNsMYSM1gmucuAaachRln1F27ZBmN02Ixl7fiOZOQgQyIQ04cFHAJcryxS05AjAP4ptOWGKLP
ntM4s+sXJvfza1GXZoSHcrYqn5UHgegQUCwJ+oD3ATSjdnAmMcAZfu5Ha30R+ohqRQY/g1JgmtYX
ojQz4VxAAi98/vupBVCus0uUxTqmI460qhrooyxX2NHqcHpaRMdaJnN4xytsuyOF5KftAyvtdyzJ
EMPnE+6uVHnlFThJQ4txar5crATNOOe9nrOQnZ85YrJciWA5zeGWxx5YbwM3YB8YNeoAcTfnyYCh
uAeTE7Cm/JpsI+V7MIijcjO4mOtQRvYXT+xicPWBDA6KR904FDb8K6poakqIOFLUXQUP5xq0krEo
Ecy8dIQ6qxmdksCXePizNWCOpk4vLOAWu2V1Qy+/Be/c6uCmxl9yRqWFTu681Vtl027FdeTu2vOQ
H7igcwgCnSRTmwMuN0F0+5o+C5eLdWKwH5G/4qQ6BrbgVML4IWXaXrjJ9LERmbUQcD5+pvjVz904
B7kt0ic41M9ZEtYamc/xqAUr67wQYW0/rfxUQMT+gn2DiIDshvCCpOtF44nQxAhADVXFHSeRntPK
Vt0wfGE1jHhpyhD9MkUpx2XoKlw2mKQlRf+Dphn39L5hH5+KfNYQpQTfv2TgNBsavxmVH52o2wHn
eNWu//SIRZ8SootBgaKz7k+e+t8mtpaeqoOJar0JT+c32ky1E6hvuPXNEV1EimG7pWYUmXi7bXGz
fMjxmYU3Q0lSoelqKu75zi5tMfQlp2k04H/n3vfWzzOfpBol83cjitTH9pYB9jstNh3C9cMoH0o4
GnlRTvH+/32hjnNfpnfcKwy2LJAZixp6zxdfkWqJRuBxFBoonrkfp5L09xluAmGRBYlrAXzRP1YL
rVZhu2uWIWy6LJweur/2B66sm2YHTXm82we06fxCBeeP+2uMn5dN6UDJfEa5vddK3sPUMYVfNc9K
YmZZVVG37Bc7aeF71KKDAlrZZoOu1M8newpy7YQ9gnodAILlntBDZwafkVcl9GLWx+lyCbHoJJ/j
aMZPSe8baQeigeQrBgilVVAfL0d6sI/J1Y3ikln+7YWBUk8XSyaUydMYUy1pGfie8HRNlOqn8rve
LBUTNAvr2wwW9VDps8AnVKEN3WEq0GnM/o77bQTini3p0wtlgxz6xfR7HEC+HABjCFWAvZp7X8tI
cWLEH83pSoreytp4bONdsn9mGRBH6RBqAFN2imXTRILy1Y2EBQZmYJ7ZQ51gdvg8qyiubjgZ5GBs
fZdMRHE2I3kPG3OU4e1Jc3CoGEPY0l3TNKji9x6gLQCoSMfv6UaKccISwbENY+Hh1am5rIaVnSzt
vj9AXlLlrymFjwohWIEQlAYyK4Fcntu0fLkQ5/rbNGyyVma9UnRRwoqSu/cdSCUlHsmB0B0IJmqX
8W4M2GGR1OAppy5NDGxzM1qO7QuAXUzZU6YH3JLdWNKiu1n/th2/jYSFR9gcVqIHtGxX/8KAY5fs
W6yVrXueIZ9dy7MFm88LPkCCJwpbVbu2RCiNy+GxPEvDuOqD6cs+9zAGV6IbEsYHnxTnYYBtuKjU
7j+1dSrr84uGwytFhwnauL1Xx/feHQqsWYYbvX2pamsKVoFV/qPV/6OVwAGamfmDZ2tLdew1NlVb
SGn38Pskdv8rxKcSG92Svd09ql/LTOPaSQod9rRCuM8WsdLeJEwe2PFN3ijTTsUiLv4q8ioCBLdw
3HgpKSVaaWZoNVDOumV+Z/Q1nCtzwYrc75UIbZXGfcqz/dSGvh7+ebwYX60LqZqu04I3HWIMnJAX
uHmSl5SgdCOhnXF+7B1Zs6iVxJU698eQ3JElZSE2Qm8nULYhIUzCoiyCkOgHOwdD8PNIC8lsKHMB
AfjWoLovJVNGJZ6L1g+oTdFfZj9gXuD0k5ZmVuqcaNFNQqpDDxLN+QsQYnuHqjXNNZnII6qk9dqr
s2BlOww3DHp3Eex4o4A/Iyrg93+8jLg+dqRA42BLdyWEI7+A3MG8tdhmOS/Mgeyg9fjcfcCywJo+
47JSRSa7no/97kDOCjWHHrgcwVjGIpL36hC/8QMMRZYThvalEmoxs9WnZnjtuv4ZLN8/npFYlUot
QIPerKlfhrcPkBsMfmZaQ7Ps+3HNTLUUrknen5Dx3Wc1O0XDqsNPt0woFPHSuKY/48dwk9SQZI6Q
QIE9se/uQ9ESB0gJEfATk6OMlzQE4Y5JIvzfR+MVlyW/UoUQuXcuSBMaEg0L2lDhCcQL/C45LnQc
6fTFUV8udTA/zndsIG2Cy+LI4BlD6eY5ptpBmhcvE0FSaiipkRwhXmpxLLYDQwCM0g6eVt8Kb9Dk
V/kNgaNlEtCOtgPlIURaMUWSKRdvV/L8ML+eFiKcRZ1ECEJrT0DsKWA15SwfgWIBoJwJUAovIJyN
DDXAUUUFqcDq42EvQVpseEb4Z98HvUrpiHXEx0bVKxYc24y4Dpbv73JyEhAbAoeVOm6HPwWqocOS
efn9iQevgrgufotW8R/BvR59e5D/aCMPpZZ7/M7zrdpTBHQOOyh6OBKsaFmxQY7fNa5EzgSOQ/N7
7YbnGjmHT5ZQrQWMgs+W36Zcv0PknP2+nFb1Af1YkWVaBClLSy2wlpNUihczHhUFuz677MBO1hfb
PrThhF/ypwMFw49G+o6R7VFcQvIZJOFFlaq/WZgt9/RTvFRrX4a9RvVdL9paVL4X+pZnzCQhRkZ5
jh09Xw0lYzqgUYKal3wkXOUiWCoccTa9yJ3r4CUq92/buim2pjKrKJbgXP3VqpkKErw1UcxPW2LG
KitvvWtdWi3OuZXIZ8iZLJ2UKw5YL43se61I9OQIJKVLhQ1Kg+yOC/HtdJ1yoIPX8HBkk5jD8iNW
yah9PMo2oMnkAvyTP7kw0A6EyqjBeohi2AUcFC6B6cq2eXyhKjMStNn2b5Zz2Qm0u91j7lNtVgxf
wcYw7Hvzmlubpw2oRqLLX18aMEa45DAYtpufnyxi2m5NTNjIyRgBqj7FYcMUc3RhiUebJPofwrdb
ZgjpXvBynAxUzBXqJwiFlvmbDNBnVERIdjsG7hy1oOTTMZcVdULL462yqP9fT8eV3RtPcXzpDeT/
yOhwdr8gF1sCuuYJVzXYtbGbcMTSgKFCC/IF6iATbVaXlEHPtVkxqePEPooryJv1oiuyCc+It+XM
j/3EzWZcsmq46SHXqibg73zs1XcyX2iS7zAF3mdKWe1Y9P1412KTEIGSm8MYJez9gMOhGBM/n1+N
rOnY5jwnjFtEdvBN+benq9I41rkYa65T8LZOL0Gz3O61R3kzZVXFuEMZvw13HCNU351QBwTcegew
DWX4oDdUsw0JM7LjaiasRfaKDRAz79MfsXgs4pzucWcsxTOBVod99oZJVb0NbMJCAwVZS0BtjGaw
eLlIfq/glcMIZXjow8r+wEBiVN2F6ObkgtRXbV/po90GRrLPKdUx63QnG7H0p8Jr7tVpkujSWRka
vn7KrNLc84p54EX4NpHDQuiKQCM6WtSguodG520y+73MZrOtMMGHuNOjCQT7ZjX37iaVgouLj7JL
sSyUmxzqGlxCDgDqU6CD3FlOgeybpQJKihP1XA8aUD3Vbp+l6RoN6UWW27VvM7l+jLnEDSZmzzSd
zscnInbJjuRkIFLkeXTG4bBA6fXRMhmDCBVZNIY5+V7sjUv6F6QGm962w1IyBzmwfHXC1mAo58QU
6gq5pphdmc/2utJyscyj18nplgO6qeMOvo1PNGODcI7jePzQa2NWaXdEpC2MdWBrck498k95fE1B
Us9DhTGFUxLmEoqtnS/A7MVvsVOP/QkhdOFHf7OmSCub9uhk7LP2yy4RCT7jA2S1YIuefvLCt4by
v6gMt+EbOBsU7fGQcScL0d0GFlnca3VXykSUUy3EX6r40Ta4tpSUW/zErk+4nOi5FqsIVN3x4mnE
PEUjVJbVdaNxqrClq0HG+Q5J+Sl/311/LDhzZ/01FyYTCemMpxlgia4bUXZGRyMW0fcslSoLHK/W
9729BtTHPxQpYx8AoMjno1Habr6b81cKe2XRAZFtUTPlAv5zXxJSkTIZnoEHMLT9kMnn/zwU3yGC
HblfWReo//AwJVygGNMRt7pcBZTCxKJKsoyCkGksXi9lMLCqj0UYSw0UEy+uJEOmWaVBweoKjAKh
6X6Z0uPdFp50R3xH+L1CuOrzE+d9ObMwuGk3Ri76uK6+HR9TRaHzix1G4CqMebuy2DP1TRbi4FcA
VNWlJjuMa7kQstGFyHMDTljvO2BToCrdq4eKrQCGOrBpdLNMfpqWQjG1KYXAn7Yu/arwaacrdHsu
xS7vfSl6TR+oFCS/DxoTtwD8p1ksNNKm/Xb/JY+7/+ET7bdWXzaLOp5fVfVnyMzpIuuRnEsEmuuL
vgPLAXA6dfkZTvFZWQrtNrNZVu8EYRnOgD29qiFeY1AknxjDft6cVhKP7E2TNE41yyWEximVdCFt
nSCvBs0GzJBBhdyQfrduS2PHvkHB/0YN3WJYX/PG5GVsHNyhGlEdtRA1nSD7KAs2WmGM7IP4togM
cLu+o0MaH+zpeCqY+aS0ez+qcGpoQ0+aZD3X4JOPV62W+zkanBsOnfWbEMPid6P7BAb/JV1jsF31
z46Dw5t0RUd8ciqm2E4IMP9a+/pgALlmCsj6lvWx+qaY+uVlx2sPWB6ryZ9aC5FSDWZFjp4Flusi
/JXW8sLexHlX5bLrl9tTZxPFG7P9hfQ+8cksljGnQCAyi42MA/P5RqcjBXA6A5m05ISjYjH3Ywql
N9bny62+ZsZQ6OH9BrfO0xqBXhZL1UbgR2o14+Lu/DGjyqmP+KOWiaWWjbIpAZvIZqwAdfkDqUnl
QgLiTdseg+Ole8L0W9m9Wdx/AqZQl7rVJvt9AVjNOAUfy8zX6UYaN8hzvXaMq38PISWDAk3aGJ1g
LE8qMLbSoslrjuyPZufV3RDx0cuMNxyThFpxvdlcT91nXfyB/HU3ucy7xJa87qsX6leTt4KrS/29
3x+pBlhRskAR/reCdq5RRrcX+Kx34H3l/xupKedBHpQsE4PLc9aqmVRBLhVkpeMO3G9brIHaFy4O
m9jffteBkjJB3nh2BYTzCwhZY2fCYjW7sEpZZmq2v3woj7ekk8Kdb6fz46Jxk5bif5YH9F8gPPzU
5+WHQucN9qdL3YJJAJH9ZGNpgQbL8qZLki0LYBbNHGPDnLZ7KwfN33svBVR9jWkxfSuBkhMRXXmK
9Mrb4RZFFU6WkZs7QOvJ338zqAqEl1IUiQijqaMCcPanggwbGZXv8TS4abmmEZ3lL96YPVuLwQdR
VDwSGtqHO0ix4Woe4dDAHvx9P6LZcPlFVVLQTTO0AJVsxX+DwI5xyEnLcOn/VdXzW5isou5MhZzc
PDRYU8hj4rPEbh7jaRv/e3PSqqHSTnvSHtipv0d6tzEHvJVzRqUv9NTVnZTWcXV45yxWZTMMLHm9
0WqXyulqo1RcWJyLXjC1oYtjxBDwkf6Km1UXTe2LCuHWs+z6iKc7NajUgn+A4knLtjBAr/xa4hR4
GYw6FUMfPyj7jKrXLxqj24xp8C688NOGTbWbFCNIZjr9sqWxp4nCIaIZehKQ6ksY75CH9TsS9F/S
/a3VKDDB4FQNjpZDjOOe+QOyytuloZJXUFeQdKcQO9hUo7SyQVkXMt/FXcrMy9uvsdkYmUWan7e7
r6EK8EXTumMNMnfXmbIg+Z7s/Nbj5SWqWvrg3PPrk0NFFnlTzQam6efO6nXj1mF6O9tIw8vTdXIa
j5OGkZNyRKW9Pw9D3BmvGSbiX32BR7cNkaDEcuwwDCb4GWMFG3Xrc8nEfvdiVe+547zJZ0E9j1Dw
VMNvxHuRkD1x4cGvWRQPr2ipspES8U5HwJNR2AOt5BWLhiE6bQ9FYK//AEGByNvzdOmqhdNpptNF
Z/mJqUJBSV2bCKjTjFjHHTmN3LGj5pQdXcnVsSsYXmFL9idj2lvkzVMcgKKBYteL7IQSQqybikMa
79EVrJsFRkgJl8RZd+96xBvcUEdBD1AfYepEi9veFUotmK5/i7h5ppErpJqQi2dKpeN9vE3Yq8nX
WfCHeoIzIenG3j/YI7oePYrpzXm9BBLoT28Z6x6DAk78Xv2WXNBI/yc+5rUNlJCIKl08NLi9p33W
9M6pJ/hBuaRQv1m41MkcGM7SH/maUGNKLzcUmBHwRpkrcjztXO5CvjxnuRW78KPOAjZEDG3yT1Uc
D1Mwg8NfI5u4WEwn6eVcdrPdERWcAHC7W1QJdFisKA+ktCoRoX1xTO0gCClnSmhWW8Q7Nkh1+wZN
/MPGRW1k4rFznvsp0WmuaWKRgBoDeVQB6gWSiF4A8TjFVju10yX4ttsgXIl9pKf3psoaVTyK++yz
uGelR7wgNIJg/47p2ilzAA2Vf85UBr5La5Nbs505pmWdYfMMWN8DoxwU8SaByKn4GSfX/iQH2NbA
JjfJUAc3dCxr4ZYle7OzTDvIsV+Cucgzh4mwaKlSG/whV8iPSb5VuK3rsppemx77KNSe4tRl+VW2
DDAnXoP2C4BYxlk0bYToFVjVSCzwqG5kRwdxP1nra0Epa5VBUXAMSX9DPGp4cbE1/nJlVdOfEdrv
M/yVyNr9gmz01LGO4H+vF30im2uDiwTKwm59yd/XdFgbkZCdt2Xgtie35KBsa348qa6ipYh3O6vc
SAdJkB2/SbmrTvKRwz3XzI3ScGXnYDfIJLgizQHvaRscaL7O/AhpKATAFzJbhtKdiZouAOPxCifh
ySlQQh5hf+swBQOeAIrW51jGIMVrZ0Hk+nOskyZ0IMPuGWaIqvuQqVOOAvHlkyvhw6FHdooaO86y
+iTK20xqj6B+AUmvZU7Jw2gSGmCV8Bi9dbsM5/QY0KJ6w6Qce/5joA8AAcpS4dnc6+h1IFYlOfnW
ZKYmCV9QuiBtavwplXQi4CVlpupPwIihkrECdSctIYW+8nO4KX21592r8MbcRykozJcnpUpCYUPf
kqOTvNabg4JdIKqRHNJaZI4Pi0Wh8BzPhArfq99eI+rmZwfTZR6t5erO87m4N3uW0bsph+BuY9iC
/kmjKnDoxKUfslErZ5SevLGCS/7H8CgOMsgH6XfSmtZs/O9HitJOaRWQx/Nmf03Hw4N6sLI+dX8h
miA3eu3UVSvJheImjqQs1uZppSXrOc/FaMfah4v4C4xKlQk7HBWD3org7GfUFzTpviDtOdTJMf7s
0xTfqKL6cqkdT3XhIJxJ2WKcROtvZwlw0c1ooEGiSXyWmpD9OoCAxnewzljvKw6YEMqMW5IrEpxa
p9aTUvNiKfUAdTh577tOkCx2wVE7Y8ab3YtqEBbhKYi2sQjnraEoHM5maP6jUm5nWcHdDSn9J9CA
hryDgJyNhGT4BhZYap4SlLvcgOYb88gEPu9pIuaj2SuLDjw1dgDknJrCV4KrvCshM+7Bf+MU3GsD
TmEa4mCCVRQioEarceiXl8VIO0WI7wXM+6RRA1nCv5uESRLgRHl4GvG50140hyWPJaThMhm+JKL4
kR+GbyQNjNGtgmLpoCJq+qqxVn2MGGKZoT8x+yjP/1UhYT3pNFIq80jc7op6Uhj6cokHyaY5cNbj
M9oqpvrzErdqCc1stqMM/xH85FXRR0Vzzc3yWaNsVQLUfMJ7Ges+GMNPO4AlTLKjJAdWpYKhybM4
9rFHhXnFh20KyZpWXSGKdM3DI+IDfi57qf8Vo8XFF6vwYPHw/UdpGTsh9MpxbrQwg4J1XwAqob9s
5pHwM5TP9Gg5hqtJYp9twS9oOCK+9cvlZMZKZp9pCu87v5xE/kOsZUeYS0Fzx5NG18sh+EPbQTgH
P6rrMW7EhtUv7RxBvM11Tq33cKK1dlJO78bY42HDXTu+1dHZp4jlFLvFIrR9L+XUAgrjzg7OkTKe
CB1PIxxXmEBJxt9RGLUMk5sxnEGS4/iOa7HXvTBmCz/RvRJXQCMYcIsQMKOA7mS7n922yorhbBhJ
3oaMyppN2fbBWET1Y6iG29KlqJ/4f+gyIkUKK5Vqdzhl/Qg9nlyHTyjjcfFS7nntnlcMt9qQwbC0
X/sOiQFeaqh//4GQhvyTTYdxDH98cLIhdC+oFRarezP9f18uFrUuk1tWquqR9qc/g+Dp3QVzt3dh
+cYRvCG6GH1JhNgJeVYmyMauEcoZqtlmm2KZGsNPE0banoxgS9XT0UAYH6iLk//JS8+CkiYqV4V8
MlWWDblsWF4Im1ZzztCazbTp8JNYa9N8VLLS1ucc/X0sHtsONAhJ5iR4QFqxLc4LyZvXjS4JH8II
InYnmnkbLzSsIXO3iZUmfRItL0qDW8qyvOhDW/TWBspnfWopa21Sq8LA8rTIKEj99VqtDI5Hl1lL
y3mNBfjD0QANf3f169SJV0+0HMxfpbjnUBi1UWs27VPbokVKVpu7+4uF+yJCK6M7Dxck4LLE6ms6
iUqCaqxUdgw7OJxOP/0ZNGkc4NwGDrreBXNvvAeb6/1NYtWivlQcXv0jD/qrNKErU4b37VL8axu7
cha0YVES7vZxPX/KeCfAp3HRHzyUNUZe6w4ZO3meRamYcs4MJEEgkPytcoOI1Yv9pqPh+jHxEh2b
COB0gvpdmgujTML5zaVTiysjMDZFScPUSgEwMXOGdYRUiudRornmonfeOWCnge5LuN8caCyOLa3n
gv02n9+06F6NnfMKiY+4mepc3/0rgrw5AK/nbc3QiYAhNkdyoISRrpMmV6Vf8csRfaaqLxek9ECE
9In1bKY1duLdc7pdnEA5jD7dC5Cgp7bnPhVXrVH2OOpgQQ2CC474l1bTKpQmN2zwkGpbPMZ+s05o
2W3COj6T1LDQQ5PogUAH2ZM2lekty1oHncIrX8BYWF/k1q6vgFQFHdPxiH128l3hoZdCacmxB/mg
R/OBcbewws+2Hm0ysOU2IAybGYmPuGwuJcUA/qZY5Xqy/wJ+Q/Pkix13XC72yrjKLMGjA2lCS55f
xozoOKC4aSFP+EQNv2RLj/Vq1wTfh3RBNzTwvCpZksRnhT/LzOqXLNcDa6UxC7XkSS2anioLCzte
VnrLcaZRWBQ4SdKEOyMteQX0HXV84moQSe8wIHN32xL1gUqod8DDK83Cc1ccAoo+gcBnEi/uYWEJ
DOGGfwtI/ZzeOTYC0vz0ekiDkpzQFkYvlHaEBupIbnwnBZ9ATL3BSOTRwCakQcagC64bagPfAcdQ
8S8U1/4HrX7OX1gVnN45njSIVSg7BfZ9Rx/uMeyzTHYv3k3kqQcI+rK4yIltmufFiJjwUGUPfzSF
jz8qtZmz/gSmZIBfUrGx05iy+Ph7CcVs2ydJsMbg7+EQw+seA8M8GA00Z5OyiaCoTPnoBnRCot/U
tqF0Dds0A0+UNgYWQvwVQ1Whh/lxIZRZPgqhZDPWmQRQ25CZd3aRIjy5r1c9ZxYwmjYe6TWJpRfR
t4fjX9rwgOK7NFRvKV77zIHK6P9L68j4iuTJWOl83+F5FIHq47RfFwH1nmdcPZoeSeyjh+kZ6vyG
iOiS54cNfzlLOfruomTp5bNvXZUMWGr9vzd0x2HLh2AU6ZjiQfO/l/T4OsCptx1O0ptR3NJfA9c5
ZT+NLmUtnA3u8ZzcULjH+VwIqsWOLacXS/mIFMj+Lb4kOL60tEiwfDutETg19vNwo9RCkxPW/79C
oiLKJ1itmQR4E4pqe/JIOR1AMZPh6bvmRiqQUBywlJBU8Ln9qMAWeNLQ9Jc8NYt+wHH8A5CpsNmn
SFCwYV0Olb1f1SdUlds99V6+d8m1nvSHddpVCsqtF9kBKIaY9bWeSpTgilf2jLduBuT/FEvVB+4+
ITlDzvQoaWJvP6JZf2gFNGDg+K17B4+6vaT8OyRDh2U+fFb+fFwfDsHfwlTL9B3M2hhevyMG9PVC
4W6fV0cGZmXgYVlFZYadRUmPNDG4sxGFr01+wxo7AjwXAMfYwMTaI/DBPzd6lPaAmIBKQSyBuO8E
pZ8wVwgy6AzzKDBUTR2+rjVxOqcgKC1B3rB3KHYLkOAXT2FEQ4QjazdBtULWim3KD+2A25mpFrqA
bxARvzbfdjimUrAlaBUz9GLl/EaJ5xM6BpdZQXh34eS5b5qOOeI94VlVXS920fw2iOMOZchm8dYH
YpLi4oEsjenmUDbjyqkFPW8klCRiKw5VjgexJqDrURRy5NgrW29vYiV5FbC0nZCnOAmBobwuSQSF
1rIVMkIGXTquOv+308vPRWbM0sO01nPzkm2HbycHBMQ3H/nnBuRjQonYTm+eaDWDFrFNCpEE8CpD
LzOYFcNnj4G+jg3yu8xyV5TSXJIlIJNcOBKE3L+XoaVp0I1ndjXjD4Mt4UAQFGLcUQay++wKwtbP
XB4s70CRNsjL9m/gd4Z5YMUd7TMyCRXNQmHNRoxpsSmrabSAsqCttOlYinNHEsndQx3pJ5YcKQyd
I7WuCIDopUXmefy4FGSnTQHb6UJdvYC2aOApBH2G3XfFTSKKzBNiBHuEv/Qc0LcNQgmYS+sJgOdT
SQZbuEevwkixMjWPbM7C1l6mQhMGnaL9FEbvAIPdlx47YgmVHDfGXoWlR2XHa1Fmtv6ErHt17EbI
cuVGh3Fvfgc4yhLHKzED2LSvmUoy/xVHCONuhjH9HUHchRAdCvy0bjgRU1qBLW6+l/VE9JyJYBRl
hmnWWWcj+Bmvnm9UBYdHEONv+HPxAWao07o0/ng9Xh8UvkWu3Bk1KuxiwoXMeb9fQlbBf/xC7cOX
72FuUdFPj9LzSH/FMW+otXdPgdiJjwoSJK9l4EwmAKrUs+n08xIg9u1bYaj1svl1ZDnI8FEN8+2d
3PR3vFyFn55x37Mwq76qfnuSTTTP5urR36PByUKw584RoYpZq7TQ5rv1M1sgrMhg02t8k33mfYz7
iXnW6qa4p3Ek7mlgVNNQoqhQ0NiP5+QfKwJMfvIlYNEibcL7KFMNVeS6c3VJLSWXMZu8p+27/I+w
rb48exbZuR7Ma31VCkCwBzFz0ePoLCp8oOcpyKrqBFM8gJU8f1wkh/vFqbTteGvmqz60es5gMCt2
R8+KuxW/a0feRuJR8pmWeXSxoSq7FKx9S9Gv/rUQJTjAgiOshVZVWbGl7q51JojPzOb9uJEzd0pr
2XlEKrJpz2XwxEKXq8euFOGQmpSJftvzEiX8m5YeGoMkiRPwjLEBH2Mm4tq1unEIPtORK4PGwAKh
eKerJq5jEpGb4ZoZl4GIHt/1UkvcHoMKy29mawr9ocqroGfvmM3dAirrckeilPJ8Z6vvNhMb34ki
HePyxfqBl2RJybgqWxJON+lJKSLykWq9SO0iUYAsYHLG4TxP3xfQAEL3ZIpzsIWfdi6WxCqshXZq
Cns32TvC9gszEaLvvfqewEAVyLIRJNevfg29UNa4WL5DQgkepbu8qiE7WcxEW+Ak14+Mtc3P+OgX
gy1vG9a4jDOVoc/AjpY0fHqtul6E18YRNiFvxuGG175WQUZHvdKOlON50NHapDuZhMcTbz8leFHV
9z/wR2AiXYiuPnwMeqh2oUcQ0i/wlaC/+rSnSm6+hRgQwodEElQoW5H9Ef9UI2wUUcne2NJkqNsV
XkUlM0cjlVHYVvakTOTG+/xXCFZGzIuMLmEgPrDC6K0xeotFLwzQ+Xxl0/XiHTOr7oXpw49UNRHo
+sTuXfK6HCGEdqLVd+vwYHBhHckouQ8eicy3KtGbGYuDmmh6YoYhNjPEk8mDnJA6dTAtqMWhVztb
cxrpoUKs3OGWlJB5u5Wl/QSQjnNsBOInjIcxkdpbA0ruxLUD7MtehzziDL1KXQq/er9jpvmB4Fym
kAw+Cy/hzhQuvJD3qUV3Qwj24UcAziwlH96aOywAzovK3nFVCiiO4l2bZsUXHThDE1xJtQRjXShF
0EQzhlSXnPkUQ762zezOoGH21rImtNJ6cmNSpur+a4XUI2WYIK/h0KZxLTg4UNPeXA6CfdoJllyt
H74phmnaVqtws0QP17SDJbn6nGQAk3dBLj/KsFBCzsKEpPf/D08zLwIjZZTQiV5j2UGs1moGoC63
Lg0CXgEeZ5Ii1Y9YcXYPwb1krrM22i49V0ytXAJE6W8MfHDEPDOQiXHOrXBNtbZwXNdOrmZejYXW
v9Y7H/7O27iP0K8dACi5iG17dj6wQDDPJxdhrF5XqeGUqhl5/mNHIUQIMWBZgShpT7VSunxlzT3J
AJOyWLJg94rPhUAhKDRM/AJ/+Bx3M+iNqv1TCqr6la687l99oMf/01UJ5FBeovEFwvQoPWwSkl1d
Am0im0ANLiUYoL+WzgoQQGDwz9JgdHRTLmxjtPN8oBHWa+rl73USdxI8C2sW4v+9WT06gzlhc3Dg
pWLQkvNKUMo74Ez14QkANZDGfEco66rSAwjjHfwaeACv0pUGBRQmYSLe3KejGUfcNWzhkYSx16g4
uIFni9PBk3XiKp7Uhrj5NDVY3RSu5ttSNRBVylQmUp4xRUNAUgTfLeM4q1dh4a5LbX6vOEenkAQJ
Fjf+8fmosFrziarffth94wGKqh3xRbX6/dLNTY8tgRGSrtgeCTw+dW5OhdQDrk+RsOBuTflyObYQ
vosPlEzDgOe6ClyXxZfgmPut4tJTs7fXMR8nZB4N4IVV+Pmn6y8bNNfzWSPwaV9Vs6JuUCJOVlLb
kqilCVG6X54Z0TSga5kPMbciiYf6EBhOswtZCHxkYf33zsss4ZCA6mzhTosBVJWWbIUVvCKE/+60
Hm4NVleuclKH1UwpjavEhWi37J8MHeg4aF0JQ8HXdcpcGiQzU0sHhIxMcfjvJwZttm6YpHMkmE4R
+iyjLNXQo+bL7520MOlIKN3817WPEfZUf1rBwYEtFN2NPTy9g9lXScLIPJ44j89oGQGA0XUxLR8p
Q+oiXMrDI6UGW99VwJ8wX4Mzk3bI9AGFAx9cFKF1yjvtzKd0DVL8iZcbhG7DvG+jRpjJONUE5ugD
fOt0u1u+EHck3YxYta0Y9yJaRNzrLaY+rNxeyjFyy33j21puuLUrlV2VmkpcWdRNEkJN9FcU5BuP
OfMX1wlOwk732p1sMMC65ESemJ7ctniH48WSooJ5uzQUUxOc8kqAYKTlJ611/RqUHtRVPmLnHIBz
SVokre0aXQYu8ani2Yy5Tbw5GN7yAF3acKgqNL/jHtNAxs20eqPHh67zcIeMCDhelKECK6a8IBTg
etJBGHaSgu+kOE4C8Jn9mm+UTOHFkuqqQE4DMeSQFVUNBzwkmEeYstT5WNKmX+bhtbGhuTK0xHLZ
hhiYNpN/mfb3nZ4iUwWC2EHpzDEQqXIOSoB0TbZaW8lgnJyVyq1JsZ6srSHqPMUOWuStRABd8cLr
ag6ba3dhIH8XDOvqRQ3Qi00feNkeFgT6HrV86m1jHfQcVuCc7cdpRP0TCdYvSO3P3NwVy5VFx+Vt
K8oEG/xSX5iMBgOUmabb3IAU/WOlWC9LzWS8L92HkpyLIyKB2HTNQTEFXThKMyjagDP5EwXC2SHq
NbCUkeNkUQ0Gk8O2/mFfABuaic/olnR9hcaLxfsZSuL281GYXj3Tu0t+eYg5v1syLeddtvaoCDlb
IBFyUfKFmWEO/t/FkMqOTqECxVZDuf8P1YaZY72/RmmbZWf8hn2Y+chQxB8tTr+wJnvIyMoolDj8
6QKPZ5h7Ontpu3ALHsAle1ZrAeTaOxkR7Z+YbsGWMAUTWhRjIT5ZdZLL7veLYdxQsKUDdQtJ2a1r
1wP6x/3WHhTHwirsPsZuizb9muQfXy4ej2xAb407mXFeShpzGuGe8Vfi+DCpUg98LZZDE56pwbkr
dVXVIEblMSQX5sWM0DsIBS+m8IChLlHMjoISuznIt0eGzUCclHdD6wxRD+LxW/9QTWY/XD1maorw
CJET3nRMfF0D6Z31kCLFxWO8xX7Q63p5sja4rANeGJEbq2smUhALBkNGfQC5dMPHwmiN+2lPM5Ce
VLZXJJqCDvtsnzPmVuOYeJsay/wBd5cDXIJsfBaz1yqCncvRxXXNGruO0lTehapEfPjD2B/5SlVQ
lqNb9zjFD0ukkAL6iuVLt7K825KsDh8bYzoXtGuPDu7lRwpDtYgJ9sxR5NVXF15hmiU31m6cal4m
xzEHuxypIOuMrmajBLHuBY65ozVRpQr6QEXu7OUXdHR9EbdNg+uju8YkIN+wkqb6Y4zu69TEjDqV
UGxe/aVep2GHeebbLzk54d7IUQlFT7bMuWPyUlj5Fxr4pCFvRk2mKviovPrA1y5mdILV/IaGywKY
aPGs5m4CUAVcDykaWVpRNkL8HoHOGlh8Xc+Xrik0ysNz5HX0Wj1yxECXbp3OfDr397LC+ED9DZpl
1oLAtaHGvZSJ8WC8ra4tvDquOp+2RjQTJSQRzS6oiC/d7uLL99+XcUcYZbh9lD3IcpjI+t/NgH5Z
zuVisTffheEJsXxmxljt3/G6885CUpC29An9EccmzVaX9JtYSrGkpwUF3dAfY9gNUc4RuXTcxioO
yDcbbgMJZ+4ZGNciLQV0I6Rpn9F6vfuTyTQUB80FpAjFE/yG2UWcF0EHt5Y9fuQMvl1Dycy5wJU8
h235eMQ/1lrgvOEs0Zf70QtKuNIwLQng5uGuplhcYTsXPoTfWN/Qyy1r07i6uMz6F+g30UKuB++H
HBFGMhJZzsga8rZqIKrJ3ajaoQFqBNdOi1XHKdZWftUOkTt2W2EWDfPUVQoZNf41NN3hSxGAyPFk
vRNlBGUCQVEG4QKjVFJ+TjivChTjHPqszyPMiebDCCsNRacOhVCloEICCLndMjlLZryxi0Wjm0gr
W42ju5/GevZ9CMMjND2jr5tVwxAIzFfhv04IINkDO2t7jn8ycdHr5V5i1Cj6UofxEcfebMZJEIDF
8+to9vehwKGI+vb4pEr2TIU0MYxN47LyVj8gJonhWEGBtsXuE3QuLYaNFhLA7u2JtDq7AdUFQrtZ
W4dwV9e+zN68WsWGCnyR8uxepCqmvV118/tpOOWC/ccfxzsgXmP9aY1McWGcnxHLufAbnq7GK2Ek
8tPowLT0gfytTcC3zZQZBDMk/P+lawcCfZW8rdoxDECq4hDU4NYqajcf97PqmwVtrEMpk2pikp60
0CZiQ2lrpSI0GS+sSohbYEJwlsCHwvKVAAx+V6Lv3JHHwOBi2b8OXUVezylqKNPF6pGmkK/q20Kb
WmGtepe06AdZymGw3U8IZjFpihg/+/ylrvGRJNjjD2fT7v61gwCgxoYf/db/Tgt3G7zrinbRfdAo
kIQBklOSZqe0YYmIGfiHwSQ6xY8SYE6Y7tykThshd/64lrJBFwSPfYxTQWxwDQz0OoFX76b2BOKM
7TZLu9o1x4VjJ9iB2KqlGL2t8Zk2NUg9RHwvmvYf117PUohR1Rng67HIC0RlizSRxT4o7PCWAhw4
yj6ao3D7vonJxL9kBYk7kbkM4tBGWWN9veZ5m8/q8r8iZ4L8P4xzIExMmwCQpNAmS3R+Rt+ZGL1Q
ginB/Pv5auB3SSBIyaVEuN+B/ufGyfM8NhCDMFHdDT3QC8SiFBJXG1ybBuRszqaqeAMnpX66ROG4
67ms1zdtY2sWnCmL8/Hj85ffMfj7x2VDUB9Mki5GRLhcRaKWwKE3F/GXMMD9VH2ORI/slUZfSKkP
nJDyGwGfnh2pGPc0hT33/FwzNhHRrNOM6oHypCiqnm7tsGhM7oDY4rWVcjw4qJ3s8dPrSJbdZgQ1
qqLJS8l4UVj6fRiDBC+7gw63+NVaEXFSKtJ7hRbB0CGpYMmLnTHMJQDt4yMVEMFtcQRq2trsTOW6
Q1Ifp+FXzXpOwxn4OyyIVxSeo/QNhT7udWg1i/9STGCxJEVQgLi/2QLBhtYDE85YHFJBRul94Ipx
f2mPHuFYPIXrz8p34BbFm6odZMLpTx+e5bBqjMJ3i4WZBGxiy2U5P6W0LYd2GhixWqdcFh/69BFF
93fJ8+1dVVPT3AK08bInUuixQlFjNPeRFjEIbY91PbRxnIj1Xq4hkVOezNoWNvfvS5ELJVeVUwHp
XajqBjJ3qDD2oT6BvHBrVVhSR5Mt97lm+M+gZsAlUNZzP7RjYbUOs8sMXBOiAY8RepR5vat2Wc5W
StMUov7axx6pENd7ABHRmYtHuiGzJsQxy8VUqxL/WnctMrHfjODvODZS9We5rw5KOoYJtZ+OlDDs
mkmYvds125ovJW9YuuNZkRt1WOgJgS4lqWbHT/H+VFnYKM9RG+0xVD9+rv8iMr7BogXA2IfmLb64
h1/K+gO1EvRYrrrjVgiAQbFieNujLcaeI1ya8XTjj+VWrq2jT6FiQrgzEokY23pBBlNkbacW5lPS
38v6wyQNb0GTMoEeMIamhCeLGbiaQKOE2ufW9/opVVo6AiDrOEMutt5tHK3Tw/rfvCRv6/MhYM52
DhCcZgZ4dx2FpzHEAZI3SWAUzAopwu2z+Lsd1P0zWtnaHTCPQMmiiyaZcbu5lSXnwkaUyZi17CP/
7jej+TEMfGWFZjcVdN9kuiGM/nSNg3QymBKjy46hpnl7+CYZTCSj4/OUlPfrgBFE0W/4x9kJHE5d
o/jOEcmAZjDkYzt3PGm9Ugcl2UvQlLT7pWvfkSYpZS7xZRJfi0uGlPjoGJOiWId2vzFJgKTdhuXM
8dMHV5KfwXoIswmHcosWbbgv1qDq7MBEyaF2er2cRRS/JR2bF4GBntQZ1FAhjMv5CKPfVlm2+K/7
+lvmbwgxEYolkaQhPGhcdihLH+b1MN6ojqFQL2/osMFP99d5gDpaCZqp8+2ZakUEt9KtL2pTeBV3
oPdufF7TUSwZd6eMLVS5OWdO6zs2Gn7vmNr+2m2TmSBhf3KvMeQhYiM0J3qqywq1qGPF80DzOai7
IyExFaIu/tBcVQtD60EanOUlbxy8EnoDsPP4MJpRc710GczNfBBfvvRl7YDfuYFpckpWtYGn0x21
Zp5Tcc1vwIaL0DQlmQ9Vg2wOulHLpyfgaqq5GnjRv4l/j6BbloV2Bt/LgxPV7ttM4OqqfBJ2Pblp
YSsuVqcQU+dYp4d8/yi3Vwv+J29GMi5gj3Oj3q9p2tLM2Nwksx0+wf2OPtkW28lWMldFiDVGKd/7
PX0U6cKqQzpKPNvawpOG/ZNbJDzWBzS9dwsQepPdejKGjF2RWlDabfKX1eBmpaPemMEek0f9VKTA
zK9q+aqcUjWNi7Qewr6uxy5Ew53Ok8UsaHREbJK/cdDngQBIHTnJwDaWt2JXqjomT5fTlArguoVG
LNldLs4lw/hBSURppQRRqPoYRiEuk4l+VQWzwnOP/BSkrFm/ld7nAE5PJ3WfSluJM1P1u75EFW2l
mLBnud1pgX/Hi4UI7kQDcPoUbZdSSkapUsKOrDTJIRyRF8zSX07GhwHdbuJ4vjGd+gVYGj6Ev6B/
OvCZbBAvEfZstFl/Mp1WKxH0joCcQRg7n4JAU75l4L1BsgLhPR0LjFtq6dyejPPH3Blun2K6CqmX
JRZXRX0Wid7fY/aCgokFUep3OgMkiDMTB7HtChs3pO8Q+qYD6Vj0c+a2UZHxyBTSOy0hQJT/TAuX
2F3BnXpE1lqycPkR9tvwJyG2SmPQzxZydtkYCL5s3ms4Dn/07WQxngyDFjb2KZcfbta3ICB23cSX
aJpfMQ4C5H11sP/Z5dssnwIWKA+wFnomr/mYRRXab5X+njYrEmRmNMSgGVLEynvEGbEwA8h13teL
mP31SoZWTuiAHbF5e7Pv7LZ/iHl2TDsFQvmVXm1mAt7jLqc+YF5vD+7R2PhrCTRuqQ5VvBj8RE33
Ik1gFQsZQYNw404gp/q5AsebhzoxvrkIkxyT8JsflsgjKnZREG8LAxWBB0Yn2kGwwirGeKXGC84k
0Vqj8HQ5RzqikqfB7swKKCQraPT/TZTT+IOzYdfDU3Vm5J7m6zCsgIQ5UWR1+k5o1PeNGXaSKjW8
90kC/YSPrFay5vto6Ex8OKD1kbAfKjoL4v5yc+vi9mzAZp2Rm5gItXt2iTmoOwJiHlkkyyWRCW1T
gCockjAZ1dexKF757DK9TX2Mxg0cgh/K5kzkzoo3T6guwfmaOc791eGHeij1VSA8lrxr0FN8nS5N
7h/PagNJjNONN4n+NiTUAu9LLZde93HpFykfLzfD65A1wD9Y82AcLPsVfliLT2OO55RjsEdAMOUE
C+w1nJ/26wvSTPKSdYJYlSWGn1Mc++553q5MM3YwYSOZwrpWS750EgYUf1sUASyvb5As4C2C1ctE
5n9bZRfRx3xr37d4+Err1nMV10oFWwY1KUmnwyov37jePpSg1eurLMTX7c3I+YbQly6zfpI63daj
1aS6x6ZYJQ6toBdXC+q8twSLEqcyIqk5SHIMYumaUi1tdh5iMwNZ3ba69rOAbaMWvLJKtzQVuDkv
C7CQ4lRPMbJSK/x1WoaHI8oa5F95k5MAwxHtWS0c/aafmlQik9R60M2XOrB03o1jDIfizIgPBRM9
pWlwYeROpFYDeEtHUwPMYxxC2k4tDp+r33/+JcZTkFBBRhEVwBVG5dqlc5oSOqtdxfbOfTJTs8WG
uyHLjPzIglXcGp64mf7hRj6qR9rlrnq22iyy1yeZ+litUfUmHRe/tgTXqgFbJZ6lLgUZ2XLsjlwy
xIuLiQWszhPLptVT7Pp1MUsY3RmSyE1HiysXRV41h8DnwzOFbUyVjCQdqDVtXCTCdb5olxCjBkpn
xBzP3VwYvRUAf0luTFHNsaHujavXY+jJ2yOvJvcEQomTN9ZspXVGXFq21HuF3mc8HHXLUuO3wzRp
Fp1aftxQihFz9USCWKsijgv4rIRoy9qjY+mK0yhmGllQi4KkReImSpcnCMVGReW2VpSSqG6/WEyl
Fmcx4P8YI0NoEvuc/41pfngeBGCYA0EGpY57ikUiY6zFO+OjrOR5RCGYk2M66nzKXlmQJIb752zX
OuAkIFM2SchFreI+ZNRA6ciXkSId1gS4t2vUvcGhgHFLb/JV6EQBTNv6aIh9wvn4xmpc+FB4LqyZ
NnKJcCH49PmPXVmG1KKexIviWqS9AJlk+4Rr0jc8VeB5MsFa1m5zSt8/pYy4/mXXGu0eBulPySJf
+gFeAmI5iB7bDcIHHwM06++aINXn92rBeIVuMyxsjBqJynPX3DGiVeFA6bvUnBrgf4gkVnATFZMC
LRlwVh94OeSyb17ccanNL1lsY5e5L+iq7USPPfEyV0Uqv8VzKrM+/qDT+P9fyE+YbJ+L6XJPGdjb
/YFzW5xbtPHWUZ4BcQozSPDvaAYkC11LTjxY3PAYcJDGTiBXTS1yYSXP0WpmCkuJoX0vLjf6zLrs
peBFlXZ8yoaljnBmSA/AP07QY6ja1o+wc2qKpHiECdCPBlcIvKSLA99cHlZoUmEqMlMKDv/+UmEJ
dH54xLfhWRWIfUoqCIoLaSqXTGmdZFcSCB3HTY3bIxWdXviqBvqANuPR5L24bivDVsZmj4hLP8u2
SFaa7OhwqIJSt8XjZftmkUpicfU0Agw+aREs8/k/sQGLXgPrxTZLMjvppw9q8mrNAncbcALrXr1z
Tfz4pZxL9usSuzMEzVQX7xgFIH+ByoNC0mQHREP51zNxc4MDPnWAYRqR9OZ4j1sQp+OkMQtRvK84
xvqUH7i9o+gwjYKffYRsXZfM6h2wuFL+NIlo2MFSY959oAji1bBQsDlF95orlm/d0BcPlNp8j2Zc
M+iUqfBwPxiFWK4wUVKf3Q5983H8J+kHTr0AiV/5vCvU8Ufqqs+A6R3UwoNS3uy/3uXnlZgTEema
FOnigF8kROdrRTQY6MV7X1cbYZBnE8sLj9ZKIIqyyP8hEiu0o0xWXRQNQk66M/YCbrYoF9FCsmMA
p5ZfEEfWL+lSGYBduQxMdqm1cwj9otvshV5lymQDyDPq3u5nbJhNmNCtCnjCf3qxEEvSTF08ErqP
6BpEMR9ks4fCEVs7uCOKUEmZrc/5aFcJsYvozR2ysLi+6Jkf2lRHIzix35xP/1hB3j00FT1nb/Bx
7xDuXBIBLck8UxmxhvUrtXjCgFAPiZ06FcbF15rv5u2v3hx6YXFx63U5xt4rD5Ps4/OSemuoUcyV
MSfCCpzGMcslZUKi8JMgJ4Hgjttf7C/Gmi9P4XYYXAS+vq48Pc+V/ZNV9rIzpgtj5PBg3AcNtEyW
l4ov/gtBlTJm3vsyCzNvB0/nDWzZEMb9aHNPCIRN9c6rgiDVJAGpDRy8ANg4GcNvuFG3R1EzUDEA
DOeFF2Px07u9D8oKZ/24/0GqOn5FxG4DxwfA1YcJFNdp2un/dnRpmMgINa7FvyfjWLart1XXXIl9
m3dWEQDf7+6SXrHuKNUjVLNhF3YdUgLazlLtyG8EUg+GIRP0HIMrBBhjQR7qzbG+GYP8sjQV5/Xq
5cn+nuwYZOwIUa4opqExyvyHUcrIcE9Mgp/+eLk4GK2qSAo8SPze8GmxDe6fJxKHr9ieNABoQnNG
pPemTM3pc9Rc8gjDv2cfB/ytDdhzmUu6jgnEZ2KC77PpiyXbxt3S4xaP90TA0HA3ujbR+Shv/+lw
RpY0OPsEX2labuQiQKha7R94umxChQLjNLme0r4g8K8q020w2mZCqh8kUGawK40QKfuEitnnp/tz
qKs8+xqVKWSupDy598IiuJPJBn0PvON563Ywb5Uf2mhJw3Oirg5NbxyWNzZpfhWxllU1reFm3cX7
FIn2gZ02K37I7wd0xDY6vfhxIxHbxZRKS/xvFYOopoZLkMiiL7ZbV2N+UqvJUDLbYSAKxpq25Xu/
Fe/DOXfsX/7pOcdmRCu5XFjWxaoDQUIrLN3ij2hWUet2XkVcS3pLkfzOK6Y8Cy0g4hlAVpkFFQEU
z/mPoKaAMd1OMu/JEH5XW0tp+HglmNjZf8Zil3KzqR+BOIuTCmO6PCRrPB/OWBq9gdL1ExfGvArU
Fc/89AsF+ofbW5P1WtACwowLO+E2ZHHm6ddVHJa0h0AZrP3TIkERVZ4IbC+1ypB1z0LwrXXQ0WQx
2JRNTN00tDqPmMWiLQdxiCfYAm5HSKuRBk11nh6RcxzSMttS5Cu7Y04s9WwouvWaXdmOI99w2ltj
6p6seH8wQ8B8evrLtmBTUbiehhhV4B5rZ0Za+ohaGClrMm9M2etmeVuHRvrcq5dI/QDaWJk1lLcA
wEk50c4rJCG5jL+pRc5f8bjaOFD+PiGDI6dxdJ9VHTQbBrWtEcF1eu+8Uycne2P3W9A78RgOT5s+
wE1Jx/CMcnyHw/8uGfFKnVCTZkWsd+zc2B1f5jzmXH3dTMgDIc8QMW6tFZi/a39xOC9itVHg6Qm6
Z+jkA3h/nfKtH12YJbfWy+pCF7IEFjK7ZkjgTfAAmfnxKa/xr3BIR9+M9owVUeYZtV0AbTdzx36l
681WRrjgjrWDAoK38ShvfI5ywtEkCz8xCgfG4qCSaw0iiedQpMGllb8MSGunVhXSyJ4xaJ5kDaKz
/fQSCq8fheSWULk95PnVttFWUh83jq5vnGpMUoCe/Oq8KCYM7CnTCIjj8aDTT+67jZqLNinHTIws
Uf+ruo/huyiG0hydLk3FxQUaFZFRuy5Bl+XIMccqtOH9BGYBPn/zjxBjM0tG9sA6cnC7n6FsfdXt
gwlKC0+d1GzCwBakdTdt0GJYM8o+4b+qlxVaMKIJy5dYqCDKBG3YgVAxO51MptQF9wiv3I1Pisqz
h5t0RVowfHn2UnBZYZRswD8gQXZXH8o0V0hsg9hoQUbM4fuDfac3E9jUz3xQ8NQwBnwdAZvP48xs
RMXdWj3IyFKHfjY0PAXAxb/61lQCiaP8TH3AxDrSlmrzz2GL9HE5bemPjcN9hITYoMVO8CdluMxB
1YNp3xGH8Utfo8FwzVo82HwmZIE8F0/UXrN9Y3Y+PxylLSN4et1+vaysp/mUdgRNSh/6cAJbj/iT
gmRJ75ClWU9+BRhVA4YUYQENHrDzEGsRS+L3b6CA4K40mHejNuwJ7MHtou/eJ5Gkl3Y/mxtGumEO
AqFiHV4ngRre1v2gjxqb+Qp9T1lyM9758FJSNA5c4YV3mhgd4UyZ8sJbzvr5ZfZSwEPNI3X1w/is
jv84p3WWh4+0TuLjsn8oqy0pSKKnG7NpwhGcltssKBR5fa9EaAE6Eo2qK4Jx8qITlz9wU+WekbZe
bUzQ2brDHoQ4RGkVYo9E/95TfKxK71WumSBtr8VXszIZhyNaVz5uM/5D8C7UtpbPc1BXPchwJW1K
S2tDU4sZ5ActgU1ST7UUEZLXABv/dng0zIRCvk7OWS0YN6hPtRTzarbSLJfVPU8J9pioBijHK4gj
DRfuMwI8ojoF0kCyOLgOEEG+vMvK7O874GNQYCf4zVVqWBR4MfcGmt7y0hUJNavjFgWlhDCEOL0i
Y9OYO+O/UD/UFf0IluhEL+lS/owd9CAV8Gi9hkVOvcYwL5RYNkhnnNyT9GTjJZQGjEQgIkZUSL85
xkpyJgtcPRCRy77xZz/HesqyiFk3WicQK2gnHjHU5xSLrY5zRxng3jR9ZSHXa9zNnrO/J6lxZ4jr
JNYmtjd+8QazsoLsvGgqzi0MZ73Pw2yrlrc02FyRhMm4VDn/f2ZqbTIU0O0c8mp6wcB5608P2Ky+
1swHv/dbtfXsYnfow9oTiMzIUYv4BCOtLy3aGqfUvqVpRaq8aNGdj2xyIHByULq44yPak6eGJSRD
nIFzftO/t1cklDjt+eNwQXk/FD3olcKTMfExqUvZkMH2oVGNLQ8sE77EH99o9H2DPHSZQHTs//vh
+59/6tfYJOC1L1lOh8jSCkg0+Qwt7GlwRcYty0QhuL3Okcvli5cJWTitBIlvpPi6HVtMerwbAjia
ZTZb/5omUJxNReVeftICElYE7YgHfCbbFVPYFSmzF5QDjhWMz9kzHSBnEjm1xDK/xqAp8hsEwmsl
K2O9chzaR0FNN0NOP7p2TZA/rI7M0Qg6wHgg0+9H4KZWexQn47yf/aFnBWXWN7qczp5sfnihysCC
P0RgT+RLZbKinlUoYlKPTJRjJgJhmFEKxtf4BcbW81Teb53oRrPUbKxGjr6q9t5qgr4LzLVm904p
W/OioML5Dq2YLXsgrfHCY94+uWTYgM6xaK2t0Gpmuyg1JKdIg/VvQQpJpu6s74AsFJuhVmFOr4w2
jUHx30NRByuDi+Kf2wQwaL4PILvfDAQ/PuCHIWtjVCqFQIDQaZikH/i9iUATbl24sEaq9Zg/77ZX
dfS0cUvuZzQYnivqW4fiJVKsZf32iPVhtaC4pRL+g9mG/aEQdXMOrZ8pr2mI/dSeRPiqZdHk6ptr
xjjm9RmUdjsIp/b2HcGMX2Snf8XIU7lUs89JNCfALpmLJgRvmajymq8ifxLmotQtJLwODAm+Ship
OyzV7JsV/aZaCRPz3qjDpYAHXoPq+mGWDelKx/P1IvjobfhF14K3mGtHvOcc7CzWbYg8sd+BLLUB
1sMS8wtqZI4SyTNx5FbK4Z4tlE1JnftVDPzWTDYfqlyfdEUDoOHbHRbnqzi1c/+vTTTM46BsbG7q
4HQuUaePo/l0IPSu2hlOYJXP3sYWydvkYa+tFFNzJhZRFE9dbURI9KtQwYLNoW/0vCEMOJs7C2KU
NdsvvrjP/EwqpE7TDngDfLUN07/fyY5JzYHTzcvqxFd9Lj08WUxVMVpB6G4JRh25nt0jP7/TqhVI
Lp7DjW7OovW8twRMhuE4yI6NxmiLA/2eyksECALvssB1BGN58h6pk6s0ZX0r8azSWvMO/vxZvNYL
5EwUPHVBLK0cQIqbkuhPHy+3eNi7DPdmHYcQNhGWERh4h2IyWkcR4MWWm8pFTwgYQVvqIN+dg7SN
5t6VA6RegrFia9Q+zJv51AoiecE5TrmlXpisuWlSwqAVdzRKe8zZcaEy+HdrWu+JD6k4nvgaB2V4
iihu9T/D9CugHLTp614jfUFWVD5QKgeF92hrpbvq3qw5YW5uXYkqe3zXnfydmDC7SkK+oLsdJMMU
toejFVq0aWRlECNAdtjrXUqgXP8jD7JcSXzu07xrvRDKNGYLHpeb8nd+2d9DAcsc0NGa8lS3Y0XL
UlXUhFG3QLh1TcW/fw1c1lJgV8g79x2J8Glxrn0GhTqtFoyzLxfcbHsGGdrk6aMyUBRqJflU5Gyw
Xo1j01LHPMRIEV/W4U6UPcA5bsO3HnAya3XSix4xNJRfR5M9zhHmZw/UnVyntYXww8RVVfE1POMw
ubv4PM5wh1OnvdsRu7r2WDjpyzc2rKtuiPARWlhQ8sXYMGNf97eRUUYtF6vY3f3gmpVvZUtBzdR+
ce6OsGbLJQnrfK+i7cmsKM6ExU7OgP2bLJdEyZ4LEOb0xOkm7jpNRoWr+rZOnolONdStBUDzhBU9
z8dKqCWd+fjWIdctSOX18+V+1XsGbVm793v9Vo1lSNXDl1VBJzrn90sm3W6mnbW5/HxFLa/nsAK+
HFEfb9DLmBk6us1xQM+JDde+bqJvqyuUAExcphn9O5djr9qTAerZQotDmJFHh4G0drBRem/P0n2V
9ITUkSX5OXK6D9bjbAWG4HQQP5GO0g51uKQvSFGlStPRP3PBFBVGbPS9qSMxs7nR2gbGhvDNA07R
CVSTzm0oXz4pa1G516U6tzxjNuMwjNWdz/RA/9o1XqagaIsgzw+SShnDgc9fQ4Ma3VmvVEvekD3N
UIepwmDMBn0KSxgv5wvMrI5MrvAO33W0WRtSPMSGl2frx5v4bvO8tpYiH96ByhazQJpKdoMO4ciK
ZxU1vH2TTdOZaLfNn1RzeXf3lInzr5smGFb2P0e4tsiaRWRXTl2CJnkofrYtKrnpu/6izmR8o/9w
KTpV+ljmSz6UTxJu6542S93hJfmRDH8GXphfme01qkgq8F2KqEigoXIXeGaUlVmnqbHovAnmxkY2
1iW8sgzuC3sHikm1sMJYg28jmpglj9STD1ncatWaS2rJF/I/9kyxQFxJeBSOsdlLfRM+ai4rhoNN
BieQ0hSaSgImuVS8ZZmNjcpxPavMHobbytM3Bo3zvVG4XuU5Rc2BWM0+TSBI3qTTjHoISR8SNbBG
iXJuT8DWtT4PT+lMWY4Ht5z85/GuhLGzNCnpVvnKoKMdCVt9/dPF+LogiO96OkXYuSerNfKylvYZ
XovmwYQzFdgHuQoeCJ8GudrxRFDh9o5KF6P4XYiLog6PvmPZdFPD82Bbc14/FJYcTCvLSexmWDnr
SaIm2p/R+Q8iltNYg3xnGXxaNLd5fL6w9X4M+YlOQTF5mtOJu73IWjLPQKEV/k0XoLz3vVR8NR2b
aaH9g/1uTdtwkBFOpwyC4ZOJSIjPYmiEUusjjvN2MQAI1EtqN6Da/0YtN8094wEEg5buku2lfnDr
AvFpjHLvX4ieJh3L/jjDBZvFMbv2fbbQ3qUw66Ed/LmbPMsnshH24bisyGDJQyGR6Zn3z5qAWR+F
ymXffm25fZt3zFZwOIVdQ+UpMoIGu+6L/Bs3PT1Mbkhbj0O5u2MC8vBporHI6O65P1Aec+WnXiT/
J41M/tYdmugwZfPv2w44Qcw85NsfxAXWqn65JBJAesGnhHNEEods6hxAWGWneO9Y4XjlV3hwuI3P
1UqaKpcQTF6RkNsfZ/ZZjwr5fesjSQBK9qDdeezU8zB4CcISP3Cow4w1nI/LMqoTVVuuqu+A0cfV
JvDYhn1frfXHKvt7+3lL+dbJnI68Yrc4i4CzfrSMQf9e3bMInigUf+8Qc8u7941mPvPDcndMi0Ad
aCV/OUxqbpfIl+3JuiMh1RNvQJk8dRvz78NT7cwWGLZ7E6V8WBqqR5mU4S+gh58yrvfa1zK6xzHm
yGsVyGM/ZBO4Jkgo6oJSrdRDb+TRk0sZYwlSzISeese4QEXtNngvVBWLFjoY5cOajH4nbiagbJrZ
Oh3YKSQqwOniy1R8+y0dl6Z21RMs7VwDDi+QxM2parNbXX+rmf3msyazP/iawj8FjHBa2yzgu615
T8uaYvanwFWglKog8QvDy5WddYd06/o+4JK7Z1ecRSCuLnwFcb008lU03TqlpLTyxZ+jhJny0RHO
5CcPcbE5uimt/5oTu/Fm59D0EFkBx6fF6WAHB/4m1lpenPH7fibUpQPl6nvSOnEv+Tb7kPFAOb/t
3Xs0brtSyeO3mbQMLnUiFhNTFcg+UO7853ZE9Tn3m9HAniP21mvFxYBqGlm6E4UQ892ziS2juGEN
ytkkuLxtJPyDgXiWZdVHshPOH/7UQj4TDmf6+YWRex9xKjJVhRhRBHoZQHpNGp0vAUJ/MLIYks7d
0Jo9pnK44wzVxvNGapFV5E2cHGHnkpIhj5wiVDeQTXW+J0o5jbiSXdmf3/WZ5i/Ds7RsY6BuvRwO
yqxr8p9CUHoCBcrgasRoMvD/xtI98i2ObSHMX3nHYX0jSVQF53AXdzJBjkwlZ0voSqQaXz837Zif
0IE2AtzxvaX1Hm+3RB60Kj12Jxn8Q6IERvFW1U1i5YqJLTUp12oMtVgoSceh1cyRmjTe3OwImpvj
1lABA/ohx49accECnMt3wwiqqHRNglocOcys+90Icv0eKG9/0PbStVt+WIu5QZtOr3yJq48/rgNe
+no7eVvTv9dHtlkEc9t669iKS/Pl9xSQOk1DyXlidP7/0RNpgZ4huq9xyDIFvl3XD8APFyCIK/sA
BC5T1XGpADxF46OVXC5P8kJk4+rntMiZDLPbqckqlMGaekY9gTbr4pKajKYOUBVSchXDe2W/D4OY
qRRZLE6Mz5KrertqdDlv3/Hj/OWn4oD1OvPvZ41pjAHPhgP47uAg2x+HQd1NHty0RLVCiACt72SQ
esfnD5JY9p/7dNdl5j5Zl4tZ6s8Tr6Tj7fSLJChXPHmXYE7ec8lyLavKM+1iTgR2EnFzm96W9dUW
mfbBEho7QyqG1CH2y606A2YiGn2xX/KSer4qufMTOYMGjYXQZqkRBJy2B3a1urKRS73GcEhy+8Jo
qE1wwkFrE7Kc2gKuBsXucQa34O9mJuV5TSJkNQP1Lv7HQc3Xw5QrO/NkLH6Vcc/bTYs8X/BV5q4X
rXq9wP2EBMWARgk2U3E+WcNTpfbyfmqXLGOmapvxMKMIQpeQ8aNcRTgUqNcKBTRt+9GUuWbfXxoK
nEVQ2wtxCs3yXA9/j0MkBfSHRtZu1gIYX6CJMHsBWfJTXcXt+LP32SAtO2Dzn7JqSeM2fx56N7OE
S+gzMkTXAykdVltqPIW56Sk/6OtSsnIQ2A5O394IKy9HDyMLNSgK56O3M7Rwy33EogcX6WzT15oy
RKvdv3+PbxpdCN40pBektCcq72FkJY56vSC9Ywy2e+TXQdm17jhdvqYG1TVf74He9WepxixQkxi6
m6TPO5fiZw+wnRv4JCYuGl/GBQJD6h9HZIDmfV+1HrRANGX5EEJ+OQl/QYYq2itl7WAOwiQFPn+4
379+9zZ+wjwBPax9BdtBSyp4vGq2N/exW61Yo7xNi9MNzp7tmFohAyOToJepDOgJzT+HJnQ8lgjr
MSdv4RfmHz1NQOImmaKxbBoV/OFnUGZmvdvgQQsERXU8fuS59BwR0CyR0JbWZuP+x/uqzWqT0VpW
Dc0OgSPAaNq/i4XJipHGyUfT4Kdy7JYI8mY0Z2TfYneNXDIQeuF9+Eu8Y9hlWo1Jbdcw1zbbSg8E
whtxPkdLgzDOPnUi0C5MIh0Ew4CmJ5Caasj2yI0cU7omFAiMAc9re/RjOv8TKuCB/P/BV4yzsVKd
AhPThoCFU/YuW2FdmIEdSjKVkfEXFSOETeLzqn3L2aM29Bvf7CLvBPBVl6THpQ83IsKsO3b+wrpu
gmVJhYRbWF5zAJwWavlMDlCv/UpEtXDOnnO7A2KSUwdFo3C7QNvvCcpqesai0pgFjyQHl6ZjSRjq
hXeruoQbNJaPT3V5wc7dYNO+ctw5ivAm+VPtxdgDPPPDfMcjo8L4rWuO1YjT4nzd+YsfEyGgSHac
+GdoYc2ziZbqP5wnToTty3IIais8L1TDZ7HB1+TO7FhsVLUPQVPtb3XrwvIogwffKsBuEHT+Kj7S
Nwt0ZCi0b3GIgljcz+VIt3EWyDti2h4GhBTGae5PesjaQi93YPaa3PKiikH6HSzTuKtbIs85SfEt
Q2C7wa67pMwrDsZSv4L+apD7Fjabu7Pz8ApElg3cV6rb5kkkFU3VtsF7axxafzrSxJwERjqx0G+k
jgcURKWpBZFTsXxKrWMVjZM2cgRU2xj9vFllQpndw1O4m8MHaVFsbxxQYQ65jWxfB5xDqwyEN57+
Nmsf1L/qfa+J6GwQvlkEL7youCP6uibif0oP5+QSUEBlgrF24jKHLuwghh9RMgc8Rqw6+LQHPUYj
YoezOaZsDKEDNaA0LHr5xYqWAUfcm7QVvcicbxcBDfWCp5M9vb51yatYX5sXaUQnjYtipU1B4S6b
OKpacUWuS/uP8pOp8zagPOhz9D4DB4Ex00hNYfXVKGjKVrJN181q+ax8+XCXH13s5qyZi/5E1Gxs
iDWCTIzW4epot37MEighOvdBcVmwnfsh+CQ8xXLmdqdAs2zNyBiAULvXZrwCFIhFJF+mYTZEgJSH
PFLWLJfGbyGHR7tDhAglv0iu+eks2epDmGgerI+xQ6JYFRYVjkhTz69PxCgIx6HDWEo75zkwuujh
h4HZ4kW4VI52Yozoyfpy/MHZ7pSGD0n8gpjPoktxkWVkoiRudXtDJv60Hi2MZO9xqtfQi1ARDTEs
PWcciZ1aFIFAD1VdfnrEsffFwEdMnhlHZsVOrLFjb/D5PslyqmHay0x6a7ZBKKyadYltzkl5k791
Yx/cECc2ROGmnFPcQhtfeCuzyWHzjwGzobg1b9bPIgtmZ/owSXY5NraurtRseepf/Zb89gJ26Cae
8bIFhhay/L6giINsfJYOklz5ahna1KKwRBz5J2hminrp3Chy2SFN0zp8/fxeWCQTq5k1AkmXFUOD
5A2CKGsgpbFWwzcrBVMRiQjVjr1NYFvySpUMTDV7IOcXeQaJ/+dKvU9aDfBr7bu9Ootho3ICrnXO
N5blhihfA16C/wB/Z/cLw1J+u0BSu+sIE99aUy71X1sNmmDygYyBAjraFQRkxuanQ+BygxxjJZTH
H/22zfVzhsF8iib9dbSzFaolUJASqsWzywq7PZrHfFcB5vdBw9I/hZAkUVAvz5oXZjyhJ+InYZoq
EC96Da6DDSb36LMOVPglytLJJOXGurgmaLgCK01LWNzUnbtPTrmQuMVm/JV4nysBXid36VtGIwdI
vQbrxJHPG4lGngkmq+Mikjxls+FkSSdlSwTlVigyFlpxYcLm7VGxD8KBoGwM5EysJb5BW3niwlt+
fWekVneEl/ZBbN18rnhgUuvGoS2LjMWCZdqDmB0vV7X2pa4ma5pLMl3Vw9tWb5Cz9vJk/x7GetzD
hDEWdzcwDj+2mXADwcP1YpmxICQmvRwYTYsOOecbR5a5eDnQBYGI1qsZ/RgtjbW6e1dooKlDyi8V
pVTxHy4oEgmRvPJEKCCaXYS0/P+163z4LeLPRQq6F9RvdkHTeQ2FlubMjSDABIqSw/a9bB3u2jtE
4XprMP42paiHfAn/ZhZAEqeRnyXIij+RrLP5gXrQGtwl20lEb7gKSCHZurFuTV1ueSmJkgXCAiQk
annYjpFlnGxPU2o6qgMZgWMKZToXhZdl8sH5rmmvWJihCMOar6QsQlgSw7+DYA5k52zB1HLBNsUk
cfdsVI938cYjFfCswVmgN+T1WpT0IbOQFfafBQH4h82Cqcp7pX+wimhC/VkYKzmF8jUOFAZjDWo6
dh+XJm6nYRKpcWREK3hRumIUFR/YuBeUKUHZdzejrWb3T1WGxtx9X4qgzBQPdp6G1F/HJNfAzN9D
XDcYFUWFW9PawliyWSOBw5Q7qki915v5VyDJDr6iGC2+1T20pPZbI3CmNU7394+54OM3l61tYzFS
QAM4QaNpVo84DpxCTCAhHK0PDhthHUXihcV3lPpUibUHWhpVmxZcx4BAsD/vCGSLXtywyFcNo53q
y5N8F0gq2ryJ91kZjwwoE7h/8wl0cb68uES/Apgljl3tvqD3cksc64dro3TBAVCiCLk2tdSfFuFb
i9GOoDIQ24/02Xv/g3DQaaMbCfj42/8sZ4tPkPDuF9sfeGeNWpX2bILCsn5PZjAXqPlSXvP6+D42
4imItraf2sxXcrEQPuB7FyPqwgOOKlLJS//7p1VkDprFTsRbgQug7sjWFeKWLOmDWjIKxyHP7klN
x7b2MJjG2PlEX/3MCpfme9ziX16MjWVZTfQr6uoPybRxFaQIJhLRZF+IrkR4TvppC7RXTsso1xuX
NLhDdE1FwmsYuMjKrJ0joJrcolblhm5zHb98hzh6NEufBxz+1jPGg4e6lCdVBsqj+oczZvBmSEb0
xYCmUytAcyNlNK9nY/RN45WhMJtmsD4lPz0VRB+HKqMHczu3J3HlzQOUR/Gq9ceGRTNMjeRWIKr4
GhGStcJTqITf7t7LzY7Y4pyDtjkDt6F1v2z33dvsjlGGDticsL4EKmbhW9Z34orRuvbtuHP2ptNy
JDa7WfRiKe7U9FTgLnLH2GnOlHvNySvuvs0UpTBMOVVrN8b3yAmHMgRD+gG9HFYYlgdyzbGzhwp4
BWmNH5ByBCQZcGMW/tGk95TMSwY3RapO6RpY7H1b6mZkvArFOcEIbYTTcN4icvAfnE1IBDpIh0M6
igNzS13afV64u+C1OvWfWQOf08UR43d5GL8nTE4BjZOL3EybRFQzNCiEYLM2u8AgYTrJlov78ayw
EBVJmMglBipRbkMRGYEBwKXP0td/jsIFw91shEIm27H6G2cW+4C3JJDBPif0L8tLgA+/GMbgYQYy
QCEheJycbkFnI0IvoGmR7vS6lQ5+Kr799Vhf/pEIiLfwL0WGFroWZHMCSwVOJElp418lsRXtyFPw
qHKRHSUoTxHqKTHp0m1r1OcsQTqQ4rpG2nGFEn2YnCtxjxU10BrDBgjx+IHj9jiyyfO5cfpCABUg
FsOf6CLfDvQIjs2IGHkTfYh4PP/QgRHhzfrxP4nxoxfktA1kZHhlyuHSbrZjaV5cLi8L01CSUSxJ
7ZnTEAL+ZgmnH4rTNcZLlNGv5EcZ8MV0D1lOmtKxz1b8EqUbVAuM2w3dEK/3/11Dg3H56n6S53VA
fyppSoUSfOOIS++wSd5bMiUjLda+trxnfVvB8a3yh4FCxVVN2c2m+MKJ+rkKRDKFznqVLb8YBrUW
wsb8qVWVl2v9Tq5SH6FG7MPoUp3tso7+/ZaZSU/6SRDguXApHACaWuPxXtKwLGi/BKzHcNdxwf8e
4J9BPrf4QKB2qlDZA/PpHJsJkLwzmanE3vnNrs9B5yj2Du2tvT1TBxTxGLicoYzqBJBlfLvlOigb
0R41i/oX91XH0Q5CSjMN+wqD4juppoFOljY1AqTzqimC4jRFR2TeiP6HkVqElnFQsfliZZlZegkn
wBYI1BeycICz+bBJFjsh+hNI/WxEPmMnglbTInfbtsXK3t+hdqFvgYOXJJeFWeZz2+oy2+Q33Y96
8Pm6baigqShVBmNxLYTku0fIxtfuSsU35d2YTf8WxgmgOazAWgb7PKaE1FwvTU1wpatCiuMbsN5L
YgMPgjE151IgcWc0fPiuU2Q8hEn7SGO/bqjzjalspAUwrtD8alaB555thqts3+ZzJ/INfBsZKuvJ
GDiIp3vfSb1nwWl/jGFYgRWtXvyVaPzXS7GOBlfDsV627DEBuq3iz2zKHb5fogbeDPPxX+cz9pvS
9QsYUsD7pmQ7PpzBsx1DwHBzELLFOumHO7kWEZ58MwU22phj6T+L6DVnyj8vt0Br+dkc5XkO1JEs
f+uiwRjhS7gK/EHI/5Vik9k/NkpdKq1Z5l02AApLsiXH2ad2Xy40NC4X9/NVWPr2xvRR+29hSuLS
51OTjP03VSIjH6AAaKRCm3qNtPdJLfkFY8a2nz3JRgHAWeQpRrErz1a9zgC83XMd1Vo5rl3sJaBf
j/fN/0pC4dXDNCg1ZDT7g9vIkjKp12MIMY8c8NW100rDXj1yoTaE3oUVGpAW2Skwzs82HCooId8Y
Wp6DqEWN9LP2Bi8+0gkUSqPtQHQsXZoXx8tkcbiirumw8NYQxU7+eI2wj9EAwtxkiV3rxoWKFqIu
kVwN4/6EcF85oyZmLEme0A6FzqM6LQA1ZNAbcsDspr92wCFb5RXz8yLek9nd8+R+ZvOGoUk5rQPH
wUdvAlGVeCz/I11DTyVOfBnL+m172VqQXptX0vBe99jPcS26aeUxOkcb5vBkUNPR4WptcM92RCUF
IlVsVL6O8UaFj6pwZVV6JbJj1cgaj20aJKk/76q0Tv3my+czFUcT20Ew+g/xOLzjqzJ1PtbkY2qw
K99yBBrc1KmL4Bb2L1J7VxBCpz+B0ZJDd606/gRwZVysoHYXF/uaRpo9o+ghabuKKXjGsbV8kLn3
/GLq1s2PJu3r1ff1vQG7gbONXmn89dbF9qXTj4gXcvc5iD0qNYLM1uobEpKnP0CsGdWJPoZ5WZcN
EMWhNsunDtUJtXEEUTyPmxD4qIZ5AYDdALOwFC2Q+D3jCzyc7B3e/TPBB78uh4gVg1cpl+4ra2dC
MZ65vfeLfEy7xdha9dVx/wInvncaLRBw02L7uZruaeF+3XCePIHOrVRnlg7Giw4NWUhqGEkB18qU
BL5JoNYELY1z0C4HjHXCVvnWdpeIqWBUprpf47R/SKjOLgXWcujtxq1cbYEgVNI9DB2+1KWHGiuF
JcclPMHX3Brfeg2OyPaV5HWw3O0dXCPFmTBCJI09M/TWq/34l5kRnRMfJ21hMig40B3mmFZQO50O
wOHXCkzYFZ5QK0odfAAEeocNidk9XzHYF/kY7ZHe/yYrz0XhUfsOr1wXAEcwewbWl51dVAFEmZvZ
Gq6KGfNhRh6vIQYlgz618kChxLrne1dFjyadUsgvkQQouQHouch46089+xFZdD1mKS14PF8DWhbZ
k5CzU9bNtQDPFM7wtum//0RcvBX4l772+haw2lKsf+DxF7IMAXUYjFiVLHt8zWeYi1LpujWjP65s
kHVnGPR2AxfO6701NhJqrFCgAnSfRQ0QQPwJh3BSdZTbN/gyCWnd19J8KHiOIj41FuHxamFiTinl
cegFjUi7LIf62QgD7fDNqpsWTnrjc4E1Fws711me5X3Ud6NJP8wypilozMGY5c3nL710pqR16dwc
ZGio6N31gHT24wt7SC4DzGT1DMEzk8wOGrU8QvKE69QayoQq/5gmYRRKEW/D/OgPaBPY2YDwsjT7
ZFGQ4qj7sfi73V3evcZRVs4VQ2EnG8hi0l88pCeSEmRGezXgoA377sspmChlEcbiiPvayAlr0mr/
6boSLUJ/6mIrsCTouXXehORu/Pajq0jVezJhqbTl7NR2TB/2i6AJPd9NPYxGWPydhoE8pdU8MgkG
9zDo/i5b/5Zaq95b+jJFr9n4pXYvYh468JJirYo3lOQ4LK1tbruhnfEkX4B/b2r8P2xDkE6v65rz
8ZQpA+arT1yHTEq5/KRT4x6803Lu5MXzeD1TlDdArI2AEGPjC0HcWpxZqlJzjlPpSguLnjhfrj5y
9kBiftClQ2Q3rUaBV+dqtBjbHphmZ1ScrGvoZCFkQYQHtnUDC4GEcnlF5FaZyLIvAtIQLlI94msY
FehHc/G8g79BkbnMIn2nciEM8IHmHyb5uNaGoixgKMayLLcyIc75fAQPZRW6ND0UmxBaNlBALdf5
SJyLnBHt0smFwbTZsZZOr3JXYF0dMpzZEfXkp1i4GAPU6ycHW0MxiwbMjfNNKvAHwF9Nt19xlYDh
8e/xuzmDoYCvgOrzY97ygtMbLsVTxMfFTNr/iQEIelTNLPa3EqotW4kyrvtq0K47UWZmmfPUA1Um
HLcSZzT169tAumFfLo0S/LXCBuVyuffZ3w+FWFizRdpCMymuKxYh1fuFLhjX0j+sggUGfs03aNcr
TGRZP5O5jWeyWwCMGcSwkS2qZakZxtyRS6fjZQIeQYoGJTGQ6tcylCDcwAkvm0e2E1V00dbx4585
eIdWJ7OWMeIGRM6EMeVpYSUNbCjNqQVQAuDiaVerptC+HqYc4OkSXJvbP4RT8rJRjw9WRlI7DVXE
tEFHG62I5E9baUW8sSYbcKbR3h7GzeJx8hPiEfva042gdF04/6RBh3oK6EsMRqmyPGq9L9Nonkr/
CMujoJu0PHSzvf8sV7307XpevuYxZmg4APchEjUgSLPLSosgyhV0Syr8q2qBQTvFjMchy5efPhP5
0EZZVrmtn+aa/FPc1SlyRhiihtd1Zinw/mSDJ227xCr+PBxvD2VWLX3/T5Ix1i7E+MachlE/UWlR
yX5Uwn5mfFvKLms4i9juv5DWuvqh+UFw74egmrEG9zoOsKS+iYZdooFbHRGY5nok5Q5aTK3YnxsH
i+xCJbG8XqKxRS15XXWbm2j1zsDd4elkLDM4hqun+aS5R/wXTOslSRJA6jKuToB0JjB5Ys8dHcxJ
6nGfrVBcNtFPBS3d98KhIKnoUhMRP5JBaLRKoaYb6EZ8BG6uunJjotjZamn3wWBjHIjTz7oXpqpt
IruZ/nhwOo0wwboY3ZYPGOXVfgPpd6Fx/Rtjs6+VG0HmnNTTChasTuQ/CSwZzFCfLXfirQMMrv0A
Mp2RvXPiXK9g/rUPoSJ1vkCOGhtlZ8FDt1cmGo7GJFQWXgK7YKplFZhtIF21FSrf5GpJeOiBKH6L
/z3nTaPJ3IgSZMVAhbQCI2RMh2EdIUvK90bHzswiUPtj2IN1maPkY3Cc0v9S2ElD4b35/S8QDs0t
GLZq8IZnIwcn7bTU7vTds7ip8I76UQq60RNk4X/yvO9EsIFn88wBfY2vVw+fAvTXU4yAyavsZ4/a
/LZ7N9/DHfe7UgxnmiydvaOZnMmVIVc0rL6/DdTk1OS/EFBOXMlGt/716/YKdE4ANIBu31QW9RvI
MSmCYNiPP3pQ2yRlWSE/Rmc+ByxAEvi4nTJKQOGREsWToBNc2uM0XVtZqW2L8n7XnIATP1Pfj25p
sf2e4mHs5W/ZH8akqkHsv+MqznsFfXWWjROkLrCtSJlWqd8T5+5XyxeQrBVrjOcUrWpeRRtqPjZ1
OEUgTuZMyrj/xUu+qlXyUR8E9lqqkPh7L33sdzUz+mKStE93gTKQSlE73Mw8RbbvjuNXhlVFJ3xR
iqig+vvdJEKF/1A5PT6WZW6pk2tdTxVpD/+sg+SCU3nrCWEMqv1aW98SrfRSbq02KysZI96yN63i
OELWf6YbW6Yfl877DqQIHOkg3c/X4XiT63E6G0RB5VZC1xCcRGMm6atszX8lJfZ+vBp6Ujcf/wmU
tGwM59JaBcOEvoGbwIPR1+QlBWU0HMiAPFL7ejHbAOtznR88emyprtVeUP2rNo4OWPuR/eclkjRu
EAn1rNxBzFbAawhKEF3qJ4TvjpDQ2i7u60BgNvsbprM+ish0Dxo98RmRg85sdL84Rm8CggYxLT7S
Dm0qP+bQdV4m/Ak7gdWyZY+/zAp+ZgJnflwpb/5WmoQIBbH2maYYCREBrqJeQZ6Qq1atoWQ7QBSZ
N65VOwTCi/SWSCLQP6S60wEwhbT3EqfTsttoFQSKDNuG6z4jEVNk20Wuxd10BmchvBCQqnM7PZhB
15pmx5IxQ0H8rVgdeddv0/aTlsynGntM9vBmS7emlirDJNRflgpgukFTo7rlSk4g/pnU6MmqUsS9
knhnHogD79o0M2WZMfhWVQp7X+wyEiQvFb4BleDDqoB7deLiwW+iMtlqo1fuZXR2m58xMxsnhr8g
Kwv/VxZ/C/S3DyLvfcshDLBKlJkoQYfIZyJ0L6sUoWWD47aOI6+Pb4mhrkbH2GYDbNy3R0tS+zFp
FrsqvPRNE9aj9SDOUJgYyQ0yHYH7Xz9poLZn0PuCpmjydqXJP7QvfcEjjcp1ispT0i47h4AlbCwM
26gTcyrZYhJ6anoI6IYcJKMJaG4yu6+IEjqP/WahjWksmjn45rxVbwTq6onBKAZsNIiVa00DSzy6
HzaN5EZMf1vcS7Q/Neu3O6DFUSVWo2yFrmk5uXkAsy6duFfE6VEswXmr3MZFPCs6AYqGxOp6fUo8
AuBzuv6775ID3dlxta9SoZ/BXsDqUZKTU7qsZHiB5X67z9hXIfQGHOuudXKLXbVlbWifPhACP1Kn
wIOXNLqj2REZ42BHc95U20qu7U+TtVkIEGnqx2qh6LewaM7XblUemc3Pm6aebLErRKgYNPRLO4RP
bFy8yURwFcCecgV15kaSZX8L6XsTBQUlO+cbIrRSLsQzdrkkOgfNo7uBrQpV5YQKAHWf4+GAP+1C
GTFJrNhQ9Au958RwGTj7+oQChoewxMl3c97Fr/0jJpW4mDUTdNbfXxZIOnn6NDh0UOKC/iyTV9QH
873Qjq3FN6NSgWpKy5xPEy86TyLW3biM/9CbWt8nOhtMoMSsCbq25UgHbw19dxIwq9jwJKQCC9vr
fEkYsqevKpXCb6lTuBH1Zb7rcOYUhaMphRdXEgn6FfgbbBRQKSFGJijPQn1OYxbgjTdWXZdXYxJu
8c2aDl+ogBFHfzy00AdLThx8L/TsnefxMSy9L6+lyCd33nzw5OVQXxhYsUfpO0HCX49HA5af9fdW
53X4gIKtd0jkhufJqYeUXzfz3eCGvYdQ2oxPGQDiJeNVxUnJfBwwS12b/q2ycIlHC/VpqwnGcTiJ
svh3mU69pf2lfie5/ZKGlKFsVE1vmtx7jdhTE1o8ewnnLDA5EITQMpIJhavoze13pc/EVCFNOdbh
xmSupAac1MpIpv5nuI6KduWWA4TtaR8KrjukMlpmyDFq7gJZT5jdzsAn3cqY46BlD8cPRZ25aBdT
+A/x9gskGjHerU2ce2w1geGrFIfbjdH212ADeBdV7XhSbiQxEyLSac77WO4wafhlBC3f36uyUksk
gWJYeLGHP65M36QIgto5s2H3bd7i5oXBssELLgIkeKvZQsQc8d04sO9h/XqNjco0ucNn5q6GGeoe
VYXVSCOOaLmcoDKzeWks+UdgRM5/GH2XVBmn4lB4Gg7QYnkjExTv/a511o200gQCEKLX9GJUoblQ
3bz8VeLkKmNMhPRYMPRT8VSRnwGYMzvWDv/OpLco7xcXSaKcY1tWm9OJYenkT1jt0ZqOMAabtN7d
wxlx8DxZwwlHeFWCK4BKN17Gc/sL4yc0Y1d8y7iQyJZp+AJZeZW3HEQ5KxXMoM/kHHKDLvhwqXgb
bPRjw/C/yLAv9yjPPXoN9lYEFCVzsxrFjUuKfTORDTeilrBDKCw6Sc3EiUEznE9g07WtMJyLDkh5
O+8L2J3pmSTp7XbjBTIubmTD74DC2m2/dhumwS4v4GpGaU3YXTUD8yGuXM+3ZGYwDDLtEor3ArqV
cuaezhcUbfWDZUmDGyAy3etKbwihLnFFWb40Fy1zysL5Lzm9bET0c/+WDx/xHzwfMy7mm6Wvj+cK
8LZYtNOEUhDzEMSJLgspSEiZGDezXup81TrpzIh07T0aU09b/3ehzsAi9yd94cdMqzYBNlmNYWiq
/UlxYYfuTELnBVLGkFPXCNzMmxD/cSsmwabAi5B4pcoFCzAJQV5QBSLJveTJI7wxZjMFWdIJiHNE
0BrN2Fxvdx+Hnovb+DJK2Ig1fS0zfqB1xJnN7eijdoybPnvOJYMULsEX/B8GpER6nJWJB10fjCqw
x8iV9dQrIW9CQ5ffnOdOmeUNkKRqluTEKIlvv0Uwgrc1wBYooq866b3TgHEsX3u7vcy17nmryvEU
6TrpfziFyqhCMYeM02zpLsxQAnryuxqHKDruiRNliZXL13hrzA0StirKk5fJP4c8wJheA6Goq073
I0+LupS5al7VzHv9odyu5YPeT+Uh/x9Af3cGtXuzRwN4vN2WQpWCCUK714L6082SfuW0xPtHuXSQ
vrYlbv2c2NESdid0vQt+JBUc4zf1DomRl1QgQauNUf1supvqi6eRGjUjYTRYbAvA4AzWLdoVaXcL
yw3Wt0+0RwsPqc5CzoUK7jfdr1ftGbPSU19io5Y9aV/4ep5VxVms0FXszLeEBeqxaDD5anC0Qzq2
nJRCQRhmBIdPic3vKNICCeBynRoAcEXoVayxe6sslPA2A14Rg2AVdbiGabE6Cb0x5kUdEZe40pnk
x4iOPa3WmmRphzb6ViPV4FWiYm49tEhJynNOz6ds5QCIeCJRKuB8aygDF1mAzM1VMsZddfT1LWuA
+bQg+01mnQUWSd4rPmgjduyRORL8pk7mEdb6x3THXJNx17zjCkPFxXdgvBU2zQDMhUOEAG53/gDT
fz/i0/5Y5EFndVdo1UEYx8mGZpmtwEKCVX7sRUSfQQ5Kmp8eCRGc4wBEkVRAiQnsc1m42NIefig/
wOZEtUiXku1Q3REMpSFlqR1RVnT96iXNtxJ05Y0g/fow6JSwXnxM13Tk2klmQ/qUU8AuGlfUVUhn
Fjb+mrpRq6kVULLpjZ4Q9ETqSvvK7b7P8DEn4Blhw2lpkR06MTN+5Zl62EQ/X8rdoY7J5OT4Z3Pn
ZAI57zg8RJ6vgeA4M67XaHc0bpzk21MP6vfjAhK2b33dKJYSfGGwS6jeRgHAWcfdFSWfh8q4hosg
ZNzlgV2lImnGMlxADXFhD59ZNXBFPMOu0c1aXaMNKGQdtlwQevG6CxYNKdBJ4zcwzgsN5f8t7g5T
jnBE8w94eT7j4R9cGdeT7EJam7B00leOuJUCzXWCgYrOdFPAjp+aIsMYxPQHIbi3d9tmDL0qcZ/I
6OH+VCdgIJkx8yWsimlSg4A+0IY7AZvDDEzjjHNouRZm9ueacR7XPMpl7negYF/c1pz2EgPy3+M+
1w1QjK4cUS5BvtwFq+keijJYQRDhwcoKWBAmz8LwaOj0u3lwwFhvUrUFy72/zWn8PzJq3zvisLu5
+wdGIc872c14ndOLOSSXlmmO3CcEFlzpH/u8o9eO8W7+LgaAVf3lkqkRDUfW8QThO4/vDQdN+5O8
OJoSjGmyZysiavr1Sa2Eo2YpnCffjCMYpT4iuIoHQD5+klcdRpCvtjmUUmLsSzzt5mgv+i4HOpwh
TQDkCWR4nhmzVYBeCdCD/IL93FvNfUAdSH9acit7/0wGdmpnw30vp3jFN3vk6pzJFJvN+9PFn6oy
G0oQSfbirJK3/PIO9rvRKFwmcYVD/wKz6JIOItMPEPyetbhm2uDBbpQJJLYOWz7cQUOdhMyQ1D7g
ekXPyte3TUnTF9VqaZqij+IY10uxOl65BuSGDvsJHhMySbFp3ZGiXapOtLZ80fv8xIpphTKDpmVm
1aKUPQq8+exs6d5rSGR3mG5V9jrSOk8csM44j9JuMQ5E7tmsDhJyvJoEzXTzZHDpB8uOxcaaqq7N
9MGVTOWVfWRFFV3bdC2N2ia+AW2iXu01Tgy38PSguC86TSmo2u446vlOk3SI8ZtIhzOmgJR/8OzN
kx1zxi6yqOX1+CieeKrfl4kijLb7SEti/cm9UDkdjUIg4N6TeePrSCY41lChKobtJ0O75gJGkTdA
o4zWa0OY9yi8pg+dY3nk8/35J5USdAMsnTBNmyEkkeORi41CLKTOLiZena3rzouaYKq4NbTqDc9z
sIMoRA0C2w6vZR3AM93iNQ3GP/4qSGe3mwcGz31u8NQClAyoEJVUVNKqR+ls3TxAeZv79bB6z4Vg
t1Okbn2QxnCeEBwGzqINwLJhcd+pDAr/FaV5Kw2z/0+ziGu0agCYx1icNGXyeFAl5FBVDpXz6tOK
gT6xsmjUwGGnUmxE9vIChHvMKT+DvssJFIcygyRrf66WZiGm8442a/F9vq5wcg+qNsqLnyawgW48
0NuGkbS5PKd7nA/ZYBoaFASKW6ZyNvdUce3GJnCKXiI4YKhlyE1A/UXmLuqMoI3qUm1vdoUHUTFT
b9Y+sRq7be3ZI9csQWe79qI18jSH+nYbm8p2NncihklgSPWoZnq+xv27nJhqe6rCryjRb3SBoEvT
xpV8fIEdCX1hup5Dsz2MOq19A86JvH91EmtmPmR8QQGPrVcJLYf6NitHaYnnHJNerONryBLGdgpx
caNYgRRXT9+Bwj6iraDPtW517y+3PA3aWc0vvdRe0UPa7yMVJkAXXrHI78U/fhy+ZJaI8KbslhQj
lsP4AyiOt94FVlv5DL4jBirRVTkLJJIfWq4TOfOmLIkqIgWoMKknfSqw9A7tqsxWQd9AkAyEOz59
ZrpPFYnVpsGlJ0BRBfUZro2NjZes+s/vQ+UPdhI7DWSk8Flw61Ma2vDsJBDGXWdAR19UgA78bUsE
+Y0VZRT8ROWYrWxryyXQKI06M4Hs1S3lb1nZ1lsDvljhnV8Np9+enEUsO3UnAjnVJaAHyPJM0kwQ
u2I20iBAnen701hg3VmgASKzigQVlTaO7tVrzFwCO3Du8uk6N+Vx8v+9H9xom//1C6tzH6o4LOQ7
wT041V8I/P5yH/kHHGZhS06ZyvBoRtasYeZLIq9DlyFa7LAMLFikn/Pt55dcWX9DiHKYmN/5mazi
zkC4y4Ud3sgYkOyF/eqW+JL5dIu2z4MitUKpxi5/EHTQho1ofjpSGUlWcM3cNPKz+F5aK/G4cBBf
2uQTsKhrq8gdYLYGvqbAuVnblD35qQ7LTOrrnZ9EtkPc5eBA64YzlojHSS7MUNhrMuvuI5Kbi1oq
h2W2SIvqakS1QqX4hIZxqH1bZ9U9WENYsrUk3Wb9NcpCtFEK5/EMp4SNeN/WHXSVq52rWP4zTy5D
26UlfKEXnKGTXxD8RA82c6LOqNmwnUFaJfefi3hqbfJbSMjvlxQdMdq+FYYyo7Z6UjK7r+oOCKLV
rMgHA1fnY1EaLcF0sycMfMzJyc2rknNU+yZM7qQWAUMKI3LifWnh74qoTgVRJy/WmetVZg1ywfXX
Rg12kwhy8k9kvE0cEvvVn67mFWS807ioUDkkX11jTRiFdvQ3kszQ4Ks2xbVlJdOWFQiaJNXckUma
R6gxChg2KSIg8QrwdCCTb2GAafi7kG8sP+sZl47LQGyMRnjCmEd+6W30pthTsdW474wKa+wwm2EC
tndA1MDSWE4bad8Nx3Y6myD/KDfsMVxbwGUz7ZXqdaxzBBC3n/O8ATqzvxNsg0mZhhoXTUe5gMuI
Yj2N4ZcYayjy0mDhC2UIIbsVhgzP9X5keTU9DLVowq7sH67Ixg8UDdA6BnsjSH5hGtsYHEz01G41
c6WSCxnLiVxzo0iYO+dJFZHTfkKEIs98r8xgzIK3Fc8JWHfzKRqrlyE7xWv+v623Uh78lebe0mJr
Q57ILZYm7BgzJPTY4efdHNhSToFYQ8IHMnCjyc4GzrWXiREivGjVhe/RzBLDNMjsj1m7HTjy35Gh
F4oQdxwFTU/GcEH5UYcUhbzcz9GRzXVedjZlpBNKv1qDl5GXJ1Tm/SEQlPAuL0r4+CY2nBZ98+2U
rt2CAn8n2OBYhqATXByzSi+/IFpAN7OncHWl10hmm3XJNcrf0em/SF0lYz9JipZsfoKiQDpjUchM
w3OkupUD575703Q6cI0JKcQk+7cYT/Uv0T/l6yD0L1U0a6ivA/DGfC5Xxi4A6T3mUZ3RUu+Z3ygQ
kCdCNN1ULiu3/0IxL37/AQLcX7O3mcsxTL3wVuexP3y2JrgJNvy1nj7+xWRVSn4O0lyotXnCVQSh
1SoslIuG2pcxTipLExGb3avdxDhEBLWJBGDUlMCUafRVaNN7FAJ3ryS9xOkAYgAkxFulBe3WA2I9
l1l9gzesea4t93FDLR+P582V+gBUCeRAhglCg26pvRC0lgOgG5Vz8gk/t2WObdadPYexC3LAFfsz
kDKJ3FL6BbB9YurLr0VpbcurfD2ofYLaoWcseL0q+HIvuLU+4RnwZgYrFDzz8Ij3FETl4qoDnWwZ
ypuAHg4UnIaqVBOFCKdu4L9fZQud3MQb5gGgqjMIc5HOAybpwWc9NN0TFhLTA2H4RJWdcey/aFSq
TprA8Q6ynhG58oxMdCYBUWN0E9fPTQcQC6WlzfEcsrUrtyg08gsm3IhsykT6V7zgJJYR9MyFlHvp
NogonT8L91Sl40/c2PtlkmSGBOuTuHZTodMvvLGykduvmUja/AVLxcMz+G7c5HZABS4u8RIx1uRs
kNNNH7HIgqPoulMAeKZwiJd7kRpz4jfLx2FsoBqanOcXroq0xBNci9E+XZsD1Y4vtXDfCfsPUiIC
svL8RM54SDca5wXpvsnomtqVt6aEWTgeefX4ZUSyfMnxYFphRysUic2vPHcXMUE2q7O5j2UG0dNl
3h+zUg4xoOKYcK/XZbih8Ki0NhJwcYYBtQLSBDacF8JYdimX1EP7XitZAKWrtLnDvUhxrfXycdgs
5TD2q+q2zmIcuzxJEbwGXvSx1kGeVW2q1Yh4wUfZFwT3REOh1CH0Jtfq+5IMe73LtbOljurnSmak
f+DdK6aih4p1sVpNrd29OB21z4GVK2yYxPSKGza/C9ygmIwj0mbnGMBFIps2+yuiILchRiCbh4au
JWzQ5McH80sQx7ywyVvV2hCxxcmpM4TVzYT6ryogu4mPQXH6YTaFKZ7S1GskeAa5Bj/xeWT13ojf
3PB2kkpbWWiH9Fn5U91o23QSjBqyFJYLWRR7mwXPE/OZeYnEEordiG6gJDGfkKchx7aIUz9jUSTh
op/xiVfwBwuzcOZLesJYGGyPs4gT25iwPNYcN0KCCB+Qw03EjceDvhFSTI/vMUZbhyvMLvtvO8kG
uEgL47IApvvlqsV3ytfXtctOM9KZWC64hvpfhGPSiQQKTzVK6Q7IUhkMXqJBgDKGzq2EBG+hHzXz
YjpKckaWJ/UQhJI+nRu3ThbgSqDwogM1Z+tpPNpnhmtMYnLhnqaUiBguzmqTl+3+OraZGmXbBWh+
SDB0QghH9NhyajG8vBMEZiFVVN417HSIR36PtRSyEyJv7oxWJG9Fgx3+XNHKbbDu2nVdHgFY2wSa
z/657rMpwR0tmLwezu8LH3WgINIMFYchQdXABlMcMbW02IEqD03wDl4C70pYJ6Wqol7E3e8EChBC
mADxcHnHW/y853Ui4Qjh1bLooTJVBflF2MPElQ2XmQJJcAtyDV73EJFBBdbgZwKk4bPQdD2mIIHE
hTZ4UzwJMZMHXs89QTv1+QjAntrOUsaUjcjsYWNrhjvSfGtm0UKH1Ab6tjcAHeKtNyLaEsBGmvVj
qAHV1Fsg6PdG28nRAsg5nuIKgj2eIG3So9vccYCadnmgS666qD8ZRm2jrQVzY6aaVYx1uU4tf3sc
K7mprJgEMBzzjy2+L3Mr6yRe0fyOVb3vVRb7Vb8lSAPf0zicVW92HDJrKcdMYpul804uYVCUN4tI
a20SUlXYZ6lac8LyU7DMsSC+MIuMvDwKxv8SGHFXfR+k9lzdQQYmGc8LJGeEWWcVm0uIOJu8X7Yt
o76deoSrvWUUWkmgwWbJ67TaLIbp2wv41RlRDXhkEpr7cw/U5Zidizg9sWvYx6rPye/NdvfJHdqR
XHO2lCWMrnknfL54U3f9Lsq/RqBr5nGXAAhUr+D2mU72vdp1uB/K/MqiqsLhkOp8CpYib3bdBPiG
u8qznC7oE7janazOZUWFQxw5B23LAWAVpaD3ei/riPd3TrZ9JaXX5IcRxQv+YnqWllwaPtAD350J
CDJiWXZ6dr/M3qOplGmswOhYz1HgkZrKDhqH1E43+EyVyhQMaA6QpPQ8FgMwS/yo1QQ95SZlFGFi
ojnvoe/OFEiV3qWmCUaB4/ttprCTWoKTLkzRUNVw4YbJNvMMSnoTtoRT6W/3sFhwe33q5LW8KRBk
FRSvkVJzyPeGMt5tgtCkzkAsqp4zSGQ4F/BVRZgd6ECfDEJpdS3dk+2v7ci78iCCFRTtys+C4nE6
NWfhWGCUXQ+Coh2U1VG2lYj/847wDAeZD+i8mWFmJUZe8wR07Zw0QjNEaCbSWevSXfKM/MHOS2qg
CtpXjH+qg+YZRwxt/MpI3AB3JaxQ6mu0Risza7RQKfhmIo4hvM93EplF5P1fCfz/F82PwXJx0H8j
s6GpH7wr7y37YMXsIU5o5aX/5cw3+1v4TlWhVhO86POCo0lSIZE55Kntj6zVYV8Ua6TTJI01Wf3u
Ys667o/db3OFYKUTolF6YNz7zsVFDFprGoCAdsnNTNbVvBb25pmdXPuJnXkHyn2rJ2jqX5Vfprke
egY/u2MgqZCQYlhumkpXyX6xe23QkDBGipQU9YLSzc/NPKtFLjLLTZckdq8X2gaX1GO97r1x/KdS
5rUdxMIX6bEdNyNtzL3krjKP46/dCAUejmUhGy569sMa9LPgTJvA+njnhBVJ/55QgrVSWa9kHdD9
JnNJmqaEUSAPGEfjfDrgVi+Aw9w3nmpkP36Jr4LmlTEjAO9eHsii41zfz4VwYnRxjY2454oUwn6r
K9B1HzuSeSSglAEqFYPoDi/kb9H5Qj6gqIDEIHBE8SBTWI5Wqn/8i303JoV36IFF2Hf77Dkh0buW
jLNTTEYtK0cb8Fm/thHjKiiteYN9SxSMH1KZGOB9ttfnIKnk6l2PXRaN1ePVy2Br46wWy74risLL
gVwD+BWxkW4Nd/UUNbUIDdELTkQHVDRu0H4F/f3BwALflK/WXDC+z3FJfrLfO5u6Eh9nBhilyFMv
A7RycJjNevneu8U1QpW19TMLgvf7r5DEg6l8pvI1MzxfTwy4hkRDbasbHYn0yd5j9gQpWmXPYfM8
5oPzay6CCQA35MuL9ROBR15L2pkJdHMPvK1h+w5prhRpWjTdQu+ScLPOLYABuBU+Ph5kePS8XqaS
/gerd0pxevFNjQeegANhOInSUtRdGIlw+b+vDLWhTla78iMmka18Jh3AnLhDmQTqtihMtA5HqwS8
WcUTFtZW9orRdhG3kMRFbrVZ9oGlbDHJGETJ/Lf5pVUT1enjCs/7Xj1SylbgpVnokw7Kr9FRRhUp
MykwLeYz0Vx0Ih5w7eVlDpAdQdySkEZ82G0t0IRc26TDz8x/jM0X91bYsQyEa5hau4RDh2WPDRxL
rlbvxfGTA5u7vyF6hUvnV59lBG2vu8flc8wKw8KOD+aPJJZV7asg28Io/xmBa4mPLz9/0c2SJOn5
IeW/KrG7klFpNUZux/qafmOwAtmQajtUmWvVZl8oxcRBUXa0Da8X9wm9AZji625fOI1l7HZm8nvi
w80SYflILXFsRAnH0SZ9Hmu/yLf0jmcKH5aNT308O4u7nsJScBQAqe16mNLumQ/uxlI4EbYaRgUI
hQg2Ywf8BjtZ+91LSaSYJD/SY8G/eKPJUV0OcK7MV17RAz2suvJp2u3J2VqT7vkmyB6RdczumSNr
6Jb1FYMOiZG9gJxSi0nCf9qREb/t6ukGGaM5X7ZgTfrJTRFOIsmMc6tVpG7nfWTD2jolcTcyclY9
xVHSPMm2l2XOrOHgKtBjYVvNbS8dCQbyKADgdnQW/6uWA1hH4cXppASvGnGQoIJgQ0uqBIcYFk4W
v/wevZdFQwiz23BJ3HdZq8t2niG9AnbrA09iwVfujZIyQ+HYXJpHQhAP4RUxs3X/Tsdy2mVvsd83
YGwFECWZuQgc08xDGlW8nyOF5Q8+Gx51tXPyCQESqS+1QBWAW93xVztfDvpBSf3A5UiocygUsZqo
CD3cN4WvK5ZAyDb5CI1+Q7b7cms88+iRsrWCFhZsa++GtoTYuY5It5Z04MyJ4xM1RkBcXlA58aVI
7puWJFjWzVLA7zioqVlYjCqs9zOT1PHqylE2c7ZjCYeiRlA0pcoDslJW+pwBOxQel9iEG2Nulj9A
OyWtd78iqQfqrLjjCgcukA+BInDW6I81USPOoIoP9qTdAw+y5RNQsbN2/MDVbbsKNR79uZozGd2G
aGaqHAVobF512HmD2rV15C93kJgnTt9MHhcX3F2M2gQ03tHwG8aMXOpxFgH7IowZhIU3QrSYL6QO
j2IgoTJWKcyK53S2NcoS9Oxkaw2LJGj50ZWJe+qxi1hXxPuGr4oW9iB/J9RktxDputEYDnImnzBG
aQI9+kwI+EjxOG0H039oRJwsNh8TCL0Yck0wyBLBKEu0bGB3Qx0UjYrQ4ClIdfW4oUvoXUiF/cTY
sJQ6UivySF+gKbJ78gFktmWF3qZnWKUUUmp4tJZdHhUxReQrhSgEG3cQQAQloEErjvID84Zb/l2B
XjVS9CXIp/UBmF909PaYtsnXcY9byQXZmmkhdd/2AFum8b/XSJi/uzQTO6nDsK7dcUV4adSlhINZ
ARUnEPQaVBv8FUAcIbJu31vEi+3Fstzmplz+7nvMxlt2pgpLhcSXdOz8K2UHF0/S+zHkRYM8Zi6H
Noi5bb/wYqYGSz3VP0aELmBUFt2HD1aKhWRCbPOeACa39+CorT8CL2EYJUiUD6SukswH0sYakhLC
Q1rpauvlD8DiqbjFKzyMXFl/OXRRolmsfSu0puDMndgN+ASd5s8vtw0hCPX/HgcrnPL8eCusok9a
oJJZ9rNgUYftut1xEplxiW8MDgF+93wKEt8hOTkdqvlSfqG7znCNhJ3GSFC+ja4Q703E4i7a2hjE
ceol16KT8AhXlknFYjp82YxSiI3FVD/5VBdQ/yyn9CdlpZqnfayWZMZyfxmi1nuBt677oTpaRyy2
H9LLyFb2ePrukb4YJuNXlSLEbcm1RHDQad8LW6xlN9PkrT+inW6zxbUQ7CQRgJ6lOaBv0mSVU9wr
3+3DOjstwPFk9QhqtNevCoJmbJj+L+ON3qRyZcenix4KRCucwrY01IURR73X9k8nCV6b2O29wAhr
THAoEAOg2iUAbkHw5ArYEz4r1jtKNJoEhiBwcpQg7QZp4m3320GQvEboVw41Pb51wxwxo1wvmcei
FutvhfZfi2wVoo2Nzu+7drOh9L3XI8Wb0Uy5Kuv2R4+YknVMxvL5ewZAQqGjSvPzK8/NuD4TRckF
Cv7Pq06IqEM2xPUgzX53BgcQtpz8lZ1x2Ym5w1GHGjanhEKaUyC9/NrCd/R+LNxb4DY41CuA2916
Fo4JJkeuxv1+KaWgcGj4gdVsIzNGxB3QTU6PCPML1oSFLn76QgxE8dhrSjlNljlzQ/GlTBsdbSkY
dHwpqQfrF83Qgu0C3COGLcXiLhqMlig0fP/WUhG+fBl20lrBE5MENX8FHwx3gjIF2CGVRUvSbok1
FrPVgXT6/T8Gv7dnkFeWNzln894FRbXwDoBZSVIU//Tx4vZ+rwBm1lmpfiOeKJpxC9pHsATgCzju
B/D+0BWhy1dGi45pMTuWHv29BkA4OqBSZJOkX9dI+oeq9HY4KRQydCbDBprbeWrD92ahJNTWaH8X
1kZHcxYA2MIFCfUwvyzeDN33SSteHcmw/QwnE9HGtBr1qSW7rdDcNnbrRiHYUeJU35mdSxTm+I+c
CdSMBy2v7ez+zUseNhfYprDw2ftJZIRHuUE8LjCtyVSo775fS4jWndZdE/SLr6wsX0yYTRpn45Nz
KfEjUVcupVunBZRilMsVGKbgMuUYXlD7qXgGqR2yVVNyk9Pk040qXgLS9qcrZ+mqFTefuBglgoey
xKg7mPvcxNU+LAl40YaypoevOT5ogT0oNQry8qGtcK1ayTd2McMc306yRxhvbpkhhEBDhG/PIoDI
8+X9K46T3jRwiSiDtQVfp6RFOz77S9rvjCsNuYkOuiU9gRJakem2P1O2kVbrfaO48NNXWHG6jVZm
6PNCzWmRRpL+VdTGwydJYpTUK5g8PUkouaArCWThTWT+KgdrPYS9wkyKgmIEqYC9KmZXHFFf3ETl
gmKMNZfD+jJjmDWofAOG9+Woar8tRB2Dvdsrub23Oxuqks4PkbysruB2motf1SmRTajMRNOhYrna
ZQIkMDvL/WB8CsHV0AgYapTFfpVtInel9H78qOGkgB+Ydqtntq32MyXJszOg4vDGfZF6hEw02br8
oO6yEzwicttsuG09oR858z40OcPlw951uyY+hCbVhdTjbeorK0WXhQP5Faa5ZRQWIAga4GA1u4kA
vpPRXGum+IKQonNuSdcedQ2HAlatKr0e4fExnm2CZPgkv5P093yN3oZz83aA7buFJiPG1TAKpXL8
YIFBra1iiDmtFjsQxcQkV+2+87Vd70ffmmxO1P0indz6MTvqRzhrUGa9N5RHl5O1+eMqgf02WFZ3
Ukx/ju5K8vcPD5/9q089EzNuESmY+cjOpSmxugXQtbtzErORGnLRVRecsLKc4r1v3eVm33T9PBAi
ZNbYMz0ZGvRbkGgh4KFL2F8N5uRSsCHUp7I60q7W/cuhVb7X6n/cSJGQnb9VJ5fw1kB5AbngNKMP
MEGxx4U24cettkhOkUVntCtxNy0h0o60h/3MI9nlim8+xCe0cAvUfto7ULIL1nt1ACz7FbcLKV8U
fZp9x2FLTYivqKkI7l8NsJ1dMQNkQn/gncys1lPg4K/Ke9ulGdiP8/VfT6O0xH/2hG2Uq46XUu1F
hfcArRg8Hd8ibJ2eZHIoHbSlVhoJ0pN0VirnFi0EjDrydBTb3IQC1bLgI7IHhPm09sIUaNINfCX9
AOAAkHUONz2QD8lfJAFlTBWu3XYLtkKdJInyF5XST8aGtAfk8YVrctJ/hAcT7MfZP657d+qyy5M+
FS1wfHowEpfV/yB2xmPTe0vtWLo78SXFVp28+G/o87x6CAXjjMmwg5vzFjrJMpAj0UWbCWDzVTtX
N4kJRkyyD3hty7b2TFdCvUGKx9Ow14iDlXOnCItC6XmXXJSp8wnCyhdCKuHpJIOjEuKpq9XrvqEp
LdlSBfJSJvYW2uxeWGCNypHWx2Ox7FqQv10Hj82SwfSYA2COyqdc1QcyGqviKNWo6+VRK/w6+W5F
mfpzjH7r/ywuTX6K2nYG85VvzOme1yuQZTk26OmAluyviBc/0eiMn2B3Im6HcIoWIdqHFQEsmncV
/gKaQqC+R4mSlyN4Zl/RCjxTrMhtFHUjFhHnaWI1D+3NDDEJv7nNaN+zvHOIGBjHpWziat6Fk+F5
e2uEXNPPMYKXEQBI/dCZXVQfRbxKvkTM5rmoW3CS7vetYlzp5UDxZnkbS1u+uZEys41GzcEalgW/
rDwWbt20hhGZnkvxJb+Ij+cbvzjRfVuN3JEYuVAl1IVXY3MyE6A/sjZdPDuTq9Rw8Cg9oGk/LHlf
GF/EjwycOk3LW2/Na30IwA15dOe2ff/lSZIY5sY7OFBH3HwLoWWVjmQSTdnT9aW6kOpHtNYj8Fcp
meMKD61dT4wF/ME1keSAfl7eleuj1Jb4pILbIArCU3zZUQ/ksypFLkdmqE4tsSRIl1KNEsNIfCGd
VYJ81/RYV7jJF6Df/B6V9eT9+L/OAOXQipOrwfXTJiT8G6y4CV2DLAXsPH0huU+Tej6FNMYJvqm7
1S/H0KiWNP1C0RWaAqPlU8bhUXC3l5uxMQ/q1BWa4O3AaCXc7fVui8Uh5xYxj+18HiXsSyR7BCrv
uJ3uZrqz/J8wk03lRI1Z0r/jTlUU9dasZWfhGAnu7/HnB4WZdZn2V+u8CNqJ166Tsmm3utpYXG/g
u7456zm3xH6jfz4M3AosRecurmxhhp/28Ph2F0Acb4+Nu3HCczNHyGTRDMpr0H3B8NwaKB3pyG8M
dG/b7rg3yDGyuJIlMEXfQc9cE+TjSszANLjOCoNDzh98DqT8raqSqpGm/iwESP4UvzH/ueS3uXCb
xKF9LIeLMPK5NjWodT8LtNj1Dll2uTxSz6tIkGjv6ytYsxtEPJI4UdemRJqID7FQdY4DWwEU5txm
a5c5JM46RX/3VsO+kGS+CScw0E68a1r7zzfF3AneptpTHjhFWgdPdWdsRsFErKvq1r8UkjvzvlUg
Ir3om5jkn+9+14DbfV/Yj2xYt97Rb5+zcArmgNK13v19fMza2GBCDbSYmD7aawpYP0u0owLZibez
3YGp9ByIUn1KyJTdFZNaGS4uwXCXaV1ZQrcbqv1c8BlMdhfACjZzyn0Id62wKnLwyuXWtR1ayzqg
ONq1wgtRWc9Akrn2euO8KOAS6xWa63t+hcpsGemHmpYfvkWue9dWTqQLo2SzLQ55fzjZwu4eaR3i
lnedii4Db4x7mYU8kFPgl0cv4YBy1ROVMagjqCSu1vQxwrQYbfnhksNNNBtZnTatLwsShPyrDGeg
De9IVGXPoHRu6LpaAMHqBZweUDGzJj3nZ7pjHkun2pndHWYSb2OIUYazhCL3ZitVf7xVYP23joen
a23MIoubl+DIvT0EHoqotYC6v+9A2DCZ3lSv9MWQAu7KO7P9LEjdlu79ltf8IQ0OJAlwuT1cybGw
KlXkBa4EbhpgWL79Z5pUimGCNm0Tu0VvbqZM3cZKzlpi82il76Z6xg9e9ckG7zh1hUHUEhPwi/X5
3RVoquUCqIVKbKehegO02DXQG0WHKy9gw+fhTKxzZennCUA5wrJ6/yIQjApUq0IwI6BUNCuRvFFq
CbTBdFyszEOJWh8EUHITGdXzmDznj1h8XXhsrSoW+/lz5vyM5uA2Id3/NaSWiBaBmmn4pv1Ii8Rt
errbw1DaoAC0J5NZh49EMFmYQWWtmsEiU2YYKKy9MMLeLCSYoEKTqct+X3wcw9vLAnjKYHiylXYN
0MHDvf3JvEJTIYcD6iyFFz5N2ozYr/1REJ8IsvvLLjgbdHvzDCDscsqdZa2hhPGnEhwVI0imDy0h
jxxLMQzImZq7YkFaX1gdoIj6LnKoh8qH+h4BFPIdsR9bjly5gLgCL6MPz1+q8wVnMvVWloab7pef
avgmFDUH1ZScvbAMSDgc4nSw810a7plxEcytcEphFN5pVBOY7bGZ1GcTqri9xNFvho0wRs3wvTED
rDk49IjUvV7fVp2YYNej7C2S5U3F40uMEWTWYLdMGGHpITaLJNI1SJ6/p0SDY/Ozwxn4IP/T23MB
CiwmwBzDMu9l+6AUfTXYoP09PyXN/fbQ39vQhO1mDR6vh+XZ6v8IVGxEbNv3pluWTmaoz2twCLx+
gX149Pz8NbCJSkXy91laEe/QH00PUuccd0WsmzpX6imLLXCZRPhIV6BJyy6bCUdmnnhkNZxZ0QU+
u/vqaav5dsmVT9m12uBm5NrYwXEc3qVAAQnT1FNxhzGzK8e+QD2QqjNjf6MroA6+U1ADpD/G3Qh3
BmfLvd/9R11i/neY4zzsbIxmrXCo1+qBa6y4FQ5qW0zVBs0APVqMUKy5CBixUym+BOVstwxaJ+Y/
Ju2oH6bBwgimhuNlpwrdQ2j6rYoT9ea6I17n3lMcU8tJ5h3/36iYC0GkUTfrormup+X3FUQoSHaN
YluKmArmwURyjl2IjgyHCu/WpnLfiddMQg99MPtRh+F4jo12XqrPgvV8C145PsGBtruUqynk7ua1
wKrXua+Kt/c3e1QiK7z+sBTaJ9WgWn+RfH7EOWC2wkma3no4Q0CtgiyKoOeY4egN0ZD018Xo/5zN
u1W4aUhC11xQCEgberde05/WoIGUIDa73N7VMEAbkQCLiELhbzuqzT16YKh4q07tqL3OFnS306io
NzJzl8YDiJmLVsZJirC6UXhoFJCtlWRXrSUV0fMfjgh2T71k2ikSmsS21YYw7QryzUxnRTlhP6Ip
n35D9u1iCC16hNZaJyOThO1jY8CVzyOr35n4dgJsXi0lBpTsmiKg801dvtxub6rbPBPwEfuPfwro
uhBJOF8NQu6nC8OuzaCQqh1M2p9ikPBWtKXk3EO4XBJhH6l+Qsms7e53QHqViMQza993F9a686RY
ViX99h9QF3jpNHOBfUCgOE1q/+pfrwrji4INjofwlf1mtfK6J1qjOfMSdjWkR7BACLNb+MNZYc8C
9xHwPaJ7PXR5gDWJoWnXekYrKqNgwjXNvllaoqR7WRd6Qk1d88OlO0xWri9jrrG7uk1Zf+9tekDn
hsaA9NpGxAnUdykLIki4rZd3o0IKt2s14hxLVafUYwpUKNgghAXiiPv+CWfD9HTyRmByJF4IasrG
m88WXaRxkmPxoWrITTkxRVaJkui+cAoOXMYT/0t1y3+9PobMMqKqB5zUe14RzgCNXkbvyytvFlNY
qxTS2ItYAHGLbr5eyG7vZtbP0pGMicyyl503KIZ1cHVYFPgqr7rRz/t0fkzSCSg7A3y7uPfK9b2f
YLQ8KBjzZNMWcRjKuHRKdP0/JAzwzjcbuZ7iqGZrKXUj4kthHS4JKb0EhPRfoqsT55mkI1dZTfcB
d2pgnXiDYdJJDffz9AfCVqqAjiAj8SK02Z8gWd+y7uExsOrqdLQ0nR/UF3tu1IUiIpj/EpM2ZsID
F198lgV9UH8jNN5T1uCWYCrVUAXMCNzSsRjduAbqPlmIui02Ywm2bwMakjj7vItpXhnYEOt4xwM3
y/gqO6zq2Fchc5GGteUWPIESxP/JaoD1jHgFnWkam+2i4JYKlm7auw3qcLyDuEoFrhODr04Na4k1
31oLvzoF0SP+S0/nF6pvd0k8/xDJoQX38iM4Jw3sjATpifH7qGWnQFNjno+/L7PCOR2xtewTjl1W
7qD7JoOVquPW9Zh90eNdhsDvnVY15Nz4OQZ3QKxPjlLJAeOUkIlfEomJIYk5z/9/lcx5sTOtiwuZ
P41ej5pnD4lMvAR13h8vZJrs0Z8SbrC/nyYcxP3sjkaV45/iijcmNCvzWjNVCbrU0oTH1QER5O9s
yOFv77mKEAfWdvCKZdGQqGj/1A4Yt/oJc+k2S2NejVfxWdeK7jKWOA8T+1HKqXLTNxCJ1LfhgyIO
XTYXgHmlqv3UTcQbcCLkG6ilnevDrrs1IQLemtm1KFEA1D6TkGBevU8+GQMG8Rp1oXQflCbJq3Ig
Su7crVj/4Yzo1CrDkTuXezCiH3rq56jJx5b73NdMv7Wiu7zSOTwpfRl50sNOK8E4lGXPjo80EJWW
4f+p+94qXCxOjoXoKNpRGhDKysTk+14998M9BJS91dWylCUWWzATlr5hsrjeaiV4v7TmyHOAuI/T
lZ7dWRU+MNzIUpU43J/ThNPoc/OHATWCqswas/eaEBID07a3NcmBxhYJfMb3UZdUOEPam3CTLisp
vBz79IB7AzOjSbPGoPIkvR3uLPgH/zgYsygih7a222cHWkFhTjQLA0hD7aXnW8vY/TRFRryEQzv7
+CxZ3S2XKaf7yvIEBo+sQaws/WTZphKceezvKX/j1kJbzmasQroEvODh/JeuS3uo4qYrNajdv7Ve
P6a+mOP3MbrgQb6JeSHipm6shPwhDFoGGsj2NIA0T0DJzbMQI+gIc3RBYtlLfV3QtBR8CVx7oe3Z
3Jdrpxa58COVQ9jCUFV0Wrzd/2v85NxgXR10Zudz6ClOnqPODWjgs7eIfKKvxAYBU749nDDkPYIe
mIfdAgie8KYsf26Evfs9UhglROy6+zAjAseKQH0L45bpx76CuAzahnSfkHaRjNSbJltV/XuEfwxA
TFzinjxbmJisjvkw8i1nrQpy1JNVa1Yd1MfzDqseNJN+Gcy5jJoZU/HW8hAW6l59b9QsXYftW4pp
Iae1ATTPOhroXj6Djy1MtOAz/8bpMjee0kgnDne8RvDWM9IKq+Z1eyDTXiwNcIm1sQECb680CRW1
a/c9+5rTX1Hgdcm8HnzDTyC2HkT9RxqQ0ctdfEnrKvPSpJhktn1e0JPDZUuy8mJ0u1R4Ggqfchgb
PjujcCa3B2/2QwaAqbxpwNr8ncJlXAkBU8F1fq7b2I+r94/Q+1dxLHo7MPvU7g3SDl+1uqYrrKUy
/jPAzURlTN0CGv/Q39M0nSAK6jBr05HCK4pBuvpFT+TywcKPWweJnaW+hZd0l5rrvwSQKscaOesW
X7U2BX18dfL98vkwxY3yQ+Kkat8FHnJu1xm0Ex9junoeAPJtotXlw4bbC/zlmKczpTD5Kcxqwm3j
NJ7TixWP9j6egE7ZkqRoBKo818OcGoYW0KVBYr2BNRY03lB+A/TI9UxFTsgcRMVqGIWLbBkcV7qM
T/A9GVFPIOo7M8AkpNVJJHk+qyOh+Lnsy6qgH40MwbLeUlrjSHJIz0+M542QRdZYzuxiuBo2b9gb
gxXBz/I+MqVtG9gimdwr+zNIRPCn4khsVwy2A4zFbRxyuNaZhvcowHEKmI7raqbzswa3VxkAZV6B
De2D7M7bf3Y29V/HBGZtxOONQ++jlY/e7mCW2GG0RmtPstMShmXcZgznEURvFgrnUVeB4KY1eRBB
ZMBfkF/dFR6IlT8a21VWhviWma6FpR4dIUL/hf2i5/l6LHWGeEmaOVtw46OnllWu0CJ0vgRWfOQt
0DCiO/S4ehU91Yi9/TFJva0OSVu0eb7Ib8+MqLTbOl+6eZ/ja/NEUb2YyUHYCgGuOpiQi8ZtagVs
mX7tC8PP6DxKOQkX6MvSa9G91V3gLHA3X4Vk4+9coGPCVncCwPnXPpcZ1QfqPDb+foMufCym3DTq
pMbAkqOKw3ODdI/yEvldrvSNMm8i+2H867yJs9AjNj+PhurcmM/SH813Whk35/Gutt3degB7YYRR
+Ol4pNZIBFxPQBcIRxH5QcdFSGlor6Uj6+a9yXPPrtVBym4ymnqghq+t1ba4+A9V/WFiuTP0pZnn
CUKUi1g1bPgnNJ1wRzju+t7QX8p05rZZZ9TWDc0a/uVjBEjMXrkxZo/SFAQ2buBS+QtX6c/yyDGv
hosPRLBNNBLYzMuFAoqf0b15hUqTxG9wJE1RxMf+5nkMBqsta0cEX20VlIeysJSQo2QATbfIbXWz
lIoSD+6gZ+JMi/UDLv3gv3Dpvqv2N/rSGpbqOyp/38kcCaoiDr67tYKfMa5wagm/rw55Ezd7u+73
r/M1G85a3em2IoKwzibZfbfTIEAVM+T46NL6FYdns2dCchjDx2hn0B9l8HvwT2aEQEbRaaDy/pOq
6Hl+9EGKTrSaEzNWz7TOGv2z9Pv1w0tqQ5qHAnJkexeU55CMfVQcqDXlkxzyzIYe8KI0Xo93ay4h
lcHFDn79aoLB/kmdSPuZj1HvlluUXm+xVnDO3MUoZGeTUjpUtCFaQdLULteANpyL3+yGMCk6p3D1
UwLjF9XHnH/ZSurQMQOey8VohU4QpIigIDy3N+rTdIDv0Ay3Jix79pHCK+EIz47FsfZwgqsjanyc
WVRdRYD+BPduaiBkNuWA2aIOLqBuGgQglCvJ4LMCz9IW80RKJ9p14gKrzHm8zqjDxrZAd7tZ68Nn
A/7idrSyBMBWfdzySvbRuHA3RUwt3o3fGeaxQUukh8P3J7ScVi376e+1zqQGuS+jJkk4lTJ/EP3y
jBfpCjFK03E5I4MUF5NgNyPI3Pzx0Sj1p+bYpRXNVLXKJkEDhEM2SGgPUUKdyV/Rp0tNL8EHDuTw
lfHFwCphtWXze5GepWOgf7L+AlW724E+3NkUlB5jm+n3sKGihK3nXHbB+ullI/tS3POZNdrrKKJy
s5L8pM9LUez76FMgHOVK1HjXFC6Gl6aGk3gLYeXJY42Zt+MYZM7leZ7JblH+5DjCJLZw1lyMCr7g
PlYOINARPkRYHLO1RWZLHlcku7oqMmDu5xQbC78nDJwhWLptIfV85vcc0o0krqVA8/jEb1UDUXvw
LrGO169loTOLdXeqlcHKLuBRkN7k75+oiNyhAmWV2xjvmhhBX9YFf+suNmaCt2U53d0Fu3qu4tlI
3l+w2JzKSql63wfoCguy6A3xVVYLVpaD3t++MyIXn++Ep7i01AK0zmPGknwm9U3BTlTyBt4aoIzU
GBoG3j5E5uemAcjniI5ScnSSfjAPzabNroGHaiwxcb8/Il/CBQByIBQ9eTluNYCpW6g92rtBO0FJ
NRTHeNsgP4aZPbjg80OMgLSL+qUSZgnxYX86uSwopsfucqsfFQQBASVacCTo7lptR8s1j4SkIIVu
FdvTo1B3PlAVcySp1v3jiBpy9mjX1zkJJ5kFaArdLiAhChBQqgSJINpJz7vizJsLVDTY90wvfCwP
qNDkllgqew0u4ZuLaD1qjymnNpYixAhbJXqDA+YUURbwa6S++Vw0xA6gpMR36qwfK5H2vmJRmLMd
hX1/1i6hpmJ99GEkTk7yBDD0OG0XML9Z3mWXNLJNNJgtAq082oGsIUKAq/uOjRBB0hjmI8EWC9hX
BMwtGUZPur6JU6lkCmlRVHfbnEWlWPMbsVoszOLG9QKtfv9lr+REit7K9O0FufjgLRWgiVmD9Vb2
rYkh9NGM9KUlM6uIbBYkkc9FGrRsOPfimRIX7CXclDRpQn5cZ8FuMx0YqgoZ98vL/4HacCPWacLi
UcZy+jrr4AirPYxCQZhD0eic8dyj24nrr9PeoLf1S0az5Tzu9+GAjPoUgfDWoUYf8ppeaLfVYq+a
ojeeDhOmShKesIjF1ceVkOkR21WB408uRvdiPlaMr0oJOi3tZvvIpvqHR3HkKW3Wh4HrbuGPAx/2
DxJ8cCbKKdjhRrA3cdeNiwrj+d+w5yq7gM//b9woAD/+Yv9ImMrqLsnwBUXAnD8PlW3ria5yMdN3
CLSL+owxo1tZSBndHU6EYTFdyjubEtqYgsPhE2kBqQ7VuojznASiTm9t2lsvEG8u2fdqbAaaj540
fPws9nnoPlkQ53qq+CFx/HSSqudKRdATCES4/tR390yVNDjkzl7nRdWzPxapmDo5/OOHnPNFJY3J
Ue4tvu6Ht9kTYoUUopCH3XKwYMrKZdQS2b6d9kEQlf4NL6nTMm4JAzX2tEf6qDVZ+ezHuQK79NkH
U2q9HdRRzyXj6TtPvGVcz8wxds+tcnicA0cCTZbIPNloulk0MzF+A2OwIrOpXE/aCjYKOKhoQY6B
lLwkCeUsbHpllFuGEIqrI00LGGrzYFGtreBfOcSaV9DjEkh18vRQhzvQWVYqrBGaMcpa4k214Wlr
rWUTavWjOsJ6QqIo1/icuVumDMIyM6lnQYxReh0GJLqCHMK5cd9VYOVm44hLdsoQATjs87sPDWgr
0qNTzCUZ8mlVhfH4uvxbZRHVDKO4Rpkm2ELJhkn7hjWhNripB8r5HLEmUiRAIOxTGz/H0oXFPWI2
9FC2ELj3JnQ1Rcagt+49PSv5LPNf43ywuDX7Ffg/W2d6xIAfXdd4JRyaQ1yjRa1BCha/b+ZGTlMb
Qv4U/g89cdDMEpJyTphNEtRPRY58ZXtRJOBev4FhmaUmuuIbBEB6eq8bYXxCaTcY0fEv+X1B4pCV
2D8Rer7f75ZefFM98vnnoTS/5MAIO7GfJLlp4lzkT/Ff8Guc0p6f9kKFeiSxxb2aSHL9FqJjB4BL
ZTUhN1UMGKXe1Dy6cyeir4y6AG5axgtCbGtafURWZjY6Bk6JKFhSAtmXe7wpnAOG07tdjJ1KBRpQ
HQRwYoJehZU0UdTM11qhUBNS70z0BoAS2HgHw54S4XParh9rwhDO1t1fvXh3SPMXF9R83Y7YB9Bn
i0qN3Xm21Yt9NxVyxiHiCVqX1naQMXoP+ykz3Gfk6zRAAeaBcs4NS5QDC/FspeRm544wSevtFJZu
wIqzK9IOMen4RmU1kMmNUEMp1+HalNVGrZ5EBsthKI+A3tDSl3vWUeIHVgJqKmQtW28NeBtx8wFG
4DTorQ/BY/yJRzuh8JznHfMEcgAptN27vK4FcwxHMUOqB8lqenalJOIiZZoIEGsL2/arSJgdn4Y6
Y60xr0KC+1DFQ8RmOBvh3WhpAO663mKbNeTV7gdX8AkOWSKYsQcV1XfT/IrzDicIpbc30TivpzoQ
UfdHEA2evqQZm6s7hFTrh4zZxWnyXK29Tc+0Lur2YTpiLlj/1rej/45ILlTTXuwELz2RVuFwcirK
kSNVDzTchI3qQDakgCCMzxKY/oA5FVrfaLQhcmijb28zPEC0PZOBxV69UW/KMu/hj3fBj8BTTtkD
fP1UDjveLRYdjU1qkTHt3AyD69nSPdilhoJrN8CAARSQcp4iD4eQ4IqYFCiUK4QYpyfO/mhk5HEd
cMMIWLEgASz3cB8YvhWOr1ir4+UWN6Rg/fIdRKP+8m86b9btjWWEKN2+30KYTzjW6E7mm+N3cdS7
ZCdR2pi28XJprhqWjSnIZ3msdUO71zpFsdBHgrQwC9yjVbtQfg7mh/phULfdkxncjJryN7wgFmbA
o+/C6Sv6YF72pXc0H6tu8x8Z6UlWNLItlLnPJaleDd26yx/UP8eg+d/H5TLtTW9Umwm8Ge1Dkxns
fDjD533+rceeZTkrRp6QsjT0yzFoz0xlVkaALPu2k6U+/SjG2VhxqKqD/DG0mDUasvcJ/YxlSRes
lhVr9IXRizE4nwBuUcGkLSEZtsOloRit+QS7sCvslWNDXmYpj0BRrwk4c/VRzGxLsXQ66K6pa8t3
rg7m5pyBwAzpzNudc9+xqdNHmw7IQhoaq65Fpe0cfD9Koru9qb7L5u0Z2PlRnD+pMKu2lK7IcZB/
+UU8lr0Oq3QGywiOUhBv3iBAPR9R4qOnjganzR3HPeAvz7lEF4g5a6hK65+DlV6HsxbynxiraM7X
SGkKvN7GPom61+iPjKwHyl8tHJbtgtqfa5AOBFQ96eo59SXKpJYTE57+T+lb07Ty+py/byW7ytEk
s9X6lrygLUVwWrTmYM9XVT8IQQVfHfK0WRFFlTQDvQq3ydk/3ul/abGf0vkg/RtyRDXxWOOYOOPd
RZJipwPSDs10pfR7ztnY6BjbD1O8tRqz3q+mQbbyYLvwoJ9Sxx/zd8niXvPP4LMMbzRLM19DI6XS
Js99E+8z9ODzTOcC/O0KTGA9IRW3LqSMj0xKk4hKxNDyH3iI4N5d0/5BZbZ+NO5M9vdzWyCnu0Gq
1IeDqXk2g4AhleFO1UzyJ4IbXUbZDfg8/KCbFmyGtldFJRWqRBh+hQJfisucgR3pdn5cyibFZBpY
HDF3pOf/HEw9+oZ6Nf/ilB8QWXxHzOoiXWMHhH1Q2PiZVKqG0CmpOdy/MtZtr2RiB2opZpHtmpNB
R5GUCS74qDyvLOP9rq1CPWeGI37vsqpTan2b4xo29hWo9xiVeDGxJl8pMntqMmbbGrmcCAsrOYl7
R6cW3vFBPLcF5n3wFfU1s6r9fHqkekP4enyFu8NYbt/IBcqYlKVeG13huXdz6gpJy2hzMjdRysZD
UB7QsF0HRait8/VFL+iKWMX4ZIqQtgb4GK2ebmsoOifjepVLALUJLRvwm+aTJideCQQ3DPGwNabZ
1O5gCeD7uKC41DLi0woIcRnGQ2prwwDuFcrmnqJZOvLY9U8dQHRJqS+UiaBhLcP0joJf3S6QP7Xi
VLliIoD2Qn9H4lLi8MiUMTBzhhOhkVuzuJItQVV/Cv2u6UAH20NqOcJavDSfAwwcyUj4YX7kVp4D
I6+/fHcc5CKs4TNppbz1VxN2afn62M5uWTcwvJpZeRJTvpft4aK57BYLGdbuzr9bEww3KTMOJ1/s
OzPsyXMWKgxDPJaDG/twcb9xnUbUs4V5clHW3bHnkA75agjOyQ7kWnJLFpAkf1a3UFJ9rdGkc2++
bAY+/qWxXHtJojfxLQ6CM0xXCOj+3MWeYMIsni6IZjiFc8v3kL5ZwaunwOBCHUuKnRSCF373iTGb
jZ3oK3fQu36QWq3U/nT1DASiEZzIQGbGfSBNWernm+rT2nSoTnjaEjxAvv2ZdPXVWBdHjUYykUGa
+b3D8bkk8cf6QaSwdrObT0RGsK5drPiASvHc0cwmtYoxYQUWg1KO/0QXVk03VPbz5Bh6i+BK1kot
k+oqJyZXbDRQiMpXQswmlTOx0Ct6zMgUpecelXmCvT5Kiir1ta2sc5maaTLNM0XSGcFT00/c+3c0
uI34QsAmuJ+sFm7xic0cXc89V15Osx8fKCLh3Jlxx1pfESg45G4BeOPLyfZBKeEuqoXodYZ6R6Xf
3YlFOSBTmMbmFSmQPvsHFVw2TtDfw7Z9baWOG5Q7gZ1M9VmObqkNoDA5RlUlJ2721XrrmSqOs10B
VuAySJ7G57DvR75mfN9wFEvBApkvXFehhtzUdSsWRocxZ8k/i+QqGyWROj1Bpmctp6d62fps6bLL
npYg0+G5RNHBkoB4gIpGFTdDlWgigrL1OIbcFbQGDS7rjMiLNJzXgnt4Dnxoml8YPXkN9UMmRjP/
+NiBmn0chaDT9yNfet0ZYlK9kp+XSTKmtg4sFENv36REtDzj//LedV+NJX8V6d107kn1H1Ji1dLq
96ucTwAOvMVleqvERjDhJ523TnntoCRt4uUV/5jcF4g/lKgeF0QWZlXMuBR2a0Em4Yn4QAIEX+6a
E2IxbyFpFro8pCDYAKspDpCthu6ydZAao6sMHoVI7rCGtZBFk9+2zEiNIN5YKlozsab5mIy3mZ/K
o9B90iLYpCcFtfUx5q2zQ/qjtY5QsOrN53lqLfX8fDxmzOFRtibDSdRNvs+ap+BDEUY9hHtXK0nC
B0FMy3LKASGVFU1jr91YcXCvrIdschJmjHECP9TvYJ1xjCh7psb+bjRG41meHQTftv33HSwqHrj8
CYwZKO/VHBF69iBv00pwMwpF/jufd7EiW6buojEYc+akHxmAog2zLaFf3f/MrUud+avP1AAH8IBQ
lUg9nir3NHi/wKiAzsN+h8kFTZCPljYKDtgMHLGtOpmPZKk6nq2SrL/TZI0fb9F4L6yDE6ulnrBg
xAB27s1Lek40tSWiHgqC9eZnnXodCyw/UY4kxVmiibDblthabGTa8vqWqxV9PzhLJYKV4+uVife/
TifZuq8BxrnZ0cJ3hMGX7B+VBp47ktgBwPGW4zJ9QuGS5kf9Q+JY9yr3XEqzG6KsZOqu+zYaykux
a2Dt2NnJr39Ui0V5rv1Iw4QbBXgGl8N9owFFo6IT11GNpp5Rqx284KCvt5GhBtBC6JE1RvG6Z6dx
1U0GJIOe0lmyIHmV+e07JpJNPLNFnEL7sCNKJHIdLvpRjbheZPdSimpWcVZ4NC0ull7tQdTcfsDE
yWmMZlGujMIDKny3Er3dF0X19Wl8ayGNEPqOOOZKIySSOurnRZEZeO16pWiwWjeaOYtTgTkTxMQY
fZpZ0BLZMwS4E0E4S8w+RiTsWvwD1dArCKfMkLdSi47Q2VjtmSG3KE7T1xAsPu4X+2ajLupSKYUJ
VAkf4OU67FgwzEXFZygsSrTteBVes3ge8B1k2giQWzRP/AyElRijIi1IsnE+DUb+kSekb46j95kO
SoAVKTS0YGdHswShJPRxFjNEGwEY0i2wGY/Mf8lfYdMonfVxQfFzKeRJJPUywcPU2NWk1U22WzEG
tHFq+S/GAq6/N8nhzCuGQThQdF5gkNz76KGO12c56du/pkc/c69yxof3CaUrviPulZoWzzerk0i3
BxZKkAHjTGEs/lwdaRRpa4/qnX787pEKbJmi7lV09mtZ5lkUWNc0a1qA2J0PSSvd0Mj28cntWOyH
28uGs8jdcVjJnqLhmuprfyw+naxCW0fPgYeZBgHMcN8Ep71A4E7xOY8NzahbUV3HjVQqpO95s8U0
ebK6P9dmpCSbIZITvAY3wkdxJFFXi56Osr5TVgbLeF1zOarYeJ2krSplrVLByelb1EpsWZgpJF4/
N0YeCG5AxvNntgSuyKbQRc9SenH5N+2kT/jX2HCTISXGPNrd3/UymY0svW0kezcyYTtsucEpIfuo
B6udypX28Av+wTy/j3DdPZKOZ60JfR+ZvFgsfZR7PaeuF6+H6ieEZaNPaB9R7e+Oy4hQKsCaVApn
ZwYKfH8ow4eWWqrCHCaapI0PPTD1UNxokYU3uSGBOK20bvO/KAucW49hHwzmnp4VnhXqzTEwXEVt
GMeI0RZzkhp3n4D6umPJMtFs1QU4vPj9xO9NucmYErDnqoaBZjPVWjTMaJA5cc9jr7uO5VImh300
dooOp+ccR1Si/ACunTNgu1sETMAy3uQP7puvHgpbcioW6v0iCUhvWc62vC7ax6/kfDgznBlEQtXi
4XurIONiz095oq5JObac+Rv5etT3ADVgRX/JtyLPwOoTQQ5tderhQXJkvkV09P5xN6VG3LlUxpm3
G2qG6VSynjYVg33mBcPrh8J+BEN0V7vhvTeZndRuheKK9mGVbQK2zgevwLZxk4V7tR/wY+FbQhoi
8L6TZpilNalkewRuwsMj8++LvtDCtPGux3dQCbMfrznQKZ1/VTWLuPNxnJjwKRsvRp0+FZioJ9Sa
+L4wSt6ckUjAERzYheUQ1aBWCr2JOG3cSN5gpgvPWmQ2xDNGLfDJz2i7N9wQawD7jCDQFrFcijR8
CBEt2nKG6FxH8ehDfg50itXoT/f2/5L6ubHRbiJeBOczX2LTiyz05UOVmk/UksQnaApW4fpZPo4H
RZKOySQpZBc8HW6vhATLAFgVIes66zuhZYVv6ec00uKrlI//ay7y3eduYcdsXgodOsx8IvxmsSSL
IW5ClL/6+2Xcfwkx9DdX/yRjKKkSU+0oN6ft/pgn3ZZrODLq5dBum2mGcyhMj4FhzgBRmUpGYNlK
/bsnyznXJKJZQyRqE8no777Zmd87MZSfsQ6r12lx2XTgkdRjbrg7uhux3PdEm/lN2LRG5PioG1pX
/XC5gYzlCWU9VRVMgIUeFM02MkwTCOcUlq2fnlrZwh+VRZAHjz4yCnow/r+Qoii0e9fFIVJxnWTi
q4DjL2ElZjTBo1RjkbKPHhZd5mB7PARPt2QeOepOJ1Yef0nPrcdlgFW102uWsgRCA9TRRbe3BygH
D8W5rluV6R4NI66Kcw4hEXH/GAAYFSk6CoCIz37YyeouwQKD9n3cGSct1D4wWpoP1xgC/X/4BkgU
6MBaN3byB6Oq9Rp/JG51Xzzrqk0kvJyUY9bAaYJBykebr45mSDNCGhDRsjY0XARO/jjDNaPHevyV
UB+EzAVRbxNOrKtGXZlDu/dpT9XX6scRArguzyDOmsGjrQ9J/X7KSGeNhqf6R4MeWK9e9BBrXXLF
KOtw7wRDVUQuSjIQGyITB7yzeMcbDz1fdiJRWAIA1gVZg+++1Z7vuCNpW1t0s0q13IC94EHosZiI
k4lBtoPdC4HXw2TsqbTQKrv7JEoV0R76VD6CqKlqBAsZEo9QTCoYXFbY2TBUnXPc527dQ+IyI0Qn
O37FNMXwkX3wH1NTIy6ayLMOHYQXlFaL4NFMteCBnMegf/VdaNi4zumaNPNWTQ3KiVAoVMHTOD97
LIOi4J43er313Ry5TUGt8uSk4g0BQjR9qI8UVDRIJLQ7imaazqPEFkZ6/mHWjtv7B4oh+fBXgnbs
R0RPlMGRjx36uKZ5/jpCgEKS0rnLtUmo7PdF9ZsbCZUf3Iu80kydQ93Z1PMYzEdeK4U0OTwwEZ2q
V3XsXWaq7p97Z0EX8SkwIQD/X3xPgH7KWgj3GpScQ0OUtx0hBDfKPtTACnBSbJsfEW5WibEzUBew
Lrn4Vpx1gXK9k9aM+rxPhNUUiAoZCJXv58TBUA7tyrUZTZvTbMOQMjvJDbDGw9uP4X/MKI3qTuqI
q8bZLWovlJ8LQ8M7gkAOyPrlggRq4kAkAWbtZJe+2zi7+plVSFdg7CBtkc1gJ/0esTBx2SaA1z8h
+3NrrUKAhI8458jIV3e3SGQ9Nb3fdbItH2lTRJFbFRZpTU0nX85rzLrPzxWJgphHjUY7K2+Cs3yd
fApoOg/cZmO/uctJO1XiFvtBKenmKXkf1Tb1+wQuolKs65hjR3v2TaaTWL6KLQvZ8JR76xYmyv4l
obv6VRvVUuCvGLVkCX7Gzo22VccDvcJNPAlxk8Xy/c4pnKBpxj1HcdoZ4p5sIWh2fyMOgsE6EQ3W
6wYjd+CKnAVpGHzj+nGhQ8QdWoIlC/2mtbTgdRhir7PAYOj6WIo0fIl3ZRDi8AnicgNHysIhnAZZ
DBHo44htzKtXsoUlq7FXPFUr2VjtzlnPghjlsOUpk+Majopu+cuA7ODDU77OnMlHyjHmr8kSQrfk
EntGU5qULJGdafw1pZeOunIPPZy8liQwXSCCAWEEViWPQ2E0D1VpKkzzMYRULlq1VOF/44uwDmMJ
tIZTPk258I740xo4Kn01UHpdTPmIW/6/V0Wyt1EwBTAO59/93tsAJdXHs4d+YtTZHWBMVovFnA8p
q3fc/J2fxPIobMPVKCeAVFVEpSA+BD51ZTUxA2/44WEW2cv3nD0a0jIK4u4v+Eqd1Gnf3Lz2Hwv6
j3tNu4JD1m2eIfQbxKooI05AilGR/5mELleoN42rSnAVPBSQOAP32/1SBP8alfOhAutH+zoRsBtW
U8Kxaz+mSmAtFm86aYxxf5A2X1iRkDwv2306K0/LGCOjwIKGA0TzL+7Ri1OALwqxnedobHsHnNuF
RtUJmWrzxfmxCUpkkB5hi5jHqLf6L+Beuyjf2cR/NTCsAs4WflkUto210FncC5wtbPMkNSkJHmZr
GKy9Wbqbd1YLypMwouzixbLBxMhqr+8Ms5stmvGQsg8PwaY6KQdwQN/UyNw/KjLf/s+15T7KmjhY
wmCodPCuWnRsx2EkMqRlV2IdhQBdULVhbl3AJ3ylP6s9+ym9GhCcfxCdtpfU1F8ihmZBTo3apNha
T1MUNXoQdNSApwj2/usH7Zgaxo4MM8Jm+ZiNo+lN0TUBshvdiB3r5VpfxQuOLNeFaJzJgceU9gr/
OeCjL2zi0/2+x11taLknvTFCd7WuhUtINVZmenPeY5Xc5ca6wt+XEJDLnXY9Ov1vNEASxP/BSxgP
Z1NZVwtQJQaeR1k0vcbbYDKt6RXuv8gi3lO8x062wHlJ8J6txIQ/P1DkNZ9sAQ3t/VC2p67PyZVl
qE1owiAdhb084EHAI0mDRlcLrUhQuTzLiuwGbX4uvb/85jn1ouC5GREf+1HE6jWkgEVpd0lrRjmD
f/yUb2fhA6Tq2SW50cXmfswLj+oYuH2vo8poBXr00/alNhGPvznswba9g3nq5PTRFh5y9i/YAkPi
eVbOkGgDEsIWD93+8YXbSNINvzEdEodc1d8hweCOAwmKBHfM3tVDP3NXyhak2aRadvYQsZDDC++p
CmWy/FFLxHW4n0lsR2E3fYmdRgxfgAGXFFWCJDWtEapVrTe+nwtJvLC7chA60ObMFLhXJeZES5yk
F0ijQcRkScri3T4HENnchueFqkq0FhUyHS6DWQeoNpQwu316pOcNHh+nx9Cuqemo+fNwByfh95yg
m0l+TzUbTo7EUNm/XF7xTEmCv51K5+C0E6YUbLL0QYm+U+jvhPKu9a2kDFR39gekwE3eWbx8ph+a
0AEGH6oGGnhqm2Wth1jlRz9ZjuD3WzDxVUtUM+2UfjI2QAj/xM6CDDZjlNA5EAmHmbJ4vk/z851C
uRNyy0okvghHfgxiw0cRplpYV4u7Y/bAQt+2hxnT36m1miP3KmiKWWrOV5/waCdAhJ5TqyTM0wkH
8zDevSS/SleYXN+4Bqzr/MY19ZJon1OA/YfF8UqcCm6j5LyHwJew36Iio1teRCRazxPkwPQJOXhT
xhiL+WvK4DM7j/66Js2ncWWEWf5Kp5RYbo5/LhXLM7qyg1G7IffHHOBOa49GlUyR+Om/Hphq3sRl
Djr0o4NMujNk3BSLU1BCxV8dsd1dZ5K1r2q7hgIq3Tvpg+MR+JUK1r8b36MwsKZodE1kNRVYyWOW
/SKdHzpKoH/kTZh0SeUc0ukqnBstcBAWqg6HJQxdEy1ECAcDgn/BLjduHgDinlUy/DHqNsLCY8RB
ymhFbqJk35bEmqAfas3nxWHqDu2M83BRN+lgCqK0f7Hmg117yeVwVD1M2Qy3oYxEmiksP+9DTOAs
W4aVSiQKbLyy6tc+xLNeip6MsmWLHu4F1TPuDfyaDtzvvoUIqC8Dd5BDzYgHYswk0ul3bTfsYCu0
xY5RcyQSJbJc/ovekm85uOH0kGHnyPJDrCuPb7HJm3FBHWH6vHXeG25fEJeWG14c8qNOIINcytF1
JRQMeMl0tnAQBNXvwujSi9sYQNFxoh0xqwnY/4m0+AY4cl9Fqe9UyjTQm1zXgB/+dqkYFiJZ0U9p
JVtfY51d5L3oMC2N0z39Bn1i9fQ3vwwrDw54nZpVSAqAAtgljwkGakulKHW26uX5WfBRIToKmtmr
9H3UWlYHV7l5dXC+a3vojDm/rw6YvKCLc4Ln1h4G8lMV4efns+iYZuHEczecsxPDMCF0oHnmLocx
1ymPC9fwwxDA3QJF4W6s5Yx3nwnE7VUvg/NZIJ330UM1J4tC2l6JzwOWwVWHYu3PRA3ZcbIzenHO
I5F3jW98mU6C8SSm921JfhEHZyzM6YYuzOU4pNQWCYinUUkJjT17V4RrYnFfZLA6/3mfc9oF6sNf
OaW4sSnCvUTfcwgQDGGAaN0D49JiMaiWuzFt7F8HlE2LJz2SZjRfvyYiEwGq3o0L87N2XTqJ5wtn
s/zj1CgWeWA0KoKQb+3SLRZkhUys/OR7qSsFsnJzDm2muby9dgJuuhajOFBfFJGu4VDMOkMo23Jx
fOZ6u2WSDLJou1yARYQYCwtTyfPts4mfTNw2pH13CX74izgNh4JsBR5LLkhqO/pY6H1yMlojzUS1
ng/wTFNdtmTEe52degl5OOAq7U4uaF1FrMx8gDSUbXIPGCCzbKmwa8LWifLDbxdF2N4yZilefl5Y
DHL1u4yX8/WMSO1R//W1svAXtHfcTstElo1keRBNlZgdJ2Bo8lnd6CTY5A8m+U3x7ZTIR3p1glwA
uNKQahu8xUzhP1WqrnAUIS+gF9gutBepy+/dx+707Z2EqWpaChZeGxRWsToIG3sVrQ3Yn+rcgUlr
Zn3JV7LV3q2LSyiaEOzkfgL4kM3ybcj8/kUXIXCEypQ6s60EV0XqFAoFid/KhW3vJ+s5Ija9lv9Y
Ke9nwkK27ozSnYndI/H+Sre5H3SbsFp9AKKp4z1utFv6Sv3x5zkLTxlp97JZgLJ6HGw2tjqh4XOe
qawgrkABSYFx91/qsChmrQyUd2Q1gySqaMebc5b2cVi999qr/pd/pXiak6bX4p8Xu/7FnGijOoe1
kU8Lpm28tux/rDh6vc6VkeU9VESF5v/ZJhqY1eTHu6g2CaOpcXY76I7YVHDYVEdpnH9qcelPVaSN
padj7sgfAwMVcG95zb1xsx9KuxqUqCJZ1sJeyndInu36upwE0qjxOh4fiTwvguLbJWmC0iRAIdkn
KIvT+fWQw+rGiG5w4aiUA43t/cy3r0biLylMxErwE1wPYmgm5lPYxRaHhkFfsckh7HTUW4QvbZNu
OlWy2VfB9j7lNWrtO+qUCiPYQDfj39VW+r9GePrtIkmWXDy8Utikj8VA/dcGzaunoLKmUgTe0Jpk
wfImj0XEFcMt0+oESwd1zt+LiYynt8TUpLYFVc1Dwo1xUBQ/HbAWfIlGtPNVDzpIVHLIuLpLV8Rg
aW2l0LsipRCW5Q7MP6gHCNx6u8t7pwh+ChbY4usKeBMZZghjJenLtA0k9chk9oHOo7WzNVkB40Hm
+RymyA6gZzeYmndB+YE5ifVScaCwOPrI1qPULp4bLzAR1XSAP9rzE3vTUD3DOLqx3XkiGqxLxcmQ
7/7DjHH6FzmnBDM4rs5+84YqMuxwsOK3W0q5+SCS+lQ78H3f85EiIky1floM4wxI976Op1ZxxaqY
lqZRkIHH3aaB5/fvbboI7amUigAAsnQO3WxlmBeDKHkBeOLR0NUXov1gFo+IfrmiI9pCUSvJAHje
ZR3FbPIrsqr09YJT+A+7XRGHzF0XjojBUhV/Yi6kM5gqweIB8f0WDx/LFOmZ16qUvaG120/78Flj
fCeOiVtZdBxg0epul+ADgUhiXpDCHuKmglf9oi3QEsPHd7HtaNP8QDXxft168TxgFXAe5tz3nvap
h3WBrLRytoVt4weZXHOOvcg66y3wNV3ywyvN/m13T/jjQS1j5zHMy+TUnloW6y0hJ4xg+eyZ3Eyb
GDqNGh4W12scS7oQUCKuKym8aU753neET+7GdhL4nNLJMZ+FW1Bu4eT8DUmR91iri/IvFiJmFFAB
yUQJvS+yPg4fssqTE8o3mX4t6sfIOJtmBYpWnqA2oEbctPwfgGvFeXukzp7kFLgParCndujg570P
B7ktojGfOwgAi5vD5xGmogv6vQApJgfDB5qbl8Fj5MiEhFV3oJYxw2HrsWkyRVXvvVWeAx8yUV+C
grHEXh+ft2TK4HMUsihGuKXhi6rOahtb2hWA2qlnXiu2niQOFJUZOQWisjq0XkBjYITuh+8mf+4X
qKlYzOtYi6omeQPC+K5DAh/e6Ghvu93Zu6DrFWJ19xYn0qH8XT4kScOu+teB0PoBjyVVXCjWUQiV
5iWajn4VPW9U0eO0a4GPoD6/8SxzVJAiBWFwBbfG5r9brOhxOmMJcT3Ly2HKFr94f3mrLVf5Ptob
EF/Yt/B6n7wK5UqSXXu6JGJO8u5AgF9WYuzALC1+J2l8SXzWT5I1YYlTuKYc3OCu8lRus4z/g6dI
qHNy/ahfGDSe39N9kDBvD3lT2uef/OtzqyEzp1VOHiZWI7ePQ9s4gybj+EkX8yrvcSMLfDnRmyqR
1DSFjZRV/nx95ks9QhTxEJMFNMBb5daqgHp5JA1Vm+XulBBqmBiQ8wnMXOy9AIyZy7TBdtz0AF22
M8TJ0UtixeHz209CIP7fKQAQFfuXy9epB8ClmQPFbWR1gIH5A4WtdUnjYRNKOPNhOaSCQGNHALl3
DUjijeSUGx9UHpx608Igk5594oX662GJwNqvlhj7+Am/nnVrrbisD3eYZPkrX6HaVKFeEUmB1eZP
l0NoFBKfW4G1VBswAy9AgAZbLOFpofz5cTGtZPtnIgdLqwrXSOvNV+y/9Z6PU2ZCBRqxvKh+tGwp
FWBna0tEw0QPLbN53HFo4ofvfx5mhLnAVHoCTsyVlkHZKzLYfbBwVnUD80AMGcnvTSQmLHx8vnha
EbBr5cpnX4rCIYqts5Mow9mQZUaUDrX5LiNh9S3E7i1rBV5IOxIL32dSzow0odO1HJotTSQxw6LT
ahtrSrRHn5LOhE/eUbjkF3kOQ86dRFt2SRummttfHNGKL0F6mc3RfNrPO29pahGb/GUVSTAZijqx
wmdwTAThvxsxB4HmaWzouqFCDV/rue5Mwc2aGVRU9G7GJVDMPC9W31z086TxyI0s2djFM8O93T99
9fIkw08txUU6IrS8gKZGOwo5yYsXxxR2xDyoC+YjY1yyziVl3cya8rpq3gIjSgNqv/Yb6i0Psf8W
Q8KX9rNNf7N3NtVtuqz8K8KPLePj1JCGgzX8bKC4TdufL4mJPJQf9f67ptmwhiGDlJH7QFvPwbW5
RzhHQ+FMhwOiyxsqxiuP/B4JTNOfkYuwNIlevRbwCEPk1Mkq6jUx7ur7uSGmk3SLxgRHW75UsEo3
kXl0732v16FhNHsEJYYN9cfeTa1K3767sZuG/HDLKLcWNnpOmG9Mt7a0WqJy1MYLtbUOd883jtr6
dzPy9VV5k0VvgaXiUGr19dQVqaPlaNhYr3ZD0pWDBHpmMuVQX3R2zjNtvchs6qPb8yqFklmJVQoy
LaYBUVTTbmAR2VRe6bVwZZdj/jkvBu9VE4o1fl8+YJ0BU/iGxNrXGUYAH6Ij/YMGa0jOmNHLFP8j
9mzyKX8m/VA6BTOeH6G1PVdywA74w94vDxQLjU49qAng5LM1PA0TFxS5nmQWO7eUHLURZyc+CLBf
6tQaPZxtpBTfui7VPRi64qeB6Ci1MUg2FK6hm/c/pGFAAiE4gwa9NxWR4d9fZ/pPzWfKp2tQpENh
NyzabrXsZaB55RR4Tbbl5FeQdVly4hrX6XwnRC6S/Hu3Qj4E1sEvDv+tTCxjF+mkrUIFik5UKRdk
0tM1yz53qALwb447DgxZDr7mQll1U7Y/L06c67UFjZGaZ7zzfPfUh5NUfQJqOjZmfslcv5TJD6jw
IOUF+3g3rCGyAsDDKDAoOaf4aVULfyDIMTzF8rl+06wu61fVZrOqUb9Xl9hUiynDuWA/z0eYwrPL
ajgU9HK3wvkLAFpHmtT3KeRAnUGqVSVW2vkf8Mb1yrIsvG40lMx+wHquqF3myPQfXNI1NqX5aiK0
ScJ/tSZOJH0HC24SJRyHNLkB2eLXbU+OveIRBmD/J4TTW5VhWDg52KxPHA2tq+tOgSC5JJMfYqpU
6xezjno6zTIkKuUugO+DoWpK1qc99umD8qR7pasLVucs2ybgdRrD3YFTPDQyaOmR+T57fh30FwUc
7sVpOUHAom9YrR7bheG2NY3EjGhvviVYK+hPgKyv8oAySUFXNv0InX5W3igFFOeITjclGQrxOHQ+
2fCNM958yY2CR/8Rbjibm0mALK/D7rZCRvN+Tc87Hr/1tTkoLFm6tSdXbZWgufpqGrIwtnq676SP
ampRk/uSqvPvbQVhign/Pt9WRg+fG6XwQLeax45Tn4iHn/5qZEPdKMAbKIrB+oqmdPldyZA72GjW
FNAMe9pmkgiLmnaIJZ6rdKUgdBGCdBEcdkn0hQ5HRamearIszRItISkbCuuq7p4ekJ2uu9v6XLQP
CEfYx+C4+jSdUDA6NuF7xdXvvFFdbkv5kUilvV5+Sx+Z+RrpEOiBYDOj8IWR+Fjtxfnkw5x6X73y
PgMrB74l9QpfrNdr//2p+ojEwd2L8x2xR8MXRXJX8bG4LPv4qi6geWBMyCFNprYkJvuvcJ+XeU8P
R+c9rQxcWL0gDFHdgcEEL6qUsjhj5H/KSdWOUweVVyHMiYj8Vz3DrAcQBN3I+Mirdsl0n1pGN1Hp
3JXU5ENpxpjuHYDzKzlYXz5l0KzAqKMxBJQiDtrUHrJ0rntq3+hgGPcqcju4x3gEDovGa+xe1Eu2
MiIJ94M40Ci1LI6NzZ8VH9JAhA3zDvWbUY3qV+NCJb5nXiHCSwSO5LQda2H8FwKFPZj2Btg41lHh
m+12um121TShRXF53ihgI1xsJL9RHif4Ttb+kNK8vB7Z2cqjOaUWO5zuwa7IQONwlvTgpitMKCTG
xiJ0RuHBuO8gTmqMfvNdiBWM026e9kNj1F0RE85M3YQWu6smYXwre10nZCP87oMUKnusLoTWUxYV
SoLGZzPvjqK0w4DINuca2BgVTvObVJzRIYDyA7zkbIfJGOb4NnxttovLwzHj97guM+ZdHjfKQjlV
L+uY3TOE6B+m1R+Pg/F8dfRt+dIyo4QsZFZZcmcwAJCHLvK9xoyqs79A7tYViLNrki++HKs2tLfq
5I1H9coYvgjd38yQ/ntjiasXs344V3IAdmWQewUErW4Xn0ndpMZrWU68Egr5T+lsa/sFK8eRs4Rc
oLwoAlSBIh3D96ruI6F/xs8JJwTygQp/3JbW6ikiQo86veYQx10+Onxq3sySzS3pCzP6eF3Cdwcv
GiXFtjhxvYDWlLkniImWqYJ+hQLX9uuXz/ra1Okm9Cna1tclhDBQ4/MaSid1QMlsadchmikiAZvk
8exW4WLxqXfA0bEz/28Rfqz7kPSb0Jsm8GVFdoFc7XeT/RHbRjQEIlGGs4QSenq+A6l9KmrV+/nx
5hp4xfXcn5v32TCMCORS5VMBRP18jjJvfsrCxyUlzRtrj+0Yho++OS9FknfG3XeKwca3DVzzlKqS
BQe8cMdJCuaSHEzrPdOpiDImCdmKFGg6EtcQzPzBgOKGT2ZuKbYhAFQfaTdMROesXNyKS9Wo8a55
Tdm6aLgnmAnHfIWY8a57Uc1ULhWKcVy9FPlItyQ218jv/RKsL48CWurDWMegwcUViOJXQy3y3ubp
rqRWZERS2Pm6IZrZiWPuEwB+QKUf0RM1NIcSJ8Bii4uyXHDx7o1/NUxRpYUHRZqnG5IElM9PzuTk
0OHVdo/++zJOW/J9sIogBeS9Viyr+vZXZkjhP2n7BzweahuH+bVLDzs0vB7EncOEvhkAluu52TQN
hD3zFWvSfHdeHL7K+F4iIsjN+0sy5p/aq2oz+99i5PHq1DktjFyY1WflUO73SBCXdljJL9jMQFKJ
Mi9gQx+mmGdWY8Ho+tg8TmnO9s6FbtvhWhUpYqN9K3z1CTUsNHS4p0/YZ1blqoXKRPmjCxsjGRlz
cnNjdO1AVwE8P7ZvNIeYmIS3bJO8dXw9egAsibK+nCD0NndIsUy5UsAoz2M4brn3/vuioLGBO9ic
Tvo62pJZz05c+amQE4b7ee67tgUkGi0V43Qsml4S4+ROB5WJQjqjAk61bWo1DqZXC8Mol0Y=
`protect end_protected

