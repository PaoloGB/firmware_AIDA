

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fPF16TcpNgM9dNC6nyb4WjUK+7bY8P+I62AEEiiM/KOMhIKuPOHBoWeWL2UjxSNO68WLeYIZp8lA
I7rHN/CieA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E6OKJxjnDRUVVFwAhrQMAtoyRVVpuMKsXlca4m9CcIt6QI8vnYN0tf7gH3uVuxZ90322B7kUeFw5
Pu0UeqAoBaSyysHuDqXazxHy7oyk4BIWChvcrp7LULlVLcL76obtSwsXi1ORVmpdTi5b+AcD+WUo
OP1PSFj5jpodG+LwXm4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x+agogSsgbiI6PGyBpMY8RQCDzLctIr3EaG23mH5kJHlNmNKNolnP54yJ8Y7nIFi6yl6tlyOLMoF
/kxU0pyFmIj8QM0/MArMxPTiemXbDLS2VKtonyK9dDH7VbjFnRWwzK0Ngkas0+nbW3TqGPAY98x3
251QPjQoZCw3A7W9PDc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KNs7hA49BKKrboRSEkqIGldOa3ndCnhjRkSn8lL1xFfKUn+p+Wbc09ogKV6YYnPU/RaF1LbzyoE4
udPSNea4bST+08IjO5GAxXqUugcig44J+hzpGKmh7oO0TuyNbYq1CnYcsZXaD9vsmNYz8fBDoW2S
VK/mYa21mBKTOuTdQ1yp3wi73aJ1G9N6Ngt7ovDUrjyd5oNxxNlvWU8JkJDinbEnci0qjZ3Wu9Wg
y44pHUXf6xqwFYJpZ1ZcGRKl83P8p74+pLzt19lw9TPlTfKI++IowVjb6wo36ztNDJS0QjQE5Riv
hwbPU/Bt3S82MVCY5NAA6bKC/8NnoWMbmX8Wiw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QaRubtGbYrmCghuFdQuTgTEtoVYYLcPnD5z0C7mo18fwCG17qy0y8mj8xWiwE6bo49IP1/JXSIw7
rTBwHFOVrmbm926sWNrF1r3IHB83C5cstprQ1om7vnkw9XX87SjkscphhkrHmi08jjzW4qX96m61
/ymclz5TlAocMQJGz/jwscvIMOrrbuH4SkWQOLQnRfx9GIOv5Y7PM+w/wuDSeFXsAXz7Ahq3/qmU
cylNfSufW7/zfN4RZB4u+d28AXsuFe03aSF1dpW+uBK1xtNZccvj9h9NMN0cuwxt8ZUlLJw8l6e2
hqRfTTZl1F4qnnrJu6w8h8uEGrmgnQG1AW0epg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XXj6Nc59BeA5Kznlx14IKravf7ohERw7h0fbO7pT7/HsiPDCWh2DlTGpFUcnbNZslPN2RfE0nJNX
WMzLQtaHK4Bm6kxY71OsXEKm7MAIjEdLwOMtJTtlZrbm7chBbSxcW6sjWvI36jk5De3Yct9Ao1py
DpQ9NICUtRTwGG8SAiRkAXRh2Jv3rKvnookQrlVxIkNRSBMSgbwuTbq1ze/KMUZebBWwJNUVIC9r
RV/i9wjYXBOeCCUk+cGDC5uSpwdLXYV9ZxhQUU6C1ufAaK2m4OIUeBqPc2ski2O0qQYQ67c35k50
ynO8H9PTEROPEOn5c37S7feU+36OcOOAsVBTBA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
Ee3F6/2AhtVJEAdVw0LWIJftVQ32lWqZ4euveA+nZYSRa77E39rAAGffhNK77KuWD+Bvmdvebpq/
MslKKmF1J1GlB12APgeelFkH6EQm5tU/pnqkGExxgcDlKGS7z64lfLfxmCZZ5j/4uLU2CT7B60jr
s3sPJqieI5dSKJiQ/HbgwYeq9nbXxESdciVzrIa51GVLdamWftfIn81411vcaWqbs+xEqaW+Kkh4
+xCexe2GyAaQtsKWmlsGgparEB7iwAKQnxvhruNIx7h4RN5cxHNk7ZAm/FpaYCDnmdsQwY1JP+37
m5/uvjYmtrLqzgwhy2S8sfH4JgnJ0prmEgCliwH4EAZedOSxmNby+n07bCJLMw4voqZE7chQxpTX
usT7QMg3/9p/RQMbj/TfN4EWfEAF3O0j3P969HhPjb00ipdhdB+y/W+o3JPE18bVYgzupSsVVLA9
fx0m5LxNxl5owqrjXkgW1cCACtcvrf4JVQNI4QuX1o5xYxeGa8YLa/RVJUzIxIApe1iUtzbpVwZ5
xTrIXH6UCvF9O5YMW/jqPYWmc9MGvig3dJzaytlOa1CYUu7dIJgftDiKYF2nv/wZ0Ms5lTIzIZdb
oi82jxLQ1EjbtpmjFcFA9tqXjt1TdhgqPXKnPXr38B8q9nD6mnDIM1Qduql/rcfLtpzBviU697xe
9nzDUJ10yKIgV8+d4ODTb3zGz/+AlxNyH0L8AsW12ovAUEuAQjIfFXGjCocpGLluTZ49U+mIUfYW
9wvryRgHkth6Rv22tBEgMByivL49WNu7kK60JUXeRihysZGF/PrCZQCw+j/uiYg24HMy9ANiZqtu
SwwBcKdzfzM2e8CLOSxYRJ7vVKpo3Uk/el5bgWj1dH1D2zP+knuptQYB3CnkXPlUcO6fS1BVF+Nr
PCCFN5ddcGsU3f28f7RGDNjaP1Z1w5PZepr8PonB1jJLQwMd8Pvmh94AqEe9Oky9GwW3+aVteh8P
MSK4Yu7WbbuvBNlUbYYk26cDGo3GdH/aJe/lhssHF012rbe1OBt09crENxw3y/DYyb1uaH0IrtMZ
SYLAAGCkOlNTW27JtqcpmyY5ihhzB3i6VEE9aE1i14cnBxotVeVlCDwLTj2iW/cq6nftDC5hbnQy
Rc13Uz+KUjdoj7kaXlMA9C0aUYvstWNedX2AJrhYjw6hg74WWvoKqGmroa+nROWU05+1W+weNUCd
OPbHXNcskR6uK5pTSruEc6zkBAniy3NlQalmnzjj0q3C9Janz/eEM1BA58kJKBMNDOoG7PnhftGC
PtKEtgj89jpKdAVhtYwxsyamqbzkdq7BXET5L3YgxpYLCaJ30chpzYjftNcOsx6M+iq1ke6Wbzv+
JejND/QTgQYv0fJWtH6bp7RZf7xOl15IbwE7rFjZr38+YMp+fMzvwYq9fpdFfsIWK048WW6Zl0re
ABoKVUgiicxKA9as4sArMVYqGvReUmBXiXHwZOx7jA4f+XuoJch2bNRIQjBW5XrxYW+MJfEaD983
tm4olIU05sZH3Bv0nLqNx4y22peIiY9mRYr6tmnLlBZ+fNVtKG92iRdo6Knn27MnQLYGpsV6J0YN
LtmJkrEMZxMrfsf3CrO3q0cwdPAio67fLqkpRUSFfPYPzEKDCAUplYQ2JSsV5Qu6oUikijxESSjc
YZaAwapF6gUuqXbIDJyEP8oyGNCJw90m4Fa1I9WdRBKpCkxgrmIHi1UIeSrpId7nfCbj19pCCQSl
6W6+0cUxbQtlRPDKJH6vYBFvSn2ZfOZtuM84Qvo7FoZrGtkma7n5CVqvIPGg61dXklSJqjtZ+Nrx
9D6hqei502keuT45sRGiUagSJaTFI5hZPVGiilmFvd7eh5j00xCWo55iYoNp292sxPJWo4pf9tSz
cyW7Omf5qtPI2xKa5qi2NMSrpJxW2dTvdRi9eNr/6tecIqP8f8NjnC5LGqxBWKLYTsCQ/NKUYkT+
EaLN7IkD+GRi3+NuOwUxOrKehY1k6Z7s8ARZbfS088lDCwgj9oDGlh53BqFd5gnR6etIEljYd0f8
Gg0LVtTs31wxWiPuG20o15sBpNLjjR+Dlm/+ocalkNYBEicSW8jeBdSxpJnwu8J701kLVuZQBPRC
PI24wi8zNYUDjPcogpjKGze7xFrNMiHzBCziwT7Q7lK/u9q97Jd72TwTC2Egoxn3YFPJTVtjB65M
IdzqoeVXR+TdzEz+TwGVCUrGJr7qGy1FuUN8erNFMPT6rIZ4wN9smj1POgj0iovn1j0B5t7IUF+f
qQB0K2YsJ9D76/1SxI3tM4y0ytge+2Rr8O4bkGyLwiKYMi/4DSRvkL5jc1QAvndQ+h7jdeW3n8ax
kYInuzcmsUWq0vLph2+Q9n4b+EQxm/NaUd7Sk36VAt/b6vd/SDhQZLnfkefrdpacxD/FuM2RxOBX
KFqGJ/6tHYPAIUXPZLrKWFDEWBub8zvDN0jsWp3mBWm5pU9IXHELd9uLpEHRvgoo6kfeWl063rBG
3aK2tRRiMJ407tzcRNMZaJIncfgyeqJj+6DXbeLbELs4FhtD4M6HlQxHK2Z1OjSpmcv/CcFyOh0W
LEvpzwBUKy43Y/0FYDzqjV9GvD7yUgBibRslDm2yOiluXHE6YuRil6MVIwtRrCIX+LWNS+AMc6jW
Y5MloGcpxD+FgcMXEzxMc3dYl4/oMkAUKd7ll5Ig1MEa5By+MPUyKiXlI116MK4hofNtfC7dRr7a
+006QhNzmaFFvJYm1SQV4mopXw8wIs0zMvq11blC8A6i91nxKkKQKu4bwh9jDf+XaIZGWtxB1vMp
dzeR+GFJSxHlCMaH9PgMNpdMHP2e/4XHsEA/FhRY+eeOtOdgV1ilTsksXuPZk3t2rf2TVix2OaGO
z9kxeZG1CQvFRi1CJOhyKbSTVRG9QnARjG7WtG2JeIy1NnuDaAopArMAbcFFhDwivJ52mEHghW0Q
AKb2+Kz65Jw6WGkbZ2K4lQnYFMwvdK/3M3R5bqTSxFMuVY9x03SZFok0lfmWJcA3zJCtJwzPRNJT
gIQqxDy5Lzy088A5Nj8unNh08gPk25tsj6IbdAYjK7QYZhPHaL6cnsF6jg0ZyMs6kQ4ZnAWmGUzP
3hdiwExtNO64gnYt6omRzOWwaeMxefkIeq5u2OihHPDn2AFTReWFUOan3Uztf2697W5tt5BF48Eg
2hx7DHBkaE/EyaqdYUbYPaHefakjw01XVJlyE2Di1Da6dthRj1HMMpKZilA7wPETPfWjf8dpMEXk
xQyTlSYjyhs1VXRVpU2iufygZ8juwARj99OVbmpzJGKVa++7QpO62Yhiks6rkMk79RS34NtXDjjz
lH+oAWGn3yAGmdXxDnFaaFMxSdxxJSHZMABTUAB1BqsSeBtRenRqROwc4G9v2rAf6HnTHQyW++HR
t5Qm7vzinc3BJsOes380uAD60qFliQ8zS8zVxxJkH/kLL+kr6oqieA8YQDn6dVgrywx1cV73euaN
pwlmtlmEMw5LpO1RrXAynKFiEBABsHBRn1/7jgO9vRm01sz23TkG5SRCwMYItZcaVlGS/ecqic/F
XcLKCAF2uHepNjz/XuaphSfEo74QlV4MhN5s37g+O7uEMqSjx0J1dAJBC3u0UQC1JUVIYkpGld5B
rPa6p6T+U7WDBiZfSSZQHTuQsz6ZiOtka71diTswsYThsymwLND9VV/oleGnndEq3foNJtA14Qdu
bMRCJEKrAy+rCfSMA1y4ha/MLjCadIf2dH19H3QX4oWLOijZ/chktSkAuwbwxoaxzwZw7uvgEPoC
An2BFgzNDaFTSOGy11xWbsdWJfTqNBD2zX+4s9fH+u6LWXJUVFHDJ0ioQdeEEMXfLA3cA63VfBWQ
y4/bvhx5mNEwpZd6kJtwaLVAPsWciSBS1mkf0BId1WzHjdQCivsmbPKq6gixc6hGrNNpirxelEbl
vcOt0SBbN4DXStS4BNsHVJVE9LeimAq8PzyEBVIIl87Ugz3zTrwrO0KyLd7mN5EE73J2CRh1pcWE
VK12jwEdnLaUDgkce5lbLMHDZTIJQrlH/6HEquvVk9UZsxdxwRc5W0H5fwgyEf7UdLutb6BW2dDd
gdRrlJIn6b1N3whR/4hONkKhyxPuA9QinIQPJjV9aQckO4QO3w9nHKd0F9m2z62qPD+oRlUzhDfx
iBnSF8TibPri7o9R3ZdZSlEEkQBzeZsuqA53Vj4PoqxzMxpOn+0/ESZphN7NigwzPCNIl17Vx0zp
HA1+jkTZRZBLE5d+3BclFSG0PS5Nq7hTfp+68baeSx9oJkHlBjX7NoR8vp9518aMo7p1j4EFSDqF
kneISeiXw0QXXUoWGxJ+M23VJoCQ2RDalMEslySJNEhYFY2VqZY+V4rHiVxgGvTcT/UEuPFDtA61
FJG//7te8wPDsVb1t2ALBNZzxtiDiGF8nP8vJZBm2SZ3JSub3sFyWmQNAs3au4M23xT/m49BBo9F
K9nO0n/z1L2tCwMRzJcHpKjLslK9ugQhCQOmEoTu2gLTnxfWJj85ArBXdD3MGcUuTxh/01kAfFwO
zJYmWAp03H4KwfkowXaDH9JkkwAbQ7HXOtF15Fa0f0mZJzvGIzhdHCDMEUv59M6BGiv6sU+gDh/p
F15Zo/NeEihmU/kxjxnlNoPfimwSPFxFoPcNpggGwKGKLWdEZ2WdopuYAidiLvp2qpO0d8rVHpJI
Y7puppHqBZdHqj+gJ25llfdFlN03H81sILnXmf9zlvuEtTmmFBf+sFz/DqzMrrSmB2du8ZoFONTT
0Nu583v9c1F2Z/iMw61ujdpBUn2uKFE76n7fkEN0P7rd4bp4J5as4JND7vUrbnojwAePrHvygIgT
/cpGc1yXKwHwc9KsdzivlCssvXNlOKnNVt3jCUkOmVA3q3+RT4tZZZp7YV3u5FTaZjJOmyJEwoR2
MIHxkmZFIbXPdfCbZqycG4gZJFSCoQnfA2zm32G8sEgztJyzab/VPq+uxcqJIg372wK8U7kMyrrK
mnESvZaVyYCefL8bcrPY+CYbZbipTmMvAxW3K2yku2WEVYDf9yD0PdaK/gGSBvno2q2zAlfTJOY5
ZO0NdUWZ/S8jc1obPsE67QugLYnTGCr5DVb1Gp3x1ZCc/sOVa2Y3EeJRJFHDaNe9uk5mBv9vK+u+
vBFl1scHi6xzZyXTFWT9NkV3s7sq+pmymEqdfpzme8iE0MnMpzfpsdkwy9O9f6t1EvbbAO6imF3k
cy7XmjYhA5gNxKlhlKToIBVH2GiQSpUxbfba42IvI5C+a4I6cckzYyLiQjxZVdTDveHyzkqDTFMv
/1/Ux1s0IUgDHcC7n4OJUCV5VXfYOE92//aXVpl9OAHCTGby2FV5UUh2jA2uELrPRO7cT+DT5Llz
HxfQSY8DXSLMzbw0QNsCrvnVEg16H5ollaYTJiSk01PoVCtojND34WyX4DjT9Xtt1lMJmM8l+aks
gJeLNyqyjlocH9QOmqqERpgF4ooZA2b7ONRlPGgZSAGHZaUmSGs1bFJBEQamKtOS9gvH5gihz42t
g9pnKjTns4u9kyKPK0OKmeF6DGoD9sd451EjIlHTVwMcDPleVFr0vK16FgWPTvJUxJMC/h0CRMnv
4PBdu3GeudlIJipqjzf8f5aJpUnRE9ia4qzDKj25AKsXawcBIOB/G58lZKalZm3FrmwWlwQYyu6n
V06xB9DmdKy/kgiLWBlZ/pPt+z3jxNtvzxQeQ4BIe4x/Ga1qRxT0IXC6kMe92T1xlHwegu3XQP9r
DYoLIcF98VWlotr3EctSpen2F7Y6jlCSia52yrV0u/g30znX0ib+EJ8VNldxUC44UrduYTx0DuEk
70b7RYhLdG6UkiJ+FXMDnjwqkv5h1lrHI/eYNKl0e4L6E6kJHHVM9I3YyNb8ZnfhL021ElVYrhFu
iR6dJSodOxm2o+nKvGrzr5vxM2UR/G0wwhAnQJp5+tj46QfpRvGLjBZA0x9vihikPJpDLeFTyv//
giGQOAPa8SM6ufEGVlLZ8UGaVE8uAlwdkJYNT3JQBdq84cFr4iN4gzVEsXkQsFxhdCKjEHE6KRvh
L0dorPBSPAfJkg1Vr0vCzcq43bVzWtCHCotCIcj9JcH+dNwi7FUYbLB+AFUVzMiwx4wScvkYLNQT
vxkxy3TrnWU3Vla9+lSmOjO0/MV0YS018jPQiOgkBEdsDmPclg5eCuTZr7EMXphxV/b1Vo17QweV
JPDnNjO2d25Xje4FUouVk9ktjKBSSTlR92qMmF3n41Q64uqjBwI7tuT5iXu64iHh7WmDl8J7nlp3
7jGc5RAtZbMbh9oy1X6efEzZOT/hDKMWFYXEE5rr1V9qlaUwpExBuOjcytZXn5AxB14Su6p+Ixg7
KIs1tDpoeSPjfvjoXsp+bnCIO9SOH315g4aHlbtmh7/3K3GtVGNL1tCWgDPWGhItQlWDZvzgrZE6
Ty2Yi0DHM07tTRyHJhKtEdUmgMJviy7O/Q+kF7mgscrj/zGxKMDE143srFtR7+faqEzw/WWtgDZM
WaK/ZPSPCyW/PQiLkZ+iI3G+fBU3Tdy1F/EKrdrJOsaq9/YlJwvvRjY5haEmy5l1FKcMx4648u1w
r/U9AEE2+d6IFT69VBKyHvxirXkRK53m3tAMXUKS9nF8p+wXyK9Sxvrxkr//XZ3zZa4DOFXHwkk1
6DTb9h9rtlGwsBPEtbMQZOg3yH488bwMskbI8CE2NkuSgBn3eotOcGiXxjDjGZ7VVf+oKnUuTx4D
9lr1LnhVn9/t+d6UBk5jwXdFoJJtvlZpQkcZ6OhlYDLew359XqfI26eDwRazbWfmGygsZL3XyNe0
nyieiJ8RrklzJ8jZmmJFwZ2DXRqvde2SjuAH7kUmD6Ud7eBL5Py2GfHgtHXL0YjM4/NlA19VV4jw
h1OEYOoGwx4u+xLHgaSgD79JujlGupw62Fl2kSKFwkrdfk3b0v4bz/wvA8HbzYlSi680SXbbPuG9
qsuNNVsHu6JmbMIkr8hWw3G5e1aPYCslix7pqVsgZGqeBicaDtvtB+7qjGbtcxQVRdYQhJnSaLw7
ySPGBYLWtZyaRui/xdEBME0h/HGERYxWhfkPRf8rKvB+mb1a/fyA7vguUFZaDP/aC+QMP5kVprB8
8JcPkzwQlmK4qo0cWHxHpgNQtvOASaxNONkKSlKovQmPdeeLYheOPKBDL2Jk9IBN5wAVXkoGvsof
LL50tula3awfjOE8yTPEqEbiJ2MWImDT3yA0HPAe0j4COb1Rkxi5/EP8SZYM/7zATH9mZD15sIHF
6AZ3cNOhk1XVtsnU0Nj7h9RUOESyX4ikLXiRqfGzl6lWoKZU45gBw3J+ii2NoU1Zcubc6nnEBC0b
WhOig1JhQoIx8L24wkfnPXxzKQ0qj+axWe9y5NadLcVK9zKAAFmeH2tFkK6B/vQWN4Xx6ZYEDW8V
fwhJ7nhHLVyUy8TTyZi0LxY83YkzimkZMIhpNHz0w7y3n0LLMmwEKnb0Hy6SAr0gqU5wLMTkMQAh
DjKnr4SQp3j8ZW1LOZc2WfbVk9KIfgFmSxpt05OXrG31dIovJFZw6oXtVlU8j2Bsdg3St8kpkw38
vNDaixeY2zG69bmtYngRuvEPAvGcMGKz6Yh+odC85kGTxAbZ6w6Rc0gPCaS09tFn5dRcu7mXlVLJ
rrYhxK8cKPn9uQAgXqbHfhPbJYOgwoaQRuwzF2QQFa9kbxphvOYh7QUhC973eDTTI3I0Q1+ajOoO
KWMw1yO12O+VgzpPN9s5QN1PVhkAlRliOrVPyHx50ruEqSbkDdwSuyv7zNpGNVeyjfUru4WrM5lo
HXAsf5cmUKN1qzhafVhEnm/wMhzRo6PYwxel/eSzaQ6vJB6+8embdw4jBM9FmI6RVqlwuXWtCHWf
n4Ej/bOxsj+ieN/8zUwUMwk4hZsvlxXCCRVkGnpWcUGqKexzoL++F3V2z4xjdWtcJ/jCcHgzZGGh
3Oj4WltofcXnbFX8roeVw6ext4/Abd9VwIIC9Rgz1SOTqo27dc+0iNo6T0+ld1wxXT9WNe+s/bWS
g/ZHz1zMSMg/3s2OxeckzIa0LF6aHEoOxqXBNIy5Ur9mLsR0WM/j7K6jo+lr58YeUKo8BoYS2a/d
QWktuWNd4XAwV+9MJuooV5USiqRKeMCALNg3YMss4gOG1o8Pf/yP1zbNxdkqm9rUKXCem2XbvYZL
WZ1l+UkyJSoqntwp8X5UhI02bLJG1rKiKLCvGF6jG3IHY0nbmDIuZM5F1ICdM4Y1O2XNT14azhS3
lyw29sE6nw3+gWZuxDD/hI0AWnykPSoKMlAXiCjnFo2VMj4Z+vySwc8Q/bUdxz+x99+u9kUdM/OX
33vw7tBA4msYHQBm03+qBW/LMFQqMJg799II3un5T0A2zbJNPkNFEia3rXc/wUm6/6Ek/Lu+mdiN
fcNSSiNe6cu0qz2InkVJScgXh/7f6OUffCPXhrF3Ir2IzNWDPeQw91UzjkpuWqNDEzdW8s/j8x7p
AABYcnyR9lsmwugqy2T8+w0kYEkkunIERsniHYKlNDd9K/rmM9CjJSp58K34gkHn3+0bQyDf5mTR
+6OhFFi1dHcJgUPfGJ5hODf3ekR6xxFBzEMOxRzWydaHzQeoBtFnmNFDpi2B1mje6Jh61bjnGPn5
0pH0PclWtQI5RKKN3bNV3K5FsaiEY8Jz4fDDwjluJw6GM+Yh3OoAlyNsdMoPJ0Lwp1PTZrV9epJI
SlHlgpR68hfNPGu43mk0NMwTdaqQYv9P6dQTBT18xzDGZaw/daxm5T84QPnNgM2x3KUrzZLNM3Bz
T7mZkLREX+f6gh2gJ5Yjii93GfJUmlqs3dFK9vaXFEocjy8U88WWypTc7xf/i/BopzkW1M2sTItl
u+knBnuFplKIcPY4GS2hnM/nR0oZVyfz8NqeSwyRcw6ZSK/G7izpOcyOWQrVv3kY+Rlhl66M6hqb
3s8lr/yAcVI32zoGn74ZkdDxgXnefSilJZVPARu9kVQbZ969KdlxWQF4fUuI3IJn5Y5Zmz321x2w
Thdbk7B9cl1U9uGFgFTflT20+Vl6c1x+OR03oOrN871KK6PQ+RupQT6qN3FOg02AnM/JteYyHFbN
KPQbb6QVl0SUlTMwSliy0RLDOPHArmA4QXR/VGYNGVOfbtKSNOikiQrsVZwKuH28mJ39oxq2YWEz
4eknyNngdObOWcaYSD6jnvySdIER/vxT8fO72UcZSKkIIzsnadgF2+L8LkfkL5ixicS75TRP+QTi
2nbSane6v6QIU56hbojKeqggOAvxN6l0ZGdAnxT6muX6uR7qxz34lxTEDxOFYBtG1fS06VKKalT3
DX7ikQHYQbc+zt3Ke8zDgeYuvvip33tuWoZBjxZaqJ6hAOybSJf+AgEXmkmH1MmO1nDpOy/xbWIe
0tf+Ve/+MwGESZuMQph0xpeehGdzsrNObWBE4cvzn7C17esI40aJV4c9YXT4GJ5tYxTp9q4NARg1
U61zJOvsB/Dkn+9ui6yrPyML1VecSJNczzMIVwEyPJqVl88iJn97NGLj9RvRwp87DzfqitMzuibr
Tztx/rFUS1yWFJA/+xSkANESY5b8gi5Sl5B0HZGmD1apxWU+Ax8XutsPkyF7NDFolE5YG2Byh4ID
DtVZmQTD+Ve/lPEsMcoBZ472MkVxUUvrW8PMBjr7ZZoMQrtgo4hVU/YFx1vTcu7Wgu/ttxsgMPk1
YyB8SSyUhDp6AZCeosyGUNsXUk+33/jbqZ6MzBSA2+ZLYKLeIvEBjI3HE7WvM73sHBWgQyDtO2dw
BMGvsQHfuL6huIxBl/2HZ6ilc4KhXJ/OK3CoYTVqPZIN9dldkpZJ5eUC2kKkFzckIzCiYmY7ITDv
57URBEauVp/3wWDevvknSHmXTSYee/ER/j617HZz6bOEjF0uPaAdG+EFQhS+vpDIp1bZSamW27ZY
bWzNhhu2dxTRxN6f0T/+1GGUvx2i8vdFglPrWuF+X8xr9KphK1PmFL20UP9Ln8guYBGau6AXy6Wr
j1CXEfswaUYMSKZzIS+BGdb+nWKPnnysPmbaDhJrdC4fA7eIJuBVdcDp6VHaZWx1tb7+yBK4vwcQ
Y2d5wH3bwGuEdtPCHtDt5S0rWHGVR7qN0yvVI9zmxkKVtdB6X1Sj0M7wUDE0ds7yt8S4ngCqCyT/
Dm87cFJYBCm7D7mwvgM0qpaS5+wgVtVytSFL7gi9AqnaQZioOgkPWGZBeLUMO+UdIV96AleAGueG
1KALWuFkRhrlQEt3OpZ+yM8QRuAkIAgqMxN1591dWw1cS9nHPYkMey38pn7DBBTwqP4FMAJj5aFM
DRVo3mnpgwqtJ7rmA5yfYPz9JfUMOt7PooIAj5t9hxz/T4h17j5ez8/463kk/KjEKIP+DKCS+smB
P/KQkF7IDfc1HT/72FRK26IsSOcOXEZDNfVQV8bRyXVvuy+puRG2DPTEt0S5Hne67f+xOxAEoikU
lHTa5J8nNapvltY/hI0twrBFyQR6Om0iLgpNVBHFi6F81+/aOcuuW1l8tsLpUBbSAcPtU9MWRWLi
JrxkUstilxYOXxt9muHiGC2p77TacjrteKq1Dsr7PsdKArQsGsuRzSGR2YFXAo1AmpPKHRmGiR5T
AR6xoRNMT9zRHEfj/huq3v30cJBCCvIfBcy684gCMAGhBCgUapVM1NfqLxR3b0X9NAPWzLkEDNB9
URQh8Mg1voUMIGBZJP81jABPo/r2CVeD5h9MNfP3oKASU2qE/Gs4v6yCUhSp5773No7I3CwG86IW
ZkxcVvZGxOlRMnvl0IvktPmsbvJeZwgz9gB8+7a5PbTJStYkzArLS3xuNw1EeR9ws9+HJq5wEX2c
tFYGTP2YSpYCYpG/Vuqo+8FjyS/FWdE+5z6v++cUUrD1hT9Bt1MhFK2Er3CSyX7CQgFwAR//7TTI
Rh0EMosJdnAWfG5H9s0zbx2jrtTiVewCpJGX2mTw9+NIcmMKDRgvDlw7t5M55lp0fFSjMhwLJvRz
FGMvq0qTZqMr+5/Q0kxuImlimqyLpc4JGlZviNoHAypVD3bTzL/qV3SkwFOn5ExG0QiHNwIM1boq
zWeilTti6lG0/nKfich54oWgrsIm+5h6webXhZydf1T3AgnRww4vGydeVY40z6yJ4Wnx0rdw+ujX
r7aSnFINZPHOcWAppukPOXiJIHXh0fDcQDjsw3co1bm1ZIUzmE+qxi/pLv40O3au0qq0QrbdqjiB
bH9JEwy9wLjSlJ6Si9FV+n2f9Zp7ie1pK/ROR1kva+auoSOD7NncVq22Ro0xt5a7RM449uLiOyYA
CmBNzsEX2duLhko3iOJARX2V5/pGEwXpbm+9I6cEhTjil1Mwkx3u2i8lxXWprkUYtCFtcA1BBPxB
m1poXHNZFeAaGljVhxozocwiNtZedTt5xaRvBRoyuNySyjMP8gBjhhJh74kCFkMbUoudOgO4qFUB
72qfgOdyhjN3yuIax8coDcjeO7z7JLoEd5nlgXWFMQi6l5rcQT9zy9J2YRjxAhH5obLxE+XgzA5r
EPloYquKyx+K4lBu5WDWeCx01LJlJ8v22eLUnudy6DKfeEYWJsRcN5sLPy2nD5lHL59bbVnKi6n7
b3GmArblSiuVwNjqOKDNid+oXqpBPu5066i+50X9U7LY4fk1XxSOLKyTOqtuu6Y+SFwO7gaFyYkE
awCfmtxAQdP9VuBsyh0kcb1FqNh+hq2+v/A2e7ksKaxdV3tF4sOmIkURDWvGk9oV4vbXgYQhMb9k
3/ZT48C0q6wzBXjjn3H7qFa8/BZUvOBC4huyIistqIxufnCuHSxn5LNEbEwL70CJp/SMXqtWF8gk
TEOhDW5Z+71v5RvDG9Dkthjh0tmTAyfdmvTsYo2VyHjF+4hN/YCaQLJyOE3nxUDad4OjTgiG+v0S
NtyOjdo6dH278Nn4gDYPUVPJYxIh1LIyFBWHewITnLaajPbW6AsXdZOZodZAo4URgGTwE1WR6h58
U604VGhp1sTHGBanN2uUoHuuM088tnFLZxgtwXhaa4sAc0383F9wVOvlZK0wgge3caFi+O4wTULh
5Grq6rIy8+NR94zexpC764uvmB8TSTbqTQCDaJ0RChAbPnKehmmulDXnJcC63yXTsaFUrnd/8GrG
OASvYnLH4osZiGRnxe9y0SDNMgYp0ajxTamZdGb4phP5eXBeQCBd6T+fYfLp74R//zsy8Dp7Smko
7OQ5hEgjRpTb3gf+mQDqD2+q53oVxojFj05EUjPMly9APGshdF3+lfskWCs9hEa3eaGZBLtSCQaD
axPuLKRI0An3yJSPC6CLXALaNPGWM2zTqbLf8PV6ei/2hyBAZSf8LCmtfi/F7kaperHSvCXkKLgq
6/E+rGCTPEW7dLpLr87ATcKfBNQwKq+kNqexN7QNN7IWIE3pBr8y3I+4f641iEiylLagxS9zrBgF
nGnFfppsfWqqFzO2Q0UZqRlTryxFsmyz6FKapqTZgaJ4dJYZwyWiQ/2xdnHz8hi+TpRT9WupBbm5
YcWvufC0w+JsBETAArck3VaiFNtTiV9z4lQbZ4DwErg3VMZfAz9bHGxgsi7E/NB5cYcIqGqhhbc2
iuHH6pQuNg/LADAx1D9xkNu90w30l2qZlFjOGKu3SEASiuKCJ71n96sgLiYRjUhtpByoxMvueM+h
cD7JHBIvJNjyIIISpldNfYd5Yebucu9YW88DBBkOub0uC7FaYG/j3XICe3femHZLJmybo2+tp7Lo
M03caaWq1UJt7TFns4vuJAGVtBoiXARcy3MEShDg8FykebswNzHAttHAkx1bBfArhh6QC61Z1dm5
83S7JXc0pnQIvhpsjRIRcnG+u3/mnHwkaWuhX7Z60RtEpgForlTW44dTdxY6yNlrvO4huasHX9CM
jbFiUbcqK2bfRB3aHZo9+PYqFkdav8SWzLPtDs/HaeHbpT2OUCvz4Njytk5iSqWg1eXm53uiOYQo
4TGZENSvLyT74AsrcjK6SA4cT/8TiDzkoWvbr6Q+kbXREOefr4bSIWpm9JeZ7e5dKKsR+vWejPgD
0FMSnjEO88o8qS34OU6HSN6Ea5oFMZ/wv7JewhROBZB0QcWFzIJLsQIXEXjr9aFDjsuROeJgctll
N/j3ehFAy4vwKfBPk4Z09zSRpiugSLsO2/T2syLZp7ZQJcCXu4rAa+DhQy1d6Qp080BmN0SwOhoO
xqxThJXTc6L2O2prOWOEi2Bz5y/CcPcmqWVHCQKgDh/lrw6cumvJu8f/wCeZ1NOburfk/FHVuddH
GYD6kvnTBz3pO8I7RUIZkIoUgyfk3oNMyfWH15b7y2zXsc7Z1h1HePwoD/BAE3kC8Oqay4vQP9gy
VNkycgfz37/9byK5gUROHU0woY6qK1wQTMRHFjCnc1vrXweZAQhMi5iKLRafcmxcBMw7/3k1MV4c
nV3YU4OBkQnQ/1+Qos7aifxieTrEWldXuJfJwBZzxiEqpAecKE2S02UeIX2kJ3wXZ4XKxKnlHt9a
9OIAEy6+J7VpaQdE9AO0m/Ij814lTPk7Q8f3bAs5+9NRvugKBhStLMOsAQJ/89RXRHZ8fBorse2f
gWYTdAsHSKA/wglBrWXNs+nYLCU5fs2c0oUe93s3w/2MExz7CHUUu+omBF00TBwpMmgoyEi4Llck
/GRxpSC7XGsqcExPSoifBzEIKmuLGSUAz+J8BiajibFrQGz4dhZk/EYKvvcAWOiKuUzQDcy6y6G7
CTamd088OvSlSdJh9DZG7QsXiGwYZNoN42Q0cKA/zzpTlc+dCUX4KW45y0/920tvVl7OPWmnJrSa
vuX8NjLndhnrOCN7YkGsMSLCcoUN95Y16RVw48yrhC+o+ocFpg7OlkAW10MQmNPUPDfZKn2I4gwf
zPNABnJsPRbHzvHymJfU/LKc9+T4anRRQJH8+nJBg5PFDc+qVtrL83vCN7wRl9KGgEZbMP1vOvV+
RU4w/0A3PabhUY6wGF1UqBQy7G13aVkyZK3zFpaI8oEdsd+DD0yYP8UPn8WKwu2Ai/yz6I1pzWc5
qcqts69cOj0bZXwYW4koFlyR2mkZSVEyJX0jNRzejqTBndD0fRcoZ9Bd/ap1HIRkkrDHC+GU+oFE
uh9zTnrF4G8cUc+p1APeHsg9zMiWGl9+hSbB+4MutZaxTx0CZfHvM/iYEt6Np0WoCNBSu+ANttaI
mIfvk0qth8/H0hoxQc0DFPnYwlenG214YrqYcwiuL/Q82Xt3OqDailChsG20JQ6OsK8warscWxY5
9rorEq8+gXM4uCVyYwPU50M1iLcu7Ge4GwVy/HwhzFeapRta3ynreYDF/8oLI4KrCjrgY4tgH9bW
1FveQgk7vCEbcdSbplw1bYOO9xtPYsXv8fudua+EM3ChbfYdEGvBq+nZklNVWi36SL19Whe/d+Mp
kGGDsRJW9MErLLdJ/jfGTr0evErItbzhFvEbKueTrHwRk3JELYfPRt+NfrpTEiw/y1mmg/ZCtPUZ
nsq6IHEGILT3D5X9+rcCcspdOWWO5WxXrJayL6azuklfkL1KXuIEP1Op3efiF3GYgHyWEzgWTmJj
5JP8+mhiFqmrvK9of3VnXBU5o2zta8AEvokMobz9+puowI9GYjS2ZnkkfMom3N0Oy6aYlHnp8XsC
NcLQTt7hDCzeR/5GbauPrDEZ0Y/VL1lWtlcBvftJXNwrEhS0y2c5VQBrGGEVNuIwahDd9DVfsMQF
umKVAkXgLwK0EEMoTZuUTxrrhiEIQK84joqWkP+1ejgn+pqHbRoErQOz6HjQ1ICpFbd/hghrH8n8
wnY0veElcgjCvTnI3C7miB3JJrrsat/gIY6d3CTlYQP6XvoJSCM8ZGv9I1wPwX+Ts9Ae/dM2m+Gi
9XnC0NKGeqdvIcX6M7XW5a7/qIwNShzv99kVHWutjVRTxcw7JPBVR/t0SermQDWMSL3z/nsts/dJ
X8yP2vkDcGeuEo6YINlIhY8muM5GLWw9sCzv3IK+5o5ZLAS8nGu1mtSATVzz/liFSrRwVJq+hfyR
62VpN6DHodHkz5ZjG6S0aqtvcL3NECbqk0f8iii6k7n65yJPn557bisG4FdzP3Z8uQp81Zf1tyBl
FZ9Jx9JjTAVeObgJ3okqdbb/UlsreqT8lMYPSzVi5FI3jjbZiAaBMgiSqbTc+esy2O+y2ZvpFYc0
CHDWe231jxrqAn2litYRIbPlSTMhlaaUx/Vw2o5XNfPTTkIIf8LcdKh5pPNnF22w3vCK/uqbvGOB
tUK9EysqCaw8qcQKLgu4rXMVkuiqjDbEZciYNYSjm+rPT3AaHjEyVTS45uhifA9xCPrCf9t7UWwc
ycmdFCbV95A7VZBYOZ9rMIN/eZXTvNMVjhvV3KUrobHLpp0dwtYknAB21WkgxmhElgOXWUoYX1Tq
AIl5U3/xnxr5wcF6XJFuV6W2H6YCuhmrhu+4GPAcxsIj22Mh9l1BSMBrAqhwH+R6aJZ3tIyn9lBa
rGNy8Q411iPH0Bm6BiFzLxNralUwdq4BYDIeDOP+82BJ89Dcx/DcEJrMegq7QCNWCVCIqj1RN473
8MrTEBhW7k5xkXg+5yIAbSpLfdxXOtYOjNNNwE+yGe2J8Gv8nfuE8owl29p0Css2QgdE0Nxw1WuC
8/ZVlOcOODcTB1UeUBeCF0mZo+CL2FPynYjLG5X7NOhVDltzdss5r0A/k8qHY1cU9I8vLDiUMip8
B2HT5feMbIgrdDKrp7Bw3OBw17OkdN8eo+j79tsWiajeJ7moa1uMAHgKoeAGIW7O4JQj2R2OESS0
wYbXSqnPaJvIMVYuIQo5vPO0c5hK59MIz9EToO3tCLZxBFD1PfvtLhLoYM63T73RJD0gkL5b2JMv
Y8Npd1PJjwnbt1qj+ZRF6tQPuMRc8jZdvUjMa2RRuXnAWJiViU6LliGTwS1TDeDNHiE5+FdHYyom
lTFwTdIGTTZhhXY4xkyy5jZIki/gvYHKXRfET/FfJz5wIEjdQDc7UhIC3My5DaIQHStFKA4WG2US
mrAt+g8ZL1vts0G8m9ulKs95f4UZj8z9hXsymSXutO32GfvMv19D999+QcTO0LMS8zimPf2sa3il
ToBY0nkxh9JMmw9m2xse7XYpa2UBXxI8OuvBfnqcyWnkxUYcMpz6gtmY6AqxS9gC7syjfma5repI
BLYjsxvCHEMtJ3S0t2/tV79VA9kUeK5aWa29873fybSwGud3v5GlKNlZgnVgmyJpPNbii6/jdtto
DlhRwsiMRuU/Po2fZYmrgAh56qP3RYDw4mBLtRqJJ5cgr9Kkh3V7Cqp5BrZRYcNpZaKwJd32SopO
6OnnVpYDAEtQdel6SOWAMZIouGpy1T7PhwVtA9YcoRsDd8JMRLGfaZxKwivIJnf8XLEr7TuTq5M6
CarUi/KWcRkM5F+EMr2i1gNU6yK34bTrIAMhoHnp4/5S3CBCZ90wKSMu5QSMnmaIAeuAjBVPlWHk
79iEbLQeG42lzJRy2tPNN29+wezWk4nccFXSVKNcH+zX9uCPjXMDvB3qGuSLm9q1AVBHA7z8hlLl
syrcNhaFRx3Tfr6W0v2GxU4h9XesKfETleZz9vlFBYEAcV56CMqSiooxbvM0MuetFUAlSxHC0VnE
dqft4OrLqetdKf5U38HNl/jASdjwaXBDSDJBw0wnLSCQjOYKd2u/YkMOa+kNmfl2tOxROF+Wo8xa
ZAL/kFKYMrONUvdKjDRimu7FI7y3f38zM1yHJaj0bkTe6IynKSV9hMzxi0tT/B0jgj88M68GKdbR
G0meEPhN4f1EsSFmSUmJLL6GnGFd03cHaKjoACBTFSz0We9khzaRBeEQ5KoLeEOKvEfewN3VlAOG
JTqXl14A+RnVWMoz7QmXc6spO4qZ2toUph9q0qycsccG2HES2IOq0/Jq9HtE4TJdWiIqfdhFE05C
1C9PBmb1VAlsjId2jHXgRa5DfpootikyeA+X/CWrs4RsUtYXdrAP1xMnB1evDMsmOcw2kV7ITdNt
9K9jMCWSMhLfUNILsb396eF2vOEV/rGh5ZUfs7pMj17Vx7IIwL3/R63fnR+XwH4PspaXKlRcX8Im
Q3KFGhbY57OcrMsgUU8G99udZp59fzqSHyhkTkdLp4UNngAZK2MC+iRNxjHNvvnENxB90WSlO14A
tYRW7Qicqsg+4dT5e8y+YFpzxu4qXpmmrGc9kJvLGt2JSIn6v6dYg17PyHY4ENyAxY2BHlq2//sF
F3uL6g+CzhgoA4vB1VWzlYgupg8/aGxDPzBhtnQuBcn8R16Sr+XiNHjsBBaikwmMjJAqBaZ0rbtM
wfftfoFVZmrAStBjd+dFkuIPIJaWLLBm1rN0+83Vm49QHpi01AEjSAhQmB11EmPPquWvLT6XCgJW
tfZoRzMaM4fnNaqTg0aO3uK170j+EP9MXsj4SixwroF+wAjQELAszUAeyVRr6N9Ef1gXo4csE5Vm
mHc4wt1MNzi3WULxgomrCmIggWL6f2+gcEudmMIxz8KZOOphqWRTPisoLe/2C5Plv8ms/Z48n5Nj
R1WNh/YEzvCius2hZ84UPT9ITttbq2u42OR3ujA936oWbTFWxqPv0t5FC0RYWfyd8bdKPf11Qqut
RTv8Z7EzbyXudnj7UZsQKy68UZgSZlosMvWjCS8zejtv3mSQtBOOngjersMccRiUwDLCSohNyh+8
5LRu/iw3IbzgInSCCDloowo654efCb9f/Spc4KkuOV4YntqhlwJf+wfWqW/635iW075Eo2LihIS0
xRyWcSezX/7majI8yY/XeX4sNMNSnr7mkll3iwm/k44vc0SVWA+nekQtDhxp2N9g4k5MOvYif5W5
BCDVt3oZnoS8JGNIZW1jW3TOTO+uaS9cpEJSDmvYIS+M86RFfszJbpE0ZTzncG8oHtL+MuEt2ROl
eSlE5qHHPjJkPrVX6RaNOTn6itB1UeIyfrYQ6z26oMHAFzCNSLLH8ipCoDMbbhUwPM/T3KVm2Mzh
6JfzYMrcizxnFLhRVaVTrpSf9xAXat/xwqLeLNPTnP5EkqjIX9jLDB7Q6qxTDNhZOy4rd8Xo+25p
gvn1vhi81U6g01G53D0VnbDbAw9Dsx2/kbZiCCSgXHjyqNbzNSe4vMjHbKgsnWmLpxrdylSAKsb7
qdZTOuH01xqVuwyK+G+9X0kV+taVBQnhCkLjVBQyQatHEbuf5EYAf1jwZjDRM0ExnlRpdbV5AT6q
/iPv33Y+6DINdb7sNCk6F3+sKHxStROGQDmnA4ryIZxHbNMAj4Z5HZ+iQKW3O1d0UiaYtw6vjVNm
JVAbgqAOCL3hxzVgiEGqXkgHZ7V+FCHdaeki9CHI3QZ7ykDFDUwq28N5GJ7Anof1cSXZ5zdLx27Y
NkA9W3DoFzKvB52WUsCWVZQf02+95nLiJIsBw1GNiQnAgnbqU0tqdDja2y1Fd4aShrvqx7HaWGuc
yjzItO6Kzf8FE9aIWUZYEn+AfIBJj7GymzXYIcR+B0syMKSZ9QWLGBJPuZTOVntDn5VK/wvkXWIQ
eTt+6bzTsGDISHkVDb1n2xvonqG3OO8eY0T9D02YCXHfnlAYvZC/IJ6vVKzK5WooyddA/1yfKZm6
dmlbNYuvIxiKK0NmoEKKx/byIjXDcotBBg7jJoKrMG5G+RfnAHyEjaGbk8NBAVtcTimsjn8AllSl
FMUbMTUqPJXvDoT7dr6mJCE5mfc7As5fmj36LvL3VdUucbBDL9yJWi68ad5q/5Ian1zztZoWdfmJ
DIAOEDaOjmN9lu48pN/7rBRXUktFOGJ2W1+xKhh5dFyfKeYhHEhw0KBCQTTn+RcwV+9Bcn31zjMU
V2/A+sYEcrNvVpaEfBfRfLke3suAM8i9FuJfTG7zkpwAQIipUnLdv7LG/6zG3MIdbz9u8HEIP92D
gDCZp0D6R3ELG/NJHufN3qESR4iw/IGvh7B5cPv6EPqzJZot8nhh6+I+vUbOAhva721kToD1YhiR
PMCWgRssOpJNl2yb96vQQN9ysUQr8yiOKHIKIGL22Jf9x9QabPWGfFY48ktZ+gZ9j1B6oOUVijIP
4jLCnViYiM2aTbx7Y1OLZ3rHoNd8Vs8qZFs/gbAg1M8yIcsXnUAKin2gQYWvXV3NYUDx1oslK0eO
/G4T/sVOHSm6y6idHOm/TAWv2TnAvjRGI6N+qTqzrAOnny9I/mAJUq6H68Q1KRWW5+A7IHjOS0QQ
8jD5nnXNk46+yGorUPnTh/UpFbX3lErvKQoqmJtrUFNmKwsterPEUh4p1vW1L1HJlehPbG5MOxzV
KrtPGzvozMbIElMHSjW6EDBRUSMooq22wBbb7JWU/2a3GeZwQ6J7NOwaFpbi5E/afjUIgAWIy28P
enVIkiKV0cMxwMlX9G/yrtJvGwJbRM24RtROoVUJDq2HJICYCh2tDPZGqEZhFAHlZMiz2A70nkjn
8Q8i0UO1jiZuI0DPMROlsWmnBdPy4c0VhIV2tAw67gn6Us+mZaqtWmMmdeEf6aBFmm2X/4JLzhqh
VVGPyA+gSAPtavgLzYe9jmdRCgFgyCArf4P/P/na3MCuJmJBhOEH5DFCB42VCTOP6AGJ5hhHe1uX
ih5OcZdI/Jsr7M0vY091QliiOwRWrQ0ivzzf7cVl0tjz7o3tdAgpciAAnAVOLkSlcKkr2j3tEJTh
8MIKNS5n1JZoIGUB2uKtdOjA4uLLrJxFsAdhQNIDB30d4Bu53zxQG9XBNvoaXOcgNLJPPsWIMnPm
VWhe7oQCiubaFf3k488G4lhquAkDYnb9wKqNgPL1uNhguOD2uMsBUKWpvyIcy8h4pNODfOz7JO0a
4VcOwDIF355OfS6IJJq3PBRU7vGQQCVbb/dBoiXp3FuyrIALlDpBK5zavLOwBgPMiJZ+RCqE+0/s
gAvZlmzS2VR5WfqnMFxJPQsutebepMN5k0e3015wcZsjneuL044ZSVLl4TjkIzIPlDpfhRwyiO0B
fVbGef1DaBTm1dG6buzXnbfzxPMxSElshnXQJqdYXDllFvvGSqd0eLlg4isrAkAT+6tkZ1XMndCg
P/hT/ueVQNnVKbVlUiG/yxdSJklo95J/4TTEtMpuyDRp+zBfltAq5zG2BwZM/vjej3SRjGfMId/l
6fM8o4I6T5H9FkanNJ3zGX0s/WT2Goqs2ryYzZVIaC3eEsRlz5CcyRWf8+NZD2ysGliihfWOFnBi
6JYIi/vZamXnN1uI8ihc6op+2L9IOgEdV7b72lrXHx7zoIetLlC6PIYe+2pzBdhxKrVfTMabHiSM
J++LbDhmqf+ebw1HRsqnKoF6bIEs1fOblXF2BxFs2JHyhZRvauq/ifMt9KHdqh1TLECmOvgVqjzt
33B1MRpOY2mhRN6nK9bbG7sCWsWtktdX12Hc63eupNFO7SBSuv9mJ2xcKJxfj568xP3InD7vNs+v
QBQ69raai7GuNarjk60ge4ZLLJY+NZrW1KTefKQdU4hbVxrwQUggcfyH0nBqTNRrtQKwRF2JVmXX
90nLXOWezNoD0H3EdLy6z84xCEfv7RwYL1zZ7zUbp0c/m0c4F8D5z22tqvJuyEmxPJ0qkosuJrtn
oq9TzxNu5D0U0bpHqffLZ0tNXAQfK+znDHB0iMWnWHUq7P1KFqWNhTpjTRvzgCdH4fUMuuegCYhw
YX50RXwDAyYVMTb4YttgMCoJJcrAsHvhraKstbb914RmQ61eYJC2S51lNaRwqk8cvazOoRWuM7RG
30bUpjSJOHpsrYOQs7mgwSkeiy5oeeEKSaZT6Xdin+Dt17ox2XGKOD///p061D+8lw0MxOG3pPZA
3xLqXpUbkqrxjqu18h79FfTZkzm5qy8MaKwRobcdtgY6AR3M/kri+crkFEZvWzJ0EUc5tNHcp/zB
U9y5lNit5GSJYZsOANgbAk/71Y4kOPlahJDW1EUFO0Kj7EU+Szve3BLpzaopPSaoRrFZjFRT0h9O
scX732Pr46wFYy2cpkXw4kEAxJi4H++gZ/NzPMvwl+agrMg88hosxnxkIMi+xPiFF1L8zSLwiagU
b+D/vphz0JKmJhWYDZQ053SAg52DOG9BUOArHm3Jie9T0Y+4KhxwWIvIZxmxJvSMWhdNKCUtTxhs
Q4YyY+SLi2JBjxRcI7wJ5PvN2derQxcLZWlMisRS1nGkXZWtex7R3M7io34JVhs4Z45jojuerYJu
OxSFjvf6+qLQb9hWlUMCfrYjf0uyoMORhHFNtAI02/pwaBNm3g4z23Npmxf8DZ//Bn9qeZjkKn2P
vqpfh6hhAu/75bz06CKuRJbUQNdFywdATbhzoudReGUWZan4zR6QDhjSoE0UbyQe4gZLCJgZ+pxL
HNhqu+I0dO0IwbKxpFqsNx8sxvgGY7XmDXqxlMbeaR8k5I1956W9xdLR4uU2xmYVRX7zMwnN1+GZ
NB+Eh/bIgOfa1YAvNUBcPnIhD4ENtPi7S20eyvbCiO3Qpbg1b3aebiafnRoagTwestA5LWeoqH3m
Ek50W6bFwSfgLAj+qabBG6/bX4CvmX+1QxooTZ8et6EsDtJPwgYyvH3MXVoA8bQzIDDqrNJPXm1a
scySgUAcFOjT2YqUVJ4aHXgU71eTwX36jjAUOfMUn+0xqdT6u/W8ysCpY22/dFCH6gTmdTDB4hSv
UDtC+fJMoarbH37B2SfLDJrxlMMa40memCj2QMWrnU7s97yBnvEhf5KfrNWkp1gBG7hcX6fc7/DR
iB2oPCPiOEtrCG91rdKmAKpMTid9gyDiSnL1i7Z5DiE0BAWhk7p9Hl47ajTQVrdJd9ErR14apKSK
nqT4Zr4/ztoAi2Q9ubh7F3ZFsERRVxAgW/HD0W77jr94YxI1q2BXSpE2yRNmY9Xl+9gPTDyyCayt
44Qn2Io/0CsvPstnptC7f9Jy+sDpBBK1x47ofqSGgBvbgzSD7fzr/gQmwun2/ap2H1/+fdJmKXAC
ZEIK3isluFky+m6VPH1eK43Xvv3mlkwQt/jwJD8u7s/+jZ4MPkbhJwmHr2/m6GjW2R49of/qU3CN
f+yi2rq0zHPMxMujGRf30596huUde3OEg7lK+nMwn+mwVK+qYH1PLBuEV/9pyLdGgGZKJLrd9Agy
wXTUZa5UcfhCLqQZNkKB+lfakMN6+X82Cmh/GxxR8dEiSMk+YHiSTUJJoHjeQzwoG3y9+g3MvG/h
7sxpw5seSi4LcYiyDkwkwNZ6LbbwwpaaWTdrSDJxeIS8c4KuREJIJKVACUMHP5PJPRMQ7UFQD53J
Qt6QcfXCDDA6atoFceIy4CSodzqalnVUyOJ9M9/zqEgGkP5RM1dWCc18Fv+ish4Ya1ZPrIrWCiLn
qgO/1OkNXLtqducp8QJeoUjU0qCSw5f98asIw8rM+TxN3p2vpCa3qrD0ZNjPuiEnSLPy32GzbVFb
NvNfz3K92zk9Z2NefMRJM9FqaufKbqfnn7UGB86TNGnk72PcTZOxr3WzolfE72P8QKfAre6faPfc
sRPi3prFrUGyGg6l7AfOrAzTmd97O06/x6LG5/y8z3qtOhkAd2TkjYN8xQ/lEV1rp6Fc777kGc3N
KMVzQW8FIOgMVY5Y2T6OSUSdldYdO4sNkpL5s6q1L6SsUokq9uA3VLHnCx7yC6PmeYCd4QAInP2O
zjQmQaGSdRcVXVYbHMkmUazIur2IVz/PBDsc0yIj46qgtChymNAAcyZzmH5N+dybKVIILpxf3M4B
1oKeSxua5+5/KXxm8bLyWjM6cPVH1bYrmrGjOorEAEc35ta/SJ3X0XPu/aIVxRjDUdBJEBg/WPRk
UKLO9Th5CJPxJ3RJKcAuYGgFJN7R0N2Vfic4VDsWELxH9XLcXvQqA+ecvYPo6tzLE0fME7UmTwFD
2CFJjZOxxd68VHwY0iJqYcsZ+uJjQNk3oqCez8W9AJOqnE/mRixn8YFmTpe7VtIFheDkP3DqzrRX
5fDiXJicNp8kTHUiUw12JHV4G4v/83DUXkt/yzWi8f1lj7FkWhXV3DtuFF1sb3/dn32Z+av455z6
bncjvUDnS8flIvpW4TkGCExmazeyfaN0PGiGFvXug1NTJUYgcrSmaVUAmfLyeeMgO7N+QdhuyFwj
2iLFATRYP819W7hbwBxBGeX8p36Jn6m6rsOTj+VLFqKpfBmnjyqaIT7R4GA4+nLxGTQhLtrnAe6+
qh6y2OxW3tiX+U39pFj74VpDvgndIIbMM1acwRfuko97f8ukuvM1OWoqHwJLEot3JCHoEDlNlCMO
rFgwUhp48gohR64Sqbyxdv9b/R2GV3s2cUwiNVpGOqAVVF7hApm+sr0Ythlsv7P6RU/iGhy47rxK
RTxrLObzFx4Yzf1O9YBCmlwiNr4O+PPuZFClVHhN5NDbxSS22eQg0k/L41o8XG1dBH60tuBC6rII
NhbhGeNeZ1BpIToufMiDwduQUrrTCznkgA1Am5SrLyXidODAR87lrLRfzcymaq8KdMYpqMtBBMKT
RJVzDzLvdn0o/C86EspezOuffeQp+Iukf5gVTDJDMtfHwGVr7P6xrfJqlRGe67GNcx2CvP2aAAPa
xeTQW1H4qHtHRdxM3R2YgcntmlT1ZVbewAcYmiljHFrMapiP+e/yqsVWpZtf0yx3rQmhXwxfHGbk
esRwaq5wI6Zc4CIgXszyhfPdjcE+TwdPHQ7rr5aGmdNk5y5oRyXaZSockJyQmZjF1+dwXNze751p
6x0I8RjYW6zxTDmToU117aYooEtdOOsj8TNtVzTGpUjDR56rXMT1eBw0lPIXkdBeKDf5KUbbkCle
qB/9p46CQ3WseBy2BwI751gZcnrRk/ELpDJfvHM7Jwa4Pw89MgYZTC5dK2wcZkNDmTTV7nPFlFmG
FrOvPaIavhg1I+jB7pS2EexBEOqpo6UOt6OvoKFhYEmsLhk5tSq7ehNQvHUYInbnUaYFrsuOMaMM
TLH8aQAOHbCk3dI0z19muvVL1Z+xSWBRffkAhfTllDLn0s+pSIl1h0G8FJ76oH7vvGDlznLMsnCT
wAkB/LOnJQT6DDvyIeH6/9Z71UJ+sEm4zeU5YUNJnF79++AK4Vs+KdvgNZrttFIy8wgI/Uxcr0wl
vYAyJ3bQNSaHFkGu1XSB4vlmk1TLlTnBbR+V4bNpbX41dv8GYnRa37VWPWnN7EvaZ/yTFZ6lSULm
ft3Xgko1qJGdHJtCGnTr+drkxfDSvnHr3ZcKmQjcBZZYirlwIMKNstREUidaz7BvOJCMtv0Rp2c5
5NlBPdutZSJanF2QoeAMfpzEgn1VqSebH+HJ05sL5sl9fYLLmwjfexxGlSNxL/NoQhv1bD9FQVXb
mZlhIWNIIOmoeDSd4Qmwavd9+lWhMMlVl5c+5B+akMnNO0Hov4RQF4w/WNt12grnpfws+2mwBsIQ
P8DxS50aFw9xQapzZG9xY/59pvi4GIZz1PwKdOF7dFfZJ4f0KHI1bhT0vzvebUm8awZGEWFO5zYF
Co+rMYL/ulsR3V7ACpIO5+x8tgBHjlmjNNoP12F/y5lP7BFMlLo74GWNCZEgjiG3fYbgZDnZs51g
R3/SGuSVl60WJmNvR8wVWYLYDU/ImStTk0efZ6ltmgZi8jCwwUw/t4kQzkFpBUh+4k4nCblqi90k
Oi3HhqgHpG6IyPlQ6XU2mtINaQ7iL4kk87uxF1Mb2vFQkH/aqV9hlro/1cx/Sdb0pbHZM9XySFxw
5b+rIG8esB1BRoArgVZ9wqZ+h0iaLTlGQGZDeN3niwvx8e2e8ucoS5RQOgx6m3KKJPLYkyKVcuV0
a4L+RMTCi4FUt1Mao/Xg6C1u8tbJdDYtdrmXndxuLxFjhAokaGI0E4jwI+Jzuvw+jW7atbMFKosr
C8WdYe223RVz91bD84tBWS/MhpOPWYdgJWG0RybU/0uOo/br4BWY+MM8hSkGP/LVbIc1fzWcdC6I
tPIfm6tJ53PHHy2isa12lPqgYjRfH9Z2Ruw/Z/UqFy0q31BQae2rN5emzbohi18ug9q6x0t6ff96
sIM7JN9bpKkjqZq0tGe1R+vauVgg/VnzGYENFrZiGxHEO2aZfP9+oa66Sz8l50tZ7pqUsH7f7CCC
/aAnrlxRoKv3Q5TtDMlnjqYtDMTUoIvgHl8EnievBAkM21pXSEVCRkgNRH6ZN+1PBHMDrOJFiVEo
ui/WutTnrO7f4ta0uhHlFzsUALRjXuDiqit65VgX+yzqGzx/Bt65TbEcv8NTj18hMUTnoPSW3NF8
iyq96WlnsPtenfS8lDAVEI/Rmf2lKkMVWG34wIA9C+b+JIOw+ib5enq9qL2f19ak56VR72g0MTX4
CeNp0oRdUdGGJR7taEM2+biPIGlvJhXngAKKdB3QmW8CsnxbUhilwEVylgWhuKPUO44azTtRRA6k
q6agt6CVWEBboBDZrVdPBiA6OTKI/ppueo14MMSrLdFp3aZiMSML14qBYtCYmr4PbM8cQQr/mOLI
I8oNey6TwvEEXT1vcgBLG2v8MOnbhxU+WzlNyXwosnwHz0+XNrVQgbyMnE3yHX9zQbI8WQV6PNo9
rnYO7XAGfqXdAu3c5+WGG5ZJmy7i0+OMwV57P5MlzO/+fzIo9tdVgOrSFlvjWoTlSe/7YKdaAT3n
3NSIyeCMyLQoRg+G58yNDE1XzWnFeagGvwdS6UEY7COWBPM4XQP/72AnyWbgArm1W6TmWKygBliH
m9i/vHhAywaFEQrVj9hy1jCEFX2YfyEIfQxgp2djBfZ1rQKspxR7CQz1QqWlXs7MSdZpAZQZ4iQB
T1Sjbr3b3GMoLKtkIY4PX3GqBV6WalawTAAoswgwwIewefEOyq5m86PfBPqLVU5uZwdY8KUBy4Tu
6yj2H3g+ukP4FhhstyzB5SL2UTjQOnOqJ8V9wDj1ytiyv2Dv4awTLm2WBoSnfMcnzU2vib3Ge/SO
jx38O4IXjY0rqkL3nlTCgO2CIkbQOivf5ytlQNtdgU3ZGr6NzodMVbhio4bUwtV2V8oamOKyu4w2
HeMVrtH6NxmGn/RSgG1Fuhd29x/CyOl03FUtGtPQdkMDBHpWCONyUWBL5XxSlFrX60tyLbDj8TTP
3kFkToGSP4HCjhLxCZ9aUdH4kuz6Zh20/FSKHmN84jIX/YbNFlVipFiRxoBI2dxi515lGK6DuCH3
29ws26PIl8pZfyfSMT6ATogAMVWd0da2gZQaev1KVTftaDqwqf/XIZx6Tl9fVZmHm8icK0DrlOAD
4CxFP2DYSRr8SvyMEtwv0YReSnWzcZdb+q3icyhYGoXXbDlPOeRhECeB4Tat9B1i8zAv4d5PMHfp
/wdYwVrCtR+Q0yZeqOQpIx4NuSJ3DsrzVgYjg/wEbe25Q17JzqYz0ie4T2QUA7a6gv46LsnGcP1/
HJ2a7lsOCTmqAIWu1X9Ttr3jxXyx35ajREzLpHMJN3GNHmrZRIrCkZC8huJG8/B0Osoji1asNn83
T3MhwpBgBMjt4SFCWjJ7F3n40ufUXflBvyXZkXtTCJAvk3Ajzm0omkQ5biyukPRKc4TeUtLDSF6L
itDloFnRy3gKhJYu01RNddBlwCiIfeKrC+4/CHkhuxo8ljbqo/5vG2x56KgM0m7frjiGlQYV05rC
rlE4DIohm1Ab1RLc5HtyMYR5GiWTig3D2GK8WWEoE0L21fxxJFn9civBRQQqTWbY8qbp8kvImC6V
IAWHwqzD25xU/B1m6kwyEg2gQgPaYHypyAtvXPR/W0w1GvQK6mVTXWH+NUE4p4iUxTtV2J6KGw7y
6uaUx1HMbm5zj6WFJHNmPGkosPlmYrQ3dFffiPrYIf7oz+jirbyo/TnlPcnLMT9zpjSw4bynDOa6
FbhYr8ih2MpcSMb/K0s/mWIK2CC+nM06rJYo+FwbBZRGqhs/kTSjO48OHsDuyeLKwsaWXeN2ijvh
H6QtX1WMO2rzsybzPXBZ+O+ZhHGq38brbkdAAp1mS1wfAW+aCqowt7zPlGcOwVPXnWVL4RH65Y1+
7MgGArqVYXoKGYCsI9g6DaYOpOW27U538crWoWMRdm2y5fgagNRKeaEGFpxv9hNltkKjcZHEDEuu
o5HnpTXOKKyKCULzEaPDubjtUqG26YtyTJKJoQznpRt5F41nkSOn44Um+hJjRxpBdFDncl+VfQy7
V2mzFGzsRfTI0QQVLGezzQpPDsOvmQ7sj4za5mIFAjirNpO7uXlmn9V4L00rmbFXVbmTAzMI6Tol
FOZD0FiJzuPfiUON8/yRg0PdnOBApRNfO45lSsOt7GaReLG9uAqfCU22Hg9mzXOCKpP2mVrWL5mw
T6qgdP6+Du9OyE42NeXcOoKTLTpvenF1/yLo+YgnKC0qEJXeeKKEzLIVpfz/qq1+z2H+eFFrLcwf
k5qm8TGLzoBeZcd1xWyopvwLl2uXwO/rbPmj3qB8aI/G/0KPDSyt/didKyqq4ZbLL7X1+BjWwvKZ
zWlFoqPV+LxUE93kyPyF3vt1rnjyF5RMMZUY6h7j2BdqsBceduAm8oHTOQ9poVhdkY8boC6YNIts
vWFVRHA9D/Jko/vRJSZO0npx/aKS+XHR+8uqZJo0wkRazE36qgDA6xW5o13m/QIhmQbKSHHjthYV
xaJhffv0oIyFVxecBs7gDu5m1gfOas2P/Auh/bzIFRsBufEf2DnQLSwVWFB3uOGOUh+LmFO+/x4S
1AcngntpMpujBCwCVM4fqfAmssZKeNF+au8IXWcTquzBGWY2PdydAeEXUZ+LtgH0Tcl69sMAbSW+
F2SGQxcr4oxqWjjndMbXTzxXQcPv5MvEEsb60XXoquGOanNsygizKIWhAOkgh0PLH6233AxpjwET
ap00R4Kw2PqwIAnsE5PkWXGZWngLxmb3nOCuFF/33BZ3GGrcsdpWf/fjFdRujlYXBrmjmEckNPbA
tlnrfdtAJ+P4rj6V9jCvjqpqIgwNNiJoguGYHTiDobekkbGMsbExdawF6EDyLmbq0FFOr1NHAdHA
Pngd+bD5myuHugiC3ju7A3KNDTpcGz2knokhMk6IXy1sM82vOC72pJwGe055nFenzP/Hau8bx7Tq
gHs6Ig8B1bIo1SY9vQmv6LzCliDZTvLi8U8LJcTRqpDwhURzuradjcDFo5EkDOvBgHQfTsJsOXYn
onul85gr84vvKljZnP5gmIrdmXQh9ZByeOrugZcWEfarDX+P06WpYSrNXh5ixc7uD1tgiRnjGbfU
BjGu09DJZIQusj2r5e3r+CjznvzEghA2J+WNxClOHLRU9WLW2MqRf4dHmQZNEAg8n73r49pNZRfN
8KC5tbUTmKhFDzzqglZBkjymzeaQJf7wIUHWpX8tQgFZen0C2AcVSoJFYfni/bYAVkR2GP9kEUDz
+J1HY0TA61v9w5AS9FM+z9wcya7PDrdRwhu+jozLFIAoGYJ3D1nIkc1G7mN61tO09zwHu1eNZt0o
ljBFLfFo/hFKJ8IGFHvVDNJ2GsEPyByYQQ1gMdmqZjYtoVJmDSpFjj4BRXSiT8UXoNaqkWLRc0Wd
/3+MA7d0zE7hwiRevat5U1jBCH8SKddfAlJpf00/C4/11YiG4I+UE+YJMRtGrcdF0PsddDtAGGMn
S+LDMHXeCyc5wVVRx+OfMk09M+YINAltvXKd2dx7YWQGKaCzjLJZo8ux+9pdPR/yLqTiuOarHKlK
QhPyge8FetqKPLccJpqoF9MR55kgAvEgOaTJC2+rQm/jUen5EXx4CqR8y2dlMmQqTEDZOJiCqPdK
FKX9CGXLyEpjnSHDP64GGei1ABU6K8OylU8TjlCuKGKFIjZEDvdVnBNX8ujqRmL/sQ7NBPGOBD6Y
Q3pboRJ4NY4KlTJewpaxMZKetXB9LJe2UeyBotBQY5ORIbqZWLUAfMVJjy6bRF3MjLZNG7OXYoX1
73qtQuexqjFjRN4sDLQVDdGc7HnM3QGam3zb6XjTBqvklj3Raoa2qnfdpX9fe+XhAdO5CqXfpAjr
tiZGCCXTYRAdsM6sY9J7vd1FJ9R224xjEHYnFVfo1IqPTMEa6JTnd3Osl2hmBYW24mU42bn/K7vS
1KvQM+cOtFxrOKCAU335PFWtrs8ik1AAi2UTPzxfIMGkO/NKUShuFDffZ9wRXZpbhNlR9hYYNsl0
lGdsv+nqiTqIpKvTZwsjWpjxt6kY9ha1/webh1dWYcJCDW4rItHpvZl5Tsie/1vwAYjZGOe1k21E
yAHrk0yRMSiXN3LbC74CmLX5ktXH0fBcl260Nub5um5d/g+luQNihERJowmO9aQCyeWR5AF+bhcX
Gq7H432Lsc64DRjDSDozBD87FJbMaQM7pQ6AGL42cWJ5oLP7J/5PKeDYu+aITg6oWQr6Ov3dyAEQ
jag4q5gclFWsdrVrIIL7pF2kSM5K9F7piaYmAeyLHDIMh8aD2evJjZBfPhD/4edvmnbXA4vS/4n2
RYdf7XxJP2BsDWeQhKDaOH9kv7K3dR0vxHMaf6lJtnwXB+boEEW3jXB3ccQUqoZv2RDiSix3V6jm
mol327SmNWaCo2JDXqxzkCpFBSmQ+GeupgjcTirwvGv7uZuiLIM3lN54VztgpzqOyjekVE59+tT5
8DcHfZo6v3Wo5PbkQig/DeNP9EynW7GrTq+HXNdp3S0ddMZIqanwNF8EmK/lp35UUMW5i0rRM+fM
vE/gX/MbRc+8zu7uQe6aAd7HWMB3vqw4UepS3lVbYxxwkfTcPCZj9xNuwxo0HOXgoFGcJ9bsoMaU
GqO27K/UI8zHF5JyN/Bktdkj/GcSjmGfEu7FB5GrwJqvMl8zVfwDx3ozCgS4UOYvGOANgyguQGcc
1l6YbF8iyzWioySBq3eQfH9S3/IPB62OlZSodzKqjxSBTLsx178g5L2k4I6PIRVM1OzLOi0sP88L
+xkVoAMt/emG9oFc32AbOw/+EzklX2IAKJe2Ti/sHNYPViJsFCaLB96oToK6nTmKXYhAnqSDr5VE
uSGLu/6BXuZZUimStRWvMw3wPIic+OMJsD1GBxLgDZpPXMr/AUMRnGAKs2NIQYWxpUVtfeDtzwyk
LicHIkY/Cx1iYctimMjGGvTLDZrH6G3+zMWVoUMjw27Mb3/R1weSfLcD5fREXyi8vO0WbGKb34dS
CkoPtLClAfkd8wt1gSBHacArMlbkgVt3/Yr5A9KVjGUNmo+esOsSnixxZQyLeTFeszxBQWgwFmvj
kz6obZtbPEaeVMEE2lM96riUYT8umwHLk2t1kNf2kpnZzL3SKGrRy3iEfsSyY7QhX3uUcHreci/J
cmp0xwXu4id54Y+HcHjA6qN7ig+u8+wH/lzq95wXSkNsHFZkHJJ32G1klWccAx0ytARK1r3lKisP
NlsWbhDNqzvXUlXgTThewXKdT+VtxpgM9DluGr/dK7QRi71nsVdZhSV7UW3e3XeuuIgHmSkFu/W2
+RwI2r0o3XJ1+YJkHD6UnpOg7tyOHFRiWXGP7qYLUXhjpWTmFCKBtglvJVz55yuQLQpbi12ynep5
uL3fjCLpT/nQsjcYW6OoIploI0N8i7FJrlcpdsh9lnnKAFZEM3ulSpP848a1lyycnJVmhtbCsj5/
O4y9SulbRjvaBQbR1TdQR4uZMZsrmfuZCvvIx6kV+9NRW5B6ewtYWCkEZ7HLpVpoj+I3VXsQVDtT
5jGweOLqcnx+Ai8U7bgPxCM+JXnIWs1YsyPK5Etu02MTXndBXo9nC1+jUvRoH1WF52/pCw1dzUsZ
7qFeH4PkY8fe4SJN99Eh1drqNfBjb0IFSa22zsKsgW8ZHHLhwDUy8PdKQexwt12fhcNgEKGvPSoG
TOlgwK4S/PAQUTfbiDkeVxWOl81R63SHR7AktE2oi2abavgjX8MkVod/52JmvKCsC9huxrYK8aU+
nv1iU7d747MqQ1exwZA1lESChOXURASKvI0LfK+GETTHC/wtjhaAjx6qsIEZv2X+e6expcvfm3Qk
FzyJ7enEUQTYU6UU98BExguOLyiY2NQt7XZfWlVQzCEEN1MM0YDteNd1zNYNIwbxLY525fvuVPHR
NOhLRP2PA0+p5PM2evJXQCnf9eTDFsLIpyfPO/EdT1Ov4Zz1a3S9C834T8nLccIZGSOfRibvKQLu
v7ogqShKICMXrYvjgDJWxNO/eoyt7mmtRtKVWVjbVOAvh/lkWFiY+xuScc/HWvyXEkPfS+plBuEb
J8BEZvGWd6Ty0HqZbcUoWahgeNPCNP5qst/6F3OQmK604GACAPUR9NkBQthwVA7dCJfe+oY4tv59
KzuKxAgW+8mxmaYYmdbL/XmuiGX3E5Cl0+p2H6PU7F+bY2fSAESqxReU3zAxbDVqJ+iQvxkEwVJF
g0AZtP4CmXmYSjvsj14PGQlCcE/AyW+RVwxsxWRiRxECFz/kyqFiLbAMUQS2dr81B5kVqfN/QnLw
EYJ86kJHaZ216dFgYuTpMGfWXelPwdOExUcvOknXjcjpu0QKiwEFluM9jvfdKpwRwzdN1uPG562K
DQIID9XYlcLgpJxezYPe7iSIFfqmhUg+atRYfLtozGr/0ZjpUpmAjwERSI6hBQIXWikDi57f8Q63
H5Gxrrn4KzToZx2IPJZB9y1kMYbbOQG8H2JxQonMs1SNu5jHskPH3DEvotQ0yMjIBIEsft1ERktb
auZAdTsKFkim9LpcOyjBK2x18dmWIwjkAU0xkVdnho6tFhut+bhoqlgHVpxTGUZxyxmE1EbLWeup
CC8cmqyK5n5yZmN4EjjX+qVrnpyXMkSt3DQq6Bzjcyy+/EGczQMrbJvXfrKYm5Hj7bT7glXSP2SB
bLTmy45yflGarzjx+9RGaZ1iyGOFbQUvtnho2tZMTH+x9YYCvHP7xLTRogesJdQlWXDY7lfH92cD
zHyAHDV24+Q9GubKAt38/ZaZ7gnlVtn1o4fpHwcgCNFSuYWt1SHAPIcpbBUELu+6K6onOUn8Le9x
cPKQMOt4vUI/0Aug8WkfoF+hvrYYjkgRRqskLOSAR76FNkI5qYxfLMfi5jNg/Em20ZoAm8Qrd4cf
Qh+MMvXwcpEkgq6YU3mehgia/aI85Z39lpfKdvvDORJb4sg1Qki7Mn01RSc1dImnBsmxEO4nA8en
CiMQmjwRWX+cqCXRwde46ikHdMkddN9JwXwE3ZQqmS75Ejw8XKWywoJR9elQ0ky8sADUk3zyCrou
xkC9IdSB/O5GklivaV9Okt7H1C1QRCUL4q6T8+fly9ZOnD3IDj3cLEXmrGEbwT09shg9SqTP16Vq
BrUWB8E8At5/dttZzLGuV1JVKLLBkAeOAbao0RkbxzWT5K3x6dNhNrX9BxpILM7OscZcTve0tZ7N
1EkAkrr6iR7ssgZCHdzW4ESMZW5Coayx8i6IEEyMvCHu36zYEQ53fzKnOfmZufeDD5n9TBi8m8wt
8Hl7KBsrLaVk4F19asCn6y44by7r6jPQeXX80Udd3SSOUDVcAiY7IWtijjSeeCDdCjoYqv7xeqIO
g2t/MRfK8mM5ll2+QWZbax79NSdNVbFlPr5nLmhEMCCpcMEcF5lgb0akQn0xcsFW7Hdk0R1IvwJ+
ctbcUsOAoXBj/do7L5n9EaRTACXY1cijUe5kwyJBdyivifS2ugtVAi1/dTtsw8m7ZLYz/wrjXXNb
8jIGOpAISakUdCA71D6weYGvS1rJC0NVG9Q9An07Ay3J7Azcc8NJ4ZwPSpPGH0CLMyvaDndMsSPn
mwGkzZpPu3wYX3/MxadM1sbtVWYibk1ibVWlxV20zd8uaX/KDZ7MhoXqAd9rO7ItL9S0IbM4B3tR
K/Lals87NS89dLZDkrY7gnVmypDc1SoRVQTSn4MnWSlGxKbT/9rsY88T7d/Hhc4Bb/YuRMkhT4mg
6AIossxXfeBcZXPK1bofA1WsRhGBitSGZysXmJzTXuTdXd8ACZal/HKA2UNqvr3S6oo1JI+AmZ5g
W9q+PJtIKcKH39sCONCherqCPzUS0XnUPbFJAYxY+efa5HyVpdJ8bQCtf2mTSkbBAp7rw5dIlgzg
zV9rHpJnGSTCjiTkteYLpEFLDcAlzOwKT5b9lLT4aWxSOV9Si6U+LAPYawa7RZKGI63LMrAkJwId
fTmYVsLg9U4MtEBfcqPOj+fKcFCCTey6Jv4Jkmc10C6RZQlqwVzAEdSgQGJHbXUnHrK/q0jQE8Ug
kaWCNv6Y8AyqEvdo3uOb4QJZoDpdo27S4+VbM/gk5H2diniYjBAbqWxIhOYYKvrjwP6dtz2HN0br
FAtWCiP+saMYzx3cHCn1dPtp1a7O9ODWAp172AVy2niuh9cE6S+AR1KRHL9WCiajmuvGA3Q7bQCC
8R9D2EtM+2Emg+m5mDk/ldtLepIGw3X4cnLNF2QV5E6VGxtb+aHDZ6YvLuuFHcoMzImyL94l0g+b
k3kC5pP3mJm6uMuevm4Bv5H+Mqkq/jSL/jqalvUroUZ1AN3knyr5fiDSyo3iblqllKSktZcQvOog
0zMQxW6QS7Rq8fbSw4uqZP0utDX1cel3v85Ij54rFEpgqkTwxWmrNObFpHTrwp2C0WEfGszS1Vrl
O3iXcm6DEejiXsZuUqAd/UuRfIH3epR4Di5J2/aaG4ujzueFeMqby+TYfap1llBnKVdcgPiYabuV
BXqnqOJrHTd3BT5kHiySHmeAlz9zvMA8MZyoEoWsQHYSWPU2/OZT+zhHOAvsjweGWxnThTMl0UjM
yNIbQp/UlvHDgjF6DdLG0Aqf9hGg1Ebyxc/rTSg0ZLiTpj2GH4+GBZqkQIlfzFgMwfEy7z7UVuZ+
T4NS6BUz+E7ziaN8yIL/EYaAdgR/bGEC/n+hJ0Zkvh16FO7dmM56OgUjtbKoMToqo/8Esw1njX9N
z3IWxKNFxJ6xN9ujA1g+FfPOjqukPxI/zf9mi80a6IDjJ5rn3+oRLUbXPLuutCWSfmyk46JA3/kr
PDnw5vXOIXbNulY2ww7vWppSBem+zjnoC/I9OJzhN/WYpIXPBcsCdep0aH2fklgYmhvAs7vHXA8j
Sv6Qcgg8mE/RjfdSOygIkSilo6ShBGENHHLzqMA+vNrKGUUFDY4ATaqWLNscmXhLBtVpXyn2jReN
XWvIi/F2Zbnq6RMirSrzKE4boRn184YCuw4QqoHa/y+J+DM3DMcOyvk82ydEqfT5iKhGk0YVhGH/
wztV7tlSczpNLRD8jDQReDWgXS935ADJjTJ6os8gYDXNGXREyRYeVvZ85X9gB8syWOw2Ej3tjcg1
Fenjaqwqhy1Dzcbc2uCMNYniondpXNem9xpGB7kiIdkLQVRF8seHxQNZNChY0sx2vkwICSQWfEmX
RC5W3N+PoL67IdSW8qt7DCU9cDb4Q26JxYd6bSBDPYT33Du9mxgxMC5+6VgbcGD1zIGil3h96ZHQ
oHMPxuYXzpz0sGQyNBpioaVD3LC3P5gPJlpqg36AUVkuskRmNFaIlxOxmtLrzN6+Yp7XXrtddKLY
geYLdAzSkPAWD6x4nOtmZTOqKLwag6jUVD7RYFquScwOZ5SMw4rTANi6hygeuBkoG5aQWiiIDD0L
C2cE2hNW0i3pXuWus+a8GFUpO3VOW1d/U/sNwpC/EuO3hlKEjO2HzmJkzsGbz9cOOdEHiskc1EjN
Y1elfaHosMab/oVeEWlZjZatXRs7yHDUDLSgr6w+k+Qkr7MISKTfRCGx+VOHM6q0nM3eMYVAb9GL
T1lJaUSBcJf2OrysRqHracxm46HAKqjwfC7n2znkmejlJ0rR7FmuyscKXPuM+F3HVVin58+hLMn+
+3ZuJOfaEy4MpLMVAdNlGPQyikgXD/ddzA0BjOqb9yzBX/sj6uYhfhAuGKjLzz0a055LCBLDwgiN
/kfpNPMkxQUNWzwjnF4gv/iexO/jRv/Kj/9Lm6fHkXne+Oxa847KtMpteSiAsQ+eTzg05IPAfhFl
UJ1RofzgF/XcDJPpZFmsX7NXnIs10t0XgunL8fDQVNd92FXXRmqrGr7FX7OQKVsrwHKgj6AdSQpn
E6/NTNHPtelUTzMfk2qUXgLtlm7rqNQeuTraK+tnoXhfjn1oZ1fXO2N9kh6ZKFMIzV1zTrDq3voi
/b50m6mU/vlAPGOoVecV2nCpaR4F3yXlwxri7YgYkjq4i94J7FkMZ0STviWEQaFlOQceBXfmcGck
vE5ZKmifuUjJQjBLT2XnXYoVCHBNdQTvZxY+/uV6MIvsbmBVOdsoJnl8dTsGjH9DNAOwboC5nXO7
WMSyeAd80CcKeihRkVLPYQ94kz2TvepMiEWyWj5qz/8tGhOKuWg/tWqB3CeJUUmeO9HwLMgy/QH6
jAOTdf/d6OJ7W+gzheozosvcFFCACvU5jq7ogEaGmuyppUjnkzWheGNVsRaFCeRWAD1sg9DHywvW
6o4Thrqilxdz40NzKYf+KWF8Mtz4T9ryxCyY3E/n7MldcgdOoc/qgkQ2KPrO1ivNCDZhRdPV5d5l
A/JxIE06dkppvgW/TpYP9Zqx/USWUzWklc+IGD3UIX+UWY6LDmGojIh/ErgZ5XlE3XxYjqwLni3g
4Ldxdgyr+Ybob3jPcLPe8pEqpd4xODt8stqLZylgkNI+H8BYwZZ+tB52DBUu8Ai6krHNBflbAN0j
V0KHHfoNL/RRvevokOVdcKe2WtoSMn45bDnsuH7KqUUNdVqcr2oH3X3goRY/uCTUdNT0ZPWjGAme
Cn5sFcu/SenXD1CvDT3Ob2vrQR2at7hTLTD1l2agcdlLeNuoG0GhQiQtrJRgn8a2DWJnPdKmi6os
BFDYZ0WG8vhz7RhzCsuPtUGFIb8TDnNcuUpcFRy+nlTioNkeSIx8ucqBMRGKJFHVL5/e5poBG7ro
7eaYO8juoTUZf3FofqhM4YpXNWI9yRcPVxB/GuyVNCGsmYI2rQIn++rBWohVeNmD+Rk4ZGXP5wIo
jFVpTd5cc/KhDTwzXbW7DsgzAcvHA7H1xxSfADK5ZLklaTHUwPjOY2P1UiEo0dvGhj7chiR8dItc
aL0vbPsNzc3heyiP5CsOTPTYhL/Cc0CgY+rlElT26hNndEoEIdQm6g1tOezf90i5HgxPzLZw5VZf
UMzmyR3GEdDoYNRIhdUzEj27GCr/DBcf7o4aRUiHQU9KAkRF4MN1d4ni7OQPXWbRE3fsqwFIqbpM
cyUm6wEQTWR4vZOWCWdGnxTrrqKTUZC8NkvRHkv/p3Jz+aXsgvGd9UBAhXxoZ2bW5+0J2QPFCv2p
XnE4cavZFYHCjkpk6M+YZ3fnZ+jiiJp7PT5aR+gqVPFkFyKBoxYcQ1gVrUj1Z/r3YABNnw1n/z5a
9XAAW73wcoMhGALQ9hH22Vlp6jvpEYV4mqqmyX4sPw6iC/C9F7TjWN0xUn0DEiapT6RT/pPt/LVd
30UnWvguxCfAppDT7HDAiRNn381L+Gp+nHJJWFp1me4QJR+EmqRjBXWE4n3Yoh7eKj5xOHi24R6e
L4GUPmDglzBx0tDKDyFKNy5TfMkMXn1iPX8BGkYjpRK0Ucru15D8zaTE300EieXT6Ezs26SWEED+
PFvqPotFzrX/optEKfsANln1Kr0Zywqdbp1Ob+4V5lVBMntFQEt4TzHZOdzHITuMfdp50ggpVs5Y
AL2X5gppzjVk6C/8Ac1NfpLlpAf+6K5yU/0fumApsBBUKlB+dApdtMJMwrsLlZm6aedPsWQvMfFM
Sx5Xkq7/utY199WoJInmw57WPdMZxTCQbKPD5iVSTH6w29CYnPNSFMOxl5ygVHdXMzb7g2/AtFzF
j2V5Yhf/CnsuDypXidMcl8cV/ey5lYzHalFodiGd/rqSXxs8U+x/9ECoC1wSgGbDDD7iPQYWWLUy
06Eb9d9pNDe/htwmU5txh9F8tiDDVpfYXuVBqWRw/PRryTv0eTIIG/wTQbUPghC/tAV/ezHosCiu
3a1vR2j2h2NLwmHuTukEXAAOii5MJ6S+r9ejzGtQy83wPsrGD6VQ75YY+XsyPvAw7C+v+lKvk+8G
RnsjKFbXrr0mKrKRtWS8DohNns+A5BBq2jK/Vmur4SUFnQMRgYIUPd5PP8OXHE8Y5mSTZrrvI/T5
/xu/jdsXy9xvQ2somC9+hypZkBuNg1gc5fXDc/us9O7Co75+RPz+aUp84A4jFNgj9V8JzQj24igQ
cExbHQwoYs6M2DzJqHjijekSwgmiUUha71gc9btj8vuKxheEpMwZ4HhNezzxVmhEZ7wsXZEpe4SP
8PcLHp21EK6kdGPx0RkNk5Gpa23cHggkAemkW9zZ5AYxBnvwAwuy1x3C0rVt9ouzfqg83OARZc8T
j+sn8+AlaDe2qH4wfvsMEQjBKeYSxncnai/RY6ElHZ6YUmPUwzgotIU6sozyut6BpXTHrN3mxvBr
tPEZPk2pk3qOjW9ZhdgwUPQSxcXIFSWGhy2aLVMWGoLckiz7Gu4DqdiRA0yl0SoB1+CJhYA86191
QIJaMJwh38dveCiJLg8bqYd1Y1Z71puTuSDOTjvrGFlAggUl4/Kxfw4knDUMoCAQQtrpuuY1GO2k
FUyk8OvtO9WVGmFXX9K8QY2A/rLDIt8m9F7jGgIt6Ry8JGBTYuTmymqOAwH3sG3LwJl7081JOf/4
EiDWbmh3oSYBhRpXIhxZghZYI5PphhcMsadW17xD/p0uWBG5i5jcjTHlaplJxw5UMW1WVSTPa3P0
U0/12TJotfZYssryJBNWTBUbfbwrcufQd1uOge+HluiVA9FwsjGMbKneeppcLARWEI7cj8uvWsus
QhEAbUTespnnQRFmn29GJbdlx8XOr8oEHkRNDaXswR5Ogea6tLnkv9el9+tKBefiZC3ZMdusVCr3
1aj+7iWS8Tvs/pgXaLA0O7l31S7CqHbIji7735tppXKbCjXq+TD8JEUrx7Nc0Un8KZbL6isUKsSH
KpaWAGwVkaZDVbHotgoae1cauGis2ga+InpLnN5hfF8hwTI7jks6/e6YQvHr7LWEviAHUbE/BzPU
qViXDSSmPtRjOLrfAigdb4ScvUqgNmmgJ/EOv0lOfUTPVGplKoJgM7YBOwQWl0RFRHza/yBt1gt+
uffH9BBN6DinO4WU8ouWBiUnLRgdWHh50iou702xwGdlPstLvEYuaObiRM9jvHfIjcYj2+ZJcGD8
NFJhWVXZ5M4KuJloP95wRgxjDv2xLxRze8qQozOQ08C6whfm5f4clJm8fitWlH4s6gxEH2JLJtS9
AQRETTsA+0Rwibzcgh0sSc2aAg+ztJ50xyVFQfZGWts1ZEFsI8eZ9z5J51zjej15tD5GELcXcjdF
Ru6GxRfbb7rEOdzzevqpiGndoKtreahEwgICP3knrgCiK8J1+AAbNr31cJYhevb7rR1/lY+Qx1fs
eQp44wSGhVJ0OZFpcUTiD0vbGiYYKEa2yYuT3yy584+p9rRAjgGOziiJIuaAWEcP4JI+ID+lU6VD
lq9a6G+Ef5ooJU4wycrjZ3AzOLsTPDTjlr7GLa+K/xTBrhRX5vH5dBDQRjUTQs05jYiF0S6rGHwA
3kztQpRLqtb6PKxuVwmSu/BxxeAlPCBa+nG+vh04V3lXfXD1MzTqf9izP+dLNO6uywY5XMJuOwgT
6ePlUbjvHARi/52x58PM58PWFJ+iS03bHHAhb8DpuAZ2BPbxn3nAOR01PfztX3GjwFKXa3PMWie+
YuCKX8482FIIspNw4AjwLX8C9iA0vlO9Ql3PDg4UCT7IzGCNchN90HI0QAq+1eOSQF4zV7Pakyjc
yGAhT7hqEIq432C9B3jzNyNx0Y+21S3Lz1L4/mgA7OKafneBLnRo8Idpz99y7/MQ0MtYwoB5Ye1R
qCiRUKXrIw1bcl/fy718cY8OCaf7HFsoWUfvED4Ia1dxc6U7wIsvnQzO+cX/vqbbQVGjlOCUwr23
mS+PUS3u6z8dt3n/tNaPib9oK0uijZV0guFndpQ+C9pgpI6jWi8CtyhuKyuSV53E692jvV2S+ssU
zw7yv3SMu7a7XyCt2sWmaMwHostMkeSmJdDVBKGx0oIDGtpUkyccMJdtZaV5YE+EOQHF2ed4RKOU
in5yY8L7az9+xIEJCAn+0us5Mwxvpj2yhvP8MvscnIE027tpcFYPvbY0w89K94SWE/5kXFMwBE5A
sJvHDchPPFqPSMaWFPpF049MPCmzEguBs2FynQs8Ofjn6s4D9ujAn9jXls3OM41dbAnctRX24hX7
ql0LNS3v1tT1Btvo+NkSdqAZ+GbALlbQApUCpms+6mmwYUk3wecRT89bl3MJkbxboGbZjbH6xtrF
TG60Xw+rXHzLJTcI5xxj6ffwgFRl+twfC7yNmI+I6RArUvwPdHFmn7Ucwzbg99JsQiFiURNewlTH
yW+2JaBOYOspiluSNtGsT3KQ03c5QF+iQm8ogIYLITgLjKVq2cvOJV32YTtgHAoWIjbgysx7HO92
2oaeqUinpXlGax7MYb5qnEBUPHhf00FshefYmk0GFbxNdJIjN8LUpV8GhYrgpD1kjuVPtydzeUak
GeSrWkH9m9gW/rv3iQLHpah59zmUWZFJTrqZ3DKphMLH61w273SdWS5sSBXlDIVjIHMZ3iTfspJ3
e9ncee4oU8Ko/v8LnrXn4jjdtyHQRwp2f5cFbm+xvgM8c77znDnPb+qti4nBEfXh4SKRizv7k/Xz
fE8OFNjBMvk++hgHQ1p25F2iWbF7ONkrPRMmNo4qpJG5hq0HCDNvlPFrKP7F5TJ1m91/RCQQbr6o
nkjEvlnpK6ay8Vbu+BeCOMBL4NB3FnvZ5Yb7YP70F6BvuWB+zqAh/hcrchqbuJKM9MvBRnFU45Ym
l6646YsrcwKVetqEqDccib3JmVLoYDNctJQZ+bJ3XSofzH1Ny4lIxXggLmNaOmVoDRMwmf7Wscdm
HaxpWjjHXGBH3lMd3kPt6bRFf1L4HI70OiSdn/fuhgFafnlB6kX5Iw1/fjx1b5PN+fPF4PxJ1p1p
9RDxjhM7FkRl3khDioH/fSaJzRviZlGgzbwFDXJstf0mtsitcOnFO6FbCsFB/LaiJmUVm6NL1iJF
+wYkcrYvca2WW1b0t/GuVTG3SAIatzd0QKj6P8Osubg7zYjnHxX3nmbz7NCTEVFzq+iXgwFZYXvJ
6frGx8Zo3TnOiuMgvnt7SiYXQHQGHrOHExk4Sn2yfeC3ATT3jGfqAuH/T2DkPgweqaiIc6+rt4k0
YsDQPD7g7ie4BsbQHrhhsQbONj8LcxUy6cDkG29U0ShMpZMJXdcDHIZTkAVeCs9hrjdzz7NB64xp
k8v6PpfI/xyIiRUhx6g4/CxQfwg7XxFS7Mg8FZZLPm9oWQY+jD5PULoZLA5x4lpbcnFzP+fzQG7N
F0lLv/kR2DBV8BctQ6HTvdkaUddqSFp6rQ5J5Q2zjIKSdrS4MeyRJ3fHIYE9lLg9f+aKnNwh09t0
8lfVYI3pDmmIH5cfhS3RupDQQ5kJquR2ctP8pRhIVTqtZSd7zb/LIzsBugrYCitR3km/LZ/BMCDY
oRavOH24UxSy91q9KnNV7q99yP2KujgGY2IX4bPpC9A5u9FmineTN0POSl2V20XCrYa6vZrph0r0
jSVQWS5YepmRmknd1yGZrAkSFzWXyKOCp7NMYr4ZiGZ28+kZzxxuxcBD4yddzxr2G2Aw7MtfGMJR
GCBKgUPu5sT3XaKMj7gfncXq98uqxavV2KFNWcRu16vbtXZXaneUlho4i4s7IlcZyniC7rCYmb/f
mMFoXt4jCuw2JH1NrTJjCzKMFmjk6B/s8OkIuEkcRmItDYcCGgKEm7pkvZmtlE6iIMDicI0LL6EE
O18BDH9pKdbrK6/yI3MBZ+fXFKGV3Iwe75N5bih9LIDWBKMbhOnT3u9XUk6ZdtUfnyrHXrKQpWCn
KnYEerIuUcJZwUTNTQ77NyQaWqhOK5wWP7QrgXnSdtiISGIFchpyDWnKTyazHHAjjs/ILalI0lG7
MhnAtHnokqUSKu5j/83ctBFbZMC+D2QcSlHytUnMb2YPKmeOq79yMLzt13h84xyo8wBxw+03+ztA
TkP2qbrsSjQGHc/vBuEI8yC5VxPa5vnzcNOXOYHyx9fj4+ysE+dZooZSsPs4IajODzAMTU7eyo2V
jSKKqLsz/VgUGMllS6NaeWgP6eQwej0BZM1VOxlhgiRJ303udD6YOogrUz6utpnF4wl96YnCgOst
ya1ph37q7atf7HwUU1aRurdiATJ0lTke7WFsdVQfCg+5gi8XQo71pzhTkPkBt9fJ1OgwcAIkOYuL
ywvlVLtrsZXJvVB5dIasvK1U5vHYxSVBoQBglFrA9VG+1pQoPVIogydK18AgSmm+/veQZ59F1y4z
7Ovwje14F8pHqgQsZaNv7rEOV23rYQCsX8LkzEeae51BGx+smJGc4iisonCc/341Ibr0JhVMnEA4
RMPtFmWZ4gMd3DfEeB5TYvG/GiFIGZsWFBlY0cxkKoXdOb2RhylGPELKWgFKmyeJuaGXAYVJNiHb
2yMPqPrMN5igSfATy0fqYcLDId2/MUXvw9fNXYHoaRgRRa7nRjmuEfcJbK641I+HQyziwtE5VvkE
LmL5kMlgoBZ5ROVdyiuTktxKLKQIalLLobfa1/5zyFFCkkzKdT/9bR8nPiTnPkGIgNZZM9BnbydA
4aD6xWlfVvjEbBysN5TvTRtQFL/BUJjA2RMaM0oHUN1mzbUSvKJ5h1IFG8h8bRwJbTd0ELgjflbN
uO8sOolaJ45HcPFH3rR5khrTvpUmYokDG/jR1gj5EPtMlNUaB4Qr+qzrd6O/OhSKufx1sk2cASiG
+eueQV0f+TojtvZ/+VRpde1YfzLNrOOhSPwLPKCH0iusyhsoZKwCtCtJ2u/4hXKpGOItEsjkmCBZ
E1RMi/HigOyuKR9cjf9S/BNDZDc4/EkDc97s+zGOfAgTFKmTXzzXaq38yBye7jGAfnl0yn4rZbYA
AkcURDnPDPbWEYLRX9OQdmABo2Uj2IHL5FUP6XPlE9KKOwHzLTiIIxT+Eh6lrVN2BUoj2IrpPO6u
pGVB67CLWaSpyZTNgV/L0h73ixPfQgkHRvpVW2EsYRuPS7R6j6TfOvfXzRZXermD/NDTROHzL3dx
MWzQjM9vtYCmB8kGfrI7OawRfN7eTLkPDo6bVUprHIH/POzt9XbXX3JUWfPapEF4KlJwe/3VoJ7o
fi2IWYItQFzYjZK6TO6SBRYg99FsR34EwkPG4rvR6CuLoD/oKdPgDXlzuSl+7eIGovWhOWxgvJ+a
5D4YkW36h0WJKeNE81Ed3SANXsmVeeDLe9Nz4IFTdM7L7fwN4FToZfC9h1jwEPl6amn1uMM0b6RU
K7Ugl++oLBJRQZ0SomNBEK7SaNYq0TS9vil513REge+QbmNddlHJyCo7K3tXVYgA1rpi8UFH0dCJ
4G26bysGoBy0HGarIf2H5fqyobutcguO5v0U2qJjN2l7n3sQ71p8Mq4yKaKaO2GleJz4FviDgzq3
UDA7ecfQKab4vFAU5JgqGm83fO2EfdOzz4ttuURVaEywqsboFw1Agkj530wD2L8AQKZ+MLFw4Gwl
esnIwkv89Mw/Rlzx6Yy3r59P6vFRy2NCgszTvYe7XjXwMC0PGh7FvFzfhp0gRVGc6FDkIef3jz8W
Nxc62Yjm+ErV1coBNn7jhKfNpPLAHick/e4UrkCGMufcaPsYP/FHNDMxRJegJAeVvRNRcj+YVn68
XKqn+YNTOyoQnLnBorDVAYaXR+yvYq86YRffSf3rbE80VuHxejKQkVw+9u4qiaQ8NVhIqM7SijAL
ylzLxXBSgjiWjR/OTwV4Hb4CJ95yoWyiIJklBA4EnbxestJdzRyYn91BZsZ9733eew3Bn0wCAwXp
HVPF627vDRFjeb8QwOqmdrWeOYET7MvsjNh6n2QfjSDqbhZpGiOD5PQumHHsIhG4f5oBVo9Yrpio
2vbDAG+YbP7WSteDMzu/V+ikc4pKi3SuihHu5dbNOieYiAQxeiTNROIYDot9gyFX+cXCURsENJjv
xmfqUM8JuLFphyS3VGO+0Irv7BaYWRNzVpJaGV+ySVEi1oUdodmiA4yVEjtsjawCAmg0YcKkkC/f
Npy39/vAuwArGWVVtwlrx8nZj2YWAeLc0tRtWwm6aXU+WPAY+lrMMDGV4ZR6GDIZVd0+G9PxQUnI
vGFKtU9LX/PQdnorgoJ31ev6O/NrGocMJNbVEdCnv6tYkXdqmxGx3raApgtR4CRJhCPXn2CzGaXR
hwP99nbVHOYu4AisPj81D0eb2UxMfxx4/9S97Vvp0d2q/62QEfSjP3Fk/5jVVKLwbZE+Db6OSPnv
WuTNo9tWWlMbTWZoyOyXLEdGXh6SzGqUjvqSxrnmy+ZyY7Bk7UA1nZ9GharO4gpnDKS0K/EjaiQw
TJvrvDeDafzxxDdqf6PKajJEiODaWsM9dWZmpmzHUoSe5FkZkyDv9/LFoSCr8GFtHuP3RzY2k4oo
Xqy8QKYkksiZHGpQLYIMFi6MlZfduJP1DrqKlwrf4Av87ize2csfZb1KwYtPmrdjl9d4wLDjrrlf
Uc9pph1P1SJLKxxrF1rCNNPcQtNPVm+aIQO4HByzJm3DHODBAuuDUrs95xzdVoVxJ19Gny4mFaIw
/+zyKpGJQPG+p+ghO2vrrTib7Py+hz93dxYOPLN1TdG3HwPnI7CW5C1819cKs1PVsmZJFIMjbvqG
ZuhqpSl4kfpx1NTQOqZNzjMiqMDq6FRGWcf/iMVDBroW2UotSU9GzMONXNeDW8WSZ5v8dQ9ZgVAa
ta4XN276udNeHTP3Q+jFcELRGN0OY/3U358AcBu6FQi8y5ac0Vfc9BtuHmBVFsh3Mg0Jz/++K2F8
HAP3nPWuAVHFMexOTdX/ET78TnrQlUAaKBqCCmyaX4zGtjVthyprxGl2hJ/UaeMUzcJPsxrwAhqd
ZixMK+cj0Wgwaf/b09Bld9flzmtsrE7d/DZQynfThRxH1ieWA8l53aI2BXRq/odkbj0+qxwr1xBF
YZo1HpxBuhMbqzfl7VmjFfIyWgqEnMn86KMHuvAxptUntdPfKFHlPS3uM64VCYWjnJUculMeVbj1
97QelCWKVzcmk6hTeOdFSQteGzYHVKGpBogEcNNsZ6cCxJLfqMWDZ0GZD3zKwS1mD4xIrCd5DE3l
3XCx9GG4D9NYu68/xhkr6YZCdvPssWfPYbkUvZaQMZyde1pJt4e8jTRt7J1TMVC2STeffbLUlQHF
0hjrikBov99zsteTzZoKJ624ipkEF2hrhMp4laf9+5jKwsyLzA7qQ44X4v7OiTV9UW79vtMcvdAX
F6e7r6NQOPcFXiLoJYblQnZbI4aPfoP6NXeZmS2jSGUFJEnPufI7d+XH3tR8XjX3vAPD+yXll94h
lKSDrCVhstNQD+52ajq2fLYnEUk+oG9u+gW+YfBMWh+iYM/EuvWng65ZRr/GIOwmtc8Rixkl0o6e
hMxHyovvQLQmEnTLiGHOYKzdbG8oLl2UmGXlPnJUMjqtIolJsP7vH5R0So3+fPxAu9xQ2lYnELgz
ijGPO9K7d1h1hhuMvenWGdqfkWFSYJlEj4QAJfFw5j6gM/7rZk9IXodKJJ+7FnLiV/UUZYweN/h7
a5OfCOXCBgDiP1k05F3wEAtdmhzIJSaqgCDAWPFAyKprwGyM/M5rcWs0Qul3ltMcNiqSd6d/vTZk
6chddH6Uq2ej2XI64T7uaV68OnOYZvI8e/P79AWL0G8Ki4xCtLN4AYFDYHwrSFKPRKG6dzc+Xiiy
n9AWbO+z2nEDr3PnTn2aDPbIjid9+FvGSqkHUlD3AEXaQBY6N1Fe5Fs8dkeU1daT2/y4v9qfoE/h
kQTsjWl2ffw063avK4/W8oDBV6lJ/2jybGRGdz3VsDJGtX9J3xTkwkbdx6PVayplE9K3pLNkcUip
mYneKT1id93gPUm7PUIoDSBP+hNgVuW1WVn0FGmqXDpfJ8Q5J0ZlEsix+xlWzl5rMY9o6XgziE7q
+XfGRKIqPzG57tQI71ji6l1YY9hMqY8OBKn15FBDvAuKjPZx3+fr22u2QkgGqD4ho1iJuR5Y8Cfu
GDOG/rgdCBqcILaIwDxykSkBEaeeOua5SwYyGJSxJzicGXsB56o3EixiI3Fc8qnlZKc2JKnPa3Cf
aKKagPfOP58J4Us1JkSyFjCI4MJJg7C8UGSVWvOZlTHls0JD5zsxpby1FOjtvu25zFJEuxNgWDgJ
y/+s2O+auCs7JbhNRmR9U0AnQIv+Obj2eCG6mZioAmeX2ek1VaN9O1nVzBYhvl+A8bVgcEJkkkhC
pwDPNesBCHSYS0Je86J2GGmFiXwFtgxkB+Jj1RWF7vdwX9E6jf6q14HZCNJvoa7JFfeV+WVgRZ9P
+K3SiPv17ccWRmJoBlZb6gVc5Kl/nZKDVj0zqjV/gPo6sm5h2QPVBrbW51TjUzExbtY4o/OrGxG5
FwKCczzENU451ANJYSXlKw5pfFzw260C4hLoLlsjI3cb+IuTjblXDHN0plilkxR8bRrx3o0fE0oL
SmAYq/P8W+4Tn0uo/qJXxkSuS28MTlYDl56LDQIINGeEuiKY9LDqau6fmIpiV2mtxTW5uwIeeggB
B1ips68OPZ/bGQmTPzk+h8+bjiatwz/2hXrMNQkMzLW5IO9x8H8ZYTzThIb6d6uqM4V8JnCzRqN2
oiTfekFL6Q27kZw+O/QFNJxtIgbvRkz1DGkudNI9Xowaw1jT7VD1rRAWjUENW5k9NwgmP3vIZDMy
tCDTj6fkGr7hFYw+89mhj9rDTPAFsJn7l4zBbIX+lMLf1YtDpD9oSLu8beKY2zua+PG8uHaVVuIJ
5r8xnCfUnC5Qma+NumWiQnHSKTvUmWgF/ipYP17sncBRUoV9/07Couxm30MRmTDDMVBIzD9L9XAJ
zqvaDh/+wd6nnXhS8kuH8+48MwtlZZkUempwQmGr7fRQsUnC0m4WjAT5NRVyBHXikHuBYGTv466+
2MIXiZMpMFlRTvQogKBmjCzQjURfbrB7Jpn3HlfmXmiTuxYMO5g+J/hGnE37IuX++suE5KfwAMzf
AItg1HeG7DQYxY9kaAhvYmV0jQczQVreknYScezbvKYdzPA0gGOPn9fy5ypO/gpMCN/olBD+bnGN
nSI1nuPJZo5kYj6thCB0NivYfptTevBxOBLkVOdkvOvEXSlTDp9Ah+BGcM6/Km0nLGE13beAHDS+
2zw+yWexUUlrBtHp6GWuSW356WnUU2BcHQJjV/2oA48/LcsXD7HQ3HmN5nFWKjQFTE5j8RmqWAMl
o3E9t8G4b3dbK1nZIQ2BR9aS7i3DDk5dGUXEzIoAGnmGqvS8KPU4it+Mln7Vqpeev9kTrioiN+vt
K8bdIQ7j/xGU/S16Xmq9efDUHzulKhqNYIFU0n/vwC7bgvXS5wPnQoFCmdouA8SLFS1aNR9VkKdd
rRLHtzQIeBuDjVZNjuhGMVhCYQKsqlf1hL4BmKsRUKbzF7LChSY2LNBHBbz4UjddGTtVX3jA8+NZ
83M7glpmhXf3h0QFMNMJUuhw6nLoHq8kTGgDV6a+nHpfuPwrUb7oAniFjkoyoBCa9ipSsZGQ+PrK
loqEoB+9mSPLlEZByOX+bJB6CjQ/zEqtmJKtw2nH8pAJX5EgR9mOGJ45nmI0YG/VvA7FYtPmwgUE
bg9ogMIdhsT5IPSCD9UUjEmQOOvcoaYkBWHirzfZ2UnSvgEPHfoW+PiAetFd27ux6daSlw5ZUsC/
ghBIONyfr4o8B1kPFQ7+8Z34WYyJqIaJQpVdwyweSALgRhZq8F9ZSGYmyZep2hluZazgyZHrFuqx
nIlCgxRUQYyrXSHauFKcH5usnRm+VCRX/tbLH+oFTRn7TVZlM7kDZWyca4TdxOkUKk+K004+Zw78
NnAwxkmkScTMRgutGT9T70nqlKQvDL8EfQeaVAv2ncTRHAfukPA8AzqRTRiXYMrMdMQ7MArD3cMW
cuZL5pH4eBtHOAoNUS1FW/BfbTcSmB03FpIJliq0zSR9wpwqh1xC+xnub3rvKCXUvZMkDaSi0EJq
CdiP40+7AMuchxOOijh3/TAkHzVpj9N3vMPKXnMwJbVi810p4q9etFLU8AKLRx0Q+tz+bCXFterd
irnPONONci0PVVpGdNTBMiiHysJDKPDZrdsHXszibYGwa3gFdRmGbMbZXKwJiIYm570lPqGR4hrr
5vYPKJYQGg9f0yMWqdUxNhQtAnwhCSXMfTW/zMWKotnhwDkkia2tuFBOrQr0lSOKh2927ofwL00r
entwm3s3KBOBVUyaIJqu+oR3sfECRAUZO1Uu836mAPxDZft4SrSKbPeyY/360vMQM/4Qeg7IE0DY
EFWu4Pk8jczCxSrSV5SO+0BRbGskxgavgGSrS+8+VQjx0gNNYesVpLaA0y40pvYpDG8NWFJwdK7q
DxWaLLI8KH5fGpl3tFZChUl/SdiP+ftItezBP7yRGStFyzsKDF4xcajSwe0wMImw8PrKur40Earq
BygqzGm2yo0I6/CGXNE9ANOjvU6TG3EVmOneeWitqTSP/VJJ22qc9DEK4P+CTQtEkiGQbjno3Jz3
SChZGGhZC4NBnqVh9XuWtsW4TFWmQ6U33X0hl86iD3ag6Ta58cV1zthfrj3lno/qHsTPT7N+c85+
7da9tXhkLivd1HKJajP0UOykW45gnHQP2CRfi9F2112JVM0kGDv4opxkuKvtKeaoaa3bpzuUueuw
M3jfCvrxaIlGiMR2vZBIOYVSW+O1/Qh+O1TnaXSgHltPlWjo+wsOj4mRUCYVs30bQ7EwE1ESZKOb
re2dQH2x2fRRFiMzcl8bq3XgqzhHcv1bSabi28um+FMBvHjrz64ZNgU0sIvL0Jqz5xfDobcS0fEB
kzGVRdpzXAjEZrWJXUx26uynu+l4mjPzuzDKx0T/rEyHqgIxbK6TJPVoPBrMU8Uure9VgsMFZHA+
BY2JIIl6G51c6j+tntBGBVDjnoOXHz9n2zr/7kVnO2gnolopdNxlMfh2pCjDe4umkem9LEK1CDIP
xLHKW8h5Zpw2PqRPPcgIO5C3HjsTnQK5Vizy59aO/4Q2SGGg/AZPMKChpVy6oHMiYumszmOJG0aA
8WIIDeOfHOnZR60HIuL/L1c6/nSsfcXX3FHXAlh7fiSDxp7wVz/J+xnRVmkkxJHIqlIfRj1Xt8el
VH7wJQ0ng3wQeD218uAsN1LY7O0m+xANiGugCtBmRUKbN6lTZlV1RqYUg1O+/rpxjzXu2UJp2g8X
iNZflUs0LBrka+6JucxpKxNUsSWrotraXGL5D3ddJ5veTQu6Axy01kFnsiBi5AOvSUssnMJ8aHVn
ayqagReYNchQglz/BOBvYOhg6Ubs1D6Hj5mpzs6r9wNFzQzcwg98SDZ7BEGLR4qhSZcr/qEPr68a
D0XoqUU44Z6YOFHIpE+vOwb7YyB2GYyJwzGSBvaop5WVjMC2Cl5gtVcVnjxt6R+Uu4yzn8jyNRZq
ugQnQakgZz0zIp3DNlbXq7LnfSgCbFePSYoULIXQP1dU1vihIxXoecnfv2N1In4OoBb4ZahXz8if
tpQu48vH2DOezk7rQLLsEq6dcqrQrK4Npr2yZkyA6IeZEfAkS7kkJXeo4MoQ8bzJsP/O3b/ldz4U
oxE89eeJa9j488i7VcsJYlgDqmLwJaivx9IHrfqrNLMFb5xmGwkr3r0DLkJ8QxHW5CMzBzV8UX21
kgmEpKjR9Lz9Q0E6G1ASmzky6YGHkyIlTkzOAynXclZhWOnQHK91SFZ07oOKc1IO3LAQ9NmqBqaR
J6snpSv8T2k1X9n09g0cHAGMKZTkkl29jNRmeCbSDELfN2HIYz9AFQJbtM5Ruf8DYTMYzvt36dw2
QyxNG7b8xdfcGPO6DGb9TMyk1QqFOsly6PmlE9iEE3pmzL1gJAIGYpkMFu10flPTxCXbhQ0Fv2kT
FGF/AY12jKjTRR1qQl1cIbQCIKLAgd/wr4KHluWYPu7IwdAYNwJ/QZRIExU0aj4DUdzppPvwuSYi
dIXYIg5W3atBkzqrpc+ryR0VY/qPx92WHpACTfV1uqPsgb8xMS2JGnHO+sesgcDo+CEe+QzOhz+L
S7kV2ZXwszBzSD9rw8eVG3Yo3S0jnfXni4/0C4yAMyDnWBGHNKg3sCIsvtd8xew5XDW352M6anhH
dCFz7CVDpIekwKuEwFRJFwljlcBaNuYOb3+u42IUpGwx4IbWgGu+UhJbIjMcwoHdVBzdsp8VMkml
BQHOoYi3H+GWgxRcxc+z0FOKneO8ZBsJ2GZntYxPvWgH0YroqRpzSYACdVuZuFiNViYj3nX7BzmH
bTnv5x4QqixK6xW0Is5+U76kJ/onS/1xmqkUCtN3hHrkmAglyHpJz0RBjiW+4LZGwhXgOQPp45ri
c7xwnL//QfQutnVpV7yXNwvdtkcA1RAAweWovmY481EKGIg6vpIj8qNmrZ0dqmFFnC74QlUq2WZo
3GhAYl6JeFPnslgNzp7+PgNaa6D39HPNfc8keLjQo9CNHQJkPoxgujlvMfpYf/z5dh1ZY+rLxiBr
JQKU6fANFVRGTeSZ5zyq3NY/A7RBkm/BakItcuXij2WF4tSFbYc5iJwrIgeTNuaEAqahOfBmuRkc
XpJQ5WL60bKzAZWW3wY9b54Yyxlc2zIFxxl6BldHPgNy1t09WjE+7QYnTCCIY6u/knGfx4WplgHk
rJY01nNrS+5HClYhHb9b+w9Aj5eOhIPWdahU2xxz091BOm6VHmTOhktcXFrJrcdtwTCmYvdhBAGq
WgztfwZbK8gYII7rdTO6JD4Auj+m8WVMqRteQZgwWKxvB+m1onYZOTIZedkAOTvaQ6fY0ttzVSEc
63Bn3oNyIPUES1afn+QBFfRCpuilR4CUx/0mTP84CVNkThK3+UMyY37AzxoT6TNzmHK87k4b87WC
t/g/jZ5iEcBIilsg23Jmd6rCIdFt7rGfAcHVirhD0Rmwb8i/lCE2SyBbAjZJ12j0SUS67mnGjaoF
3lhmc7XFVkV7tOizZhF18tYpemi46ICSZGUHNZySjjBtKzxbUk0kPYieZqfxhHgdfDkUKOXS4oNL
nuVSvvkagSGIV+jSOZy4v87+x7W80N4JEEXechG8VVnsVFDBQKBnxOpJosMdthvbiAo8ro5AiaYZ
GRfE9Ipa5sqTh1lc2nvxdLgOeYyCH7Y+Oh5alNGuRoLM7w2YqrVuPQwroeL/7tx7RyDPwAWoA0Dq
dvRDgScqrszubSww/c1gzquOuhRPaZdu9zkRvEOkRBZcaiASmGfVtAKECygkjI3So7pb+hdCaCIv
ODGU49aaWfAV2QU5wcSakDRBhi8M07WYHLOvYQgj+qXkhuAHRKUWJCrbfNgWelEuodPY2BhKVYZy
71ETtQacbNjXQLbtS7/rYPh6AV9r3nsl6KWu52mpM90xe7GD70G9bUUpwetgJSqfOVQOoWPrFvao
qTXQyOBbVH/hrUVKr24ZMteh3ygZhQ8A6IzB9/enYcJ0PN0VG1W1mkEgx7c9oKtxsWKxRIfp9ESj
vgmszcK1gUyCw0LIWpy4M6ulLWnkdXFFYaPM838B/3r0n7G3Lu7wktw5LYHONu2B3Vgop6VXqJZG
o9iz6byrAdAoxBA74y+MqnbUx0IBk6wUHhsKc6+DbkoQmI9VuWGBbGAKQP8hf/TF53qItnZ8f7JE
DYzG8bXZAk4pxNac20qym8qH7uxXW+abNTjp1ZdkeOIBi7t+8n/oXgthgCDVXp87phW3KLoYLPMU
uNN4AD7HLtBzl72LJsOnwNn/4trS1ZgI9q2ZX3gm76qOqkBi0wmaotZ/nudP3reuNAh0RkJIhQs0
bQNMffnIhyx4Sy33FCSD3ghXBczLk+YXVXbCyEhc2bvhUf4KmzzUJcyklV7cotVmHq8YPQhy/fD1
6wg/9HfncOL77QqeIdmtz1aRpA3S4sjPDksowMe9RGYR42ug+GdSlnf6CPEpsYXZiCyPivX7ibj0
Vwhv0CT4kaQfvcfu8SVfJMgm2h5rOg58TnDpU4WQ5H1EdWHPc6bMc6cItrt4L+rw+L2RwjJ68MbS
sPRq9tNe2sF/hV2v0dBDww2j87SQ2u2griYIlSOq1QvMlmco1MblxqriI9ceRbv+pwZAu3WIjEUm
lsm1YfNg3hFetgGnYA+HeFn0QPwaqyrzsOwny6izqmbyNNDh/TNCk3Vvtgnx5eAMjdq/OVVkiX8X
G39pENvLuckMIOtQNYviwt2+hq8skqqJquUkg+Fc6qf0Z65UGZzrZNoNXq5vnnCljqzrIPCJu7xb
bLirmcpRok3edyVN+PuAZZwo0w1ESFtnzrYqMn4K9Y1YX/MssnepG/RdrE1D4F/ibZKpBF3rAODt
I1p6OtPBKc5zCa7Z6ckG4/HCOy0/+8X0nMlIheXfAxk5FUTZiguQDIQvGOR/Vr2RR1XjJORZyKMI
58yhzQYSjlWnN/dVQqsqScvapQwanv3gHlABZd8tEt43I4TJ1oHZFXc/z6964lycIW65KZY5yDEi
PbU17MDStybOP4TIc/HPzSeZC2hegL5KoGDRR0l1zvw/8a8W4ZpIbp2NjRRutBUV5w6jo19M0rBE
wzrrlRxV8z670Z5cXv2zhRw9UnxIXy0r0iDHgwlsuS+6WDp+T+GklcGZmb97Lv1U0uUHyMn+nYdx
hYMkcxvcQLoGZcW6SQuNk4PL+TNnRgMN8MbHaDnoLfnqOFwFFE2NJiWy0J4duLQiC/m0okpag9kM
WImBjar2MRWTM6EYvvRD+c5Ds+YUnQkFMoz2z1zX1c6jMnug2lOPmkqAxoW1CV4WrTpeLim9H+Im
juKI3oqH9piGlf07jZbFbpySf2T2GdIbmEG86tbKTOBUSQt119H4YjlzlI0DkvN2lEAaKhzfHOJY
qVAnMHVyn9rBnMF5AEG0jpVBSEeW0idocFp5V7EF2eY/gTkVH7InHGLLx0sJRuiByDhIMvWpoc68
GC75K6soGGwVk28NLpSny/7r2AZj55mk0DdpvvSIss0XDH9KRB+4KbLE0mUEuHXsoWulTQubO902
cX0AG5rBNgsrnKgTuyDp8/uuNmbPQGB3CooorjoIBjggkUMlaa82aX3ZWXqCG9i4amdeuNWVkqRk
Fv/yCsU1rmete/fnkxruUGhRg98bRbaGx3fNHTjHyllAY4X83GNJCJBG9Ai7rFDwn/Biu3fj4Tdd
mxFiGnW4EpX6cOojw++5DYrthbBjLaFXJ9tI/sTyHPstF1DD+s5VMFeDyTHmtlmfXWEM1z9zGixp
NXq8vk/tD9ULGymJ9EMjk8bvPMp91/1ZDoAL6TEHwe4VET+Qn0OgDDN6dyHs2Awxcx+EPTuQ7zHt
zfua0D+3FrTolfWN6Mt6+THZm6L0DXFmLJ5Pb7LTo+5eQmh++9BkSdpCwd9AFa+5wdKgwX6PJCrj
aFp7IcSSGm4njGUiZD0nj8WDfc/AaadewB5hvwl9h1tH635cpw33JJCghmSAd34wv4IrVcRCLNCi
T21kDIx8KArnfrt+c5zcyui7l4KEJEBxQd/Eb5ZJSjH3iZwKE2hEsnGdsGuCTkVDa1pTdzhYgcpH
+TuOXPH16h39sMpLjfA+Ltf/XL+mgpycgZ0g5IfAg0X+djHi98wZ30RRwR5AKIv5tlh0cYfWaWeP
YahNheUHr/wytLbWZpIPSYfKY6q7vWpdyW+/NxhUh+5VYHW6ozJFmGdsm4/gCQMCsuPLrxnmOi7C
Nvzu4Fj6SXWxpa+7ELPh8wcnW+IJdbGr99BRxcHpWR0lTB/gb/vrN6GJQOuIcPtDJxZF093k9z2x
D7Nr6ieTarLVjoAOvSFt/RkX5oYQNvkrFHmncCqx3eR9hr4YXT6kpv8MBAV5eWqr1NbqNS4P8ZVb
xl4Z9lL+uDjVgqfpSoSz1qtHQeYBTNsiviqoD+b+AYpEql9c2P4hWOMsfgnheSe0dW1YeFearHTX
F9JtBwFOdGXlieQhe4bZV8rODDYgHUeVDRujNAmpcqKW1KmG7zNcrGC377zLgXtN5CTlFRvkmorE
O/fGd+YtMFgV6B0XhETeqXCXgjdVoUAQaCdOPAfm3kd5IvKbSvELuDiSgNPYq6gHmhI3O9XHF81p
LSijqOQDwssrgroxh4qBglgkIgqcNFJWgJeomkK2hcTXSEyRsqbwhZQyCKRaUdoVfNoolvhZUv4U
e5b2wTRMpyyvgml2YRsH6gudGBE8uwR1cUIuFEf5hoOFJF+JGqYgqrGkY52PwyhXNX2H6wDm0KLk
qI7RCxf5aNP8HGfLFrMNI9D7IwslijynW2EcNgVFxIt1GujFBm6gNfdzZajXLjHeodY13eiwpX+n
qE2LlYRA/MIW4RKlrsJO/NKbMS9gL4wveIRVmJP34FsAKnRg6yABP9lLObzQnwbWNrVFlv5gIG1g
ObtIW7amp/EuhA6roFDVSQNcIAwObylV6vjMFQ+qqQOO6NDIzjEiEDyYcotSIyc5QBVDtXE+HmiO
K5wU6CmiY+RhdVqfDv4isQpYU9/VHCrr9apLO17dn3RU7Pl+6u/Y7LPuMWPsxxU6pfFyRTk8qNNR
ugz66bG8pvrkEcn5c7S7YBNu5znhu8rxtkOxZGWbCSzz5Mi3nV3dBsLIDxJOSmCI397TxNKDV2oc
au8MNMZh77ahUHHLGFxkOF4lKxKaSyvIyUbJ0Y3DZYK9lMMA+O6OZK8APCaRrDxZ1MIDRdmDuSpf
bAckGtedSuNX84CLyiPjUR3inbW3lUZd1Ur0DmofB4ZSwjqB0fro4AoFTTqvLL7z1p4Vu7IhviTi
Rv2wdC9h+0Retc/J5NLS/54Rz96MVUmkrxQKgvvsSHx2UsrZrOFP0ntQ0rElCmc9xFSpV057kxvK
Mt+cDFp6hbZHHKD8wfGimUkK+AMmWAihytzweesz7hslj4xY08uhOlKjflSSt0e/wF1jyHxWHTbX
stlCFeXH12eOd60YNzqIrslYWt/JjUgCpCqWDeTxJgjXFCJlKm5YCJ91ZB/2CEJ86bxcOLOpRjsA
xLUNtdz2J09XtVEaSPG/gvx6Ouq82JXuK9ReVANyLEg1UjM5EVaqYQmVSaIrKtvg5DbrM843ySrH
40JtCDJjowy6iTBA8XDIZnXMf6/HsvWkIYT7qYg9PN/MV7jdnMh8Djq2TB7kDk6rKsH5kuiMbv9n
zPvOrtpctftLUH/+rfxYfl4zLaoq7KgOUQQ5weIQifyb9/GgaxMNgOSy2oAZ1ysjbopDp4/1u8U1
ZUK7uibmnGT1QU0giBdpxYCUDbJZXhmuVR8V+uitgvlCagSbQFzxbiUG31z7l1zi33P0wJko5F9E
7MlOba+DLX89r3cRrBrG0aMAVBKAWIWJwmSuCd5r0N1v8A9Y21mWz53Mx7R6HgXA1Lbcaj7eu493
a67ZFMndMPVR8pgy6lMjTzzCYpVBnafqaYD24J0ZCOg08SH164OIGWf78G1p2m6w8QR/uXDF1EFE
kqKdIMnD9j7YA+YILWiz/J2w94gQ2vLOHoOL+lNl9JAoLfX1cLuFvfU7j7dGus1Li5baJuUHyzRw
6EGTQkN4Ovr7f3N9ZZ6OSgkCrsMHLiQKy0ReWlw0uKyotFk/nqZgfY75B2H/KJXpDMJA6eC2X7ak
EYGWRYIqNejZhLVh1gic3EaSr6nhiwN5AJCvg4xY6rg1O7bvUgsLkncKYpRGqFgPMgM12WhW9wtw
4jTRn2nzOCUL/Tw3Sv/7p0eRfv9BENI8vA0wAbljiirYhCAgXAo4OcMPsxRd8T8jAnc9xBtve/vd
rtsE1Kb8rbY7n5xg+S+9zhBIfcHo47gomCyhhgMME8eVS/cr5jVSUoMzE6Idg8W7OAvmvC5taZcM
VZLcJWcXvEiDV8jqV1gOxcVewkfPuhUDXhyDPlbflIk6xMbTb+bKbbDtJhTny5luaYrCPZ7DyXof
ml+M7U9G7em1XOp0CrHrOACNObjD+QUFxZ/6HlMVDoAM611/wKK6u8EPF/KIVHZpDbmHaAn0i3zn
q5lOlDW6gtHyX6ut0dgf3PtAexT4SNjgkNLFIacDNUP8dupPp0QkZ7jFDrXZaYU8YDnwwZtwbEQM
9siN4FuzfnJ7J8ULY8tQIchPIgUPMCULms5hAALRIBq7SGht/uNzwaCBGOyHezXPqnjxLHw3xX+9
ayGJo+Mg2Wkot/On2m1uaXWB6ZIppCsWMv9Y7anvwoerKBIQ550fnICNwSHRGOJPnlU1KTzz0ne1
XcS+HjKcd/BJy9RL9v20zJ/97fAiw0xmDoQGQr8Ztf/OyFCIdSgskSG740BfZ0OTdZp7r9wgUwdD
mhE4qaRh9NsY+UpVXnMarv0GYKqkCpr4h7QWE8RA2zJFUB6HpAu67bu4octm/9nI/SkFC/YxiQT/
1ho569lXSSuiGmj9Jyt/Hwb3xitZ8ypq2TCXe6hihtzrHhzdM+cZelsl97LXMA+emc3zbEWPs7aJ
KHu+oL1aHxj2TxN920O/eaHMU+swY2Z/fTFbXMN7CtE+bFZOaCU/PlVQPTQQChniyOVSM8ebZLDz
08jF5yy9QS1Qs5umK02PJgbmpk5ffMOqb8NlyCm4mti+daIaapuiFdqQvn7+KyJSH1fkwkHojlMJ
wd696DZdC5Ig8bdzmEGwryIwI0//k/fEN+gZH+1P/0S015wAKUyrukhY3GsGUAPIbBlTKc6pVv3a
YNYH+fpZ/0RplO7xC/kKkYtHp0R8AzyTS5ALjXaGFVbdKOREZUXOYiX7u29XMeTb7smSKT7WIJPe
qEQWlrSan9FD7PMhyD7KGrES4E+EnFHMSgj5yfIE7Rs7qmOu87PgMgyV89YC8G+H/PVhbcx9KDlA
6K0FXRqCDh+yp7OY+N2Iz7jRinV2DtNwcH44v1+WnFhgjfN3jvb/epaFm+TJed+oW4sBF8IVU7qm
+AxWhOKTmbQJhIBvY+pgdN1OWuFMG4N1t/ZSXcs/k3c4fqhp680bi3TvyCBIInjRqSKu2QQLwlTK
GZncbyAMsWdh8sDvYDnvvgYCgGy0LmRHVY0LsrrE8TXNoEjli6YbJiKNnKt6qe6wd+9Bktd4IabL
MtC+VGAkQwF3fHMdNShI+L8AHd6ynNwd97Vx+i2J6Fr69kXFyxr/nAsoN9zqf7qpLgm3cNQJRg80
ytXWLe8HR1dD4UhDFl5o8MKwpRvN7WF7Z12mAtLoJHXEKuu1gNprhNQmSJ4nGFDOQ++2eHJFH8OU
pP6J4Mw0hfgBAGuMUIhgwXK2kbN6Zggi+ulQQkqchY67BLj6UC9S4Ri857mm8v9qanaIh2W7km/l
cxhCN7Ql48+hZJ2Cyz6/mWRoeVNAenSLPKnIBsGAUxopr4PnPhqq57zGBDM+adKvJx8Fkh1LePGV
AqJcirQXDAIdE7boyDLLmX06ITo28S44BDo1esO/0AI1MsYbt/lZSUfjbXpC2HTfjnetaNgkFwcm
wUYxANj931o+5oJPmmXoVvClmEa4B+sCyCChoDnwVu0YFFmmDH9WD6iYhiKpNCMNoXXvjFs1+4lH
H7OkK2B8qIdebayMBl8IAhXW9FikXiF3aPm7GAmjig4UJ/El/2qOCR9Lx4YCF9bxOE2aUODWpgUW
1KPR1LSZ7jfaVkr0secSiNtigP0MbbJkwwSWZMoRRo62uKWoqVCvDMnQqVO+cRXvntyo6MaWI8vq
tJ2YuNAG4ZG/WnsazUyMtOILA/rk1ncgww3Z61injV+06kqL+GAUcz4TzlXP2RSLP2x1F8sDG9Q0
OAyqqpKycBWkG6qnISByEjxw0OJq7EtQ+4mgh77n+Y0rbV+ZS+fD0n51mz5BgJO2IjkGmiDA+Aqf
kw+UWIBDTTW74/fVIiFiuk+tbLeomBai1RgUjfMZjlwTb1XpLVf9ajRRPGtYNWif4OaZP4S1J0ux
VlBRQiByPQBPn7jBFEPcStZInb6iNmYvnBhmqASnokaDivdy/0NZmzGvSD7P9vFW/wxTxnT5Ct2P
vLmrt3fhcWvo9yLOQkSRBNhC+pez7WIpkEpEUxyFTz1eCEGMtOwE3Qjzupdequz9FbwfqkYxbkOZ
gMRovx9vGVybiCYKtWsKAmhjWj+IVKQyQ60fBBCMTyYryHDasqO9cKPc7FLAtu9bHRL7IVUTsXis
NSfjHgOnaM27/0MouL5GTwQ7Q775jZA0MNUc4EqWNxPsGSV28B1dIhpQT4NzjwWpx+UNBEjjbSju
P3Yg5r6EM9FEGQplkoMVLaIrFhOaViba/WMuhqMozwR7OXiVYAN0eriBhv+qtWC8lAMMCkgpPeKq
Ms4+UmXQInEdvAUIo6Ely4K/JXRAz8+hbMl9nJqYIr9YvQXHvTpBK232liqHK9CpROE2gqxktxAY
rYQk3xZO4Ap0jpDv+ctq2yeEfe4JFX8fnRpIB+sJfiNa5C2WTa8xDvSD/JQYMPvGtapXF1MBaUSX
qnU0KaFNFt0heCaFlzbXoYPLUSJ6NpY+AVd425tB22bHPjo5bYGhBhXRkLUBEwJcnKKdGg5fyAnC
3uXSMDp29+lcSVCaZjFt1Ua3ScRnttzKghtYxqYiL/Ux6qf+5jEl6LDM2C7awSrwISn+k/VOtsm3
bgb/1uSTDfV5BRfTNCUrgLvEMIjrGNzi7cgaPrTd/YlGLj877ahXXVHt0DU+O4yoFZk9/UryzZyS
GdJFsZB4/hR1kTXKwpwVTlOpNyhZV38FXLqxYRH5uVMq1Jqi6+7gpPpELQfm2dknV53LouH3mSlq
HlOZQA0Ulbk76RrffdItw5uCv3a0pZFQeoj5NJAmLSj9sWpJHq3dp1tsBnEMpYWXNPykkvxOAO4l
R+xs4zxBanGh02aJtiQL1GZj5gkDgckqpXzDmfhtkUhu34aAu7yP2zlGGn9yU2Jr1/8o5zrrMSGQ
09q2eQkj04ge8T5X0SSCIZAYYs+2gU+JCOhyu/K9/6na4KcjhYF5mNVmbxAuZjvs0KR4q8f7T65d
NjoV4fzcHaapPF8TAvLNZ0BeU8PETDqdpOXvSvV0xe9GZVzcB6h+b6OGgHIytaFlWQeAVz/3bouR
U9MsgBRm2HMSKda9JZxccPwWv2jqjFU4kGaR5w4hOoI6p1h3X5UOEeZffAfLaAZeZ7wCRFMSrJwD
XQJBemWw6TKQto5f/uk/YS7x/n/M5K4Uay9ZR2fYcGIXaGmc6cRLJhQ7P8HK1mZ0pA79pUKpvZWF
5H+F3gZy6njB5HZN8aMF6CRI8AGBFRi7HY13iYTjOQE90DTu4fQDoaZNnrW7tWsIA+twDIswLH2w
hEU/E4X65lMCatAdlFM2NrhSgiPZnoircYAP3gHEoDwIodRBCwaSoY4mXNPSu49B17267dV8lU6p
ziNxytf8ydpfA2pe5s60qgmAl1qpOiAVe/Feyobhniz4VPNOt1wHx0G5IAWDLPCEgktLzHBOvDxH
UEZSCDkN84v543XzzBhgiLa6COok2nZ3YxoTede99GUwJudGuneCUmgb9dEpjac/S/rdJqr+PRSt
99dC9yPgfG9amxRm3r9BNli8VuMblS+7KBC43ONqQbldamPZ/0Nxjrfnv0KXwxJ8TXF/R3goa7l+
a6YZRn7J+dJkN0mYH4tHctZ+vgrroxnINvmgKpoVqvf97RknLqoKvKqbVfN5H2kPghze/mzPkgdr
uLmWW3POKJ1guLlKHbdQSaZNbhO9TiDq+//kmmAuZA1Vy/T0sETIdCy8FSVnKZu8BjwLtbUqF66w
0a2IZZQAckFuwGhyj/i/8I/WhuD/wBPoMMP9+ko9u+RZGimj39y7/4KXdKDjeW/kfe6O5FWsjq51
DTnsupMxeSoFQd66XAnkj1uShQeXZ4Wuj/EHXhMCZgMoBgOp5rvDV7472u/yGkzLKF9hl7OjvqMF
nciE5+yaiPHQzR5VAXy5qcOo6ajF01sXlBLZwpih6HMM9mqiWKNiEYZurdl0tLdU7K4qpn9nh3bq
x9pGJeUrNdakdPn9Sl/DCYMYSrOemqWhR9TzWiOF1/5CLTnQ1NjCXV6rxY4v3LVAwPr3Yc3bIjBu
zqldPxabS+QVsht7lHT2j1T1jamowbC3myY6KhIEyReR0WEkFTPZoZPS0ChubI0zxMLYr+vm4822
78TVJFVKBZpoJYGoJdNd4iKluZoUECyl5YlKrrg8RRCAVXrCzTVCCElItjXxj7bNCqHaTSvkACKp
KSjSXGiK0lxH0gCO6QWibOUGwTiGDdVjc9tXL0ZS1MqD9Htm06nk6JnebIZ2k0BukXLUN9i1wCOP
LgX4ytr3KMOMe3c11laVMAS2FyR3zJ013Wa8KaSScVtjnvnAzuBIryvpK3fzUy5plZZNMrUF4TWe
KWD0VFskYny/+IFbObM5ESb9Bo95TZrpxlHfaSB4DYCIVPZra1WNd4FHzWq+MISiVmM1gQEHhg+t
Y8VJb7jNZ3BalRodL70AgbSTEtIIcmF/HASyDriTImaSaHsd/wXRglZtJiFPRO7Hx2BNcivxD5Js
LQm8WOeYUeGudR6824WQ+9Q12e0Xin8OCP/iB1iN7d1gdr3tPXc07H02QAiYUcZajdLFJaTRKV2G
+C4EkePMDgrvlQD7ze5x+0pCA4q3ZJlKEOsWVf5PFsP8Svxi7mlcnkfFpRhO3zV++VuHX9w72CJE
IoQKBJpxz3RK0kXLS8TzQOJdjBRwIEuUVoRB0wCzLk1zsSJ64UzTyZnM8wKrex/XZQaU4IyqweDx
eEPKi9jPRk5Ggnbw4jnSPQu0ETyK9RadbLlHaHoYiMtcuHSHcXqJj4n1/SbVxUtAyVT81o5fymcu
y03JO8HDYtlngD+pScgC8xvAa7cQRqsNqjUeD7bTJn1oTb8B9nSmazPwyz4zfYvmcCgJF0pr7+wv
2BHgfFbp22EevgSUPSE520Zc8RdI4YtigQxu/oRvEDzz4oZ/eldMqiHQGcDGtzCGaK+ZHG6yHtee
lz/4oaMot7VwBCRStDFoyD8LKZ9OyknG2PlVtYVfWNRwcbMTZC63UQ7c5D7e/oJ+TUAdlISRQBMy
oLCuU0YPeCol+6k+1/rOa6WiyS9/nWCUiIRImAptGFKngUPzGUPXuaB2oQlyJXAXxxLnbk4Jy7zZ
ft6X7sBwRawyqIgg+GKaXEYvavUXie6OsdjyxPd/7PJYM9C9XY5TAMASQsGvcdw7zPuJwk74a3q4
on5DecPkPh2UsFKLjiLpxRLr4w9kau2fQtM7F72bUJazsLVDs1QU/S1wHIR6fQ55WCjVcIcAJA/X
n/7gezvQihFplDvbRjOwe4jD0rPTB4lrOHNkEt3J0kQ2XaWO2XikCHbQv8sBt1keZJLc2T7D//v4
38zNvTc9AcQh/LdOl69FjFDTrwYa7F5MUAhU+zSev7J778uzBq3FqRfTN/VZh2C9WwziXUnqPj4W
2CHWZKHTfKlC6nyxcjl7a8g7jXnUt9lr7Xj3Mw8BW90Jl6/Qif2RNrar9Ei24YjCLE7lCc1upgpR
Tc5ScCGFNq85D4MEQJUrrWEWlkF5+MoitfBjrFAaSJMiRksvwAd6u/1n6UkIWbj3F0bDu4mxQKeW
8i4amGyWjltf6nEdT16/sXXECN3q2FeThPSQuDOBjuVU3lJubvrleOKeRm392Sw1gxl7qdHeiq0Z
Z6cdaHf0SORr/eFYlOl2J+B3sf76OYz6aOMtcir/7Nit798D1PAHye3kGhUs9Y47kaAIjlPoDG+G
Ilp04teJPi/xNcplg90L3Jd3FdbbLocgo5iOKidnXSkqT0SuYmr2z7PowV5+VAxb8MjgyOi0PH4t
pcDu1U0UzJlh5g9GVitIVGfuFaU3zG/wnK1IaCeXBnuGxNDCqkmKN3tmGBqpRn3qRprZY5DxGchg
OdTSg6o5z2alQ48x+T2hkF7DoLI9N9mOhbfgFR8m7kzwSj07llH2o9DTLHMhp/rHIXvOH2Z49IFr
8vQ7UZhey+Gf7l8ehAGO7HvuFJkjvo10fSQ3I/XshRODL3mldsS4qKpqgEZSEoKOCgjVSQo8Ospn
/DcQIxf6N0HvCNqaukJYa5DxdCDO5wSV5Wf7PUk8PTiSqby3M+1xmrsg6gwofKjLCGHYm1a4iMwo
cpu49rbnmRkohtI5ruB32F63/iIScWYHkWYZI5KzgUsp9YZJvZajqsKsVTKfCDsRDdljuitf0UX3
Zd8O9MANwBAUNwDTa/NQIFcelJQjMwz0WaKk26otytG+0UhYB3UHp+mlvSR3Z5lnU5p1DAKxlawc
i5J+NDXctSk2IBvC54a7JpkXffjTxnOg9bdI6w2du14vv/rc8eExT59aLcMIe1Zqu/9HHZFc+ajH
4Mlx5zLZDnbSVFsWsBxsrl+9M/AeDCsNcYP+/ZOypiWp7P3qFdT4/fwRejo790y64rLGJxLdIFZG
SJGAFehNopC++NSATtjATp362OT3t8FZdWyFk5amDkKsSDBJnvXVYM1msXW5KHaPjA41aSXpAd2X
v4fbSYeI33R5kY+DmlcnInJSgLvUSPGPo5WxZqXN5GdNl/9NejDK8yoSIoGyC9pG5OqjVTmt5UbX
2YM7xzMXPrX0aa1xPmUW0IJNS8l3EtCTgU9oHFt92oHXp00+ITowHu1V6thHUJRZwgfIx/dVzzh/
rs3iBnUpJnL+VFnTr3kJSPfbmJoD6dlqow2JSFDRgc+YdjVb5RZNf1pw3kW3gwkbMJtVnQPgGtti
/Oi208aT3UDTgHZJbzAS2xMpqSxd46eWZqG8bVES+N8vxLHSt0sYyU6NURcPPRit/NbqRmQIC/FV
6DVW1TaEOvuGCcIeVBOmBQz6Zw8Wpnnwb8xQKAvZD2YMAWxp/iZ2VxnCd5U+wGYO0+KVaV6Kxb6k
TJthY7NPND/qt/8+dqgM7Xwj1Vd1TkNVR9Yg8vFUh6HT5ve29m+0Qhzu6TEF2QGhEzvQp2yyeN0e
7Xnsp159/mRh1Sw9dyL3Gk/IZ8pk9Jn5NKv0wF4kkdl9gzJm6VqPek9lYxi/sBgYUbp8Ahi0i7pl
ZUJ8JY0AUPhYMldfe3kJ5gAvH02LI+9eWVaBzH7xgZw3uwQAenk27UUYuzpcDvYcmnOi2p9YWSbN
8YC3xp4P8Q2MyGPlAnzO6+tZT+tLtVM5779IfeURD/yz4jBEfUuMBultP1a/p3dycMzFI1huxxuw
ecdbjn4GtcmyMQAv8PSdFG7iQaQ9GzDJqKgu9+c7ZSgL3lYSO8RqANcaaQuy6Es1gUVLuLVlGZgJ
f8rhmxblBJ9UmEeVkA7BCaQEcSlCWrSqyUDTJX5IHDQfSE8evCerN9IQUdft2skCS+vZwRtldsXk
UyG4X7G2CrMDPSmLfFSE4RIhs1UU6RS9qNSjVmZS24OqaUebjQyrZCTYNe6THvVIdcNI7EOU1oaY
NaQY9lIIehJmt/udGw/Y1xTj0YvziGCB8G2BKr/OCNjWaFP6LMG68P2UEZjuhGc62D1aFITQcjLv
m5+jOOeuycrNV4qGZ9GBpw3NY7gIimqtanQ6hF+nBFCr3QnqzqMsTJUMzLqukCrbz6omZe2ybvrB
dd6aArqLWjYNELJDE8XqLaBFzjXUcrxEmNhImRUxuofpHKv3iCxUAalWdY71aAm2HpcTyNFvte9i
+Z7Xn475kgJrzIOlSHZXC87HH8LvwrGhSZCv3qUKS+JmTt9OHb+ECHFsy0zxcTL+eHnF3PPyg49k
F2Kl2oKYf11Fe1L/g7hjF4keoWDK5rL/u2WRkRAX5DeXK6clmmVrQwExeGtirXgT+E5qzVIcDEjz
HMTxnnu49A1zb0NERYXRiqKbZucIYklC34sg3RZVzp31af5+yGxuyGgElUy3snZndSvbPYpO8ED6
mc64dyehW3imQjzbYEpaq9JC4AMB+Ec5loQqclnEsdpI7mbutfOpuyxp3ny0BqY8gpKpbsWnQKlE
pWwORvoUzZO7p5+xTmzyf9bs3YrfZEMGGK1SN0NeybSBBbhD9sGUttfyXWoNm9/s/3OrIKp4OFdO
UACMwnBFI/Q6E7KiIL4Rr9BcXZU4txF+1EVip7kSfP+YHulUSeRia2Qsq0A9okoEPfcuXb2Ebbdd
A9mJjHQ32Yk2soWao0u7KdTcpIY2rjSxQn4daX1XkE78ZaLHngmTy/T+B1RaiETvQY7X9zzZ/jLb
UkFmd/TFgc4e0OhgY0P5S427If2YrqxjTJAJiQVWxQZs3VQiwgjFRlITg9sE9ItnGR59sw+xIA7I
YCvCftSIT5gddP2K/eB35NhyYFA8GH94fjYaf9mx4GytkyxuD1omr4Mm1Xzktb/ufqFQgEIbNWVa
V8Yz9errHS+ZktzuNElKcD0ffibD/zVGwmv3QFFtWaqykg/mkP/IN8PbupoAihg32t5EAFBUpdhA
q6++lyVtOdE2SZN3ouU2iJgcC/Xex8MSHvDJ070oq1JaeyZxiUknFvKnEF7W8u6SqxaddxAl7htC
7Prsr4jpzGE4JsJwdmzPzGvLIMTMeGDIYNwURi9dyjB3/k5oosgzkcDxHcWpRxfznqwN1MSUyirc
J/75pUT0CYASjQaXHgtXEBvreGrW0Hl0mIdSzmeNOrnF7YaZCql0IrKVj0liHDz1gbV0EjRA/A0Y
XPRqTXutfN21dG5w8nH6+HtL62rvI6Z9FYDM/ih702T5SAb7ZeM2saVNyhWqs5lb2Z6fQwsGuGk+
u58Jt11Ur2rZpGqeHcUt9lOOsSItyiNh80dgfoh+LAqgxeU5psilBUr/WPgWWThCCa5jhYQmF9j6
aEbPcNh7xSqQNWeYaNKWOtjdRBFQm67PyZjjLmkPTKis8GAIBG4ASeM+su2CdFEGKRJe9pJ6EJJD
5Y8tg+4hjubbvf79q2N+QVezNdfou+22YoaXOlRXpIefgIoY+WbB8ybSQH0S3UqbM8hT8eZVV+SC
U3UwbekE6Y2mJt7kWIRlTAom1EeWGxa0YknE000RcvCMvXdyM/5U4h3ySSfBfK1kn78SprOz8WgS
eZ/DVDT6aRh4/xl63nQI3wfE3+f6nvsX6PIairIpxcDfRg7zTomoCsJ9tu2GHa2BbHwJMDHKbEFs
GPLtghr4ChV6RnWmRAhUv9ZFvq4NOzUsa0/4HqTbjiCfEjJRPiglDP6Gai/q70H6ZnriwoWwnFZU
elQo3lug5vwSq+SdvSUiqrdmTi5VeC3C2bW1C0yoqQJKbJWMob9pjEgtp1FHN3oyRO/8V0jbA5PK
n9M6Xob0Wgu2OifKC9u5mB8nVKgUT8mLJK10aLlVDS883jWegT+56wqfkmKDXOzb+olWSKucdMA+
WPw7YCUeZcwzZPdxpalVXR2wB1v+2nElDpAVhH6LuX6m5TVk7Sg5hpvldJ5AqqEvpzv9H7SJ4qQa
EDPof3kD2gMgzGFW94PiySDMV9FUff5Zd4ym1R2jLst1WH2JGl58ePWCVolFS3UOlfTXfSOfoNB3
kjFW+zh3nl8PMr5nTQJoQiXK0IKS52XmSq849luCPZOx323+nVVV5fEnKMTD9cfycS+2zRmW2EQG
tIOEh/GG3NIg75Q8beoLVRO4LssiuzRaKE15szD0+qN8/6tOaJu2eUNua6/xcr02gHQ2Qqwlpza0
MBVX2kqtwWLTe6u+CZ+ElfLtX9TNiN2DLqbfLM6KhZp0CX2/MsqLHs17wZ36l/i+HTVJq93nVXY0
g1h/1BJ/e9945TBDeNHpEiUwCMRbROAL4Cb3P7i1NJ0FWysI7gN288t/DVk/xu2S+iYct4zszBqx
gv7hqQe4pAXFH4GlYafkfoDJp+f2qAfW3xv6fMcF8qbpxlYZrbrxiaFwoYeqVQGUk9ZGoXCDlQ7C
UySPaqYs9i7ygMYJ7CsWdyVBEhLbLJohx1SAeFra9O0NX149WkmYuEqRtoV/sV9VSePPjM8oTlpS
NIpB7UCrwzTkCeFk3Ut0JHHPb2KlMO2WaWaV+l/CNGRN2E1E7zVW4anA5Xtg1WaBlpCv3CCsLtRp
NxsIoa6V7/UDGWYMs2RSCEJ/7lTBDSPRpz2alXp6DaslnnBSQtnQL2SQXdX7dvpf8i2g3GPMAv/p
tcugYHg781cI3kN09vXGxyiD6JDujtLa/3Z42dt/n8W0scJwGefwyZ1g19FG0wE2GVZbBSxSmnDR
7PBJbwrklIVj9kMn2Dqkl3wLEwudIdKCtO98ZBl/a0eywEwcrp4z+uyWc3J4wgsqEZGEPey2mhv5
6tPPy8z0YHG9oYLh7uVPolmJ3DXco/TK+BPtKjpfbLr2Jcrna1YIMtPOWQ+nbKcr4Nz74fBA3jSm
gvBtbCwHBx6IgxOBR1xD4bzyyNtwyoLBuwgBhqjdd6UrK2Ymb8LSRnvdMmllrzSMor1tTWKZSN6n
tUtlft+9s3Lg1vyXeQDN/91b4YcIA5cmV0E0IWRhtazVEvlduPxIJlt6NIdmcRO1dVAG9iZtngdR
1dlvFLb/CuRh3ZJ8WlRX/mqhxJfxAEkmDSK2InoryqzD3qxgf6kn997WxYA31srASaTLZcPC/6+E
NgHFuKOx3dMXTvsEPcawYBFEL2UanL5Lj0mdd/Ed+Ml3/NDQz2MM8wmMwl8nWNxWAWXZcMO3lUIP
pgmLO/6Ip0meapt8QvDvB6AFkyAtO/EdTtwpwDt+L+FMWT9pHSqGDw7ikpEd4soJevpm6ioU0BsC
lg4G2B9rgEwLrJ8Rsd79wbMG+D9ro2Ywyi02eSUCDiE8QY5y1EmxHoWzHwwiQzFbPZDcuYCQ4jLh
Gfl2AvqiwIg6QGsK4GNWdtJveFdQWmoVLIi1Jt4vEXQaJAFqch5bjSkzI/CtLAk1hVER/9SA1J0j
9eEsSgbOYDO08KoE1YDedoFxNUw7PQaikv/b9FnT0uZ/uvpUI/+gbLsY2QLR4LJnb2/gMjsYxNo2
anZsA5+XCbC9IVsdNCtE3RMKGFiLtjD9rYqPWt9y2Vs4UF8XPDgb2d9N4b3Plo3dUblzsNTUS7zp
enKV73iqUpLFpvXM9jbbLQ6e4rkOp2WoU4edVIpmOfIse4WK8TTdVog9V1loNvmWlr22QuuYmt3a
VS/BQUCvmg1XFVmShvt86wuHBnRATdeWk/sMulhZXjPTdbODMuTEIQH+UdLKcRvgwfXnJ43k3l16
m7/lO27HrGVqbkzbelPrNL1e8j+cNzHY0KknHb3cm5tnWTomqvIhbaDGc7SfSPhBpZ4hL2Cu4yAU
EzYd5bLNOV5sc4JazvzhzD58NSxni1MIDGv5YsB9h6eDOz3f+jkCOPXsVWj1TjwsJIuNihrPM/BZ
c2p2jukaSmsbiXLsX7u2i7W2grIaqgC+DCO6Ix2SbWyt0xOzBhqosmq+rmEtj7ovToFecbNTAlYV
rCzerfhGfKJJ8Rnn4YWi1gk8qZyHlzOto7NsZwzXMeGLIZdaKxcjbeAACx/pVEbt8jqe8EwEfD30
FmyfAXhyw6KSUn0VaZQTIIbnHuTS2mndmKeVlLkkwskOiZtKhl6x5vdXILlqgMe6Cu1LALJZyAiQ
u1EBjsG/2uPR3EcRNZut+91dPFmRPH6kjPw7OjAixqiTI1UCNQ7wxLlHnyp08K3z7WDbQKS+18x8
qiPBJLtLQRSO8+KGhuBmUWhz/Evyijy9kllOJtvM2U+Ck55nEAhvXdW9UqAY8o+aDjF3DYG8369F
+XzkHtKKDEVI5JgdIxvyrTbEWVVCam3Uw4i0BwTr1NckY8o1i4hx0qzZt6PrmaxxnPkPUwEyNoUv
AIkuyY6d23jTCBub9sYg6JhEegpqTBILUq//1F50AF/5DH7u4boLFDnopML2SN3Hl4gvj/bNQjor
2/fTS0w6ODYsvmubcsokDMAelykeDXuGEnrljYHj37DViK5noBXjghI//E5U0NKu0qPfuqCJqBgm
nqXkIdj8ps42v7NhFAgwwI/gnBsat7PP+zmPHT9N9oT/pHnERoDRp6QbNiS+fQ34A+jgJilUBbOQ
YB6Atgrucsp62e1+TrnESDQd0I2zvemrH+RZzEsKuZQ4KToXQsH7kwNS8PwHHF8aJno4mxf1rhXF
hVGIuwsL6xgOVk8XtqycZs0ayStiZmLRcQ2tRdRiKbKa2Na07bNT5/f2Vbr3JnrR+he4Qu/CA2K9
II3w0n8voy0mMmMbCl+I/ZiSTlKCBr2ozzeB4+6tshRjnQ0yVfjLFSzITh2bBgg0DtPV4D43ZSRA
ZmUrp+1ml9TwCWoFd+iriyb5LfsFRk27bXuq/dl2t2Im7AI7MTDOz1r7MwKnf9wNGJzOXC13RRS4
1LT2SYh/dGyahilSx9hu8WeNt34cOAlap2rm/cx+dTUPYp04WU62ygDbIs2bk4Gyzqu1ZevcAfml
WeMb3k3GEJtwwE9b6P05C9+NUyBMbZIkPSq/jVic6EF6MoWF8mW0vj8LtIqyTnIN/6wh9I54n+yp
v0m1HBU6j1b0NTfSixPR2vQOvj469zyKHaeLBfPQcpkaWyzS2sx8MxStXp4TZkIoDYGU2IcH0rEM
ena3ICKwlfgzayV+EWkHsxGMqIrDYdLSXKx+5jpgHOf5F/T8zP3yevtzhCrRx+eOECM7dZ4kaD4x
s6EqRGTv1tfZkZ0RNWZlieV4clNw3MS6O4X4bRfyoxhpwsPMXNOXBjYMwp9Hx+kW5RR5jJ3Kkkm6
nihWlXMGRr8N5cPoxzM99X7ech99rRWh5UZxjjfSxy4pi+B96Ak6J6Y4mpR5mlH93EX2vpSiKRRl
NdLCcNdh+AYU3VRpdDZ0NvqZBQWgSz2xTpEBT5Tl9TRAPMQwlqtBppzD2MbU1xHCJ4SW67KPH0n3
zWjUlfeYWTgW65RAgtmJP1SErAtVZRzOWf4vSjEtdwH0nusbGO/ZQowBtWXG8GWzEeOfRpwRWUkB
J0vzw3nXFBEZ2yS1GvKD3zW9ajIzznR39Yc7ExQ1fYMBGEDbNwVOu95dX0t8moTwaIUtQI89MX6o
7wSTVxZBKvYEbDYzyTr6lg5oszKP2GxpLIsHWnpaSXo4z5Wv8XAuRgYzvqbsAUvB35QpvSb16hyX
GKnFfIwaiYkVf710byVMiE1vQ2l3/G2GOtYkfNNQXsUn9MldPeyUid7YaVyGCkJJZkrKKgEdeTmm
X4nEm452Yt7oG0+43BtsSWRQozJeAK37zW3hyxg/HoZzfWfbYlqTt+EaxMfSIh9/nSkpnrLg5C5b
wAKhQ2gOc2DWcZKrWhQWOPfLT6odMXVclE5AZNu7zhBWSUvZ6bA0SrPjaKNTzcGn51DRf1rXDqVb
VOCAy+LEpKpcYv4Vg/fh8UFtJp9au/C2WA1++ANPjTx5HSNEsYnMumE/CIgn9agIYssn3vZfp05P
M/EnP64+aRUXfA6rw/Tmf/0mjIeDtYaptHbc4XjVQ6Nw8uymXNLaAR440Y1sX6ZmMp7xSH/Pr/+K
LbDwO0o7etyEdZE9zMOV1FPyj06/DPSnGsEOEpl2fFFbA4v0NZoG/NmriEGQdWqWb3EuBg8hX74s
C2xVNA8GvXgLKbeVq6xSEDfz4Sb+nYNiDJfbgyW408gQmj3xLgmAbcVyd9Q5+wwEzU336DjsXKrt
craZrNPwKlDjqwLBiwAuBpWbfT58HelYwnk/xXaj9T3kvtI05gxizS8xNEYRr5d9zkh+SJh/d2EH
6tNL+rVUl1UbWEbT2Tm1pxLTMMx622G8klFG+BFGvZnBkxHo4/e4DLU8XlDjk0XKUv0wFBWWAyat
KifuDAs77g1aFuBYLI5TDDs5MzszG3otRz8ARyXAoB8i+sGeOLInEmrx6IYgnk8v6wdaFWVmyw/R
TTJEUHH6EDJCvVolM/goQyzIwu0IisWsKwkRqumBb0MQeaZHeV8U2wTavNQm3KzfgZL5NXVkqQIg
1bJgvkjcsNVKK7Az5hA1cjzMPAq5DuQGNnfP8Nq1lRgVe7e2v2ukf9ym4WtWdHtNNW9Zn1n7a6Km
VPh9RyiorG1+3PZow9WTviLyb4HfTRjiTrFXu+VNxi/A7HXGjEIAwFAcDubDuxoKKLyT2I4N7+h5
zcjUEVt2pgFTTdQEFGjbzZKd5lZuGxXnonbrcWjz/3ReYU2soNR0XE421GQUCBfbCCR/nGVIHOuf
I9F2aCCwBjh7HACFm3K2MdrO4NMm4FCI2zzq0hxMI2SlprFmDpd1YjDNCTCWz8vUj3wZi/BjGBt0
TMvmQHX1NscR34iY27xCsBkj9QtZBPIKJgQKkS/f5KSlk72c/hD0kaoS+7AO2kNvIESaxjw76AhD
xxPJpqZi9TufLxbWhQxt+R8f03L5qTBzXA1t0KH49rKSQ8SomUbE8FfPbgY3l7dz/m91V4hGtH+3
1IksXb8qIHVJo/GVKQ3fQ1hhcmz6pyFrBZwRn47tz2CXJSRuibM1azldF4WZLQBBBDQ02xovuCs9
xaq+RUyZ/eUfI36EaTwgKTrODWYK2wliJxnmeim8PfIjCJTFgUtxg85XAHNQCNAoUjbhfC61sCWS
A8vvP/e08VXBUvCRpCdTo+aNBOuKWGGu4nuJpe1k9F4DfMfhtBzAup9LVdTOfQegEsCF8BvH5IgI
o2cTmIiqg0tIw3zWt6wov0HwlCYyYLYTsxAgV9919f0HVZID6EuXgCZJJQ1mWDvXWR77MQ6lBHTm
xdspt2wDwlNIQ+JQl60aQu/VDfgHxstTMl+9GWrsdLPNBI4E2RopDqFrrR9x4LGqIIP9hTrkDn0S
WJn7+hFqQ14vC6xOldB3j/0ZPpeUcjR6mZQWQYXlpeDnavAiVSt042eOiCGh3pF0XBCTrKAZUCRv
0UaLaSpH0WL6yiNtFkRky1IU8vkoQidinGwnn5EcI2py8JJyhCX0bHn7DJAW/FX+iJDzjWODC2kg
A/QC6iDhXWNFd0WcxXtAIbHPE9+5xh8+9OamVwTjEEIXlDpDw1J+4Au4Qy12eg9iec5xiNRMzyI3
UHaIMgvl8jPpwDIveQgqjMpJujVPF0WY12BwyMnxf6vNUqlwsWi9jnu2nnTNxEoJFkg69CwWOHuN
M/fIm2nSQYknG1+1PLornhmQCTC6J9iJNyKWZiahirGGJM5XRi6oEvrR9sG06dSaSWmXYGREv66D
+PNPCXymxKKhzcRbPLwCmFU5P0MlpsfkGCdj8ubXcj5TsmBI4s4/x7kdxnDHzel3s+Rm8oV87Y3x
z2Z8OLAwOdHwva5tqLSbKUUdpYqx6e11Bz70hs8wtp+IAhEaOoI5AWxH9EZlK4IgcaNw4PhK9yIV
j2SzuJe3WNdpCzXKnuzpllUOyiCxg1pE2Z7bJiENYwaWLt9niDKmdgbxj2qsozqhqTmMS+CkWv71
dL4I9uMfMp26wTSNPJKqFCZq75ZmtrfcS52nWEzoPN8tGJPCihtpdsBy63YaYE0tokH/0jbvIExu
YaFycmtJSHhthioEsLqMCSXdJE6JUy4s3+la0AebWqXeGxAwWsS/WPKmVwxf+a6khwGg1AimEStL
Z1q6Vq+WmXnMVAjc5O2RQgYByoB+BbW3mbVX8fnuinUUu2vd4G8dUXvL3C9TYRD+wug6bCOxGTfb
E4xUZD4lDoAlCGOSYM7FH4rTb2wia+Vw7v2b4BB7TSMxVnOnt8X7l6aYylwi5OUv2QdgaGiDEyTQ
mWfR3QSM/IZA4SwSNC4sYJ8aXWOpxA9Z1mm7ZLiggBEAMQrfmmH8ijVkrr9U2u1sXPQDi5dkHh0d
fwwoTZGnyjF9Zq7+jQQ1K2LM3+ZdI6/XxHnftlRjbrerhGa9Yp5NGdUzdjrgSm6shWG+MjRHD8K1
kwOHdXqJlvgMCaPsa5bLyedduOZFtUhcaZaaWaZsFv96BKroD18KGhnu8X+x6qCeO/88MjegwJrn
KUQe9cJ+yq7xF0iayxnmPWtiptiW0fscHxGNG3MwUzg68WYAfnzUu0d4U4pToHBnvmDVrm5/sFJx
qs61LtMtlBTCdwbBTojz7cmNZTryjDCH+RxbjMY77Q2Bxj4NNqZaf26WUYmJ3sLAwmGgQ3abKWkS
stfexmmxv9c0JDrkD/aIn/ezDMs7gbSm65oMZQ2/zK6z2KHYjrKvns1vgyKyqxyn9U16n3qt9jnP
yG7en4t2erhr/arTjJYhP3RluiuQ1sKXxKqKQljhWoWBI84SvEiZVyDl6/GOERNcwKZsV0G1+ed4
7WhBduaJqoj2NbHVu9jfcQkEK031m8iELXHFabXDl3S6WTinat369ZBzurgBvV5vH1OCRqW3eXiV
makeORByJTBnFUxXossjZ7IUqaygWYHGZncfu/wx3kO4xBhEvaW++4XuviI9b5sOnVb5m50R2oMd
iLHs9NMeQ5UpQ8AhsK7NegpHM8bDulwbQsjc0Jgvc3hNTqCa68Zky5rihWJOziKu6NHn4l7eCoAT
chgQXUFZNw9rkBAZSxSfT+yO+NzB/CE1BC9g9wtUTp2bKin9Hqp25F9n5HSND7nVRZal+ujPoR2m
sLhwKALDaRBMfBQu2Js0mNidpJuk1l7+oKPjB8VNg8KgQ/Weh6OrmAunv+CkBXVUGy7PP9sibICC
snlYbsWpHU1/jzXCNKBw8Xkm7zQnN0QGoRmbZMkV92GSZWPH4GEDT6h0TzIqv4T1uDvgtZp5BsN6
svThroAUMAc6UJupTwOEiEFu968bUtLtnPKOwzc1afR3waRxNyC41G7WkgEAyU63M9O12EdudbZz
MfJ1GMGQBqTzEJBylo3/AMj9tBgqmI/Kj210uTYGP9Mycc8yKKgWt1HsD3waIXKgzfiUXowLRxd1
eYgQXgrAY1dfOWy1FdI5xM4wvHlr6hGm57bwl2F1KJv5nMEAu+fOITYJgPwcuKpXKNbCpB8/VL6H
IaBE2CMHbidUFYc+4dScpfPBXrKGljnoSaKie3Ct6EtNpROiZifAFDv34HrqTnivAvW7ZQgDQGNM
pRw8EZToE+cklFxRBsYCOzebjaPqHl+gq/DNqXZDzIRPG4LzKbMWq4W6RyJOXLjQqQqSePqx5g9S
H47v5nElHR/88eFt2kbv+6xXIHWn1XUJkD7oMtjIpxs9r/s7g6ts7DIwpHd1WOnTCboq5Y202izK
XdcyfAJ7fwaWvTQOducLwYUjCxNK4zFPdNT4Bym3oEpUxXO9qMseAVgiIqfmc0OP+/SnVWrdJv15
pXiZkpgbzvEdLnaBswNGxOWVL2YCC9TftIzViohehxpRkvH8XNgZ5LBPUfWnovr548QpKy3tKA8I
8vWXv76d6+dU5fpi3/O4oaguCdqoiggedhXm9jJSd9Yw3Q4035egcoHyPfBPsK/iLjQMgUPDqv+i
nh/ec1WrbnMeGtY/BeOu68+WRjNgtwCLyYLJwFfNLY9Ghe90Zo+clSb0pBbJ4VtdHwlY61+QpCyc
2hzoi1yHg8DUF4bo8677sYDoN3j4BM8CQOQ6LmrkU754h9C154KiX6ozI0+QgO1BUZ+eOyBedX30
vegu2EoLiqBh5WbKs73vSgVf6hv0FMKGQVg1qbjxKC+Q93DOrsA1Bbyi2GrM/4jiba9LYPTdBpC2
u0SCplvt+rFTSQUH6wDuKH/KUAuPlkZ3Bf5C4RBG7JrSCjNtK1pZfy9wCvItu1GnbFrdSZYZihQw
q+m7ga2BOlsUnr9Yq6hH8gZEZmRnNbyDeqxP/LLk+LE1shE/o/uC5suf6MQYugSHerstvMzaxP4U
Elm+uVXRZq/Gke7We8cj0kY1X5NRt6b6jBR37Odf7ZduQeMGnClROLalxaOy8PPCvefmiZlL7E2m
75gRPTflnESHfXQWo4ySE4SGXm6W9pK5hA1syoglrOnzs0KwRBIIkpn+yVIGTb/Z9WN6+wx23tQ4
Z6Ru1xu6NoKhQH1oA6v8PDULbq89EWI5rPs1Xj/x+QkNXHJsAHcdNCRWC/3VYfhtJYZGEF6gTqee
oZlHjJ5nKi2Pm6oPFe05nWEgGrAJeUZfqGvvnTJwjlSXPD+PR5MLQm9PUexTCzkAe7q3a/MpLLgT
z+jYaSclpF1Gj4GP9f4Fpr4MuPsnITFJnpeyQAUarNnkskcT5UdSY7srfaCfRw7FbAU2HAkcuS9J
86c/+OoTPnQ1ZgKgU83soRGSCAK8aExkKiKL5SWzvEp8EfGQ4fEJXAmYdnqyeD4KYjqBD9h3VdtO
P4ay/PJCbV9SywpK7o/JDMjGATvMSIszJ6MwJp6CisDssoD1ZW5HoaZJRGdt38UBChFe2rRnAeTT
ZJSammr+QgrFk5tUa+ySlawBcYfFicJyzcTWfGykpSlGHQfB8/LUOkAU7a9KsPWEGq2nM1jpVmhF
PBeuCpinRp+ELcFfFHwdcFhmS5rJJYQNN6oseXXE07fu39mZS6Van/0J7AchivfDfLKdh3LHx09c
KbJAR7o+UjD/WuDs9TLYFnswMeflEBo3MKycvW+RgTAz2myqYSSIti4mC91KLRqfe+qPF2E3K7xe
nkp9zMYR54sLhkpLwyMOTpzMjzCF9Tv7f8TyeINqqW2zuKmeugwm4Kuc4qefZF/JFjjUecQ3gl/6
22ip714o566vkQcDH0+9Sf14ay7uUyVS+QRd/kLri/CYomGlKRz+HXWShgYqtbd93RkPXwKWTSsg
QN/vvtSP2Cn/jnadNcnK/8UrjPt4uhD//cOHxiw3v4oKKQPSnRt5nqEOALyzkCop3NilI8SdILqn
nre2hRfKKGRNzDiz1K+M5AY0/3DkxG+CLLScY5Deqfy4dJOaZfHuZSvCmOqhifRh6VH1oVQL7xk1
2AjgiaNBOqR7LIml54zaypXPydfknAJBUe1QtJZ1M9IL67IOBQch409veDhbOqUkvmVoNuAVCnvV
ClBsoSUaUKhRihrKE7SRWnCYHT865TjfRPPFz3XqiX/fHjnRMti0aC2RowPU//fkWyEUFVe5gDz7
25Xb/yi9nqtEZ9YtUCJc74cpQdHJwfAMAi09Yc7+pIlzeqAqnr+8EKg2gvqjIZ/v6eVdLlintObx
+Hh3HT06fzen06RH33RH59fNDgTCcHEauz+3RqGNwQ9XQVXI50Y64QGNka7d4M5E3Itur7e41gLZ
WyUyrFE9toAAwAoO23cmfk9LOgA1SkIjr7CQJvUAs7ED1BsJR2GQmaeT817bZMzVWBeDQHc22zPj
Ti59HCbXSgteihR3COyZ+bkKmk+eDqlu8VDrO5iinbcquq0pv0u5TDvMr5Rd/oCPxPTfSp690MZ2
Io/JuQ09HfPxVI2/3lwRBy52wQxCMpZrEQ0+KsdwR8sJY+M46vjKrO8gScSWwgR9E/PvIiqpbfQ9
fMrLlv0vp8R6wj1sv+npdkiMk1D9z3PIe7QKAfHm6fEUrG6jXO3SkUH/6yK9APw/EqzGbmJsjE/Y
WJ4EPnG6KdgkG8BYuL9wADSRhz5Dbp0dAeHmwI2POJhfPPLgqRHh421BbycrXhX9W33GGDDBnssT
x4x6xSpiX/m2rFkj90SrCMaULlvy/YM4InMSdjZurAoGHqX7jXTQISbzyv3OXr6nSumbohF+Mzor
6JC3+uG6eJAewtoB2PfFYoqWlkR+1efd+x3NqaPA+L2Cfx3TSDAsIio6FYcfhfIesihFlVrADlHT
owtnIT8FlYfcaJDSsfEev81YWJDw2CRslMOLRDfFwnF1VkPVRos/BWS0QSZy8JBu/Cdczc5vvLcn
UsfX1tWATQQLZb8lfB0TayHgBkGGb4kakeVGeg2nN1JviTioAIeLcQEkCqp/XTM2Tx6s5jKpv5nS
m6MWuot7NTSCuck1gZ8x59GaQVzsgtMNChzO99rRsv1jT8VBe76ApsEngoy431Y6PFNzbWFRAGDC
XtzGdwzHrzhJhvxIZL97oaeEXfWpfuHBT6edBhuGrf6RdXNx45/AhmWWuXewkRD73yxjSxWWEnXL
3ApAnUcdt0h2bTWkMmFTh0lcPquIBVFxrdBPdSxktjg+U9MIiNA5CekkZ/OmoXMdS2SRqjfSBnRt
bYwuffa50fNz8bjUIy9ngZQOcZ8eM4sYtm7CVoOvjOTUg2xEkuGS/t8VYiKaM+riIUTkwCzVJP2/
hjqyca9KPK7XSut02pMJpngypmMUbEq+63hdNzyy3jWi+OXNMCrs49kIJ7stRs/C+k4+ThMnppCa
1DoeCp0ezVwqVpamEcLousWcAY/whMgH9k7CzlKvXE8fnwjBpBUXPgzqMnAGlQoWRyr4E3aob+TU
tZk5e5Wlu5redqjZHun3NIhBDZ5vzQ0g+WqEA9R9RyMQwWR178G8glZ+mHfp3529bcrC4grjaW2L
Y/1jBRURErqBFyGIlST9nIeU21I59H6GLPg/kz4jZW8amb36Vi7R2Qdu0nHPlNnPp+pXR9rH1PH4
BUnyr9qHGk5SKvZQ/7Y5sBdlTWv8LmgtUn2qmHRCyLD+WvmjeQ5e5XEQzRr6pUQ3P/NfazqNl8UY
aJ0iqfNemOBfNCsWXtagEy3SlsGaT2yrDSogXd+G9/g5pTRpTO5e9DTZwPzmsSSQNLpEvaIfp39t
HtmZrs1SZ2WFvYoewFMaXF4IE0QwSOwsTJSBfEhtIQncAyjDA1fQvVmKSyYEGsuIAKy8mic2mRYd
gZupr6XqYErnewFgM3r00+da1lrXyBR07m3NYlU/9clDFDBT4/ubDhaK+jSTjBFnF2CkUFhbPgaj
inGR18OURlxsmLrJQ5CuXqGPVIbbRHSDA9A/5t9B8s/L2NDvPXYMWp5nChxwCu5duKKX/SU+O0b1
CyRE7xRI2aUdUzrnwlt1IMSURo3vGjhNNAdzYRC7bqJC2PzzUyJf56bGW/y2YX2dn8e3yTDgB/qH
pEM3JnItvOinldphh+qTnrcaVPS3ypPdVV4+P5zAd5yG0WyWhChnEWQzmXdf9lw0Gr/X0GkE/Blw
g21uN95xXaCBPL/MwM54XaU1lngdcuJ60TuNmE2LvZ6ue6+eGP/2OQOnpp8I0s1q5hOFe6p8Gkq8
X+befm5GGV5GjdhXuQBG+Po8PKrr7s1K5n2SzC4J7E8+wZtzwl1k2QH13Z/KIuRbvBVxYo0uW3Vw
kN8mQ1hHoGYhTxacOGfYTW64E6I4ks5te64tu6EEbQLP2T+zhVqyLLF3eF9OLjG4+qefzJqrRmt+
SRadSeZAhl54TeAQKIiwjPMEfYEMPfnEib1SX4qsmBqovhC3N9Nv438qLgcFN2L+ifLDxPR+guT8
yG5It1t+QZgGIiKjbREHGKNTcjIVn7I61e0a3SRklNHpRMf01zODQNZOh0g4pdZWu9/qeXM06fkf
/QNx67f/b2rkLm1vm2hdARn8MzRMHjdNZuwGKnc5/JppcS/FiIdxQLTS3iqVSwBIrgvDd+H7UR2k
qfBP31SW/p6/F6beNaNR0bSTkQ/+BViJkbnZTDm2mVUgcWs3hSxkTVR2Vwe21TvfFQUIjlpSoBgU
TvG8AuMvCbDbRwiIgsPJQEjbPvus7eMVWMv5wwKuGAbTJOI02yIMKK0hsolyj+MPUtpbwl/6yQqX
Mo2Y3Lcg+2O+PNyPYFcBPJVn45yPdIfY3bWEzQ3g8fuHTxzmuVIPwDbucpV/A6kRRHW/O5vqVJg4
MGwd6xLsMyu4erjDH9heMjCw7zANMygo3iv0wSlmH//wqq41Gtrolre+UJs+Rdian7RSOhBCZwBN
hwEg/C2Dt8shVPehF5oehPxeBrcx9GJy3hlxzYmIGpkRgFWkPpdzn8o3thkTc97J53crrovSNjkS
mdDk5GLetgArXdT2wkjLAW+6CnHHJqvrjEpdrSaIsoBjrLfwUXMrod27e7sAwW/W1yPFv9XfKWu8
E/3sb6W5sGecwihjKzZXsWmgqXDF3GPN995hVKfHbS3+YOHWrjpvarXpMcxNpPVB9PBY53eeO1ud
I7mL3x0uDpP7ZFZ+RPac9gyn7pWh0w6alEB1LwJTaoe9sugCY3NfLjRSYGnlpfnVgBnehesIyBQE
1/CowXGy9Exm7v1od/oIZT0jEnKUE8KlSKaLpwI1fDwLjOewVKg7JtwsMChFlK/SUPgGhDklU6BD
LwixVXbD9e5RqjzthSfTPwQIf8yAg4B8HB2xoFeLcZt1Qnw2NFdsKOgGmAbYXmqngDueFRltsvdi
McXjEm7S/M3mai1BRbW6+pnqbjP6L1loHU+56iGZBXr3cxrTFlmWk1aaLGteK+g/7ElmZnDZAV4k
A/2GGtmZJUP4BcZF3FrtygugzfdF8ZbsWXC3T9a4+3h0grL3UJhTZwLL1BN+Z0hbJkUP3GpvWvIy
i7du/QheEc/E9nNia8OmmBvCBz3l9bBF37+p/gLEWmFHvG6WoyscR3DpJ4fIiTyUlEdYQ+f/UbGf
RBuHg8AtFF+c1jK0R2QBQzoZvHaY8AJvscbRf7+zMvbzphEhTTREoSJUZym+yTcQb16yI8LUu7q1
+v38gpCvcwfnNs+o2Uf2f3ZMswll1LLDz2Lm3GVjt0hmWcoOgYivV1Rws7VZ/WE/vjd2aVBSyczd
OKMwIcDWVHAVAtcg6YBz26YyL3ElXIRqpTIbPrTihk103YBuNOWsqiyr2Kqnkh4c/OG8UbAXhGz1
SCfxOQRTcYpKwgJaNi9/8N6tPOHXR9ioZs68K1S8K6OX1NcYkQfDQmsW2h6K68TAi09XfKu7ifZO
S0c5lZGNHkq5s4am2VUO8upmZqgwQr8X44b2FQrHOlnuiYlh1BbI/m+4dEdFihruOnlsgkp53Y8L
81AbpL8m2dMax/TMBMxEz4NEJ/KepLN2qDjBUlpwQX6V/RL1xJjI3ua52fUZ07tAoS5QNLw4ugnT
Gv4FrXpFAsEZehh96hMt22QzxMC2yNrmkjBFg6zZ+KZcFqyYG5LtC5gNBBNXmIlNcIZjkzfWmCM6
k57Rrf3QguPwTMtQLA+Xco18G62byUdhT7qp5uSbqIwG+XwYl/VTattzVqKbRffjpsS1TYHA+EsF
FO2J5+Zy/nPHVdV/6gE/W2S8flBCD8uWyTADYC+cqi5M4Egw2LhZ2t6lomSe2Z/9H/wX5rxthgi4
lJ6XgLYpIt8aregEOzQULJJc5mOkc7O6ccpqsd/RANWJma7KqXt0ARVMQ84s0pifrEVrV7UxYRcA
VOi9vqzmeoOVogiHA6tJ3jUFc/OJBrPaWSqlBMBYfJQUl+QkdU1AFEicbXUhqWssqG/MZqBs7nN8
4525nRNXAGufemwR0H+Uk4Ldfwwmj5IUHUXKAbnOeMxis3mCOhwBJfkdzBIG4d9osdc13mSL6dc/
MMTlVm1217NCFQta7sg5I5Xqekq5hYxEdvTFWNx8zInXqpJejb9Ad9XI5zvouDIZ5Yx12THAMxgK
TU+h4EXVQ9Q0hJM0W0Q4v18BzDYoSC485R6FS3YDXp2hpVHstfbH0ZtpuUrqOKiuHVCeA0M5cYVU
/JK5fiOiRdmM2vDAFmIQmuhQi00u9PbIOh6gTsWFOyFG7AqGVRv3vkO4Phyr9Pti09kAfuoeHjb8
aQo6oTsSse1igk1LD7c/TvXYLeF1ZPqsTb72mHPzWdq341Ve8diHK95fRsz2M7o2bUDDcoXhBD5s
MCqM4GXBa/fbpSnPpOusIPCuIWAgtOA/4XCFS76RH9vlkuhc2WmvniapKW/QyIRfGuauTHmPrChB
zZiz//qG/WV/1JvNhyJcXmGhALd95AjqqrL86dtNomYoSSmKOZ2eFwYgtse9vLIvI0HHH/8AsR6Z
lVoEEEdKo7wCxqugtr7SlQJxvbMcM4wXkKto66IFBlMN0HX+sqvzObX5D3PiXvhehqsw0pumj1ce
Wf1/15PSKj5DIHlKRvQjg0lKndpUTT1+LY/qyJy7zwctEHi47tTMuCf/QGt3JKooT3fpkIBkd9ii
oMUQirLfP9KeOchj7xvbFdDzpoeFv3HsxrxmYryKRWK9qN+lk6N1V86rOPe3WsVcXv1rfsVWTN8z
xMbJ2xtIaNv661+Aa2RJS/l64mGbcjFCgGi/lrrAaAiLq9at7U7KhMDiFLXpMqTs8a9MYRVWJs/F
VMMDXJzdpmvvzgYQ+uK9ptojMYOF2IuIXltH47ptTCVjSghQbvh4H1AvILFiwoSgtVXtgHudt8rc
t4dMJDP4JqqRg9RGcYPhgMbD1KlQ7MPXmLVtqYUqc1pP4eZXiQjFdAWIS8rcFFrqk080BPjceGOO
ovsyS7B34H4mI3T7xHsItVxujqxKjEsrFZoV+NxCIcSb+OV84jYjB4LNxZU6ale3/Kj/TsfpNw4p
sCQ3m/HmBCjhmJiBepHKMDqhSdSl5e6X8gAUGB1t+YSIK9XQM4RR7LLLstcOy7oatyDnsjn+dinm
mx0i5aq0vFI1GEK7cnDQY1LO7uCeVh1V2f/ujIYoLz8Tsv/8NOMfz1ran+bxt1vlgxYlfdFMWJa9
abHwl36x+UlwtmNP7HjJZmbPvxkgTxOWalabXwE/PDG68t5enuP9VmwlLORSyHzOh4uXb+uTuzDZ
26ojCk5/NOUBn4YrI3c+FFl152u+t0WWaLcIWAvIIy2oDMa/a+v9IKbnii+XoVLMJigNaLO+zIhS
K56NHbBskWRBRWMayYB5cA9dzMsIVWVM6tGZblFJt9ejHnoKOTwBs7gqeBeWU50+bz3gZ31q1BX7
MR+BMZzHmeqUYnOEnwRRVPRW1E36/dB+c348jDE7n6D/6A1ERI9/Ux/B5FMyfvsQe5AOCqeKYaCH
pwyzZuRO2JSXnIedmV+iqQshTzjlwxltnTVroEe3dUGhP1hACHSIo3C7QcJtCKjGBqddth8vESJM
UfJ0gbTG/fjEMBiJde71yuVkLgC0oCfu+I9jmsUoHSZwUNrJCc1wZClxpFGSzB5nrlkja8xUEgRZ
7qMpxKZh19fud4dwaENGcx8ZZb5t7BaelE++kZGsbtN3gCfS7uMC1C833GlmEV1c48Nb8ADSEZa5
kq977f3C11XBaCc1Lb8NxvMSG2Mg/88RMuQ+H8H18yaZWCbHh6PRKAZXxNCAmd4MYJbpMiOdgl1b
lxi3wU78K3JwEMReYIuBJXREx92VCUQ8wXYIGtzquYVL6h3a0Upf9wdnkLkJxwpy5dKRjPwAAqA0
qmYf7FNGqAwBNrwaXrmLLAAu78uJp/Vetir6j+BB4ursP6IOe3510akLYVEFeoDiPYUQ+s5sn9xX
kEWCXYeW7G1tSkjGcs2DgVizPnQds2iAw4cam0Qwl/qqmMpAY4EVUxp1g73ljNptqxFbMiY/s5zE
+Viy4prYTQy80M5LRgYSqymf0HNAC6y7+ztsDwxswhuhyFHpzn0RbjfmqRZmFpLySXMuwn7DdFDa
eHeZuzhaG5QY+/AYOwxYXMKFhXYXoNHLY8dkAHI41sZYFROlGNnkKbUG88J4vJxUGGQ7EP+5qiM/
aLYHWi68rhuPmOl7lfyVRqTn7GS6P/yR5Ny6UUC6ivNd3B/lU4dEDxHIhczfNw5405D7y7FoXm8r
Rne4T2RKm3WDj5Qct9b0ZwErMOB8ac8PQbinLoclpNtkcqTSdk/sB2CFsNlfymh+ZhDivuIA3eE1
k5AZw5DWdCfd4mEmn3XNHCsVgf0TidRzmtsAp3BFYHIXEIKZynBxiyfLJmN26LoAw0wptuYsqI1w
7tg54A+WL5bhvDjm2I9c+8ge3QQV4szjxcPv9ntHyz2JQOwCrMsKlwCC+R7wC0wQykk0Um9l3QHB
mDPjeb6Zy1pclc/rOLv9JyZgepjhM7pd4V5cXgbzPFiwYeYJKpcYiLvrdqwJwW0qTIlpDyaIlLC3
e5xHkVc0DZCN1x9wWAlUn6RhQVTbfDUAym0kF/BvF01ROpAxH1+7MvIQXsTiYYtIAf6MwOMJhCPv
GiwDZhAFp+nnjhLDAa7JREmSZ2IObY11p/Q7zy+0pi6wic4Ii/399VAr76qo42araehK6lx5Y1gT
VdScT3eCZrPQ/zKpcJbF5hGV8H85aRyRE78j/OBLy3bOoP4dR/mj6RmYEz/rxJeuK77QQwL7SSFf
e42pik1NQGTfpSZNA4m7dG/YbLBW3W4YnwKmeJ+8zkzjroxf63KlV9qz31UqVOylp4OC+Ss/beOK
SXFbiPuIwWfL3d11T5VHsAm5UafIVgIc+Kt1GB3BF1W3m0Mo57zUVrBtECkL28Pdz9EjrD5cLd2y
32czlqtdWYRJR54T2/W66V+Z+etSBusYf4WgqKRK6ZsfahqtUo5NA92dQIFBKIBD7CIis0cFY7ic
K7of549uYo1lB1wljrSWKAQ9xmGQDbYjQnfeGewWMdsMqgZdV9mSe/fhICtz0ydSe/QhjOeWlxxo
FSTmpnA/VVveDOcP2TzapfdA8ry8dYrYg0tda9o0wSFpTI1ngpdvtIrDphIiZQ378+5M8aefHuWc
p7raOXd9YUdivmxS7iTFBFdDchZIvpImgQ6dZU4jJPmXDO8Ek3StzViBTRU4maHMgHCmLEFkju4I
0x7ce+hck12DFCk4ZXNPitfBwU34zxEqs8AlgjOLiN3+1eDxNG5FasY3GeHZYvXBjFLKvAIjMWQF
mQRvysEGxkSG/5RK8Qavj8nGS63rUKl/HjvGcT07mVMGgDvG1dZkwEpZAwrNhHy+NfHTy+nGWDgC
7DLG5klJ9mXRhG04G0X06dUFC3AyTqrFxFlL9/LR0/XCRnIDB8AWCcp9bFmGNwbDk8wT+mdLgHym
lfgHv6evYwwLZV0blpAvNElI2G3GCwSwmf0SyNxqPHbQCb7NNePydHSD6eCUaMdGeISx2Amtj7fz
+MWNRpFl1pd2U3Sg6+cPwZdKNbaWO0Ebyvu6lbQIggz2QHRxlyz9167yybmq2jq+7rEunmL3nGEJ
R9hulQ2hrzw8X1DBQ24gWezzB5xA6Yqs9hz9V48OboITRxltzI1/0mzj5x0zjjgyJZL+juc7c4MY
fjLG/Ndm2H0Lj+coHJuF5MkFfBMartO4zHDSpgc+meCNt79UojaRpMiV+j8SROFIaQFiiu6lCMnC
KPRkiIiSpRTANYuhLJIWQQvRrnDXpH8csJURyueJGU+8VKud7zU3+jeR7oVgEYq3NNLtxGU6puH7
3+dBQuCYDwqW1J1Z48YbclcwT7VSd3YxGH6BaiyUY27yoqNiOq5+hZlnZzIZP9rXzn3Guyu63uUT
HcwkZ7TmrapXrQmWmfxNWJbssLikUNSappqLK1+zEmhEhiH6YMTAiOwPEZ1B5MnNAqeiUqAm29oX
9pnfqrAMO5Lz2m/hT0KeIG1xEB1hf6Y5MMlCKRWzs95Tx4PWMo5xtQPKrWmzhNXN8oH3wXtCyHNR
7vL0FwaODYz8RWy57aDJ2wIZwiQV3yQ+P3eLuSZ7UtOXxwCh/l42PH8zP5ZNe3+FSwPoHcW33kIA
g47ObNjyen0qPziah1zP9Q+5N3bZNz/lWYY7E9vxirsNEtVD4iRDZZUIeHdELtkESgeTth+GkZBI
/g4I/XEarEzJI9yBpiueStHOwpPpTwT0Mp2ByULTfIxEI4I5usbHVBxoWqM7oUunZTWeMbyxlGnU
CEc5F6cKprrAf4p7gV5b+/PffbpQ4LZkS2XQjcEAmbYehf5zq8LN/eXD2Ald0KIxJNU3AgSgQVza
YToRy5YWS5mogg50sGOESgqgVdMUY2iYoCh4+NHBGx3bSLPUtTTtvHtTAg8MJeWywOJWVsC80cWY
oYHRcaECwYnbYPmbGA09im7ChBLBKvHuqkCl/l4VRmLdUWFctPhgzJKkWuEYYawbrwmMjmxfjzlp
vh+OkTRD7GYdYvz0VhvH/v3N5Toe7UQPRgcR7wAuigpvyT6nm2eFzJntA3XtlXTS7wlRwERQ6Gim
UZAS6w/4UqGy7K4JtdDPuk1TNm0XrKasp3ZreVXXJTJCEdL13ZdwNL3ZF3yVT2hh5C6xVB2hrdLC
fYu5nc3ffm/K44wtXrPNyOMsFH7aLpRv6iSbBMrslOEuFF5TwVMIPixQgp6yXvOPZS/+SbUarl3s
5UMeI//z3MCfu8wtjE0pBO9oGeU6Q0I+yKmnGPJAuWQdLo1wlalccnDMgjPRBLBncIjgOIkQQvLl
1jyfSghXf/9i0Ddx7UsnZzA1ZOFuJTC3Y0KTSiHCwndYUdnFELYtcOzyjr/l6HY5YGmQfzhvItj4
pC1/Ne+O+exTMwtHEQvsDXWZhV33t/c3oCd45GwhVD80o+bOa1zkPZPhbU1cELQiW+H23Z+JmFu0
N4+qY3FHJ4uqdcYeDjdZzQbRgg022a9qJQnWRkMcDnAEe04Ep7bbu2T/K/AvSGThkMgPZSlQkH6M
fC68/jheG/ayun+KItjp2qCM4t1wdC/VNiL4uFegPiaqsIDzj8ao5mdA2hQS8eNVLweDzhn83k+P
5qHOEbqfwR2o9jiagvJ3Yvuk+RmUUNM6tVC9WQBqJvVZ15TrSrumRoHztUBbxszCd7GADjFbqMBh
3vNC3xiuX8G8DZfU/nK5TZ6FFPJtlWAiSwcqZwbcpX/0AsyV6tLxi89Ne4i/EIKt5RsJqC/1WMlc
qziGFmzfF3ZEedsVJ2GfX4rVl7EJlBr26EY3VWm4msYuDyULGhEPfMYBaqvM67HvBD829jq2EjnY
bHSxJJYxcONMGqdWHueBJa/qOWK9ikPCJIBqOd09bBeQHUQDUTssqIeTBiWwIdfHQLP1jStEBY4N
akSGC3Kb1bV6KdI/6M4MRCxbVYsuyqwkKioZjo1aar3zR1bfxUA+cJqujNgud0ypiDMK8LPw8xjC
iM46OIDTfSErWZeMJ1iZNrCNVmSMRqv6nTPqOA/WxY1FbZPVGiG8bwxGGujzus7mNrSWqy5io6fq
yazzriG6UWSgepe2SKYvQM4us1p0egGwgKsbRph5wc32FxGaa4A3Q+vj0aI12adjyPlPuEVi6oIw
CfdTA2hIVq4HXXvP5Kfjy0vu7qhF5AjZZaphvWWKVsOoTB/DJyV6NosDEzfeheoYXJVGgIUcVvkM
eESdyAYjKycV+HK1Qu5oIQhuCdVh/I3f/I+YB4Xqak877H1d9WAdN2wfcA/dPFjNgVZl4ZQ7+ttH
Gk9CeLpFgfYT7kKY7JCaZyl9E3YO8ktOFYocEuaDUQFDIxpAPdH+6cIz6uKhktiY9jHJPZzhSdKG
vAUaw3VnJOGS92S2ewtg6R+SKwYBXJDZyZi3tTsb4Scps816RND//k/JWa3b2vbOTWZ0e38k4Vz/
oajVmxDXlz8daCtY8FSz+09yxLMWlOn2s01gD8yHz6ydmoBKcJa9kfRlMrTMhitZ9zZ31qhDd1AM
ygSYqiOqDlwOZmc5KcRIFR7P7JPY8c62dmXBKUJzKnJYKVks/WRXlAtlfARBCJWX4HfMSbl6cpbu
yjrIh6qQybecTC5Sxlshyt2fkjJpcFgQlt24apUwpcLelbIMLb6oWdw6iIxfyeCtrTDvyi2N2fKz
4oqTHt91K8wcB3vLDkEU34bQTBccXc8nFFGZ8KpcygyKf8l180QDyud7vxnIFZz0gjTE2ZtNSXOX
rfvtkvnAT7pLWkYMmqQH5W1kXaUuk4k+T/Qs9sj+k2Y53kYbumbTrG5EWTBf/urQpNPGF6UTJACo
zwNA3DiKbQ5KY7s8llk2mPOD+DcFLVJdC0nC4uGa4kYBf36c2Rl38h088j9aoUlDKgycWzKYsJgB
yR7aidvPwx+h6eJOm6Jh7UQehIJKv5OBWgcqVxVP07S/tbXM7fcNejehJuX2bD31FA2vtFbfcLzY
0BhQWNP7CFvKSg7yRtXfGnZNYk4p+l7eAsLLZq9ytdzmT6Sv3BTN7Gs/9tYIAjk3bIR9EZOB8V+q
LTeRKhNOsJ06Obgc/3YNsdg30/TopLJjl5BX/8HzbjnpgxQ9EMgprevyyPIOeqGgh7ONE7S/hoRd
efipD0p1hoaBp9591pOIphq4wJG4VQQ88owSkVifqb8FzpNKx9ClVCBkc1e6HZp2DZ2I8Ip/EKlX
X6oGZb3Y3wxdeSeZn09YoJwQtlYIL4YuGvAz6HlMdNrBYU+u81GfPvHqYhIXHPcV9XfVjw4gJ00w
a226RbxZslaUcSldpNg7KBL2XT3EaMTo1xXpGGVxiX+vWldYjvvmSWW/KKFxRYiFjGqGIZIdMkZb
iXeSWYq0JuGCkPl3i5hhEN4pgIGPs/8WOUpiE9W6p39IUVEOIksiBAjFDNppEsfpg4JcwdgQFBSM
pOP01SOCGyCvhStOc6HwRKvsBOiiyIU9JoFkWEY9YSnMOvL9g8kjJV5qsCccT+Bo9LGTH7TZecmJ
l5U8LV5CkzU1kQKbrmtcKBi6R3DV4k9ILvNFe8fYZhPrn8lP1G94m0H9DpL1tiBRlF0Ru4ncugh1
A6kqj2DCltTrZr31mai+G7/eqZFugZYt4jaqDqXhDScGn4pLpJ7MGwL3tKASIt8HRli24skJT4p3
69ALtRvACnBZzA+i7SkcTJ8wnws8QvsGWz+EgZryqjn+FsO02CD8eant9w9Q5N/3xWUL8I2JQ7yl
gN8xtP4bSnaJHMsnKDfrtn8LBRbFypBEiHc9c03Td2ZpbhJoaSzdnm0lmZZl1pDzo8aBTMxOza97
TS8gFBaDbRqstO8Tb2Z9aH1oYGb2UCUvBZ38MqLqa6x96qfW2510A2mWYEH+0iVwr+qlzzK247Ew
/EAmXs6Ns2U94WwA8sl6Ivf4qn0FaNdE0oHqBp4P5LOxzly4AOKy5f7TSNkTYFnw5iPCub1M0WEk
HRnl0Z1Cnvs1J4xVJtm+YvmYVTyPfs3JHS6SlEGSB6y5IVYV1PpqaJ0TjjcsJX99WIm/4RoO82Dp
CrHsrDEdy8LVdvln9jenP6ULZpep+aGYyRCMwFMcHcwpUzp5heyeNs+PDZZzJ187Et0044JttNmp
1exBAXSmpbqcGAJgfQZ46ifP75Gm8glm5+6gyskQNM6XS2YiKN+NG6mSiZP3mRmwBdkcxEpFWAbD
8K8Z8ZpYldRNGtahzHHNz94Dj5DHfO5krfn0LZNyZHRTdje++Lp0usx033Gb7/Y2LO7TbOYwdRHD
07XgnXrQm8VSAaSUunhRwBpVTU9O0D5MGRSOruQq8pcGs6VrgcxwLCkC9VTZUsINGx3Yfp66DK0b
8M8QggOanfE3lpHP+/tpTcKZjtonqxNcv8S0CMkxX2zEIUJWr5l3wdJP91cIUDuxfXuLgn8f4Vii
LBKJ68XDRcGJ9mP8R95z6f75PJm/Rw6DOfeqxfblFK6CH1nAjrN7CPczxr6c9coZjs3RKa1htrIV
0HfgtI9VGPM2wOdDAbKlWMf/h2blYBBM6LNyTUk2prgIOcQjFpfqcy0jj6W9mW1veKGI9MbtZyHz
uSdgNFgXguCllK24qqfnz2QPeZMj3yVIYGJAQcwaF7QFMuNg3X6hTJZ+pBmODBWBvqto5FKVOqFH
9CcgjKqsJOmKZgLQEq+ZxSYBu3u2bQOP03YhU6hwmt0Qk5RwJVgK9I0ksOl3Zik30rZlngccwNSs
2PAp7dzIW0ejWclYuUQgERzE7VOGudEc9XXOrBps+3YbUoRee9VgEjfIh4Ogb3xQ7gNvr75LmDxN
mUkqrpbvAi/asR9NlZEjAuCFp8/NhqZwfdKWVrICw8QamlGBtkqD9zka6dk2YWQbQl8ImVRI0dld
3UcdKIfGGk/TnRcuF8ZtOnXyNdHlvy9uolCggOa+MC/XQBUTfgpVuI9ZDpIdYsDx0kj4l9qZRSM6
kRoZnH5bziTXQnpft5sPqk5e7i9yl0izCuOUv7QgFf/Vz7IXfJUeYe9/4IOWKbB0B7wdOT4P+eqb
HTwP2cH+Kuip4liF5grPt/QzQMmTo7mifTCkB6OPbNXD9NPzkTLBqXE/qnBGuWBo7TLe7PJmQrnX
1hqGT4bqXoLujhlpz9i/vpLauDnxGcLJL3zCIhZbbmESmLca3rhT2IRs7tDjcna3sw90MRftoLam
vSgv+FjxfXa4nAZtZZs0e8f3yfHDxyzGRaaosOBik/+eWdCsJlnGXnu1u/iO0y4MlBrMEQ8nbMcr
SjzUnFA5zcndJQSZmuWqFK9VQ8J9r0zaqqVAU129E4nKKDcij5QWZZu7Y9nxfXDzA4nQ+O+avJSr
40AMUIKHhY9Izi36FtETbK23GhsloE17/HqMckIEZthk28eXXYwsOrflhrVHRwEp4UVcW11YVH/x
heA031Uvcc86Kw5te1FMnpr6vNvlkiWMuIi6jrtTRy6dxTdFJ41rqDEK4sy7uAARbUGsiVEbOFg8
JcLtCgBmQ/DpyENskIkcWRjzKNhKg+Xnf1VWL2OiVORZA0cb4ROoChw9RXqcVd+az5mOEDYaq653
VKE0a4ixIlzJEn+k5Zg0Fw7Jg02/LgzO0DGRrrvtI4e1gIKJC7+5IaCMk2xq0wqtBSmIawOe0jDA
iCWFiL/gWFaHjMtBnB53FrSa3Ur75uuUEu2EVGqW5vA4UMZHBjTdsjZMRTBsJe6Oh6Q9o03hjLDZ
bSePmNzli66jdd2YzjDOM6lulP+rTQis8b94wauDUERog/K8S7A5HceUmGh5T/WffvnhVxXTaoW3
I9M8sTpiT2+DoQp7RYYLUdhI8YU9t42Cnn9qSX3mSS+Fpj0Yoe4kJPuEyemzDQdP4Y2QSp87yRkP
UUJJtctgjMdZix5Bkg6YkED5qLkRnaujvXqj3gDm850Z2IWOxVbpgnrllegbQC2QNf8k+3RlCf7W
2i5fWj7VFBUI5+7yCx55C5ps0m1yERCr4T6DrJOK7fXjCPxg7qx3UblDJVYIXfu9bl6ktCQ2e4gS
lOI4FdQwvmlpQHRHhZhEwHtkANeFn1kDi/g/ByEUAg71jWh1UFeG7UVST9NjAKgf5xFTYw3Vp2I0
njE5csvVWcGIyn4obQVkqslNDhAG9oaF+IK4ob0j1Y2YO1Z/NRNX+H5ii+sEU61rLwi+Wk/IqA1+
/sP9zLRwYkNkvECEsCW0zI/ozzGA1uiaJOdt3e03DhTGDQzGN7R1Z7uDOebS/qaEHSlCu7PHYRiM
Wpbnu2nD9W5HmaBXl4+I0HokKUgIxvXM0CDKhQjHtanDito44sHuilgZWp/p2rmM5yFvFYRiMR9h
8buzikFZm1uKapcPkGc/8AaGnNlzK+qI5PJ0JJgueBa9qnmm8QPdKoPWouXxB6AJfdelSNCGWRnc
7WsP9A0XKMK2LXCyo2bE+FpCfK13aQ4x/tXsXK57ZTKeShtCYFjocCQs8YGUM3CmvCfNl8VgUax1
wwIruULJxHXgKdCP94wvJl41+10GKHWEoiPkGmjaLuF9GbfuABAJx9Ei+7alYaYfYKLDfB7HZJa/
yCSbYtUhquTVz5TQOnS/zVCjmpEGo50FCi1KefvPB0MJE1Ol09BvoqK9XyYY1H6uZ3JEVICHx8Fw
AhSeXMH52zPOet/MXwWDtbgYqqXq69P3OoLBcKXYWO+5lq/vPiaLplzWzH1NFAQDu3iLT7xzYvJj
8IbJW/GE/kU7DXpf4g469thXtIVFgmU6V6TDjmFgvEahL645Yxgs6gdcbKfo2aOu0HxOCpmM5eBV
j0sStgPgh+q2GHf4zaGLkrFE7xSyxRDDSXf/Qwo9c5XNsEMpkaT1rloLblRtFbEcaVLyCX3s8+NU
6EcdzmwOr/1IYtIMrjxGQa6R7F59uyPaO+1oGcjbsxIsKjzMqp995mz20UGnRJM+oLvn9vUjJMsk
atCoZ60k6MEBVVWH7MaUtow4rt071QUeqgCDOeq5ghitW3i7fv+Xli+dWjjgoEBpHUqKlgq2edno
9Hs0H+zYixbLuJiqVILM9gqmWG0yg2CeI+k2Ok5pDlpMSKKZOpav57GlNQL9peqbljNrBs0aaJIG
SlIm30vL2nJ0RtfEkxJObmAvFeeqK2ZXz1PAL4pk7rAHF5BMjgLaSBWUlARyP2oiXwkIMRZkZ/EV
1c43WLIrkXVdCujf3gw2I0d85KbTmAIkuEXMHGxJCdulD+duTiEyA10VRFeAKHAW4Vod6G5/yQI6
VhgxdwmzNrA3fPLAKWnyTj+vKuk8nuNKpHJzy3+3bWw6PIN3JqTTI/hispadtwV6undtQh2trlrf
yC3XY+X2tXam/TnYwnBkhTq7Zbg/ZY4Nt0E9rJm2ogiMPi76SgTzaoPU9cxTqZcJQg9lLbgeLLBM
FD0Dj/KZVYFc7/LOEXJHgUAmxxyLAJX9Eq+PHJnf3dotsGEzI7+HSNJMpWXYL8EK3mkME37H/jBA
7t3v3HBOfej0UrgVhirU1fLhBA/sphWFU7uUw7sJMQsyTgRvm2usBsJv8AVJ37gIrBaDhUjcwaHx
XQ1Sp2JLjtqjhLRnupIrMAUyIGWpIKHhlUahw+DH2bJLT7oPxqgovAIM4iStO9bguL2xMX78hgid
UGpO3kJ++HCBAbinw79RjIqCg9urHv/yoqmh/tIqWwZE+wi7E+3Mx7ZAm+e1GXvR43HVhn9X7C6i
4YGmub7iVbmtKfH8XwtXw2wem5nMxaEvBT/jzG+GuOBzs81X2sq/P8DT9TurLg+hUjxOac8a+sXR
t0GpLLZ8qg3FiHSkZAHjZuCCRwzcphX+T2C+aCY12RXfJhIRO/kOIekZZHLG3teZtPXv1fmbVJOU
t7w1WY4qpZgklmoDsqAdUo9tSQut/YQ95fYWDKv7iBQPoABp2C3ZaLtZqZyZD6s/MezGf7mGLCIR
DRSoXpw6Oje0Zdhex9AQmM1a097dVBY+SsL8Har4hNaG08rQ4F/FP3J1RlD584ObkIePGMFgR8Ru
GbGewJ2NrpVr64aCspo3QTY4FcwJPaTJl7GH7E0RC1Gxut+AA+Kexrp8ELpSkr98JaPvgi2pm9d5
hexDx/V7f4+z5twEciySZvJOrR2kKV95itn4C8ltmDezRM2ehc4TEun/0qFhjTQlKNENA7ZqJyh3
/nsQf0q7tFnkCzws7TwzE4rCmYpraCzwXJHVaLDN9UTyoPW5UB48OfJofFtbz76+lWIjtsC/hKwt
9G2MOKvTOjJzRfd9NRXi+cJ2jQCnfgPnzXH17c1Tr3LPcj3vEat9bGfhmONM4zao5PMYs4tc3CB2
ZqTJy98RO6tBj9bbX8pLD10yePyTpt203S/GlJMC5iG/eqhvzUqoJLwP/1/DP9mSqHV4TYooSt4Z
yrMWeYwQkSZcda1Wjyl0FyCQHFm8AAjKpQv2HNSsRIJDLW+h4/0ge05ln8mj1MHqG4GvQZWCCAR+
bVYiGLsxotX8KdbebgDbQFN1/MjEkxmlVm7oziKIsZ3H+RCjziZy8aUicE7LalcTAgBZHkHssUy+
6ydy43nLrJ5ypJfJ8XMO9b8e8oQ61rZAtM67c+t0duP/afB/g5jU9qHUc1GeovRF45RMzgXKuDZO
Z88zXokWmR0fgBv8VvOv94f7QReUQezTmIHc7q/y2VbuoEbxYwfDElslRtTa428x9Y+q10oXX5A1
IWamkCO9/44MwXZJKzrsbgID3wT/ChVsy9rLVkfZTQYDJy/ACH3SkuSUAKhQ0vmtcxD2qbOLp8H/
isw8XtIYD7ka6a7HBYR+CzRqHy1RSs/LqPhYIJ++TlcuPEpCSo4eHxz9qSBwqTnNyvV93l8rkHEY
u9T/BJHu5SmPIFXS8kbAJUeHW1sOQZInjUTUUxgDf9vm3rpEMfXM5ae+UJysgv+7SP03w3Zh9FSz
GIlmmDRnBAC6b7vjfsRSGHzlZt6ZrRr73r1T2S10pJ5P7Qp4PtYA+J9ut1adk10B7uZEv5suHgNX
Tyiv0lMBCSzMpVli5kF2lRaJlTxeHOA5zB2keRcWnP7ZcIHwIWhqxDwBfUhmhMa8wuTK174bO87K
A/iGo2wenFPcACmqzdC0p4V56vGuHVRD23XWuL4trL9cLZiNJ8Wf7nx9ensCXgCxGxIcx/utDMTk
o9s3c0GKx7nL/n7xaxXWlZ2/u4U0iCm1AskLp8a9t9iRmMsX63UAtXDRMvWqUlFRwvbQxdNlpciE
BjbTaYEQ/i62Kw7UofuIauokO2xLjxelbRvjqW88nJEWTboxr7Qar9omjX/iFzaI7xo87HzYPFlB
VPA3X7vJK3IbAShgQNucCqguWIYzdhGWXnUWx1O8kWeSHejzx/bqeXVeIRoZsaSElIgw7Ei/0ASh
ePSUi0QE79yrHJg8tQ8CBWZunAEaNqXthAPlenbgYBjGtlxKA408ZCC976FeELuUoRfDjqhon802
/HOfwKnHPy5dr08X08rJ4IeKYL0SOYQvEQh9nSin7a+65pVTRmRkIAMqququ+XXi900j6FKLfkvN
Oh+KdFDsbc+hc7Ekw3ACEMZD1MQjIIgH5Y6hKfXVdZZSVTPecpiCm3lZSi8rYjiiRdNNuXXebcQD
FLKDGzD7V3cm8C6iaJeLxd+xygLktpHA5b7yyvenc/2rVPMk0rBYpD/vgMFL2KkJoVyMG7q1dmB5
6WBOoVipAbUblrpUqpf78ZAAnsykysM1vqrXmHN350qPK7taUcWZTBLHaIqgFR/zJxG6CC4Mubva
TLw5GaA4tdNfinozY1p5sRzQS/wYHP2PvG9xJT0ie4WbDrvA3zU9zkAoQNf+aECOpx1xn14NV6Vg
mIGE/uFyfninbkYuTv32ZQZLGNsG3LKDx9Ygun8r1XoJN7C4kvARXKuOU0zvTLANn5eTOXfVGY1M
14xjItqREJSFmCMVsqr//O8tSVpRi58UYhjadfoj5maZaBOnsGVm83tyVmHDSGM1MGdZU1JFh7OO
6GdcV3VIekciNiY/Gik98EOAT6Jl1BC8PXam2SbkadTEB2zpwv9YYJFETvi2j4FqLvzMCuKN4JXk
4lu40G6Jm8zhtxHYT2t0RHgRjk+n0cwlwhw0ObRyl5PQBBtK2KY9rijQNE+Lihzm1csJZGnJfgxk
2LQoFZhuT/jPSET0Bv52/seCGzyVGcht6pbXrIPw/OXvtFK6/X+9BEPX3lp80G2IbNIctOQMO0HF
dRM5TAW9coxAKeMKSi6oODAS2R/m9sRrQnDB+wK2XNYeRO+QTTjl1KA5gtGRpf2tD6vnULXdoh+K
tUP1c99lcYYlFVsI1hK9oYX5DKD5rgkU8EjiGuoCDckMC+QxKEOqlk0c1pFqQy0G+ETK3r3cuugi
e1vIoKGS1V1GMW7V8cgTEvxbR05a8gOMDGYKjffofQgi+g/jU78unLap7CoRrpP0LqDpdi5fWI4Z
3r3pd4JRm3Ikc1MxfMy/Q5ah0ct7bLb6IqeGpEP4W/hAOmWKB2kZIRH5v47okICXffVL2o5J8M33
steS1M4OUL28MsN3P/orxvw4/IN0dLWdCPAQWZpJBXzCDIsDbL386xWxqdB+H0PHyly5Kn8aFVhN
aKsCkOVT/eCevXhtZBr1L61PNo7WyXauZ5EDA4JttQIkdFIWf7J1OibV11jTuBm1ES/5mc0LggHv
HO+WyssqFwo47HAgtVD6TCoYB1eeNkgrym0iy1rjPdZ15tVyJ0uZqbvW2Sd6xo1iEwrNu68rQ2e/
USANvhHgMWU7LiJhj/kU87Q2eikpwKEoSDArvJ/RER1atDXvfRQ1kr4gHVwb6Fh6Vj8KdeBfyRRB
HGnGBTO/FaR9gQjWqqFUH0+lz/ltyFPwcpLQdh6tRb9Ejl9ireDvs0/ltsNfOBB1IXK6TATAUB4M
noIW2d6cmD6tgUiG0eYHY2bFU58sSJFGnZDb5VjMiimlFZG7vo2jGVo/1zJs8wCegg0bARI9S26D
IR3soNaelfgjyj/vMatgP6ojlPzWip+6q+E2jz76klc/K9mpSsuNqvc4Uh1KSX221R3NMQ+W4DOT
WUp5P6p32J3foEFfLhDhuqX0lyXFqnMXFTmrca31MWT4isucAJ2UksVRRzBqN1FNGMto04cEXGJh
khFTrp7mOLWrd4LyyuhdZLAJCvejPADObtCrOtXEFxEipTjazy3IiGICsu0aP2yn/DWnFKei5weW
6r9xSLAD+1FsRvEYl9oXeKMHn1141N8wyj7Rn2cVwbWaMaqGPWLCzHTWppbiVpHpBwncNA/DbyNr
rI/Y4Ma2loTWblauCEh5msOxhu7fDCR9fUaTuygXdjHrYqn1azhinJTKIaLqgryLbac3isVPHFjJ
G7462iHV+/a/MtPvL6JDk6n8f8Xr5v17Q9AdSa/hA8EKQVMaHiZ/CqhIVegbp/k4QUh1uTQWh2/e
G4W3b4MEvKjII7fv7ttgWLn+IqXUKi181zdrCmj/5CupSWbEKMD+Sz3hvvHUu+ddBP11RnIA+qdS
a2GSZDaoCIjhkRCpXuLnDllaheigqHjxyLGJMvjVlB2qq14jWHlEkGbBjUPXIuor46DJ+hmDtbAH
l/60cdKlcyYUE7eDFDa8o+5gGUbhTWddpfg2ZQEnAk0sWVRpmIliXBo3iWcSBOlwGhUAiba9U4i5
D1595YX7ij7OJ+jUHcdFuZv5ihrKYCZw+qpmOJVRAdJvaZ2owwBs3X1sldmOR5WMaIeN9igFbQLJ
mV8CHEieLJQbT2wxVoB2twyxzJqrNarbx4jzDlEnhyTSqkqEdICpj56MrcvsOp0h3BeEsRDA7Rxw
qgc50o84yp9XBw+KnmKiDhxVCsegus5KXVaoTYYKS0mrgIEUUfwMvtUDlv850zQ7a1uqEn+ypgU8
WlZZR+edDwvHHSVNI+NOA7l62oPGXNl4t/Eb+Boj/kmeuNESGbmuSBK0iICxtPlx6861vVia1DI5
GGD01DZszJAEWctyW3zETi2aneHIlQUqP/PiWayjjhdr7sFrOd8lOooXM3khTPpwjGwwqZTgjRQO
r3RESybphHsLZN38Qxrsrlf6dzWz8QBiBVM4CxiXq7jqAvAHY+DBxTAgUVngrahOySg5ylro4tn9
rbs+lA1P0kPGliMAdPPMDK4uD6Bw6MYQzQopxCwykzV2TuPuy+LVAa8QZd6yaaiocg2Ylq9F2jIl
XUPBWyLasQaGmLybYlSEP8aNEDoqdyOWhLEXvahcaY+sJbsPKZkPSiCnbI4QfXDWSfR3a+QlsrDK
Ang0IpBMd4ckai8G5sAihDOSoVIMETeWvSk/hdpPSDIO2kHc7oGXV36af9+BEO7Ll0f7kaEQenFJ
uThKZMODSFOqPJk/N1pLX5LFKes1qQ8hgQGFLpT5/opOyAXvyi0V8B3ZguzsKf8K9B2JF6FY1w0f
g+UMhW/DaQsbmG9uWeC3fRYtKCtK5t5LpTdnU6UT5PkKWCIbWk2sI0jKuotanm8nwmkzT6HhfHvg
Pv7hif63Sr5lY+E+p4NHNPb9DZKdnBM6lul0xmUKShyy4IbE9Bes9NME9fb0rrmUOvsujC4BDgIY
gYUDqRKiiR6o/auC6NlV7eSutlb+HGXDaPEvyDvgL7OICJGxb+M+cbmh2rdzYgKI/S+9ZnBLY6LI
QkS+yEYVv5MNUdHJVumWGOq/00anvms9BaDvgZOb47WHMkIXr8nL2z8qB129JaSv8HZEHQVa/5xq
4+S+EYJY9bst27KlnsLvN79tnmui29mlRIKUc8RVnzG/C8+NM3VStB/PG9JwqXrg9/62epolibhX
CYt05s4D8gnldzAyII+cAYW8YTf/iHOWf9FFe5Gd1Mg0639drPf3dhlD+VBvMbesxw+9ZNpP9DqO
Dv3zq453AItUDQDAW9J/39+FeD8L+9ylIgGDXOhpA6zKIKYuJdxlslmK0pWL+qh8lsCNB24uCpBh
M0eRmS7446iNJ7ez/KI0t4q3B7MIIfZ/TrNyTEBQWA7tixNV5zR9TaY+9nI7SbSd6CJvrqoyr3T4
1Vi/Of+s6dZb9VEOH/w9kPuDez3r1OGGG2E3F7Ijb3uL4U9kX/E5NaEXMy2sRGCJmAaveU/UFmnt
+eiKCRP43AuMcz6/xD5TPcXsGBS/i8UyabVOUzlXK0OobI7fLNT0BjBxfKFPUoo5VJi2xT0WVBFp
XmMntJjzwvFKXj2xqr/J8gseGUapXw5/Br8xxUGvkjBmY+5JM9ar3w1ZvWM04aq66gvJic+BLth5
hhx4nc83TxTrD1u9pcTE+7rj9iwTBcoToXLVpEkn/MgdddOl278FxZgxCb+OwS4j0yAeKckkEiVA
wC+uIjhDEsvkIyimTGWxQ+nBAKZjPVetc7fl3YPkJOypNumlnt2/C62+YIPH7jvVNmZSpTe2dyHo
VGmOnmouzjKzU61f9juUhMonlVq38OiYflKeQMtNj4ZsaodTlO98cGG+yfYxaG9bMCPq0Xlg7cKQ
JQ+7HIzZnz/4eRJBNMvj9iorJmbXsFXbDg5zyEgr9qFMhqNi2dw4h3bd71foDICqAvy7iBDyVHex
W6oye0UDvzfE9NOfjEKwnsY0lggh+wHq1DAzXyNWfVM9xTiMKCN0IIu8KbVgNQOez3jKwC5UdQMa
v5/h/BnH8GTvl+rTm4r5khkzbDN9Nqu2EYdO2UrR85feX3zK+/ihgTI0W1lsI+79BCxTa47fSzM+
i6HSoK4HG6no9+qt2KZsgHXvTB1kXVJEo/d/5SFokYzySVCaT7NCEBwNEIrPSHHqQwqan8V2fAMi
i0YOMUhFQq557mqSkooA5tSqg9w2NoNQOuU7v8R0/GVp0ZBM5lh0OU5A+4N6bOm7/WnwYG5y7RlP
6k+xO0RsF7QPQ5bwEX79JYqN4YdmuIxCJ7g9EjGqCmwnIOaBn72ceac7MjXCp4qrNJoHC6Jakjam
2Xus55cZXSd3JsycsUSie5X+LT2DEijRVbWtigq8D+73h7fLo8zQRpRuzC3WFVrc+FXfsNhMnIY3
J0VkJk7hSHRbd2CmSfd3/cXMXdkt31yEndF6UcJH1HzyQ42qojjzwVXE+ybLGW3D2K7mFOvx8Odu
Lmq7Lzkr0zWw3dzNPEyjQSFEr9MvKUj/SMPfrUqwgddQRVOByup0IYRgsCQCZDJLzoLmX+EVUA2e
T8hjzwvkAjJ6HKkpcN0F4qfMnrjl4kveh0kfEBqRyKJxzi62yCGIhU+88QZShX9NOddErjEVZxeD
CcAnuysd4qBXmy2g5hjV1x/+pf16gOmnbPjhTcZ60PtPTi8CUlirDN8W3uyisnPxdCMAPNdEKeg7
Qhqf5eHp7z2vLMHdukD6WHxSkS89aEtME8+rg4cu3kWjAFxqNxTbWYYWkPNJ64BLySmjHA4+a55a
JoN+79nkaW5XyvFcWftiqZuRnTwvilLiBfqRUrKE+qMq4Brl5IrDDnVQuEYogj/Gr7wp+bjmKcZJ
xs22StJDwAQh4VjZcFr32P2IS1GNMw7He8qndoY8fBFL1eUfRlsaC1ZXPYc3PiK6Zcou2yTvPozc
ifircLo6/a4eAeJxdFPlXtCOmM/nwgkR+mV/JHS2V26sSzs4IGXAaCJFj3WbJJgD0bhbq2FwvbRv
kc8gAJQTniKA1ZdWo5AXWVQ+qA3011T/ySSn9Mq4HZKl87ejpi0hNK8NmQIJBFE0wvT70yAPv53R
N1crvoe7xIgCYNVrrup+4h/lhqja4s2yhLGBrBBvEJ372WshoGADylLVpudVnqS2bfVDHMxag6GE
OJ3mFWAbEdzOjqOwlocmqQOzK01LNS63D6hcFIESbPhs2vCLLRywpNwoId2tE9u77yZow+Ed51tY
cKzZ6pGcQ1ST09DUVRk0A1x2JHXPTKSg38kLts7MKJ9B8ewa53nrWjvAcuat3WYM4gj/A2BE7UEx
grgGpBqtl+zvEXgGHxlQProl/vlh/NWE1XKlKlEytmlddMHc1QpczXTZGIFAkFF8dTJSNf/GFgS9
qG9VVYI6URUxKmL2J8RixUsqymNTRBqy1f/G2VWO2mY814RPDATKcNR/kJ8OdM68k+TKyQqtyEo1
ZhAC0lUHtLwZOBj/UD9ltZw1NWccocumUUg22w65sTfOb+qunzk4qHFa+fmSc2+RafAZQcW/9Lc8
n0FNLLdUmPYu4XIjZ8sFDGdOikS9tpZHnPhRtXmCOxYnGULgTEdQV/l8/KUEAPj0b41/0FjY5l6k
InGs/Ty2FLN0KwRtzrEMjMEQuG+TMpSWbW7thZ4lLlb2ltZ1HUpvrbQWnFAzoMaEGmXSzTEN71+P
TD60cTOvhhFpnImej7eTgjjTiEqhuT0p445jZw2p6xA3EVaI6aVDC0hPNOtCRBDy0kcQIwiYUCG9
Tth5nWgcM0u8dwmcnOg0LFfr5toxVJhIvbZH3LZ+7wotd87Yq8pwVPdtVLw6dIifBzJ6CtxIM3/D
D34ox1tcAg8tRrf5Zfh4QtPkPrhlUMpBNHpqb5RwkoXIi4BjgEhWYyz9wcoZj9J7zbJvK+8PhXIr
McWzdjskqLfvrwrLADwfWFC0dDFNc0PrdrG0s6ZzH2x21seykCdpGz9M+PohWMxsd9QewdjTquqq
VGWgD2/88uC/J44e/8Tw2h8ZVzZjuaMddbPrDtuKkSFoEUkVuFAdy+osPppaXoxLnCmAnd6KIAQ3
qvklHIZ+vLs6J1+7K4p/8SzYiwZUrAtnLkzvBd6tjULohx6TukYLapjG2nL8knLDjegDqMqn2LCw
1TjDGSm3W/5zgUCcthuGsTWAOvKOPIeXnhXq4bzIb1LeYKIrn1/Fh/doXBV7tX1y1JDhnUaFtmJe
l1hAqlHqIyg3vhQ6Q7V+PPA41NIZykg3g8HPxujl8+fFhmnH/KonZ8X4KuguU7G+Iv2ZBBhFik+2
A3zFeaYxsMu0diwRMR8B41cU/HCvgvaEdshsfZEHNi2PgTPR53djP6VE6NM6KF0yasXDoo00MUEs
uGO3pwUOA/0TuylVW8K+YC5iJdjpNhW0gzkmiNDmm0a5taTWRP/cs8KeqAlNmT7cKrCIYUI58CnR
SWjooortpOu3dezAixa1gW9E/QeHffgOFDSlbv7tqX1g99++RACkSB8OSCRxDDS1tsMzeihlzxUR
p9IA0vuubAefHbaNisw6vb+jKEBVIxj16mnLbDVgDbiaQRgPk6rAz7aRNEMhT7TE6O+gZvQGGJZz
zzPN+HB21nftp1V1+7d/Y/Gu707B8nUifq0SGpiLteQKBKnHKA7qYoHY5x3yQlcCwq7YeFnPI3+4
e+80Ifx2hgWNQpvLtRTzEi2ppuU2geGrUh4SSsUFIjzv/SCan5Vi9y7JFr94j/V53/Z9Kglzfhyg
D4JXY+0p8uV+hgUUmhy8tsf7dyu8a7UI37OFXt8idO2Rfeu4THJZlD5zucBaYRCct/6M2QnTqv/7
majWZvN9BNyIy+B70b0emM0ozqFb74FHdwzPTcJu+3oriLMv6y19tzvoc3mNWmhgSHJAhgDC6wfK
36BZUqmy7B717t6iOmBs7BiitX2lLROUv3ocbSUcG+IASREcYxo8F2jLvsP5RrLCNoBTCr/fuX6e
ReaxMAh7eJG4B6t1xYI3k7ZgIi9UzjpYnYcNsM16JVdHVXH8RZeuokjQjI0rk1sTuDctFMlMlbYF
rLnL3tR5En950crS/ghwHqZlBaMmPg2mi6/XmjfU6eZu4cGYWYnCWjX09LrTsNPhepirsxkVxFq5
Z7UyeaU2cEhFa8rrdPu9rU8luNqaXxN2OQKiwpzLRZY/Go/p8kPSCNPl2kehBgjGHsUTZYE3neWB
TbsDFi/kvTi+NXQp8R7gU86eKQkxcQfa7U+yBS0oyMCYXYQ9Q7tumGMpeHvjVUy5FLelttQNynIB
Qtx6sg5qAEFULGh54goLjESESILhNn3TSQc+iH5g78pB6PyI3Iz1q6cHoc5GsyqAS8MUggp7KdDQ
eQb6tah7eCHtGjQBMkbrX9CZIJUHJO9zaaLmpef6kYOhqnREdnjjFO09qmmGABGOmcfhZIiiIytu
EfY/1TrB0IQRtLdI6jUKbizofR1fQKtF1cixwxW/PRuQf6uxYyYh5gEN8Cng4efmxVBNxSTOtB6N
55XYd3X53Sco7xEulImX87odL2MAogLWq2P6vvv7x3tOM0oDpRUJ7HbvKvSsS/DvwWfiMGlIwVU4
iT+ZVqfSvvgji8lyOZ3XyX+d7PB3anw10rzYhiPDrp7DsajOveeRk66FKlQO8KrqmLd/vjGzsfyr
1qjZoD4E3eKnSYywI585eSgYTbfGIjTZBn7REdwEOtUXzIWE0nkeuNWQV61LfJtXryQHwQoIWohv
Bs1R3rz1Md98ikDpILVXYHV04hRO/RYpouSF4G1HfF35pIpGzw3EQq/2tQYQ8tMdwoap4mnVuM1W
tzWtWFkvvRglf4pBbum0zujVs756NkDX59TKDoYTRAEi+5W/0o5gRZ2E8bHSIFs5gjL6cs59J7Wp
T30SWDjPos2X7z8yYy/iXy3pmne43a90wIx5O4GFGjrbWiK3o176la9gHv6oHUzR4GupRvx6z9v1
NwuWMSJNYXjf5+KAwzg9tZ5Widwa51w6TdTbpYHumsEjP8z7XE6an3ROAG5MUzYOTO3OXV2/teQM
7k6ZJdZMDei2rNh+xKLerr9oA7R0udZZYPp01ra31C/gxROaqKgds9/EYXJKu9Ru9S+C1E1h6K5i
xr2EE3XjwzIBwblWpYOpLZZwmY+pQFvrjFpkkXAem9NNcuj2vXmk5pfJ5b+zzJKXhjMPDLk+omfV
y7zn36LRmcDnaaKqs12a9CeHuOEuvxMNZw+yal2XLWMQOn6eBC/2u/mjPLohTmeiT/lAlpDbJRNF
OF36AT2D+zZNxoFt33gUvc2WOGFLFimbBUp5FGAzfx5VSCU3OkBqU/sEbWz2ov39H3qp7InAD3VN
QOdgTD08DKmgKx5RLeW8w8HPHLw/WakWk7vr7VubMPCyoSICsFZVoeliFEYDVkaIn3BHtSCyVtA/
LioO1QAGKwayzWtbuAGyvHVoN9naJAR1J9UhD+zcetKHnByPqh3OIgu/N6ErEp9U3Hze0WOr9zRX
+qFUi/whja82A3dFGVD/ONRgnlM/8TyXJNZUy4h0OZD/wMq0+SI9kjb4SGlnoNp1MgKeUGn2YHHt
sq7uH/tBHHn0ug8xIVb+xO/vLt57WBOH2FhULWsz9aaT6K+XG8QeO3WeBSGJac4/dXgynsLZbMUf
h1rT+mhYU/SDnDBqOWbxEAhErs5nYZwOVTtNwX2jJAxhOtgQTdx5RthmdqvoGimr+tCGR72GSRI6
GDI4Uzj+7DilIzbaVKyIFphxrSw2E8mZyKRQ7y99qFsT/78/SUWYcVNavIVgsY6SoMvFYz7u0M77
KglsYbpln1IgPKp80FTikACCrllw8mvlXhouRKaueIrWFNyi9szZo6EfNQJY/fNQmfGez0aA7xM8
AYAnbOP71semAfQozzh/RICp9BLIrBPZCw9y3Lx7zlXiEp2KHJAhaHZNoCItw2xS51CCbFH1Ok+l
bfCCQRSvkEQddb2Wx27RitBZVM7tz4bX2rmYPCdAFHPHikMfY0ciw+HTeSo9eybPoj5BzsUiBOMr
VAH12QxEzdoZxfTc9adXWWOPYTJAX//b+zMTQypxeHkQNP1Yz6I8GPOjnhZz/FXJTjHZ1DafV52j
ffOTP3wHLViJbdpBhjqk6OP06jhVzPGcwLrSrdmKxQVLFFaOBPs7wfcJsxsv9/nvR+Dcg1zG/f29
k2GTOhucwESHlDcgd3ukpTMIAaRiVOc5vhM+XJFacLayYgw8CFqbjqXPa+zyq0CPAnHGxcRmj8p6
ouZiCgwvE9NLgb0sG/cV8JQSYNPco60ZJT/XjNOlzR/AaSmbgBgEXFa59g1fE0KJTxIwJp1EKcWN
JtcVIin8Z3zTyzfqODR5977yMkxpkEEdkQIE4r9aoCB1+qhCqq36ufghNX/Rii6kiPW2JR2VbRTc
mkXjUWW4Gg8uF0AMCj6uvnrqnXTcC4Y76Cs7TFZwX5IWIfkZ1WqqPfmHKLNxqn977x8OlV99jrDN
UgmAfc4egzgRbsyb17I4q1bX4/AmoiiWkwbDKNJG7ovUk2CQhVgzlIs5sX+wyTcB3NeoXC4P8jaS
hfgpt/p3d6VlRSU6x0dNXq9HunlsnSM7RpnxNgj++KGEbQR5YifUVuQkirfsh8csK8YgXkBvacQ/
7BwI8tiTOggbj8vSdywVEHCIyLkwNAQN2j5HyDI4lF/JQYmGY2hdBAvvCbHXNKVwIJGxOf9Ka+7E
gGjxyvVENc0GUsLfj+DIJOtRZ5SG8T8LHcM6+Mj0wjMjfgxqMAAtnNxtGOmSvfNMdzwIdVCHwnwR
jX22sQw73m+aiGrUgWH8tqriJi2rw7gZG78dnJIx3821nW17dVD/88UpfIrISX0P+NTTEZp0llpi
ETIr4qFlALF1xNcuSrY217cPgEY2or5MUPzHq6328xN4BcQ+um40erdzFbjUbjJTJYSf8rPnq6N9
ikIMswuudeWs2YRLsk/HRhQ2EUPLqNscTWu7fNjEsUcaGoeOnwY+3Np62ZqETp0NsFEzmOgxOby9
Haqs7drhU8cf4UynxfzmboVDxpB5IK24jhmT5pP2V7IX6qaC77lesmCKQK9DTxJh1aCmPS1tDHrW
JH6AdRR3uBmfvw1LxbH4+7oPUeyEebcRZVIpoMRAkWO2k7sA9CvSXyH8Sj0m9bqSdu0oT5/MuGsv
rENJnaRcHSVSE/0r+IFqRkVrMJNBqxNA9n9shuLhb8hA7MrmTR1XyqzvopxedKBd402yangJd0SP
bYJxp59umScVwSn7sQHmz/SJG3TrzfySj05LXeQqQjOkA+3waNFGlhN/oC8IoGU9yYk4jupHQoFD
AnMk57uij2FOC4bQdw4rJQd2mzCozPQ2bBUGMunCM4KRiC2F4tPIumyA5nmdChNd8GC9hT9cuQZl
HcvEovXzJdCIb6d6OODR/966mA54krcfFa/PblJwlFazfzSXwRHo/x2tn2r+fdn75DIdY/R82Baf
28ONG37p9nuNAuM0SVveFmZjIg5WywmcyNVysH6kAMeeoIf1Va0+vfcy1vP8pNUQh73Q3hh5bMLW
LwADM+Oju/XYTFJsLOPEFwHkaQw2RosiDsNirBM7J+Y8tjBq6NuTAgJgd29Fi62gWYEnDNpM+5Bh
d8UfIGBcELTkrC3vdmiHvvkV6TCZIfVEX8g57CxsUnnc4/Qil7Wa9CqtFGJFQ0ZAG+qYw709FiVK
miaSIvqLiDT4vOpNvh7OD3coVZXhRidieIwjobGWDRfnw4vckdQ2qSo8fzYiQRu/ABCJf2RDfrep
tQVBFGf2BF3//Ch/dExYNhAZPEqh/3nLwdmqpZvud1d7knhoixlXFq2uIKLyPP/24/2l62+pbeXu
gXfcRQY8oxsRk4IiICsvlaxZSiTAuGeFqhKKQKdHpVnsvbePl7o2wdK1xRP+JxUxom206h/vt3J2
shE27EOvHvykMi4P/vkpgkhqU/1/C4+wCUbd3AXkZlcLtSO7P2TU0+UI7fs1FCwC5JNArN49aYRH
gT0Fll57KRFN5V2W54jZOHyKrqKenOaoqHpKimU3nC/2TVAPEJN7OF78DDEW/ECNrYdwBgz1HppN
3YdgsS0+EP0yDbHB3I5wKaac79a/7MKaLbZihUCB1TkW+/q9Hlg9fqQ78XHeEWqRukti/9ybDjq4
lsa0SFveHQ5UCl1RL37gL0QfWSwCbEJTKBdfiXzB07j+1GRVReIg//3gf4jr8LjSc9ek3MsLtXH5
fxo5AnpuyJU260kt/H9gnPe1F3zNasE3MZu8M0uYqTevF2Pz795t077oxuHeryscpYsdwZKGob3u
/0PfGlOgqJsPV7/isgkHvQU7ERHZdyGNwaGgpvTHFR9xJn6YTSZkVlQUgdVTK+hBzRZZBI+6pQnO
gIKarAbWpj0/emIcewCL5WuDN/kDyqmA+8oqkBqp5MhUlQrPV/95578HsCD1bU6yyAZArxLfeKdX
ZhiiMKPAEg7dgd2sQd7hqhVHfLjZpwnDu0HrCG4DfHku3Fi0fdkMhFktcLgkTkNzxB7Ob3EpIlNT
M045m1OWS/Q3F3FuGNwONNb40RJFEqQJqUQtVIVcR09CUE+210BqkKeYCHDC33Sdc0MG2PXAzo0Z
LeBlwyWHMfjvOVZuAxj+GaobVQITrL/Krn10F0BhXvnatCdeBdOyxCFWD3CWdnDFzIPB9CNTt048
6WodsimoEnpJ/DW/4Qh6bE6ze9pGGiUW+eDORimbbSi80dp4UzispngHVHWBuCCnnktedStNdyAT
d4oyBkwMFoaRncSYRpSVOUUnD74tdf+BuRRwO6yWfSw5Wdh9RCzFKnxDOiIiJczoVoEdNxvtad0z
1JiIrdG3r2WrFMiUejRGX0oegXCiRauAD/ZIppKbAheOIgWU7pk0OdbGbgc5WVVLXCI5nOSX69HB
6qRqMcrAFl2baeYnOhgT9jGsOPtMF1HwKv6L3WBFDZJ/M9qBECh1Ltz5B9sMDurVPX7JGkdBdss2
x4nefZS47PjWzJLs669cnKaIMJJMT+elvrTGjDU/lBGcPBK295Ibx65RAsstyApVV6cwCPGI7KFV
6V81N0jiXlHW70AzLGBGlZrhPip3pjdcTwpGu3RTmvoiSgeehK+diXRAEHsLXrg7RQkEHebpTS2D
yjXzilVOhyZSSpzOf+F14jmel/5BK7qr0doP4RfaijazgMsS8ArzWF85WTUxnorwToNLwHXTaMPt
rXUBNPzA9xf17oBc8o/jDykXVCNRSrVSgAB+5ACY7y8BTv9ctoQxF23Syc6cnhLv+AsTv5xqr9DX
JNDL9EKMfMg+ngKCHcC0iLW84EYvRCOJ88Tbi+SInM9nLDTJlunymvFYdjk5+3RGUMPGaouXQSu3
nTeBCx4ZN/ANeJLti/6aW8pSucHLnXkzAabd0X8uT0jrzZ1wB1AyBK9rmW5SDbr6DRbag7zx6ALR
KfbI5944H4wx7PiNFMM3TRjIIrUSLEKGb0cKUNmVaPZV2mSr5ov645TiUF7FRCCsfZlavlfbrAGU
MmwV2SOe9Fi7UcL6xpZQzSi2af9W3zMakuh5vL1Xo6aS6SiFMD3uBZdizxLiHx9bL6HjWJZqe1y/
UcwHDJYkLO1dZp5UnQVeYVxDAAqrcVzg5/UFXAwJG08NFxtYOHsv+3BLHfYQLMsBzCrQw8POPXKK
gLX52bNpJphVPITdUKaVdmHJ8sJyLWnzyPz+nKFGgGpfAWjblADGSxMuXl/o06NR4XZ9DBjGAXfl
gAEU9MQIO4IyL/Mnh2sHloQk22HzZK4jb6xVCbaDe8Cp8jcvL+l+LQRKRU2JfVl9CgYQ7GbA8tNP
oqGUFyuvFIpSDIsVATljgXijr5InmX042nlsRSOnEN1dO3D+sH3dc7t3R2E1ruk0AVL/YNtMKFqq
m04GxbWiS5bZBTSQAduu2My1EpWxAJ5erttu1ml2Eg8nnkb6R6rSSnOmwMKSa5nSeb0cQH42DUgN
k6AMP3jjkrabUzlKajUocEW44jq57e6HiznzvwKqZV6fcbG0jrbLLAtZBlk6nFbxmfLGZpoGJQBw
p2sGkHY4qnGUFBvJoTw7lhnI1hmDqMpHOiJ1I8IQzn71QMJyptn9eUdVp0OziMgxFHgWioZCXaSn
95xqWPtaJtJTdPi1dQjUAGpN/9PhFw4QKOxafri0+AoYvyvM+Fv1Y55N6DYI0RMg9cB1scnPciV7
L3Bwsh6kShvz6HQK8rav+fQzOj/fuV/Qs1lypdTBYqBR18BCS7LAmB5Ski4s50zutG2DNUWXhI5o
Lq7XpikuwgXDrF7nPnHsXvsQVKavMpWFXviLEOSpMEfpTO92A0bDgA78Fqs8JXptrs/KEnibR8cL
3y9LsUMjCprp2bfjUL1snAoJ7ne8KhsbgRx+pPO49KDQV48n1reujR7pPcMQ24jIOa5eOStqBDZg
9Mjs6KxVGdlsy+pJV9qVIIWnxReIiD0qg3y1EDDrMZcd5tDjfaMqj7/BbhaGsJw2qRn7BwVv7a8r
ZoYGnbypfKR15du1T36GZsyir+F+GbmybAY6NnZc+zLRph16zffeb9wac0jCNjbZNkJUf23ZH/lf
iYrQyGSSPg9TK+f0uxSzS3APsP7Azxu8RmNCt/AW0/Iq5yTUEGBnVsyRn9iFtB4Coh5LZwTZvmDu
IgtHhOlaEhhmYa8cmjTU8RxMySa2aUY7UUmqNiTWNmqNos5C/sc3zG01CPFVXLt1zwqI4G4YHWcW
5tDU2SGbeKdqV49OujgKMmx6DkLDf5Khkkuj4WkG9xi8KH7u+WHqV8GLg42V0Si00w4nbDDkpXKu
GxXM4mcItG7dmbtoDHt6zb8tPmzRZJr2+DCyZk8WIuNhS4I54zxb8BAN5hpQBMvarMj8vW9Swflo
vVma/88ewgOgxiHwolcaSausXZ6fJm9S0D3Wff1soz0IjM1tlJKztnfq0IHBjwAuqjzjtygXsSmR
+b59bYXNRYIljDz07dh6qhYKDRxwoPwfe7ZB/HjZ1fEVgFqOZxj83243z2i0pgSce3ZAOCFZZ5BK
NwCo4oioKm62B+Bcd+suXUQ2Jh4YaiH2dQuEd+zhPoHdit6fiEJsHcvggwc8rWNjs/a9CZ5aDU4F
YSxNaAcmKjProSu39Myzmc9OATx4PzsmtPFaTSjnYWr9EKYixezq4E82QPeURsnicsUYWVoN3S2a
NGrr+5BJ/0oinDp3yuM2YnXPrswnnKQ9+UGlb5zc4HyDy0v8RlT4ntI4Js4/soG3VPQTK0Ev/Ayn
IWY+n94LkSnGRRX0GryQEYvLcQe5JBp8QKuvLGr42zQOVJ71pXWffgDjgqi1qXfaKngztcjVvBI3
tQ4pMgedy9tPI+TDQ1TiVgHUg1upD9mnhfAyXXDxhRqGCVIYxpFdkIdmM/JtaK9JoY3ZVgeFs5pn
UqlIG80TwA+nD6VkfWQMJ/VRic0ZyeZbCKX7JpKWTgJPbdB1nfnfAJtVH/xoVizN4BYQhWjyhZsv
bCMEo8bHU5V4tJxWPWUGPfsQ89rtfbHbkxskp37H9cu3lQ3+ZIDny96nEmq7xDOA6k7BFd1QMMIc
XugdW4lunfx4437c/bkFFycoTHKWry+2Le5yyYJGF4+/fdl3Jk4ql+h5YfVQqXHbJ19SuhNvvJ/S
aICXDcMcqebHwaj8WF7YwPdOQR/pFAM7IVMuzaVOaWLVMR0RC00M7s4ERDpPnhmkTVUv1ruGbABz
ScFynFtWOeTbyPZYJKAG9zmh+zwIz72AKgkxyKssFuT/8u4qmEDGZzBG9uULSQCxdBqQjXk4d54R
IHV9oxIbOEbNa3jlAfVeo3m6bSNJauSQqHk8G3uf3wTkngdj7/yD1Do4Nc3BMaCob+KW58RZNVrE
524L1KToT/mF01HpW0RAV723DpDjSzciOC7hwEQP3CKxeQwo2DwiIFEkxUsof9cRKLDtSdZCGyHU
gaTvEn24ekLr9jtbU1f29v5PzAlz/s7w0tl8/i+qOolo5KKAxD/7AQVYpJPy6b1Y3eopLRqiNqju
so8ar9R98/RsGQ5pQdemsi0EItiuGLBuwBzxp7wy0tc73nsraZ9//MnpW3T2JSebrFBJ2Jc+TFt+
A2C+HfGANYj1AGy1ER+Nem6FlJkukNkDtYFqPUFsdLtifXYwy+mvvmlqiEcaCzda7f+uTr649avC
YfUZhE74lHYtG92rLeJYnsYTVBWgopL6CwmdpxoZPJuEbx6DN4U5q7WhwMhPb04OfOMDUW5oHNxT
rZh7j9wmjmKzY8zkMUFlLNarxBu0lTKN6XtqkfWBx++iuqNDHEEzYWuZp+SVtHmwO9VxOZ3U5JxF
kzID59AhSezzpddJlLB0lW08kfn6zbEgxgWmfAHf4f+g7aPYFMNSSHVTu5i3//owaRfuA/H50Uf2
nh4LHVuW2L5PWxlaziUphY4GVWbzM2NGzObF7iSS+4yMbTtmLuSGLbOncwOR8ro9pq/HSaXSJhKj
jkb6CPFvEvR7P2kLgMWqJqMLzeVE+Lco/dgNWAoKuulkDVCLIsOBIYOJsCijXs3aZxn0W2kiumNn
KsFOXBmu7uKHDShAU5VJpqPxoj1m6g7uc71QyRGhTXqxGh74MEr4Cg4VawMZXdBp4fhdjEVUNnMI
gVIjypWw3dA8fjf5F+aVpZNhYne73qw0muHKrwOK/sXZxUVnuNdh9a0ch8X3KyJ0bOoqV6oDoopT
5ZAexWWHdN4/2vhnQ7G6ZgHs/OO2Xh7d2WQ0S5NwsULeUH/RU//T9QSXMnKCYB/LCme9XrTfm4v/
3r7DV+q6CyUOtLNTq8PgOks2MrVA2oLNOuIG3fCn6tNfs1YsTUxHZ5nOm22saySnp4+YR6nKummi
MUSIpvdCmOkbrlfQ3yXIAS2w8otBcI//C7tGmZ4VFDXfxOhYFfCewFqEAiIPd43YUYvS4FQJWk8J
cGx5pq/1agZ2VdfLxogdSDCMAyY+SR8DYNRZ4xHcHXVFWDyDWKD9ENvlmNZofu3gbdaduG10kAri
GHoM937UrrvdA0ZzW4ekmMemFKUZjKM+i/B/WCHmz65+80f8i11v7Wu80mOdAYgJ1tpc5ejv5GuL
40gIRqD3zUJHgyjBjCSd6A0/rIRhWeTsrO23EzQtha3E8AdJf6KN3zo2bQWKF5zteaiyfGa4vBtE
VMw/Gm3f8TkIUFRuKtSwORc8P49d3S+uAz+5BK83p9v7IZDUdlth1ljTXgGHJjTOSUfHFePM7G/s
t5tuahZzXMZVYv5VftNxT/sCBRJMhpMAb6HEQeyX3czy4aM9HJyY6WMnwsG43SydKGf2IgsUvwu2
MWZ5IZBD/WaPmO1JDD73vDo0nXl2MXFdqOau+j5Xuc4fWnKVBNBwM3DYcZxNprU9dhjvsuem7xw6
WcRX3L7LvWfZW9WWHClESukBAmH+v6MVopmBmsDgUMHxo+n4r/LnyTKgsnrS/5zFvhufHrcXScSY
/so6lQ8qsFveySu8B0AQtLDuVxB9ys7FzUzELryMa81aYDpPcEajTAf0xtJMlfB0ZY04Y9q5DY2J
w/j6p1fEaHCq5tiXDNwNUbY99NLv9vDvbXPBbfAC9mOp5SWMmSRaw8lLg9xywBMhsW0H3eCaGZvH
hAmUUqrHl3Frl4M8oU69MZE/7NarOUP+GtNPO1WKHZPPqOdRAuJdw33ehSIarMe18OIfMRpsLFbY
vKhG3tdc9/83qS6kHaasTAOaluiwtr/XpcczmudBa91eJp2nmAOYOnB42YmSydidRFKAjte1lOfw
/EDmGPYeRg4S/AgRUHPygkfsSjMDRs4/uaGdc+B1u5CuKIPCHEDmRea/4+cLsvmR4H5h+tY6ptvH
wyGnrdZUP1MR4CYxQRYypQ0uPu3/OzKGG5Z2+ck0b58YMsViTNuKs/Ay9YEa7C4eODjsjB/MPaqG
9jMV9RWv3x5QlYmiUwAp8s0g554QZqKrpl+ywUMjuxZJC9YEliTEmUZw2n9fvcrpL0GNb7YOkKGc
423uoKM3KQxaA24xN5vmjCCcNKwZCCVK7zAUVI6tbEEF3STrY71HbdQxViUqC+TiCOMR1sGUXBev
YgTpt8dXv/HYpnqnr/u8XwESEoVwyf+ndfZ07IvIsUukdwQLQOjmIAftqquJbHceoMkyybEqNuwt
auVF8VpdUhgmE28ClP1tS9uQimGF00i49AAUSeU55plHiluSDLzuAjM9B9zqgH0mdbngVrNBCTvl
uEzhgeS1YzqdKBEn3nPpc+wKVrZBaCiQfC35SSykrYObIulbT6XvwbTbLZ+ApOkFrM9ub97rY/YS
rFpnp3pMsZGOkqjMlUhu/4WR+RnKgRopsza7E3EDeGgUsYd9NMY7XiWny5M8+z1wz+s0LH4igNfW
vpHoZsAYjkxpZwKUQihghZGCdh+Njnx1/2yP9/CnQ6m5g5+cCXIL3usVFM+TbAqGmFLT05aIUZz6
iJmrSLDcpX4SmwjO0C4VN5ixiyDUZfYXcXwxo2It8UzVYYmnvKCtDKXEEKQiMiFxZmPa4Y7QJqU2
gj0IKKZ8vcgFDIdTRJnFzouz4sjNohP0FZrUqfUG8nz3s6QiBMNDcj1JdBxOdPZHIDBrEm7RShOs
bvDi2PNc3gRHEjyEHQwSPdxPqQ49wziLYWAO51xVsT5WFgVxcch2/5xuF28+FVjv8fNGrbTDD5fa
9hwMa6l5pxO2WRLAvjmCetDE0+cBHm7zsI5bgPqu4QqBljMvSKReWrtYh28RpMFP189cZxE2n6FY
pCBv4uMnHxodgsgRNWeghy+13/H3MQp1K4LFPyY9IwHo+YKZ0stjCdZYF53HGWwgCjE68DKOlfpf
SYhYaYw21IGoG+IkTiNGoo1ljPR1+zF7fNmu6ZpZw3XirT62P1zpX6cNiy9ufLsVE3ZDUpK6BDmJ
DFJJ4Idi4aW/L+OfGtd7nxQvn5Cskr0LuulYxJY2kmV+i+Ob0oQ6WoJgHzVOYLUeAjLsXNH+DCsY
ZT3Qwkl9kH8+hWHVbcmAOaQdxgXvFru6hbx+YvODq3+E7u/HKnoyVdqmbJzXnHLuFN1YsdqBUNdi
eN13QQ4PVjAKRj7kf+UzMm6ogUIZkeVagTVgl4P595K5d/ryI3E9dyGZ4MHxRzXySCtQ9VhwoSTS
Csf9D3sgZ3OsrqtoPoKYf12JSYhHVrGiXL6aTPDqu/KVNJDQnnabQa79pFObO4w7nhYBpPUiY864
7TXb+Jka2+4u6rfkx3pqrlOxTqMD9JjQ7tUnFn3mknYNv6Q1THLaPvs5FQIo6GJiq8fMMR4UReMZ
KrP5uSQvwv1/C2cLI3KENWRUuoIjmI0CtmK3PncFnKLYki7DYdkfWTGjQp2nsEpG5+niyqYiKkCQ
IQAN5MppbsjPiqwyxIwgqyQcIabiNW6gOfSG3I6B7fUEDYF8AHcMqhg20av6v2QiV0tsk20cREZR
/D7iosKOVr2S+EKFw7+a+qhAWdZn+a9iTMQId05wAd0RZU13gjfAw4Y4R+oe5jS38YUwPEWfdG/y
aLdYv0NA4qxGC1Y9jUUwAvXFV+/pZaPI4VuOI3CiqyacLlNjH5Fo/hCLIqWol4A2bCvRg6OTJtvk
oewffH10Low1Z9KK4as+JpsnJqKA2WYhZfWCtp2Ge1oPyR+W3QuO6JU/3hT/5Ltkj3A7LmVPEiNi
TW4YKA5zsloUE0TqWUSSbcTG+0PGffswZpli6lFMHPN/c5OYaM0NJRHTEUoQgu4a9pxxCHCzk6V+
P97md9FzhWRwgocxupxGmKQRPEAVfIjbhZk90uYz3Cmbif17yniTmQXuTviQCWcoW8R3NwImUYw5
9y2lXOVF4S5Sq1ARL7M7CM+BwdE8CM1OTn2ikt3xlfVImQv/IB1BqBvJNOBkwuRFAfOw+baUkyLS
Tty7+KlCxXU5gteCWrcFn75GO7XMqNG7sobWK+ObOmnYiUshwpn0PhpzngzUg2BP+Lk7zikGv3cO
a6otUcE0l0KynSCGTbafmMIBUQWAy5uLTaL6+TqHrzjjfrCYdUbuqY60pm23oqZ/92daX3+reUD6
qtgDscYXJHW/FY5z2k3hgM9S9ZQ0wRhnlEWbziyMfefWt3+0cJTobd0ZmSWKkI1QYYhS7PBAq6iw
wmoDOE0+YLOXWrBWtNc3/mibwJtv++EoJ3VmtVZUAVRV5rMwbOs2w3CX+Gdnjl9ZzfxqiAevTkBU
q3jmnvTo6LT5G4Sln4xPpdh/LmyHmAMEF/eAGnrYmlmtQ/zjjPEjUUPVPCgnNzGkI+2Fsgxpinz/
OGzYZ56HPSAqpEWM8zWNs0DOB1wui8imUwCqa0RbTjj1QQt/YJH96zawIRpj8uFy3JtvjP9DWU2t
vrRpokv/op6X8IXLqYegpk/ve5KsKtTZ6DvXAqZWbu1KBrLOxdiJUo10BKOZAp93SnX8CRjb7hp1
S6xE1LHUNZLMKQCRtGpRIZDvDAaVE6lBpVakoT9hPyE7BsNNLUm8WwOlj742BkF8W787Dr2kk1fj
ngmaU2rjp4qgF6qGBxgc4Nx5DYJm3T+7v0ohfnZP4ZThLfnK6asUqLJNv5Ls29hkVGSYuaR/6i8Z
XTAkV8EmakhmU2F2VyKHs5ptVN1hgmDCp2WgLWH4xa0gHamCxueuhAPw0qupUNU8K04sYP52pdyC
wfopMvu9eJz3dmfUZEqtBlN7uh8oh5xyjywmWpLmNpT4FGeS5EA7OwFzw8vmqcDwmrBbMmXCla9j
5IfbNLJNcdOm9wLuC8c+484uFhRjafAybvknwsEHKQsdvkw1PxuDaNIRXvNDJZGbB++isnOLqImx
41BxKyI4/de4x8ze6hcQmzpSzc/xbpj+IC35l7KCASZuQevYdDAosKorcDAi6vEr9k5yOQqDF4xf
eJHZjyOv+C0JdJko0vdx6SN42Co5yBsRkDbj9Evh6bTy8ERE9QJtDexyEPnL0wM+PLxpH37Cm/0I
KCuIES3HCYf3pvS8Du5T9WXmzLe/8NtnZUxxDuawymWnaRJDY6tJWkQ66vqyqwAO8fvRWBniDfwf
hH/m082DP+NfU4S0OWHfCS4nN3so8b6QP0O04zvP5OTRk08bbfKgG8hFF5SGeZreM2i1E1YfhGSn
MRs4gymgRvLp22I5sV/AdTvX8gF08NjKFFFOJMnKQ3oa8Fl1ATKPoTYQfqNT7aXGj95EAsrUFzp3
oRCKHWXebghPu+5oAjUDRiO7KgOOdypUlop2eXj52eBkKltFEhxMm7eBNi7dkvwr/2S5Yti7kx2q
bt7DK3MnkgiLruzDL+TkuWteo+BQWdosZ8wwxEL4C+qgmmAouCb5/jDmF/VAIJX4tx9Wz07Iy2LM
fSuIiQJwhn0JK9m96e7S+ETEba8ahOllFNlLqfzoGHy2pEg4PQU3OyQjllUJwRpIQtfdWdjAQcWW
qD3K7c+tecqDn5CXPEvKOlE7o8jUmmD7c3E3Q5C87GrtL1vW7IpXS2w4kiGhiGTZspU9LOz1lRbZ
EJvHhAu5BdXuYS0NZIRLoX4qyY9Co8pE62Vz/vO0Pnjd9xLgM6zi4mp3pu+zEhIKdwd2F1lUSqAB
P4dX5IPYLDlXE2Z7k8q8Loy8rlcH5mxsAu7ye0CFOVD8SYEQ0KM80h5vgQcBvPS7T/wXZJwa2gxl
sll2fgCFATOmWx9cUsnTnZKzU4VjFrWm42dmvhVMVM6eW9emw+uilmsTGkp1EPg1rHVeeOsOV0Lh
28CuzcBSL3e2MHdDsnobdIeIdCkQPe3sNAcFsddZX7yPJ3t3aSFgX9b/8aSfof6ddJ600bPu/Y0K
K++y/JLZfvk7w3VqmX0xy9Y3YaDojZrcdcOaDTGHUFXWZZFB+giBxWE1Am9yeHtPHK4LMk1NdTTL
Gs97GqTCvJiS3MijtbCzKlSiLZMa2j/aa1NGugEI3rYgs5OfcURuSvjfxZGbm7HYzCeOzd0cN5BE
hyv67PnwOXtBNzktAlxRgsqMCwTvLZcZfjrJWmlgkrmS6ufS4PPXE7a1Ldg8Dj+9hy5VlJ7BC7dK
MwbcEXni2kprflpaH8vreAt6Fa9EPcseb/ZmHZdtvGMADVBG2mA3T+qjACKmrO4dBRfc8rLwtV26
vPPzm4ukb617KA08K6bzms+bC+bIkSN0Htcqynze3JttPL2t0Msp1/R3zCRtE2fb3wHhBPoM4qjE
gOZb79+Sy3o5mxslJjJDIVUlTXZdllc13WUna+7pG/HhAk89EuVIlkjKMKa2xxKdA6r7QRxcdHOq
a2ndpN8H6O9xGjtOwfupDjSfXVc8TbRNtvUP0T8bClDHyTCvVYjcXtEg2JZ2asyXLLZzOVy6J+fi
Nbz8TH8k+k3aFzFDnWSwj5i4ISymJWTXebH7Ozh3/nRmNeR8HZEtRd92yXyKv0f6QzgfAqyaAKli
qJg9ioZbwbXmNDfrBRZciZbW4KUtysIgZzM64kAuyWuQMSCiHa7IYTO5DW7waVp3Swz2Z7M+aInf
UV0UbYIoRt0f+3LMleZg0H+apMfU7ksdIuQCQ4iSk+bNIDSUoXtitay2GCMMVHUegSUrHPQrd8Fz
sRtxx2yV5fkFX0AfhinNINmG35ChEFwOJeiIlVhq9pJ377OLRSWyfQ5vWWfihkzKXxfrMLbMK/ml
nzp+a0ebD2pQx+jkZN8xzAcC3mLi1PxgV+dSjHNFraILnh6hc/AoGbp1ZwkOPdWBBnpAbnAuxeIP
nJQowYkuFxXItD0SDwoYPPyF5rEmWXRExjdgCtmI5ZGw42+zBJCK1qXzr2Bmgy5GMzAs6jGwtdSD
o+NDMYbMPU1ngE1kVjziXQt8Tz6NPCtzlp2Giqx4+0O2IDim0LHurJid946JamyfP4xxJJo3jlOp
MDtDNPI1s9Ilytd/lIvksqkwnoxSQcqMWpw1H3oQ88ml/pbVl9aTeRQ2YUV9abws+w0Jhk0gfYG0
A6oT/y6X2HxBiegYLCykMwyEwKkYabMOJ6LVL1pDB9RV4jPYEkF0SKhEmh/iNk/OMvSIl6BZ+f+/
JycRaEcmdg4cUn9Sry8Wcm9FmeN2qmsdd4tlMZ1hVWMPYmkH+V9cbMYefGP1yIAJJF8hhRVI2jwl
RYt5JrKYtOMTXDk9AsfXwPhwPC+usvHQwraIkIWShNC+sT0B3QpOEH5NceUbDgdxML4uJlT5Pnh9
AS9ns8PlFmfQITRYw50dtnCTtLUCtMJm9inJqGLH8GzcAVsSttbrIDNMEBVc4l1kVU7bwtKkdC2Z
kbpWTF2Lj72jZb3IY3kKp8SMKbcxm25ckIwRiLvKJ9Favy7Jvf5TGBvBZ9AKAraBeyGQux+MEenK
oOJgStKevUwuuIFezkiBjetOfO8+u8eOIyqMjq2AYDy0mIhlXmFmcS9Cwld3ySrtQ424ZoRd157k
iwPcNfnts9D+S0RhqyWqv+LocXS9FchLGt64ZB1TwoC5j0L+gLorsAYPPZ5nkFDa042RIShcCroa
/kYWkEJoa1arF937/CupkHjo/H6W8WzmSUNGet9AvAWaHlHyGoxqhv1+IEj9L7XufkAizblf3Jez
PQQJsCZmT+kiPcLLLpxDe8F+wFDAZ+ToQXQ7HPkMC8NHh5D2XgV91TwTqBZo/87wUpNdkHD8F458
uoQ3VoJXnLNVaRW14Oyt11HY3uHxXcz6aEs1Xb19Yci5ZOAN5UhHcfDgF1+9Rz2WsmDgW7kfQ+cQ
cgW8J1iBnjrG3srSSJl4S7SO2jyPfkyXQ0G6cxWhxHRr19flT3wHSC5VQx+9J1Vmpeuwp/EW0GJ6
/tt3mleJP3tt2/X6yWjqL7uiizAMrKJexQg5Y1p6b6gimu56lLoP46dBhlFb2Dxx1TyHLEt5g/Xu
3na9kulsbxF9F7eLaQ2wQf8143kQbdxlFrpL3TFBNXlaYhGKHBVwl6a1ViQ/K1zwsDwaNopnGiEF
AznXX9KbByiP2WFrYmtIKMqY6OVZryQNN9Z+zNiScyQ/YPFzwrAzp3BeN1sTle8OFdLDRCD9/4RF
SIRkSctu6EZP5Pv+kWDZ0hseHeTTnTRvHYmpUKK6rZ5/xDRh8RV7BJbQ8gMp2DDCQiYCFFpIlQR+
QPPygX4G1Jzaze5y+/vwECG8IpfZIHRsnWtVtoPj9lRcKIhJ0J4/UFZiS7C+0tnFV3DVStwVEULu
CeUrNZxpr59KeAEgm6g2AYD7NyYYfa7PczwIVX3HfejmCCWizNz17m+AHCNsmaQuisiNJVVBr5Vv
BptrdBWqrhd6yuF0fZxlbCZFa9ILWvcezLRaJ+8nqPsu7BUw0ONRzwsPByHoVs/6ckCE6NpdzA//
3aQhJLizL6M7fhQ4Gl7wN/rflC+jP7NJTsOQilBBV4xbpSsFtdWMRoZ1S74sIq24ws21UJFR2OT6
nK/oo3NAy1hlDoxqc5j4Z3NcLHMmhtE4FY2+nBYUjk2piQd8D4LWjMz1P/gjlTlZUZjVqTglFE3/
se+MZgYNvteWfpilx5xJDYJv0Q+TklHljflZO5spiji2fi/eBhdsUvRrYHDZYEfYJ8w27F5yMfuv
Di6P9kkYagSUnDqjH5cRnUPyoEDkxh6iNOfVmqF6ceDSrAbpJtLJNdigj0snNTFBr+Diaw2so/Re
TV/m6xnMpx0Bl9TosO0m7RnDqWoniATxPcbdLpWpSkUGUxPO7bs746WZrkH+yr7Qfh55Tfqyu26c
WyvVksX99URqR4oaOGAL3Bu6z2h4kfMg+DWIap+BYFKyToDNqCCvPkHiYYpFPxuDfl1SVUcG77Hq
ztR3bzCpw+ePXblJ7to7Qiy/wFja4lvQO82i8aFpMxWmyMUeI64kwZtq08GhI2L84r1+kprmmFOR
3Fc6ZeSOuKWYbTy2auHfNFW1g6TDSqKTzswiQf/cxX8uH95ZPE3w5gmsf8gjq53KI3ztYMWlbN8o
nKcuOpEVO5lvOOxiOCuy6Cu8/ZFTg3hui6JkvrYgS6dyG4w8gHE0aCqfCW46lBHteLGijseX3x5C
97zn+WvlxKAFCxJtUB8NzH5H2EypiF6STlguBdJ0F2Q/gCFl8pEWY7DW2aEB+ES+3L44TTmVHTWB
oO8qhHRQjNHvyUb2L2h+yA/ngT3vkjGqz0SsA+l2RmuGh/I53bxlRwBwYm5KjC2lItwUVs1EC0YW
fAeyFg+TwCzEzakRBaNHJM5nJ9QMxAtzc4Uh5/ZhvwOfJl3S8NhM2m31ZcYuK6zslsdRGPwsi76E
yW/p16qdlBxolyTrMwn5B0O/K6DqN7ksVsxxtu1HJEHoWFd5ym1igUK00YCUgdHRalhEd51a/cGa
neQzfMSuVEcWznPmsswOE22bEI0iRg2K/ELn27rB0zXJSQBW1JSD8DKoYQO40lnyvWWDSngqdaY6
fyL1StdMYB33Ws07QVKGZuMWbOpSQsVVX1Vl/f4UaMyGRFhrE8m28OBSyuwbewMtJ+0ns0bKvxCQ
p0oxxhzWL0Nfw1xVfbkYiF5QlL0WBelZYEWaj7K3NmRfJPfEAieRS7XJKC+W5w84Vdp6Cfwxk7TH
EwxibN0azh5uftwPtf+U0XbruynRi0VqZBwhGjGM+SMEh/XRE4X3tNoboOfy8v/7cUbDWCcyGecB
Rfos5aH7lo9Hfe5P4hmWZFfXQACtb0CCW8h1jjhWUI5oym6PXR2y5jJN7ZlFRcSYv0Ef9iFrnVzi
J/B5VpoP1UwTPgztKDyyx+nVWyw4qQzV35EPj82+6tpaCQ9qatzHwKrZyZ18MTJ6Q5NFuaMyC+OU
kGO4/qzYaoJH/w0ISGKE8/38TmYSvc0JU1+IMYKtS1K8Fsg0oZQmX8gunTn/gdf6+ikyvdlnci60
3dMD3jrBYlBfBHCrtP8lL1KHAo8Q9BwF6fTi1a/uWespCiWsVhQkmHzdZneteNxji7Q8Sa/+6BiR
K3WrmowQH5wYvNyfUzVF65Iw01uM7bu14tVGKkJtDYADPi4QLiBWu3lpoy6ZjQXaiCXkyPfInRxc
l6CiBUuAXNXbvxDndfIcLozUWEXoiTijB6UvBP9aCjRNnfpUIKUifGNgsE5Alj8OmA6lanXU1Wip
P4sY9dLx1z7hUDl5Vve3MIPu2TPQiFTI1uNvWq7MWzptjhM22NT51lNq27qy/hXe0J23855+RjDo
3ADMc7U2xcfN3gh70qiCBAlUfQF3a1i65SViv6yMUs89ffw6KJW8U5AqmC7GYm9k7phXSGEnLSUF
9/gc8TktYG/o1CBW+98lbRkr5E3TlpBN9qJpB6cyoAcLaL/4zlO5ieWyAbqjWLVBVTi/QvsOMMWJ
vQqnca7pBVyf7xZSy2AXnWBCpy92A8OclGYN5azqEsRwYZe3GA8TQOK9Jq+U/QWOFTOmPABERgNb
tyXP2+5s4lsIeQlE0+Dk05VT1zCWPoTlRA88+uvJsW3Al37SOhdSQ0y+1vX6l4TV+PJi663h/Lb2
m4loNPsH1UqNF5sNCaOaQ0Uz//nWxAMqcBusDAgdhrWu2aKv2/dkZSAWnuqs1C4rFNA8ATHdscqO
EPahojIW5Fw9sClMevK3mSpD9p6/MOambscyIcQR7PLHephD1nn465C0qjIaMLB7pAJvqRnErxMk
dhk14k3dM/Eziv4qJih2UFEl8csCl+N0cnJPvDmzoqvZWFlNM6cbmkmHRENkaUdn9Z/la9QtyzRk
qT7Ux7FzYONzr7e0q99mNgqHK4LNXlIztTD0IHY8zo3kLlS4sKghow9zO+yEKvH7C9d8qQhMIHx3
kyU+rJAa4yaLEwE6UkdEGdvSlZ/uhubEzBHROXQUPB1zQm1V+mms5aW4tT3zaLcpyqVLXrlGcyR3
ot12KRlGTKfl7rD1uDP4tpBIhewY5Cgbx/w62Zmxv8Jl/zlUFhhF2m1RPdDiTnncEOzgPJYDyFJT
4ROV/edZ39fgqMS9FHM4fixAvfirlHIPKTCdBJaUlGUZTy3yXf+FhwZvwIrSUTLaoN3hQzV9O1qy
BDgOPXL/ZoByHfOtG3kOemewQvcWC/ZkFboj/IhXwr4MZdorevSJ4rpuCjM0h9hahrM5CQXEJdP9
rtTrki0pzKTSPhZIfnJJ+WBV8pOf7FfMK+fRB/APmEQoPxw3qm3l4Z7MYcHN4bfWFixB/zQ0Zves
GbU/cBcIVT5OxvMvk/0MHA99ejuJi6xklDgvdRo7p5jHhVWBAE3m0gHtfEW7CB9F3e9dp0QR6N1W
Z4ICm9g6Nvp5rvCUdnLgyY90a9m2WbEShYe4kLcR78ca4e4z5Py80xC+DnZGUSfSZ4cICG44nbLK
1eN/4cH9cXUuiSLEuQ69w7qi8TJG5FXjLTQq23vtJvs9td62wLr33cFRc2VxIMPzO3noyXy9vEdT
VD/aEUwn9qNlztXB+ynDw1ZYSVCUnJr833yxqwJeYpoC4TAsY+iYPDslcw+mahBUz/Jdf3DTPy8A
1o/RWuQKZbGZjYs315zbi3vzBLQtwopYyW8z3Jbn8GTUCpsm3VjP2UEf2ibxTalpIM0W2bB7nkxc
DOMfoxvcgTO41wZarv5W0UNyFI6PGuijDa0ZhX03Obp+jdUTMixFPLDI1HWCoDS0sk1HzwXzcBgV
e8BIsfF669BsLy7vAYv0Q1WAJWIi8Bjm4LCxsPVJP+1IMet34aQb3xgt4JHfRUQgfC3S//lsS3Nq
JvOzXtVmDG2AYHAW4hCwfaQdXi77ZACkOQ//Q4PjEOGLuoeTKPVrCMjJQdMjiIF3DNyldwpN29nc
0/XA21nUE1itc+EeQzMxH26D+aKTesfZ2lAix6BBZflgOyzMhcyxhtzLGuXMEcEROe6ICpHe2zjk
Uph9YxHJs27ypt+A9/g3y00Qn6e4742sqOZPJSTQmonM4D9apvZHDpqPK7d9zAremAIGipscLPSz
TUQpq7rkLvwqJVmIRIU2e/5ZLcvZD8Q7OUCTttjNfOsxo0mZ/AJYJ88x8mB982ggbL0GVXzRZB9D
A+WCHQiZmB7M5MqKZEtayff2bJ9JVBldI1sURwVcJYNyfTkSwzl3zjzRQGg4r/v0w2JKOVeCXIik
zeGb7XpFp3QxpiqJF5uILFM4vWGMLLRG7fANHykFKraWB52KFI2wUaRtwba4oogm3xYvVlzucSDd
bp+nkNbpydVwMJPIp5TTCffmmKUCUEyZ4qsvD9gl75ZICfvBSeHslKKi9eGDzgCg+HSzjLtASq/t
XUJzY2XmOVCarjhsFlGO3TG8PCS4scva3z/OhGfxI3B7pAeMVLIDUbTZtEg/9YseMWNm+m7BImOC
Y1VvD8Yg0GVRVeF/dfAOvkOTpFzmBhVXFwb23ZFcZdtN/dmYGJVBLHG5M6oFpgICWC4vJ/au34Qw
vi5FPry79re/nRM1Piz0mHuKaRg0ozuzotsUJcXZyEVRBIG6g5AqRtLxre5cM5Hrd1TxkeY6V6Jw
nOzXTcYdbibvKwye+nXvnDOe6BrywHUlRXaskyP1mLUUdZxQ8CvKG+DcgMPw09f2s0pfX7JSkS6/
tBQImaMxnJkNM8mrUkOKHY2SjKpMyHJiKcPlGyKwyX+m73T+FfvrensJq/dIrl8DWIWLMKD4AxnJ
iMRpdYcrRIS8VoJYqYCGvY9gsLgwErJpQ2GB6PPvHlREiHxyDijx8nr4aSiufTTIc40AK0d+4Q9i
ks+dg50lRjIVwB5LtwG7uHit1ECrBOXr0GfmFb2adApP6Rp59c1vfYEwiFGHSU6xh2BD6+fgERjs
UpLAFCVhALOwAEc1FxdWv7N5VUx/Cq0uuWq0YhAXaWnhSg6kraM0h0/EyMPuzTrBnAweOYIC8XNa
fCoRyy77QCO75v53vJUXzCj9Xq47gVMJ5znXCCkydDFy2V7AZUsAQGHa30VvizZheuapXuYmLY8/
F5iR04mpmzQJi7h0kTPfqsKD+cJVfsrB1ijuI4KLLNZwf/teue7aXKpy20wIH9bTGF+cNVNDRiAt
X5Aj2tn/qZoY54lWbm7TeDniCKMEMf1eq3Ylz7nZsm+Ii7edE3/UWML5CwmYMz2El4+Gfq7nT36i
GRwxnTQdXvHRDds0AEOlAxl0jE1nZtIs0JocqIwEvhNJ2p3QgGhvVCs+FmHb1hU2EzLp1z8opKyA
BccOcEtXLr+3ibpHNQ/JZS/TWOkTqC97NKcQWsRiEYzVyfTxCXW1fiuVXNNly76/1pRhsLg1TLSn
DiLrTdA7Zbo99ab55dzJ7g0Bm8lEA8u5qyDoUuLz0NbdvIngytvoANZvFaIoIxVy0Xn5m+ymvVbc
14ha2Zsp8uWa6ZjGnYsYPpq2uvbEzMGxxXFaSfbufphhIBCFxy6Ih6rISjxAI+akONqdCWeuxf0e
e/7Fc/U1OO0aO4KWg69F5llYIgfSU14+yXg9VoM0Evl4cRsmXKSeHvpplE9ufjLIL4IKkU9gdGGR
dw13SoGaCJPXPsOZkGBuDwBY/L9gBVs9Jf6uukla0l7llCV8JWPxkRZy7rBxeh2soP3eIpT1ZhQk
1DuSWHoDqAF2G62Hxwlg5wddcpj7Y5HSs0UqgLecueVwfuKXwyE25EK70NTM3mct2LknD2Omo/1o
5s2oHQYAKtJrjTPRYWhhwFKYZmzjNMhWNBXuvUGqMYeN4MOisXlz9nziSFxQ8VsEANVFKKB8EFtD
jgewPufYe8+iv/MUOJdEZyAA914XJcNC6RxY95UD28ms3ITtNGqH1iU25N4N/fh0j02dZ2TmXf5h
bwCeUZ8uRc6T+Qu9GWFRUXiOVE3RdnGVxv+0BxNx8b26yz7BLDQY42D2bL3HdHZar4p6AqIzE3Wt
oSi0WAkXh4I7Stbjd0Zl8SfI+j2sDO2hnEgAoAmKdJdSImEYqcrTFL1DilPSFJxceO+lfq43PXx2
chcGJoAXXttaUFCjXUY2l/jaW9yC0JLZosqBXrpOXwGduFsbBYSNGxC92crwnxp/XxdTIhPslDKr
hoSotZDAHYuKiGeU0QdseXb0T+rJVnHzb7k6iSJS/4KbkQwGC7+HIC7GExb9oV5uriY04N11r0fp
N3cwMvPafcp3GJfJTDQGxTBLal2ToMdQHcXM5gFDZffYHswfGSKX7II6JnzFC0ooGgyvQ+HejgSf
v3nsreIJOyTJtYoz9YKYYlFIxew5nWJalgQXs8IHIJ1DCsoSPhIHH5qV78voIsCi8k+Kx/XUiVbg
VMuwv0uSvxXMDi2WRLYZK2bA4YzYEddkRCwWdJb8og+/7fgXHL3EJyfInp5eWc53oT7Hn2q3HtyX
YjG2vEJJVNLaINNRrc1L5+8sZHuqGVmkDCZXaoBKNofsX8No9CJnWeo5bbjNzmujUbdAOH8QH4M/
Gz9zzF08sfbQxe0PHtOEeUlv0sBB8vNfSRRbGtN5rBsUjo73+tSgUdRnWeNlf8xEmZhtRtGZxcOA
LmwMkhfEPxk+/RebwnBIPstRLFReeMFW8TLazRZo+bSPsSClHoT9pDhNRjfNpChqrTQ1hIVyOSvp
JYpQMrJ85y4pZfApKVb6AfeoAMaM2vwnQPl2ZsKUkFFqnQ/lERue2kUTKA3WXFCFABXN22bzxfUu
lLz3kPo1ECjCg5JGM7ybF72TghWnPC1vuI2BCJXOO+zSu+GiqIXzOPA0MjWMIp2D8ZFT3wtFwsnk
ofc7droFsJWmTaXb5+RFosIY7ftGP994l1tAzXFJcyYMHkfcza6UwiZeqU6N8JP7z0/cYbMyXS/B
gEAHqLaO42Yt9ZvMjDjffOlXQ4PurUd9mO/K+2/MmMLkWuUb+/lFJBe3clfveP33ji5ckvlhD5ek
4Yez0dukBJKinyuXIhKsSprM2PfsEeKvNt8fb/J9YpJl12ysjz8vIsNLBSR2X3SfoxSipFyqw810
AkdqvqKoKhBZomkJJIRnUlUQlLUODQj8V+EP+zcjqZfkq55db3NcrC3SMLvwsFDhPUuwKyn2xW3R
mUgjoj8fRrmnLTKw/5u18oMpLZ5qZN3HD+HN5aVIN7TqZr/0qz9t8p8zawoXOGHAZduIaIq4vN8z
3qnrY2kA3ztyJeAwarXr3fTWNt5u2a5CmpV7usqwS3jQH95kI8LBPJlW5hysxbd+HITf7GAaAByz
7VVJ2oLUQTD+2zu48ch6D55uGYd0BMfVHcSTAjPvytanF8NwT5f0dYFxzkAvxzOaH9UZTETFv1v9
vF3unMb1uzdS5FFzncvg8mK6vtle5q5/PKE3nVoS9w/bYTQx+UO8x9lmqdFvSWTl7N1F1Q4aZndQ
foT1ksuPgyAHINNfjnIlKPRhMFHBH8WkS9uQYBEuCkyohTNEAZn7jIPsWci9aiPCGN+d102Jw2J7
VaLD3FJxVH9PD3f3CfB8SFU+OnnuOxulc0Y1VobpQaaDaI+4PXq0mIxxTfju8vkx6T+ZOU3T0XQB
NJPU1V01I8ywyQfyCEMgiL8mwlpXzmURKv8yUAXD2Qw8cUqFPdR+7fcGBTVD7A6uiJ3hJFNsPKxU
63NFiIZgdfDXkbzzvSlI9YDAu/btb8omlUi9dDNntu0aI30u7Bmi+Dw6hcexolgo+0A6/47lYUUz
rY0x8FqfhNJmCGYhYed+58XhyAhbtFOpJXo9CT1/fVQ2Cli/ovNj28TZsr6CtU1KlLMGI2TSgmO5
nrPq+7gDhttWBqBbpnuIE4+GSElxr7v0t2ZhSYxUBTA4dBtYDQiO9qsZ0rVGUFxJuK8EOVjAxsNa
DIxYRPHk2KApMhQsGBaLOj8iO0PSRzVR0e6q9FI+WbppL1kd2KOBcSI23sQaYagvBW2cUjAgUirQ
JjFqwwlFlRDUiZRlAgj+zJJ7ua/C672x8M38h2u9YN4OmOhIrFNA20jLhF+i7j6a7j0QIj1IkJAo
y07QCDCDFLTBwFNbbkNe+YLH4vkNSDiO2ws9xNYM0euhmSWtUqlWuChBDpZbu9q96ktUQ3/iGy5t
eoFg5tZf4z4oPqxu3XiOuEJMTcDsFrAcWWo2++BomAqKAffFMbt7VLYMjK4DbfGAIR4oyUAi42j2
7GUZ01LGnqHSR89eUUAGL5EnGVGxJ+vPt2W+T40rP15VLKfBFncT+jVeT4lN+0/Fr+MtIG06Zlm8
3P1I35TT19Exp+881NhME7Vm+DgkieJ9udgUgn/ImpPZlfM+xmiGxuLIaQWGxDm8DlBXNyvPb0Rf
V7Ackgn+XWej8CsdUid+fB4Zywxrp7Z0zGB/WOT/BNjv9zxgG/ydkjVOwdeZSaCMQVabKvSX552/
mvRCGA7z7dOUTGJw1sOjNJmP1ICFU6lMMtpECZsn7OAm2hGQLwguuKkLIBLkrADifbX+NEWBVESN
WMFM4QQhao7hOtbE2vY+LQG8+YdAOrsf64WL/FZ5tUMR9igux/TBxadqNWUD66ErevkIZ7tanzQK
N9pUueMnmC6B6FevfAYVQCrmV+3CPBmX/afRdOOC91MrFbLuUEIEYNeghfjNjGM2wUGX/jOc6fDg
a5eda9sjxx4+RvXbS/eqPye7iuSCGvYw1BZi3NhfiXmfEemhkPt4qORbjbgGVotW2UL2CzKIqYVQ
bKAo+cCtLmULsifmkALjR/XrgDRzye3KiH9roZdcXTEvpqolMmI7bXNy79hRF1zZ2p1FH6n2Vg1Q
C7UxgET16wDBgGRoE6ipUVIt3+bsDzj5IiNPZVAsDKyRzm4OGmG7+S9s4cyApBHFXysqY7zF/OYa
pzBflIvRxuqGsEKdKEqAZms35irXiunNhrARUt/W64s+5t/1cHaXidDp3OnvUtgOhwPLBHliWlms
JznPuDIZtjPXs9CN3IIefwTYLNqlslFVyBWnfglSdIIHdusIU235y0Limh9lqkKHN/H5Lbkfq9eo
X08/a8I/yP3rbN7snme0sHPTPxnEddku+WD/wlyOSNLckKgEHcqV08ojrFuT1lhjozsLA6ZRmXpd
VVZXGWBL8Hy4uJdzwkuVJ671z12cocDUM3ELvlYAfLFLUVJPwIn8BdCcyO9/YiQtxJ3mAS5krjgN
7hrRCUg4TX7+4O9BlTy8dSnZlLc5L8w8YxMnJUMNtpjqr7QGQ42VKcRCnxE1GIYU4yYScn7uYB1o
8X2PGIYesOoQe1wtfMCxqcz5h8lxPpBM03poxfx46IpZ9p7ZHSIV6zr1FDohoULFA00XhuhlsGez
nrAwOeaw8xJbN34ixJ+w0uPmTyKEpT4k+3PH4m0DBWTP4B1X5gqwoymnPqnylAl7MAWPCRgW1xHy
GgsPO2Pfkh1uRW4Cws7AvE9PYgeskjM26m75G350izjMnmMrJyTJNk1DJ3i2Bk8b8ZOWv2oS6F+m
rUc+MibsehCQ3bWGGlolTnlBjFWhKTbC6fk/vxwtOBCd5UwS/kUP8nVjAkzWF7TqS3AuOO9iKrLd
/I8W76C09MOmSuvyA+Ygfdco6QxtaDYxSV988v7tP41aJZGpOlb3H/DHMu/J37WhlKhFzdoEc4lE
jB5CVnXrd78Fy/RF1PFBsZYDpD8yuilmGZDdsqMobIHnoI9jRz9hXOSa0uao/tyj15SwsCjjnQ0P
B51L5hKx1F42NbhoXvvShefFuCEUBHwvoTj5rJrwI+hDbzqNXxDd6eAcoZuJeZZ7lQywgW4kheEN
phKdw6DvE5xQoK6mDFVw/ZD99h8Aj3pJIGd8XIeaM0YjmgmIolIELFFIejd/AGPUoY7heOhMIZWA
I/hyQbkgB7iqP2JYSoyb0Zz8igK031KV42uQBMcupXZQc650WbARfgY0DWvRUydlOCSX1dYQbqhd
sec3B52MSAcKIV0HP4O7XiulFvn0vT9jzg+WNKE3buSArvm+wO72VcPzHAZieUDtrOPeaScvkr5s
E5N75m/s2Qm7Z+GnhRtZ2rgdzwCHdgj2ziFdlkZuMQor+LQo+YrX0O6E3xx+ONWNgW30jPWEeaSi
E+Yyo9SOPvPHYTb79ncVXVGRrv79jb05uzWqsH9Fh86xrSPy046ja3Ihq67Wo7Jj6nownonh2Dpx
1IXB+NcN5rHwDnZwwU+8sBrzlPArZLLFIXrtepsAnIFn5jcllgUhIW8hDucqvewjYJ2CKT0shcfb
beGfIEmlJyAibsQ6hcp59hIZX5wEAX83muzycL4IKh2MG1zzGf0me3yYMMqkRSJBCXLazkyAB90T
njh9y2tu1bvsgWPw0G/4gjdLR+cb3aNHlp8sTtcwW6ErBxKI6psjnaTtHg6GhqYVRZ+2qhDu+T8t
NzmSMCYAL3phb20oAvD7Xf4taVKXZt40mCSFgM4LFpodalrixZkzlLuZ2TQ9FiHB24K2X6bbn/de
+yBgKhAcnWxcusGWbx/JTCLRXAI669vHfkTNEaYaZX6r0FE+hV6FLbnCj/pmyrA1xhehc7RlIoit
+0LrUYKclc8Q1DwuU/88YcDgYnQsdYrq+oVHSVG/FgHC+wgOyxgwhr5kaUEBDD48PTE4cForupcJ
EI2i4yeg2Uo3jSJBJw4HWh2ieilsHSE5mgZTdUrKPQ26mJuJsaho+2Itx10WkgnUaP2q+ZjqXBXH
oFzx1YQTm+Grtbcfx4YgDrKaGoHLihKIg0F3ZQcQVz+DVgq+S7ufmpYxsx/GceMwlJWvkRIWiqLw
pKvc+/AAw68drxAYJDXhZPt3OT+l3ejc33NnWcwYFsC50cKa/HzEoUMboIW8RbTOBm/OaONjOH9L
rb2oY+pnYCdCDLZNNaqr7sslvaKdESFk878Dqh9hqgmHQXoud0fd2Kir8JUyISWmFY3VK3K8XS0x
ElGpbykaoJF+Ege1ZZaPz07EdMaZaTXwzvs+YfzutVGyHaQVcPBRCaMkV2Js6cuz88UL5fbNOLgJ
cNchaAvCwIMtVPNjhBTdxCsWfgGnDpAo17dEq4M2RvRYskZT12OsPvmmsbuHiVZMrIOVMSwXxueb
bJlmN+P0yxEWf1lvpmX5k/PV+Y8GFzxHtUvci2ocd7q9g54JZi2XOTY35dV9N0u9wg+iFD3VKNWg
BZu00FMCNNwaxxTpTRgyRGCmG8szplbEEsrRRJJaolpZWZNfn390NflDuxOPX5O5snOGVD0XR94/
KVTzqO7Loc9C83Drqekp42w+/K4Aeo4WTx/8BQ2QWsGT3+AKXKwbGE1MpxOq+Za2KXuP+3oc96EH
IkL3mudHlXkWi1dWBDKkEWmgkJxPSQzhr/DKcAXvvAtisvx300OWqMO8hv1nzkyn+KKYmnNyYiV7
l6AfWSfsq8vYKw5vHok1trsJNn6dpGH9udvqQQ01BgL6glfpxUAR/epeP0MFiuBD1GzgzazFmzyk
+CILy4kJ0oQdP4gzjr4jeMO3c/VhNl95XYGqOdtYKt5+56iwb4EZqSp/3H07Fs8QXCa/xWM1SvM1
yGDw0ShPmJgplqX2DPiwhQG1CkL8jGd5KrrC5jrybVWm+v8xnld/t+Dq4FdgtbHG9Bt8fVD0uBad
6zbqybyB7H2WN5yHK8Orq76HLfVgt1ja75jf4wWBvE9IDkWp8EsQqJMFgpxhAgPI+7peL5mRe2m+
Npx5YKWf4wQ/rf0PWPiQRkT+ROxnazBy42kt1gdzcODYfJ9Jsy3XyUP9c8R/HavoBjS+rcObmF2b
LSxbTeelxyk4p49pGUCkZeOO1Aq6FUoHLf/KqUwgp6wC7bvaNEFz56zd60ECD4Qi4WLl720L8e84
Dg3hDiLZJDIEeWko8CVfv47qkadc+2V4qMVtJ7PZs1ySL/EjYY74KAEdCFxx458c6CLTvXhzABWT
iAg9463RKWZYWjk9k2SQ+bBRpD5c7NgxS2UvrMkGeKLKeLL72VIVOuPXbIm2VzFM6gUjXwKZT2wG
yajUpSwfKH0P8e9aeYu/9B8PSqPl/Hn2CjGDKX+Dvz58vp2NP3QGi63x6cd9Uwt6jbfy0zdjt6tE
8IFRIhAt+B6E8l4lB7oGSf3gEroYjxZnST/Eb7GQrZ1ZcATWociqXwYWqgboy00zDOuzuhMd4ul8
eLb7DROaiBja5ofvEEVyeLzzW3/GqX+5feOEc3i9GSjW0ZlkguclkekoQo5DR7m5MGAkgIFFcGu+
Gkhzsim/G7g8udiqE6akvOI2v2yBvhaBE7Qmq14Ca9T+f4GVayzxl+Pxus/dU6Gfof3o2MVDmdcj
lTqxiIbYixUGsysO8XQhcreUoIALc3H7/mAPYYtVzKcBJy+LIj++0MXG+pYrhVFqnruOvD2Zly6g
sqv2+nCbiFbctIKabPpa3lN27FRuzlyrBDwTgXIHNwO2jUHyZfz87vv2YAA8bPI1FIAtZm0OZzYR
Eg2CfNcrSZrZwzluAL2DMwEPNpojX1fB4JEbSCx6og090vYXbaRDooiGB/NO1HAImiTGo0x7T1oJ
UzsnN8lwZzLFZ5eJ9zw/Om2+afKTGQudjudk+abQ27aHjeDJa/KqIXzQjxc+vTk4LhDB597NtxU8
XAhwRIAHxhLjKz3wsAbJgyGWLAodZsdaGGrG8C03EXXdVON2FHTFQPywSwxb/gjFPXnU7l7JtjqI
fWxxrtZohm1l+CvRjy8M+i008hldk3G8Grb8HUnH6nfczwWM3Ud77SztEwCG09K2RcbrEoQgLORA
2cNishrU3/DNXMKoBB7+dQRYOyxn505E1g0fXCs45lPqNokgUK5gYjQEASiL5+7DvaQAjWTRQaMm
+jqNdaVrJdiJjRk2liC2Y8qpQtWn1jiaH7KssABygv3UH2OTPah6zuXBZKbVBIlGiEMynAZfzj1l
j/glPlFieKGA79riNLYFBAqqMuA+5xIOmOcMsiCqRrHAj0vJegV9b8klJHMuok/0oSBoLvjZPdHb
05Ck6imi9zVw7KI4492eoQBpOeN85HrCP83RS+pgE/Om24d2MGVKv6dCnFi2ZIK1wE07hNq0sDZu
jnwSfFFOKp4O50E79McVHAnnznsGbRZnc6pfO5qCkVGBkxXHhKAv/Fna3XYzsN0CdIeJor4IQmif
RCWZwtSDF7gv0XO47yGVD19UCpVNMvTd1a1FONnJcnn0XPXVYRcr6gKICUPSaL8BBCsTEfm8junn
xcz7JTi5fDiIc6XqihMoXtUsp3XGWsgluy7f5/oWOq1h2XLH/jahRPL22+KA3qe81kphW0N/l5+h
ghq6ctEo0C9hbQp/ffzbOfQiZJjbh7DdL5eyRnVcVNHrmBMb/IHzuuYHciXTO4do5wDn+zIPkylB
1NkC2WvVDDGRHyPn9da553eoLtgnNhuIZwngCMm1M0HxGOkieqVJ3g2W4F5H8D4ysLsbXHtqd7T3
fPmsNMIE1BPNHRmsmzrFJUURa11//PeJjHRdrdpdpC4zrSo+4cZB4L0xB0CD6QNj2EdJ0CFROCc+
xWyPFwOUU6+Dgk3+c4tIMum7C7+xZOtlluDkK0z24d/9jqFEuPIJ+jA6rMQdh8n2RAAvFnaw6G3R
yTB2hC5bsPQaPzvzdn055WqznreQFp7bofF1a8mpwK7BEundxroCx1NwHXqsaq7vv8cb6iARtTrT
1rx5mpXLCSeeudiF5z+1aMgBvvugjLzZH8WrLh0AIGs6Hg9vgjxMlUzVHa+SJH6FdRYPuI5J1yL+
8j2DJ8GL89QeNhRkjUPLh4lShnFR/PTW68kOshVNf6eIitWa+y4ay3wC7SfmMcVaF7HJ3mjYDs+3
owE/+2MpoRTZUeDATUR9g5LgVCZJy18tY9xg2KFc1cVphS9ouCWoPds1B0ig6px2a8yvlu2Vo+i0
to+CJgfVYbjd4SMOFbkvVG13ow9ZccUfcK9AgW2mXiHX3dAoX0alYQeSa8hg+vvDZBffGPDXIBXN
uZ30QtkjtxhVAzIorW5FNco/kBdfzJpEK4YS0taO78rE4Hq8N49JepKjD4578MM5W7vbJAt+vEfO
qOA+wbdxc1HT9VzyBAYpgPM0RfsIGo8sO+BtLWT2NeyH5eQPtyM98cco/txxtOoK8sxKJmfrUNc3
vwE9f4FS3z7Qn+HcMRDXugiZ7rtYPDmQbJuuTL6AubG6ykbE9ivsMWpyzzHiXlWcBi0iGzNWNT6t
VsRxRJJV9IUIYrugd/SB03EQ+LA0UQkJ+SKxM597gGIv9lFUYienVV0508KnpviqAr/qXPqmJ3HO
eax/0I//e3i+dLm0FK6z6hdpLglbcsQqUMaDn99Zqr1g8sjsoure/GBXd1Xh03J9SUa00Xf4wkaX
12Pzz68e9oOWQkydkpnG7mdtX/KQ+59v3eLJGpQ6QC9tl9DvKakVv9eJwACb+M9VIkzfmUn6MZvN
d6TbxfCQjFuumO1cXNIpOE3aWwyrr6AJh+/qhK/NEw4TrURAuBxT57auNXFYP+CNxnq0Njz3F1Qy
lDI6sdmhFYxdU588SdBCslrr4IrAh8KM3PScHB/JCNiJTHaFXdICKmCL2WfRLXJO1PyyIySKTuxE
IIJtPti5ouV9jnFFJft9jMabvKkQsexbJMRPO2Xiq5EndbpJO2XqTkIroD5GvxG6h/D24AUsIuhJ
OvwGitTauU0Hftz37HPE0I3OWiSBvXpiUCStdop9nI7NdPcTKvbVo8yoeDlwRzyP6D6Doi3RFQV5
Xt05JgTRNLvUV7N2hu3i37R02sAERvOkv2PY1/b0exOKr5PW9EyLRVyRKTUiDMYumfkCpTNH6hK3
NEaWIsOvjYVv3XB4eErCwpe9NV56b4J7CWf4+VSe7a0zSFodLIP8j+tApSIRW2wRcpSyzY/xDLQT
P4wlDoTL/8bg6OsBUswgeM9+k0vVs4Yoi78YcQ3Dh+Zzu3Mgfvn5X7x4cjXIePNMf758uwJHOx7o
sgQFLJtCBgxJvkRYXqi56jgDKq53PPrjsBZY4A+NN49CMoGNyTVuoAXEuf8WnAabwmylX21CwQWf
rVWl6pt0bcOZvdNL8MxPGiMDADkt+2fRLtCh8Aca5hYpWbvbxvFryZaATpzbDqesRi/9w5trptiw
jxpMn2si5ChF2pUMtIoZgDRQfWm3of/uwPr+KA4DS7v1peA5ThDVZGCJcFJWBwGYzGWnUTfijnfN
OEBErhamOHWW2TavNLOl0rdHnzMiSzDVW9bPjHdRD9jPevODeQVrMy7QVhKddp7MM9MJjVN39IJn
hRDSFOoGeO/hXRXWLHqZjFf4ERiMUC3OPVLCY/LZQPB0NS30Bp2MK0Mw8K/8ZaFPyXxxgN8ycvR8
6mMnIDWoa3He0Xy5gVR8V7H/g58F00/PaSPNo/jA1crCKGv+rr/4C7LIp0ESmeovq/ppu3m3bwrB
xX5ceZvuPptdqNSBVCiWHn4P9nseYzs4/EM6tbXmPDHfKvP/GD0av1UaAwpwFqIE4ApAcL/4AZE7
KpB1u9LCFQGjca9JoT4GzHlIlaTyYWlNLuQAOQpzAVlXWiF9k2d84hq8DkFHP6NrqJbEwSI6Iegg
6dgNyRbNYYXvneLmU5J96lAjJM9oU4WEnXurS08Vmll5LSltGq0CdmQfJMBOIjIRGoO+CWUeAPC6
DDKek1M3JiWFhKSpqVfrbN5IHF8O/KzVyMahWXnA3LXemAk9gs3wW7BxXoJYqKDgtTnr2Z2UkkoA
NKW/eULzZ9HcTNq4qt3tiezQJFARQ33gVQgjCkrVzLZLDmI0nrjkretOgScZW3eWMTvqYjJYjLbu
IkYxBpt402qvhe+RIjxebgZkMzJxO0WIfXJNsjcz2UnASDV3Wd5lnwsAexex+f2xMi8l2PuNwBLo
0O/aHaX3k0NbNa6gtLE39QdkrHw6eFjvQnswjiA6FZXuQ2+NnJHIz2ld2B8taKn+lFxMvHN0NnTP
A9SL3ArBOYFJns3K9JtqIrNiyqAVFInYo5r79F9EaA8NxWUFBamTRb/rmUD3VdcwshQX/7EWkbyR
2NdJOtTj9KnU2n2VMiwObdoF3S0ykqI4PUW+TyGAapqH4743nWTyRywlugEdIS51NcNmo4S5srYI
XZaHOe+bOtIUpyGNI6sdzAOvN5RTn6uLcowxMIFiwTZvCi45ZC3sEhmleHXwe647ezbtNJfkXBi7
TwwRtS+vDShozK21b3+RrzmUvY+Kah3tIVFA0An+BmnedkKJsgf32Ws5EujIBmzM3pJlD4DOLgS8
vy7IW8v0TrhukfWfpjKFkOn5JiAlWXGYlk0iSl+WElORVFxOxcpSF7xBMjvbN5/odfIgmu8WHT5p
ph7svukkM5w4I2NlFr5MxMGPkrgfCQguxBMauWBTl9ZTYSQOEyjOqfj77V+1qUuvxeIWTu/m+Tne
3oYAwo6mNkOV0nogChok4mmLOzLDPoGYN2kJGAwyDNU7VUV9Syy6nXkHY0UV1zgQXrKvj4ruR1ZQ
d5ipeo4HpjaQg4SALpVw08mcEg64fWxGRpyhbbMp/bntbMrkpGnp/U83tN/EgXdNS4qPfX5CmUrY
lHziQQzoLuH3Zg3IoCCyf5KfyUvBAyUblnISe+8m+S5RONeuxQ//RGWbXoo+0viOEFCN0v3v1fby
TWNlPz1jYAz5k6jn208QVqkH6TuF382YzRR0N5cwG2WJdkjlEWUkE/ChuIHxQtiPFBwzPYA8lm1I
M3cc2g1LnrjZDVkiRKR7GT3Z79xR3JcAcvFawSdBoi3z8CqijU5NqnoZdcRb5MdpnHfveydk/2Ys
YLGIrV5fuBk3U5Cc92sg6WbYBxIy2dKF84xEa72STeTiWzI+/o0vxQdwnYSnEbeBqnYonf+Z+tp7
gYJTFaeIbq8nlKesguP9e03XxN1cpAipKs+IDN+iYNbIl+dbXIqaA8Ldnz9qy2BRM/heREBWdozg
3Ws/aRZUr/QUp/u5AR1IuerE2OniwQ/WJJ1WHzL4ZDo8bIINyHMbbPFXu9mL9FpzFpS/GmktfROX
BXFTKMAMN0IH5/KGxPfisi+ZWFXObpoc9fJBQDqQorcp9Y6xTJiMVhC4HWONvmUepWJhRCiXTzlj
noQIn4p6e7vIcLOia1JpW7bVTpWDqLs2MBDdVIiUsCOOlgJE1gZuppIcU9YnzQOgzq4YGUjZoChg
1px6zVDZxK+0917HwpShrWOfipnAnaNpyPQlhhEB//wPYSbCi0e3VB8mudEYMpvTgYmREhRNTeyV
Vg30l84EyvuDDrQgs6pLuOYnjyTz8A2CFa5lEb0HJamgeExnGNorxtPlcN/2yzubM2RPcRd0fViF
le6fHZfAP+rLCrjBl4D5DsnG12gAT2sUk7UBHtxNXFPULBASXlkT41il3Z1k5Ty5hfCcnOmmOix7
GGEvkoRmkFzXbFh1cgsPR+lMjCDhPCnzlgwHvu62vI6HYo4zcNM5fp7O/PVuiGFR/ei9E3VoMgfb
/roBvfwQV/XElqpMu4fe/GhEQS7sbH1w70weNFbViTdf6rvzD99G/7TGokkwDc/vmIJQma1lO2Eo
L8lomptCh8s9mrbie8t5O/blHJi7PD0VhQlGFMZIHBPe24dS1VqIba1dTnlIoj+kQoFm+lAYqZX+
gtAPfHXDFJjWS5+LyOhFo4lFVDslo6KUPhRdpFehu/xT4ljS4Dd9RfhKtT2fCZp6qssGZ+XV6inq
UgECsS1hrMt4zb8QNtoEDGWtsu70033Ai7R+OOCdtZ3MICngTt6bmxcq1Z+tVeOgYjfic46sOnzX
stRj8BIgQh5iVj7jnvEar4Sy+Lj1UOxqU1skwLi9NrQt5IwUX9j/rH19IGWRMR4WouWZQmZ1NTsq
RjoC1hxbfPuZOY5/f7CKSimwdpiV90cOyqd62VjGi0gyLuUFoHmEk/9azB4IBSojgXkMgNkBeyI9
VL7pc0GdCIPrI7JH+DJCqCi++N+DH+PSzbFahmnMF7K+c7qEdsmxBfPpUlsshmXtgvUz49PUsRG3
9S9Ly/3QBPbARdU+0lfrbGKfZsq4k+s5GhmKUNsTMlfctgvZUTito6onS15K2O7gnwwv875AJ6X1
Qn3KR00ax29XcOOhwdcx/0rfnIXlAHixPO6fuM6ia0B4o9vkFB1gn+ML2aZwvBZcaYG+/BQ5r+AR
6/cd8fxyE1D5d2I5FpJB9eTMuP+nUNncY1bpfzdKOQl6N6l3oVgJALSaTD+zvSqEAGKdvUF82ruf
NJs7t0SazGz0NCW0AhpZkB21+JmBW14bWijsuwxoi8+C36DwWg9EksufJBRqXX+wxAl5OuWC8X4b
jtB9f3RMT+i3kZe40hlFag3pblEkWfzTP1MNi+n0kJ1gSscKUSKpzaTw3zyXP45AOx0mFPVgnTer
qpdI0ac38aRGvMSshSv1ISE/lUY8UPwcE5BeqzdQon3VctFQVVVA5KP86hn9KM65OWNJWuVn8pRh
Vl+aVzQMmwSD6pnqFvTWTZDfM793t+OnlBNa2VjueS5Nkm8AQeh+4yIUT/2PY6PC0rUGHOfUQHNH
wOoBla6ApmhzkPKKmBpwMlP+Gh+wnb2uNmdJU+vcbWEfeuiepEB3SlCevCZrBZ7B2kmFm4Qbz6t/
c4cnSgHipTPTYtq4VxBiXv7fXHfKlKgvenJ5CpYynBmf0kBezatJfx2eZtyLKtf6NVzqqpQDm2L0
0VxM9L1QfUGeX2Ctl0acIaYr6LCjiGTCn9dFs8wePttkJsBPABDFgCjG/Y83BXqR0atoaUKAEAx2
IgseOQ+Kk7FEDMxj8JD0NFzQb7uFawb8ryjX0Nr4XHDnKupMjfX+6F8FbH8oQ9mgpnOP489WPi9n
v03eQxDtfgTEUTR+8ENmTwtx8Pp3txWw3wul0JuDgUKnGURxFcJCKXyjAb9nXZ1xJd1Q0uvawuVi
Xnt3nqWJHUwVehTN1MIZQtdjWnd1dU2QgtIlF9BlhZiL882pDYNSBNRgi8yF0B2mUijFGhD+IMEG
ygxKVz1LXXSC2qpnMTDYf+1aGMJ8+JOL2X2JmP8YldloJWXKpyJUZL37meM3N+0hAXBimjWTrxhZ
US3Xne8c0TMUt6jDUIZUzqTdtGFUlhZR+xQxrIK/yNec8aud1eO2vGyb/TEOHDuI4ai7JCMWR342
Yai35AJst1ckVogjmCp2J9nnp/k2ycX+3cQXDQXvhHanMzPbI8Xiyh+LiRZNfM/qhZrG/pXftrtE
RQBzsCcgOOI/KXBXI94P3LtCinarUqhxJay0oLKyJR7OWrR+FnuLbhhVqU/GHvck2UnboLO8ls6M
Nq+0d5qnOh3i2rWJ4lI7gtiBpPVNHZ2Gs4HuAJ3fUe+fyDDoYW+w3oNxYrkhZKhpFmO8eWCooQbD
LnihA8dJ7W10PIkzS5GaeQMOFgqvPLykS63x7C/eCdH5FHxQFr9k90JOANkIlk9A8kYPh7iioWtU
SYx+zl9EqxwMeiRusxjJohCZPJDUy3iSX3I6Ty7gHT3z47lDwTyiNYTR50rPyX2UZ66L7vwfyFtX
AKwf5B/e9A3phtlvjWMJJ5UPSliujg09ImYnHEDo/aMcRryI74XGzt0qOaZHSeS64rt4XF/2fRtH
hytWzKXLizNUzX2sd2mU1LnbrVfeN9qGIfksafXWa3WUpKRw5XeEH1FCRzVrPKgeCu6x4DXHu5W3
znBgwUOQ9vSHh9CKWI16v97p2WNcJE9hgmSO/S0u1KTjQZD9yXeY8jWdGDWJukpPdeiE3zJtVR3P
XG4OYD9ifPVmKDckdlwAsnR5Ah7ICFDkbCvMA1ZtQjcWCNY/3Goth2Bn+a5Zu/ZTucrDkl3yAySr
Pc6FbBFC9KJRWmptaNXxfjFN6zBcPJaeUkEn5jGIXh8n0KpwWCqe3OEgjMf9cSDAa8Vh2H5qms6E
qOL+/3xiIxxyHsl+XFuLO1Zqdv/MqWOyzLYDLeQM/M/Ge+U6JfOvZOrenx6pTxWxaEfgXV9ozfvj
CcLf5jochtZ4STGIVOzgtlE/KGMrd4SnKIrRjXNC63QRhXREDrb6dbefUFbnRb4YyE32355Y4yT3
DYMXN9/H9VcMW4hezmL03D1TUkHqQlMz5m1roxLWjpBWCYl5AgyJW68mMs6cgXjxHXN+rfJNSd3K
UKdxuNQQ9mPAA1o4RmzmCrwAxtWoqn8qbiRlJUC+3/c6zogqvqtqq4RomerSqi98SaMi2ljkNnjE
f95nFPqjFplcRAXyWAzz4KMgIoWM+bNyFLepwKnweqZlx87T1nUaI/eiWZKIc+PG844R3bMOOsNp
NzHv3eFW4W2oxqbv6dxPrlBPyd2+P8LhfhmCpK3wVuif6kJB7vAw7osRqXDKyEa+zoryHKuoUQfi
TzkhN6ITIIN9MujDn6iixIya3eARTVp60daDLy8dtgk+0PwuW6c0sDBXTAOecfoX6If06EPULCpS
WGZIY1ZWJH3gSmumoR6Sp0p3IcLtmVQdRXCJsGB9x7mUSmvLqwI0bkL+E6OsXJJKPKfcSDO5rAu6
CMQ+lhtJVOc14YZdx9Pem4BvNTaJE+xW/gTl/xQOyapoqIxyDeiw6RYPtBUAt1Z+Lb1PZKZ4Ampu
D+rP6mG54FHTrBBMUmV/Sk4nsghafcLN9qd69quKDXbCRRFPb4JgsFW54OHusW56S3rfS8X0SP7g
cP7tiU5K9JdCDikCFT8TTEbqGpVARps+k+UELZTDDgDhcz5JV903p7LjG9oCCCe3S9C5UfjmclxT
XyuaP62TGUEuzXG8eloELR6sgCCZ4MlgWXF4NtN9B/32bgv3t4vZiZhEz+XB1/iOhIPgAxcWVzCO
VMIXDxARMj7j197RLeJwfyHTPmf6yIvA2qaTuf/LC2JQ1+AuZ2lZqptpnHp1Acjb1j5FrTn0IBMv
OsjGbfiOFTB0rdm9Z8QDMNnussefqefu3mN2QmOEJkmhECBqaibQIUtWMCQw0MeUlPfexrSytWmn
e59JuSm9zLDZqukbFmiByTrMQQrXY9MEcz0Y+CmtQVP0fR05vhYZyqT+76O3q/GmgrBJ44jk5P6q
xOJ7B8T3wgdTvRry76/b8UdC+q+xe8H5pFa2YWsqQlpVSHAAAhR/wdrTNUloF899xter81De8EEt
uKsfa6LQjNp6dURZAw5QJZ83KN5PmYi/wvzfFnquldqHvd1pGzW57iYw3F1JFEZSrVqr+oZxKVET
lUfR1DfVtfoJyjCRzs7phT7Dg4SNuXhbCL/njPM4kl4qqXGGA2Dbf3+O97W45L8vq/VhZyCXiFie
/zmUnhtcq8dMvpRTsEgooJ2cz8SgzQIACSWfwPjfYQ8HrJkQWUMLNAoR2HsiZKf00u7WwMTWifSE
xFztywXBook9TvwRX88PfSEci2ieHK0GquzBrMYs5ZLMcoFWOIoFkpzpa+G+Yu5Xwx2Czsgy8/rp
2VeMP1RgS84aSAXaMpXScE9vxHdCM8tyIYfNP0PJPbAFeFnBGnx9VnCBkjtBuRcfJPemEo0RSRAh
uSI8iDXQZX1nF5QHlf4tlYXOaPteNL4D0GcaFkMHcHMU3Xggn1SN27fBOSSIRZ4MKb0Jqu6gS14y
q2kwjSHrKjabcA+DlvXKoZz56aZJUHcobwsJI6qb+53NrDR8XycFLCSEl3alT/wsG2kamjJrDPUw
30RRaSUHWJd0eMyXqxLkeJswjSkpUdpj427F80JgChNVm0n5QHR14U4uCvK9AnnSfwqiRgKDnNqZ
SlD7+cHFx4NFnmhwoHwTPT1C+z9MwYI/AajgUVEiRw8s7yZLkekZNC98iugb/6DP4/9ul93OWosq
vuGyzQFH1Td9xx7lfpP6NnSOZh4ZR9GkPpMM+ZYYFSkjajDYtasno0tjb1dmNsWtURjRT69ubgsh
HPBN+9oIupeQk7RuRonG5AvOUL94U8B6S3p1R74cyrNtt5/fCFkGYvhkvWEucJIwEY6y9mBUZVhI
/YnpPYOGMQBruzmoNienDDh+V36WlbRluRnwYVkrZFNoHPEncpNv4I3c+DmqRrP7AlVL5rHt/4ds
j4EhFGTfugBFAKnt/P3VfZ7nIZ4dRmBk2wdvb3VQMnGmJPfaBvzX513cAUk9KEElVUFGp5jEPeNA
T5AikAV2aubFjUGVZBM22wXw6G9/kfWHxJvveE17UcbAsc/iK9ItsE1KvYZRzhm4aZSuNLoVeYPw
jZOuGhCmCNhLgh1n0JCu6bYQhJ+QN9a2QTi0AIJ1in8nLkalWEkvqmw5n7OS3fWnj7p/gTLEHY/F
RBlfE3RU66WY/ww1DO+E9A6VOP6KOOUeRcydNHLucvcS+Nm21qoMiGw5YDqhjVF6FZ+srTo4k05C
qeNHcHqOjYYGOXVeLGE9XQYFLUNum/uj4YqAoFks9h2L7rkVx9d9EZJCM4oC9o4TNWHUpJhuWOZc
/MRLjVctybOpmhZSo2dKazXW48ppkkZdXwDuRWvjBqHeds9PbnxMv+jcTrXCtDgQXMlYcfK5Q43X
Q6fHrQ0FFNkqgxA/16/cxzkgHD1ulRwYh3VLSHPU1x5igN4I/AEoVrlS/yl2XjE6IONE/MyGf3t9
1rgkoQ+itaHX8Jj9g98+H0jhjbFQhu4gR1z+gnk88HqkeiVf5JJOI+eEb5oZA62FagWZuAUDMHKT
CwOL2fiEFYIBFUj5aJkeQOLO7gC1666JK97RqlN8muUD+MDwv+r+LjEp5GfyofB8o2Cd2rmBTfoX
7MZ8GgifJNHLllYgW7vXheUm/xbdp3OVpQXZ4cYKspE5acSfK26EbeiDAV5OfD2S4WyaSQ/2V3jP
BCJnD4015EF00moHjxZuJaKHJfNU5lL8XBvcx192hlIVkDoP/015Y57fhfSj4SSFbz8TFXM0gOFX
OI3yshmVrMfwMjUlqW6j5d/Hof4749+b2syxKfynG00XGoUJD+llT8Rjf5sJfBWkxkAyW0ToDvVl
cZKGwiwROqRkvonAMZJIEwGrJcvE/dgpVq7Cs+sk9vmUGhyCgdxs/X09XDwPXrciEXzRCkB8Pryc
luXbas77UjPa8MYvOmroJIW4Vr0bh4giLjfwKhGQqx1p+WSPMy2N3/6ZFEGd34xZs8xQoeJuXmec
D6LBeUoGrbBJ6w8pGlXwXJozp9JUiBPIiRCIwQPLnfh7A/ugqxYBaQXskL59OO3u836lTSgd/vd1
fWsoJCkI1y+Fks9fQ18JOY4q/hLJJmERd95q3ci2i3jwwBCgJXqw7kHAaAEe7LEmwKhmPCjeod6i
QPzXWw4iaC/SHhosVd2qhtFYWqnvrT4bcoSUCkdoHRuK11wo5zHKMgNLLvrbqSzhMg5m5shnN9yW
x/ZzdlR2K50mvGNGoXhETPxnNMECcCAlmoQ8tGeJxJidYLvycu0sw86qSN7n2N7qMLvQkg/DXubR
mabNDapX5t3hcB4WgDK22XXVVkssgNcnelc5ZPXVlV4EAgXNKZDGsZ+ATRogrwaiQ/vxvCYDYh8H
xMtkFP15Ao5noLMC/pZy5pWroPC0AfEFNvF7kydG2Wrfz19Ac3ksZv+EUsFol7CxbQ/WHZLx/qit
Th+jg+7r4CJtTSPjOpJEIzpht8eWGbx4QBchQmgyUZcxRDG9u5K1hSPr6HI9qz4K/yxzs9MoG4s4
NMWp5WEJvHRWxoY+fnDy4X0Hip9GIEBfzTP8Gu1r9QhHbMMrMtKKh4dHk4mvkifaQCHiyvpus7Sx
SGETbhLR/0Q0djYjhRZfCVW3pSilvzhDYo4aBNAwdysp7lPiICtK+7qwttlN2XkVpL7RvDDKGXN+
vTcYBCLY5GCIx7bbXDvp3P/o0XQmhwVA4WLV+qnxzVu+KlksiFqoWAWpG3+yr7X3rugLpja26Ocl
YD+TAc6v5/yM4B0TZVuW9/q+VuSaAFk6EBDM0GRtDzuwwahqWGK8XerxKVu52ixw6stOvct4i2Xb
o0fygvSnwFFED+Zo4I+clLODLRoM5j74IBfApXghDS7sxgOSSHAvmWfthjmXnUh6NIABGz43z1Nw
q0eGUA8wN8kchT9To1Y9Q+nOij5XtJKGp9dyfhUDzQHBNvnjO7yvZIXaEfDcz97qWhmdm/yTt2L8
1hgI75bF8QPGaZAGLVueV+sTPkth2HDg09fkys9JwTNx4foEYmraY6MmKGLuN1/ZiQIFJsLvgPH2
hSH4Qzj9eqbN2B+xO7hkvbm8ls87ajkIGOom6hLRD7sNimorH6S+70Nndno31NTE51PplhSyNMl/
h0onFIFFOSmY5JWUvdbEzXpMicrYikJnWqglqU2ORGd9E2M+/xoMCwPPA/zVIfXZS/V9jlQCL97Z
DIYVUL8GX6dusOmqcln6fuzvvYFwLF8/BjO4gKORgteBikEM1xs8GEzfiIqQUR+sSAhDV4Rhhsah
UceTSaVdVX2HSt/N8dc9M62jHW15G0wmIBkPlv9xLIKdbEtEkiKsKkFFwfBCheKGy5+wBdaj/FwW
V0abqChgDSe+hZqKKiPZLt1WmdcjaijgaRc48x0Acyje49+OdKaCUGWmE4OGFr2X1yn0iHxyNafe
4KZV6K7WA0BiBjj7V63Sbc8Ac2EB44Upn2SAWUVZTxCVkA07uM8B4ua85iEOmJpiWtIZMkw4AHdB
07truL4zOnEYuRJXCeCxkJZ2m/99mGkiHUocN113IwfJs0DBM3+I7dEFeHQzyInnaOoxvp9+PrQS
vJSFRR7A3D6GMzNb8Zxzxxue1R7pOifHjcVTJU9DdZHqvdcYP8iJpfAAqpuhcjxJs61AH5rY/b0I
LBXMtXqUSmCIOe4OMWN2LYhuA2yK+JJSiGxKWjC4uYblrzywafInKEFVAKDPPaZpa77qEWZJyph2
jz3yG7dJD2Ztx0EnkooZGJXW5Ejpfy2kgELPbwoMhPMrWUpEdII5kBSxLj4NskLGoI3AQFpoOTPE
FQbopAge7SqJy3PcsFKsqOeruGviXK5POHJenRf5ayNHnb+ESY4KJDbQ3VKzhCUUUmsXe+8yH8X0
TyC2a43tUmR1MLmp4uOAPEhwFyRJtnSlvY11Ybddxl48jRRBsW1BrcMjb30RBx4R+WybqqhDfSGy
ahRSntJ0p/J0SQOG7rzacpeSubnb8L5I/29F5NEkzPbGqdgyuI7md40iWjIHDTllJWfwJFGe9uHL
b9xg+XRrzRUU30ji09kBI74fPEK0DrUWJ54zu32jCJBV3G9muGVL4PTSAb3DE8lfViebshynFODK
XhVdIMKJMkN44Ut7mXQGNSNZFFUmIGFxjm6R9RC2V72oD8WkU6qsAsB3T63mmQIqR7tOrsxnAptt
b7H0HdLYcE1sdh2fMfTjD2yzcYn/dBWMpcVNDqsWVbDLmbgvaprlOzmPowphsUVzDkdJXHxgaa2G
EOjSptQJcDryTMBBFS8siRPwsGNcFxe7qzCCxRu+TO/kOaDmHJvALeDN1IsObI3m85YZCibLtlnR
FjJfDO9UcA0SLehEMQ405fuh56ZKqyKrlCYyWpi5KTg0qGGtuEk7jdJEBrNlzvEGEWQLvTn1hoI1
WCsUyznkqy5SaefwEMqL9iy73T1rs2vaxc3cBI6lTZLbb/PqQaVeajzukRb8w8rVnIf9RMn5Ar7u
xg0vA/zLtkHxc1YJ/cfsdgDV/Oe7yQONcTCXC4hsHseys3XMpa3UTAQoFYb021Il71Zzw4hA4fXW
VV9pCaFFPHk9/+h5IjlJVKza1RlZWgT7f6KR4bY/pxYLu6toiE7x4g58YUd5aNH9X+lrQj7pcRG0
WoSO0l3gz7gdvmkBtNA0ae/dibLoTQ+m+TPNXK7lOjmSnQxz2udvvjEe9rlMLeGZRb3QCEhghAhf
bgvsEbeopGT9EUN0pCpbAPlcj7n0rak5GVrbgS7RWoY7I0Gf8mRfX01/Em5zZ3RGm4sV4sTrda6M
f2juKIWuixwqdGC37edtaWoW/vLrQAjPhCh5HrJoJYXVHsh6TF9147XQ56z1AcG4k2e9pmZDuavY
RRLaagaGJegufUv6NSOtXbY/uOApVOjtTmXze8IZWXIuOkXEMkQTa8Sq2QhZvlmYh8gWktAAE71h
+MmTT/cK7RGPqFTKmAJ9ERTj57VjlpuiPKfHG7SEX26RYDG4qnYxELcXY8gq/oUS5NAtGvso2YHj
0yncvH5TZge0ZA5ETF4KCuGDKVFyYqliWEJyIh/TYj6W//VbrA+bZON6LLDyQPzpaQhZK/VDg8Q8
Sfm4qDoBL7F6zjkabsdLtTy94OJbur+EhlVl50m9hVsONg/vRx6TxNwEQ1hcQtMFq+4f0vlkIEhA
dmHIsO3Kvm4JQyAfGLy3Lyot+xHRq9c0S/kt92+HvlKF6VyhfRdfhZWyaiXcTNMIzyKU1KAw2aXu
lYv40el0fWksPTe8RDXWxLHXlqEDc353BLIK1+WPITu/8yu5nLCH3d/E3l3DSlLBlqqqyte39J8f
NMutLPeOTbmqRBov6OEMCXQfuNpPnsaI1+i6EKffxKbUpXy0t0xQujqBDtJ1nSIipYMiRBh9shQE
nT2ToX7Uowl3suB8VJrDlq2DrDo2YKzfO3XxTTGhJp1xdlZxkSlC9PKnk9twj9WPCels6tkWA8cT
fipdB1Ccn0rVhCYBlcSC5oo9HPuZicrEe2IpD+rE0cl5HgaLSs23xfsj60SCk2ipx4N4WrK3GMsE
snK3cCOF5r6wC7Vqg6witejiSx1Cba0CRf6x6gjfNSy0QWpd5UHmo9Fy5BdVq1phQ9mWkWKZQ2+1
9V8P7o/IAqmWmZajMdL6oH7fIqUMGYV86gKEpyZTYOWPBKj5zDx3uNxrJxR8/i2a8n+KxwklwUYp
hxcOnrDZoogfsYvz1oOLySZSNhiytMlN6vWZUCB27ixRW9/N/5oxWmWas4a4gcBMlBV1AhAhcgiZ
Z8HAQWcB6Ms9hPAB588Ie1b8HFaN86FmIJYQOPEwlBBWs8YNGJTvlkjbwSCXxkjwEQhJjRHsAydo
G316GC0bCBDGs2q9G7xxovsNkMiDnzwQxyhu+E/1289fnEvtSt6dzPJiyAGjmdp+RzT/RCnuvAOd
jYYmX0skCg2h64pBaSi8LfyBK9Sa5WCC7esMAGvbsMIYp4IlS+PLZiswngCVOkUg73RW3fcJWSaH
977V3QdV7hiAzYTxfOzs4Nnn5w8IAyTLNRkTLhJAwxfLUvTIfTdZhnwHwohaaLMyHCJe7U9GsDN2
lfO7Fb//qQvOF+smMO+wODSvN0MalVKAmWvPqQHRn4WXTpEXKahTjqkggOgzaMWFgmv2Z2B/mMbw
R5K8P8BbrU3shT4b9b5Ifecv32GOCZ7WROhCvASyEwk7+JoAP+6JU1+PRc9+aRkh08R156EUEF2m
nabd75FveHxWH6axCprspuWOVl0iJznO5rlz9gGT8V7LeY2Xj7rxCugO+GisHBVrxpneUlKIhiB9
W9PE7KRGGMgD59Cv+37TlCivvO9NEnavWciSN21Yx9NSx/tjcNk4xZyx8zBv/mShGoZE16OmWGtS
O4PovCtfeAWlC0m4V2MX6B6ZZF4Q8DA8NdS0zLIAHe8DIPGyeSO6T4pupUIhejgZ1zOuxdtyLmNi
oE1qEUfhe3++71bsBr/ZYS3pKRGYNtte9kdV1Cn197btwN/8NA3iDe5JxPY+k47x405QHIMYrFre
6Z+KKWbC7LjZObDweNdGkHUuZ2a3Zo7jYgS85EF9QBbzKFWBbSzTJ/2jzGDTUVl1Mef1fZUsEyBs
0gH3A0lOfeESIqNoHW5sVn8h1KdfkcsfQLB4KboOYjPlkPjxDqoE1CU/LXMy26d4xdWZXYF0cJad
E1HlSo4TTw8YGPQ01rrBwD5L+yN4RIDm6M2/aFXR+RAcesS9a6031Esxw5bPZo9py8Lvh3805f/w
rDyWiI+5JwjtyiksCRAdhTeoinT1k4RDtW2vd38l5h2t6Ha37M1y2ICTsbsxyKfCiyhegWA5w1IN
FTdJiKFxGddlNUd8MFaqbKfjJ9jH/3yNx6BFp1d0miTvdvgJAoBAZxJvv44ycGPOqry+Z2dnGYGm
Ngi9SzMRH9tG8cEfWmurIYNrG/te4WubNi5gFRe0J9OoNvkWoV1jyMFzQdHPRkfC/Yb3JUecQgaW
R8ShmSbJ3XHiwsK4qMikXx2LIFbzW5nyePNanA3nDwBWhN05M215tTumWzQPjmlDd12ENlbzQuhf
P0BYqD33nRdVsp/Ed/szxHIFuhXIDyEOB1n4AmaLbdXJ9+fJIdPF2HFg4ZxKiFJmxhlUOuqghpKw
cV7U8jKwB0RaWrkwq8Kx/xwAX+XAWTDFO+WsXY533B9RY69/PuUeWHUfaTZW+xXIupjl6stWRvnD
AW66vQyriMgHVC54RAfJ236oK094pUpFif6q1YjtJMQBFWBvD7UCyF3xUG1gIwzjwAmUgf51nAKD
kUnVvzTNubGfrxEyHZg8N1uznD2WeiBNv0yrvK6tj6d84kT1IR/gbhKhhiu9eOUPOKtkUjei7+bC
j+JkQxIHPdBrqX1aS6tMu9ZbtxcGXzQ02R+vlGdwMxnNSS0Fndo8ogUXfNmGBbQPRvEUn/gun9vj
9HoTYPvDN2+QXOXV4k8z97W9NSYerDWN1qw0a/vjjM+7Vfryl3RraGsw5yvTZQMbD0FymKTxpFZS
mBDHI0MT5WAtup8qaQQvvxChxPmXIIGKb0bkMgWaSQT/VxDQFPIj+RXWprnEhE3TKuq03w6PC5g/
Gip4RgOp1nsj6b4VLnAHk/i1+XfcmtJ7I27RjRYEWrWlWvUwFF5wdDSIjkhNHjit5nqegNS2uN4P
rOD6mOJz+kpyikPlI4gjroqVievxPRkXxu0NA4fgU9WantGk5qklYjrH65fQCU2iWBfh81/0T8QR
oZwDbum4NVNEbWgeJujoacF+SparOfjDXlur1EZ6G/G3HT+ToA5Ff8dQJD8jBhwE4hQJrY3x0ktU
BgEGAbTfl+c/s7BlaLmQN58kH0fMSydaGpmRVMEHNG37pBvf76XC8/HSZZU3Wja8gK1sxKk4HYHM
Pa+Mz4g4NO6Fj7GnOnLAYVYVpiKwKxLS7AkkNOt6o91L6gRh9eM3vMCQ2DpN9vfvXs0jIX9MNyNL
implssY4Fdt9OtZSIjWOCmwi/XGRu+8AV1r9O0mFbQQWIEzuWSkFGrAcWQD5M2SSNCD4BfY+o7T1
bEqaVL6apUArYI6OOikVt+IQSHJ7eO3K7bh10UOaxq0UkjdjERXb+obNNyKQMjEIWVyEqO3YD/IZ
eLeGYMnI30f7s2W0Zc0Tej94gxnNk/mynG+c7Qyfcyrfi1dL5s+XMrAsSWdmVrWL5Ja5pZZqxRZ4
tLDODLk5ipgraYpmr4AtYun+eSBv+F/QgsoQrNI/MRRjn6oZ8r3M5BDfmtXI6xuvK4nWTkj7N6jz
lAGk+4aFiDHBN+cDm8JRQqLOgMXRoCpnx97CCTKQRLBSob5gtGWBzX/nRnIeYaBm2FB3XCO9g3vb
IRhwhlZKzWw3qetT0EzJTQ2pwf37apTZCiDatmlVOMAXdeM0+OSzcxAYhI8z6uhFxzVjjE7Lamx2
yiqXiWxB2PqZPBadTDblElHuR+Wj1aeYBSZ/JG2kJy2pM4kA58ZMss+JO8HpRI/y5LlgP0i5cl93
IuG9TVkLF8kJSRRN9RB7HDgFH/S3iIsY+vqQiT3K5OsbqUvu/T1CwdsAhxXiGdPZOBQeb3IaP4lI
ok161LSxOnzBVt/CY300j8rwKcEATWB2aevJQRz3U4o7+MUXYzV35fcENL11Mxj3zGcOO6EBFzVG
5Hg2Uv2Y4CvpQPaw4pBfIxxpIYgTTyK2HkPUdPiWcuymE0AJk909dnT1Pc96irwq6ce2ZoV2Mwmi
eCVTHyKag/9FT5TB0OecQQEHtBE0gs0M3ZjcumZTrZeoLqBNd5I9+GaG0VKXxZh0H3T/If0609Sr
Xwe3mVQDKeiZTphF/MEuivVG2lKJjAddnmIQK6FF9BXOvt16AgqZVhHuG5AdBHaDMbJjFyNAKd9n
oAnLMOUVHfwrkmFSXnfqLRpuziEplZ3Wgmv85BvlK7T2NmS1QOzmbNGi5gfHicTTrKziQ0Ex0QpX
ETgGUJiFHzZBy08cUITu7yBc2nmiXJjqWCtDXLeB0J7EvgIIkX/0wDkgatZeUGwEpbYkNMU8IAS5
1QDbT0UT2WhAez7ES0QSFg7OqrEppWIYeNvwrBxEGcyhspxv8kcdxJAFN9++OPi5yfKHn3LvHmod
P4sQ/LdxovTy+sObN5oYV5n7AlvZAm1ONHlSfLy3VpN++giq8DCf5NJNpGdV0fnVXPkhPbqNX6rQ
4V+qvzUT1PK/dmwkZ21IFIBc1pOVTlSH3CaAT9mSgUw2Fg7PmER8fZhgUO1FfFkC73HSmzMaY+OT
MjqF/tGxW4An0uijOGF1qyrTer/X1rQbAXPSZwb2zVRQ52AboezAD9fw5N/7cv8lRAJG9o0QxmgX
jQwjAgaxOV7RcXblqh7gpxyPi+/U7oR5tSjtseeFYjYazTAqKnZ8YhPij32geQE9IwWAaioE0PAz
BM0PyOmQb6svcRbFWIso7RWfyNjABQPCdHq+ofvuBGifQP9Uk1+H6TWYBhCqD/jtyL1GG84njHm0
m4oal/YmU8GPdeJqnfmrqjE++qB+mMUW4T1gbk0GAh/lheQvp6Y0bhoG+cxvfQlf0+4udDU7r5zF
fG73e/AYet5kKJY8FDVk91cEYhYfX2X8uLv9sIcKP42x+7G/HCinwrwA3c5PdQS0Avn3FfXKL1sd
SYY39NtqZh1Gdp8/J8K7TqoasEJujs+zZUXSBa+gtW7w2BajSQTKvL21HNql4fDqi8h5xv/NSnFZ
p5mjACENeHExPu8sKhMJcemQDJArHEJ/0oc3ZYr8TmS8jdPZvJgQrAceFZ9q6wiWIosxzxJLrpYU
48t11dsGIcvti4nKSWRxNBqlFsYXUcBRznXQQ3D8GKDGq0R/bwsUf+OwMIU2iR0H4Z9MKKK/XCI5
chcHx1GwHynU+8vuTOjlaMCJROoogOFjJzaUdF+0Hv8HA4DtQo2UseX+rkJBl9/Xo83kqUg6MnTE
4Skl3OJ1OOAQmE5gscGbuFYpvwC5q3GIlR4hSmaXlBkV5k1l6NyDoOBqcVPqXmZ9FUDp0lM8wD0/
pcSZqGEIszzKar2mGRRnSHXts1oAuTSmudVwbZBrvONXek05eh1lqQXjUM1YkidQSUifUXkdIAW5
5ALswzdvVSyyJig1nPye6VFQhCdHDSxeVxVp63NtxAHwfid10+C0JKGxEVKR4cATF3yAu6lI8Yli
Q2qBzDKV/fKpJfTrOMJyyhIUxA8tg9x/4EYGr7WXHXbA3Wo6fhhn2N8Ctgs9fzTqjAPRbJDz9tmq
Tu9zcLhwv8tnGhwbgYWm1SChAT8Eu9RUF+CZE5uhM1NIvFFkLIidpixrFUA3LXFB3RH2ge3V6atA
beXAQLIeYGUXdQMv+KC29pix+Ho57JxH3rvaqS48j49B7sFbHlb3Mi1S/lit/jmaHJ3nFg0w8bB9
tPp/rjk2mWKI1Au9lwUIGA1dnzIiyBPgPjEPVwFL3Ygxv+wyLm/kj34bPoVosu1UGmdmD9k60DBP
ObDkQZXdJhIOkOS7892uyLG5+XLs/CY8cSHTaTivq3WEH3zcohU0NxvF1Yg9VO3uGSmdiDwM7AiT
qoV3wcqLZnzQpoVvqo/X/cnikPx33iewMGfDEDxZwGIse1sDXjapnyxKDwF+kTR6YyKtF7Ff6Ate
HvlqbNoBaSGmmNVuUyMgD5kkJLBQfPb/Wa2jXi0oQ9nNmU84ApS52YRUO1Q+QGKQU9KTPYF5G/lf
xp9Y8JA/NMXxXlE65dxJWgOvQOT8JnAGhLu8Nh7N13yepJEhLrlqiNpDwJciHjilHtUJF9vCa4kg
nnRZWDffSTo64+92o4ZNySUmO2soAULqng5/rnu8BqWz8YvyWNYUc7qwETRF/xUUtoznQg8xI1bw
9Fis9E0AncVhjV6GvMdbJ/0g0+lv7HvDZZl4hwXwdw9fOjoBU0e8N5bf2ddZyipNtn6vSUCPYnkw
Ejh+JnwsviUgz4cknwPjje0NFkeTFVTVWWrmITovuiVJfjLkdDDFxwmHImBZfYo9qUYr9E9bEAF5
295i/TBpOpBgsRR/O4e53Wa2cx4KgPxW+zPbCiGkIPAm96ChJaBfv8BgXsQ0r/MF8vfNEZBaASZd
n/VwGMWoS9EFexyWrqdlfWRjhuL3EGKQCd4XG0eTKnhz4dP5EWc2LVLaoglQa6VuGZGEeZgHUxE/
zAEq+4r1+oZbgr73ZPRD6opZiXTlAIaD4SogNGKtqo3q9X5hwrqDI+NqSUcU3GV6cVNV0XUrlzqn
K0XK6WeqPJoZ2xr/voypuFHrmcm2PZZGNLceN1DM+azGFt851k/PKBePvkHlb+P+bJr9HWI10xo0
OAdTxsSYO34Y4ft0Nn+Jwy6u8y31awt3YybLsLYzhKBBSIA59v08cMNTC5lVI8t7iBEFJtv3Aier
Av+fTFnnj9AU4wWQwQpfVXtI+z4okpotJ2uA8J5qLtyoLZEEjTfw+2XW/7GE4ZDDTOCZIO0+Q4gg
MndCJ/rDDUk2kajU2kTZpD6pbDH2xXjHxRGNy2rxmBfRvMmO5sNwT4EmKD85Sh4IeFNvDKlKiK1z
SX/u7grbNCUGK+g+YVttYTI7TXHTfxy+zDHEfCpVx2NMoXOwa3eqdjIkPGnFKQYVmUXsZubc1hdu
aJZxM2Ggl04UFQBgfN5ekXv9zvrSBRNopMDdFetrvHp6ZCPDHaPcvgtnIw9yXwUaWj32OHeoXV+o
PC0GaWUOr6gh1Px2/2GgSz5oDIkwcqJCSqZlC2z/hmz4AsDhVcRCTrrL2t4oW1AhGIpgDsdkFSCX
IgrLzzwbWI+ReVuvX24JysnUhqOsO6UJ/GjlhnSBozzsk8XErfb3Di8ZVB3ETCVsT15KZkhBBlnc
G3ZhR7kC608seXytNJvD34XW2kWh+pjWvwOj8d50/2ZEG5SOmfhrBW9jMigLvev0a3KHCg1aITQ1
H5ugRhMIEPVwlr2RTyJfObynu4jOQ0CyuCXIDdojRch9ESPWpgK0UdrJ685bKbmd7LHVJUahkKxL
CvVpKGtsPdQmUMaK/1bjU+weoLBpnMWi4VOZ/3fqnNqtEYUoEYObw1AO9iKhjH9MeMkfk4TnyG2D
3TMQlrmjpFaPkeLqDGWZCtA2rbggg6hTh+2bNclUBTjEDVcOplkQkSBgWImxEc2Vk2ZfkcwxP5W+
2GKazYrrXSHLVbjQQBVSBF1h2gjaqF22sEtZmOzSAlWgcrpi0fF5mJMil85PtIzQ5N1jzCfzGI5J
LxWXpO0SKFq3AD8Z2fBOQR0bPFxLZ302LYseGNVdBCSzL3/nnQHalZWHaeta4qo9QIWvbtx6q+gm
TAEKm60f4Iwxbz479c+yS95BWWJ4YDda7BrPcmctWvZwL+ACFBpYaKHHgIwTIOl/7L1BrGWUOsdc
Wi6YvJrkGM4quNGckn3rZpW3qPoqguE53pc3k7qCDzKcjFvkmsgHbsLrP6zoJm3m9MWm1eWwIL/5
OPhSFLjjVL7Te2eAwhZqB0arctlwWgLj8yTGFKUUXUNu7BOeYCNsUNlxL6v1G9fntmzW6UlyQyqU
tPGzi/mVSle3UYHfzxW/vnDNrC1je04rvw4CSiJ2Db10rrD6cZRyN14V8Fd9dLgWdzf5PcVdb9D3
EfT9YXShZErmn8k84Z1fz2Y9cmZRCBALJAF6yOuqFHOevaU40phvPfcuPHcPFoeqUucUlFewCRJ+
HkCDUabXiAHNF7DMRrl1aKiBhdLUsSg9zHQQZCWtSyTK4VV2W7b/31MJsYl95ZXeYOcd6SDHeqkw
4B8yI+reu/tkxEKb3IgIZObzFiKcJ2vB/DOQ9uDAUKjTKBUnffm0P/Rq5sL50R+9X8FrYfbW8oLQ
k7IoSFKOem6/TGuqPagIL6HG5/1eLW7kjXJKUQObesxLCrlom/wx2n97tQD6wCXf87Lkk/IVYGlv
2AIMNX5TTHBOEN9VrSD0ijhj/KNby6wp7gce7H/lWCZ2KpSLyJQCcOJ6pazTYoEd3SajeKh0klTg
nwyHZCOX9lZgGKS9245vJCssrhhuk7fbZM0xtEpCQKsLkaKICOnixV4Zb+FqQUn3oE2yruJtLYz3
Ms9BoXjuMXXfQsIk8S3NnwPyvarBxQjcC04p9DZ7BPVuF/9Gc7/hHBCrVTV1tTqw77qOQYlMwfL3
duG026xrBzzvf+d4ZJXENqkdARe+tfHAbde+LgM1e+DUoEjL9ls2A8SfkiRmJ4XPcrnlpLUicFXm
kfYZjGvEYK5z84+03axGr1BI1N19xMfshcXR3jXljDEoTOGaq1rYzN6AXm4hFwdODNMyepT43AWg
gBH+MNoQfgLuOoVBGnzMJQRyR23PbZydq5LJhT3DTVkTbN1E2QTaM/+sZuNgfv4l4RB83soIkdyk
0ipKot4Wqru1nt99BetY+3w8J5TVGyJvK4/zyQx7Zk7aRH6Cm7Lftjh6qLL2RtrKwAZs1fRevKmN
FJwVwsuV2I09c2RoePxEvAgIHvQTW/xq/pxzKPvRYXLoF6isBDHAaBKOTH5bne8qjM8Yr2x+rszw
knWoiNHnKriPWTVoCI6KLWXwtcTkakgJEkfyNnF9zH3ZXzrnLUh/3GOMEApr0B/ssBIccntqgymZ
oWca28EkVpPLe14CEdACJ9/bJ4weTkKgDfbbAj3tPs/mJIyhE8d30QF/L0PcMkWvEurux0d7/YiH
nORV0OqIW6qfD7AOV5nAiB4M17Wni3GhYMJ0jQxZaupdBTo2fQ3EinQlJwm61974oKWNHVtV4elL
k/Q7nSXxdslVVmN/L2cCEtKdpXoJ4iAP9ItaTeN5F+2LxBg/PIKwGuTjjcNuz1oZUyF1mxiMG7iA
8/Vlnc3Tz7iZ+LScwqGCZv2ZsEl2DfGSSSRjQduAEoLH624eZd4Jm0p2Exuyu1X31ZvdjvXDkjpM
whgEmVieuNlENL0PyIpWf9/w0WWvOZxpgBw4W5bfT1nv2H9TKndHRU1Ladixs4YB9rbc4o9aqpGT
6kI3AZ8uzy2R2763dcSpz7iRtwjHsgveaiw02gAX3Uhc3ZqR7YoxgC+FHQGOiNa/Y6dky82u1g2w
2fBbiN6elVmijlFfAZCIJQrzNeKGH7dRoMhrUjugTdSwse32ep92xzp2hr2x3lO4ypR7AYF3r9sJ
H7Z9TOrpvhWDUr353mNvNUY6SXQvbHmJrpI3IJsSSO89eRSjQI2aR4/u1dJyaixzaKw1cv2/BAJs
FzpFJN3525UQidJ/vRO1/vA0ack5YAVX7FJAILWheM6x/KnoDub3IY64+BE/yy/HHrHFS2i3bURL
YQv1pQyutq6RR0QUEuFRKP5Ohzpsh4eYKgy0Cgq4StMYx3Y3f0Oo59UvBbVY0v8178kkkwV6MH3V
lWFHdFuqcsWhnstGs2Yb8kRN9gNyhkqAquo+brGuLzrj4TBqORog9vab0ICastTmRlcl0/kDfQY1
jNmFDA2iwCPoYOICjljmV8xeBwmTnE0Y9BEx+BWrKTKI9m0uO+2rfD6hxk8PKqzLMCIEnhNehoqc
djTiURPlI9ID1KnuoD/DyD1eAOh7Ew4rUKg3kV2A2RV3ThPKMTpg6OhdGdUgAJr20UIraRJ0W7fj
UXGcutX7A7yK/21G9MXxOy7j9ovtjPnXG1X1eHtoGLcDUfAAoBs2NqLcOIVX6G9CuVcGC4g/jA9F
c9c9UiLMcg4lm1cW0UMdRk7BRtYzd8us4HKYG4VvfUxic+xWOgCoydKToel0ZyUWy+qZeTvkmxZd
SvOfnca/pkJ46y7aFGHhWxpviNPpWbA5dobwbqSs7MRroEgZjqMJUxYmRc3wVy+wMgVU5EbnrvHo
JHlobfbUjos/55wGhe8QBlc7zfHo37mjdREuP3HHLyckJZuNUYL4Y+5PLjb1adAd/tePfQS/Pjmy
1betAqtKSNmTY5hj9B76WGs/BaEqKWCG5saprYXl76s8S72k/yzIJDGoTh18z0MhSD4dYbc0Po8J
PFKPY38NiGZoeJH/UAeojbGUtwcecmhOXQutjbIugAZFtG8id0Jv136P7lINc2jCbc67nQ2t1K2v
X1DMZSTbhjBljSAnA1pHAsgj8jgaJB08di6h07IaQeMS0yzk/MIGKlCaOiOnghWPy1eAXlC/spDQ
4uAR9sJhjkXuMr3wUtyAJHNv03J3R/od9tIcmw6MnvmGMOUkoPtjcUzBYt61XuFjqz43hIGD1ap4
cIKtwElUpfyh/3L5r/HUtnyPe/l8R2fRtmKCrj/CoQhvPys/dfjTNVIbauOe/CIeTyU1WhWse/VY
DeFKHsieTwB05xXr5jh0UTE/Lv8zR1ho9Abw8S8ZLBsoGlDRCwbD+2FkooBD7Gc9gQ6/6c27ESEg
eaHRPgZvDF+sQ061eWIilnqbsUDMicZnxscbcov10SpNfmkBCICv81jBZPyFg0P0xvhF2Ne1WUTq
GTBETSRRoRmGgkIcZ42mZiqeMViPvlvCQBhJItOH2XWhNjyIp3DIpuKIkELoLgRfAIjsUOGPYpzX
nRuajRUcX0aEVWNejhU/Rdt1MbnAfWGWJJeBsVBtWC8nqlxxvnFr8Va7J2y9V5Oli+jk6nM+sfjL
RzpczsFLi090xaOAaKoFPHLwfrbEpjsty8thmaCi2wie1GUqsMtzCC1o8nlfvKhJXNOldZAIxBIz
bT21QoGaJhQ1XauK76gW1MWHOuH5/u7ivD5Wox3eFxh5LyLdQ7c2DOu1Tnw5HdkLjzqcSVQZWYmc
aOyO1fTcKVSdSsm4hBJy/a9Vd0d/cOsPADHBVkqvC6ysFfhQG3x8wN5qrROG3dE+lLA5CjSzmc6x
XbWZVX2o6qNj66T2+GniufrmZ9a2ZX+mbV6GFyUb5P6s1O/qa6JmXHwUK6sIw5nyFXd8cHsJLAqL
ePU5zPa9vyfnrtl6BDirOvF41UhMvW/qjUq29guMBJXg1zsH6O0EWpLaRVt2zwW1PUJp2Z8AUJDL
AcYcgWEJf8KhlQ+wN35uD3so2NZ2AkOD9f8zSpKRApJchuzC/eOYelHHfHwwF8Z6KS1cfvGqJ2qn
UXv4H+D64HPfQZPaDxCusLF3YL+yeF1q+dgY5AQbc7t5ACdymbvtTwwjOwDckElNfXRvlV533nyI
Ah/07UfixB6GBWdSLH7UkQp4e29Y5b8/z483I4lEyL6+0pjFlUbXqPnsH/nYKDEqZro1SfYyJByk
wDQjIPPz9AEfTGWhdNr/f/nVEM9bSNhKg6vu0ZDuURbQVwB5qfL0lVXV26apggzwsbQim5TOSgy8
TmnXN3ZKQGZEGjtXtY4/TUSfARZVDARNrdfq5SU3uvKCKqos5IQrwJSY7K497Uz2yN87fMzbKnBp
8/GHwNzPK9/1DblEPyg4eI27pjEGqGDSMcrXnxD6vlRfTiqF9WRd2yLEdg4oEicgI2IfpdcurnHk
kvi7yAMCVoFaARm818ZYCXo6pVVp+SnXOf6N0N58Aj0mJBCqWbQdLHT7EiguJmcEEpRS+fCVxPic
eoLPH1SM+Lr4bwa/pV6YttXaaHFHuTvGU55NC8DYVxmAno8AnNJtRjhFks55McmHB/X8XcXbI6zQ
j+GFRr2xLnl0UQnvNj0iL6gb1MEI6c77/2v8uRykswjKCP3KVW9mcZuaeJyYEHE0fYWFaM/BNtop
rRJzhzSHfp0uo4CoPZj9wV1lChZJBLdCBjOdOPYKYAxNzeOkwQFMgQunljbqSDJUFX99/cJTWCeb
yLt0o0NDH4r66RgxYK0vJpvjlxxiXgzxe3r59obwuRA36qhOfsshwZ2NA8rIXT1wmWpW0LIvcvZG
1bTFMsOwVl03D2Ah5gAIydZnH4GhrGVk9I4pOWr2ioIo95c5Kiz+iT+52nEn/W1W+pRZYo12eD2O
1pQRdxbSWPjj2mDWfKfxGMhab4hIXsSDgrPaCsgPlvgjbzQEsI7EihOzxJlUHUn5TstMDADERs1/
QZFhdh9Sjct9jm7XuvNTt9JbFbfJOKVxti/NGqMCP6zuj1i6iB7DyahCqMnKj7a5e0xjo+MPvKI5
XJTvIx7t30Eh9zJ6GHrDaBxNnaYZgrzaPQ8+9Ocx0ris8HFup5X1ERROGEVGidVW2w0NSj4GO6Pr
ms5xyR3Rrt6hXI9ZPesS0qFxLf3QJ+AA1Gey2s/CiU63upX7RdWNG1hifbAQNCKOwZiVkbZqeCsN
PJys9t3i4qwgHiSOWJ8Ss9Utj5AHOe/MOWQNg6qRuNwsNcODUlT3mjmJ53gHQVqhmmwQ+sYvchxE
IYm/YmSJIoSpckoMSPeCqNHx7eT38I+Wp9FVRc+G3gHZCnUcPnjCdqL1r+a3rVYH8A7Kj+39ptu0
nJq74wGgRCtJqPuTbwt8DqbSc7gTrISbQMAeW42fb3r6mkZ2uRdO7+lLbxOhzwiGd2TUaONOfMr/
S+vlct5FAmpGML8n3O140E7FIAoIF1blBt4F91iqbNTlfGxFE6R8lZGZ4sjC3nQG4C80OYkT0QaD
1oXZPrMS4XPP1xXh5U+I6Yimdtri6DYydtM21DfcGOcaEqosM8P7lD/N1H/GdEJmhi9ZeRq7eqQm
7PP8blS2wPGd2q1Z2qSIeNouq7xd2rLJVosOJyFuj6CPd15b0n7S9YqXXAkoyhSe6kUtctqm8dhQ
RgcReSvbRN4JLVskiG+g60lwPDQvxvu11N4jbi1nTSCGch0fgHYyQKEhK1U35tBXAvAl0snuNqyI
bMTeiKS1juBBHDmELZPavUWe7l6SEa9xf1xSxSdYS35Xwc5DbMuLQr9aN68GjfhFkCnJlSfnOtOb
JN8maO515bN+clX7Odd/Cw7PraycBQefCgF1zE6C7Ux+VkUQVk52LkEaYwzaPYBJXuN4MYGEvhcf
fNm0eDg8Eh2AIBvTfRlJwBkAmHl5ZaGUrdO6hNvYqDt1epUu/4H27RUHlwUz22ZFhP0h5JY2g29q
NBYdftprgD29vzzm2NZVyCS1Xtt+dXBZ2W616IfX0fvB3GdOKkHwgAt5Bnz/Ydni0JJ0M7/8pt8U
AHewS5ean7n4emXf7YtlhAv3RJmXLXrCZqakr8ONq7hyY1hy/fADQ/8iNvapnEsAuy5hYKiAe2M7
B6A60bg+oFjaAvojHKMWiT6+O8TgFv162Rh+8liBtVfVZY/cT3L0AJC+362IXlmskUvwFPN6+4Sv
ozMslbcqig3o0ZBFqXgNwxiaSeNcjjtaoGn+R0k2FG9O2d/eJqh0S++ckvqcHyHfnFqf/Ub02mzb
UOIg+sU6fkNTiVxY60ACrPqRQvYnFgESqgSHkOF1Jz7X/12SXGf0WSRXswq154uccpJhFLcvdvUs
Wiqo9fKeK94VsRPpac87QNTsBPKLjnD5xFr4R5Nk5rlsK+SuhnNs0Y4069mO067dB5MS4N4flPyH
PmiEyYOGFEizWxaz2jQ5kh3XJdTne/57FsGQbe9YQwzx0NpJSAgJtwlgYys08Z7YDY5/3lyue4b4
jjxWhnvPyISa4wzhMDQte2uWFvLrFBKWVzXjeW/6tIuVwOhjk1aZEcypWoT4JEsWefuw00vMWYcz
Fb4SZxCzR45YUGf61t/gsqbYb0ugo5Tqon2G88ZDWEDX0RGHX255fA7NJWicaCM04++1eBLon/IK
Y0ewkPwDjFLdGn3L7uUy/GdxC+IL7r2p3kcXX9O1H/jPKB+pODtCTNoUcyEi5PxCqp0G9f3DJnhh
upB+g4g2YUOB5oGr3ADTd6od7qPvWbgAOepNocnzk9cj3JDp7awPOKHaTh4QDJwiv4s63H0DadoD
2eSrHJ3Lt3NR6W+BNMjM/5r+2OBdXkdSV9osp1sbCuB3yCfP9Pdvy5TR7dVhrYmb5WEqXYXlHuL0
8MdeZxclWdzAgLxlU/SE1opv9mWDjcq7tECDzFefL+vax99EZcOV0FUEQE9PMSP73N5g21ixJUAL
aNeK36ZnWvwT/xCTpKVaY8S3QR+BqLqbwukKAQYbCg4QNG7eeqhJSEbGBHpQsc8GiJT54pxytKN3
pRmErHKS8iEwQob55asiEO9krTX3BeXfc8L0HadT7bBXcrnGgfhcatD4TLMzkhuHvzBxpvi/V9QG
j+zr3XdT7j8vxdGR0v/LSlsY9QEKAw9BH9C9phA+znji67yf2moRn7/qW8detfITmbnzmTzbL37r
WrpDHH7aRscso65WfOfs6QB8c9lu4QRuOf+MhSa0c974bzk9PY0J5PKfWpvOM7W7YD4VeycX5D5l
dkIJJUmLoEw5a8wtjKQ8Y32uTjr1WX4FucpLMb8JUQY+eZ80juhZc7BESBw0XzVvzLtwMNvF5QY8
p3mGe/ex6KvS7YTaLSJW35JK/s6cQWgkeCoHnPpxQeebPlML+aBhWq0XhZ7JjSH7iCmrH6H9cl+S
uONljFO5m8BK9grfZe5oUbR1bkfPJwl0w81SC5TJZk0wDccOx61qlwaifE1kpZwY4QG7DDn/36ty
Mq77R0qG26HvySQ+WqVOy9ACWoNxXWAqfkCJUwg8WTeiK+WomJC4k63eyq/4Y9GM4skXUt4FLBvG
Y9rtr8Nx5EDxdx2lNJuqowHmPLsgAeUatAyhJ+GmjHy6JWj8UJA+iIg9nK7FQxDrHX8zB/9Nx/lf
wU/dVRHbTEcndQQyRaqOwrjRXMZ1EtEaQWA/keqXco/BmtqqHKqFojpp4q8fc6Shwhjumv9kzoYO
yw6PyVKwmNY0rrwmrVMQYT3iRcccfCn0Q0psUYC3HE485zKkQTu4p7S//yr3Uy1qecqOlRoj1eSS
10Skh3ad4L9RmqJ4nY2aJdsUH9Gr41qC8SlOGzlJCPkOEKNiAqsbiNSNooabexv+lDp6qInAWVbG
7IkkFqPAgjRm9ACPNA+mkXQOcitM54wNhYjQk/LXuecYEQtiLHRP6vDlvanuhyg+dm4GXAbWQpaz
BQ5YGyLSanENR0YDgyDTGFYd5FJ51GLEvZ3nOrDaGXEGP4AmU+D20pJWQ0laU+VyyDSspbWKaM6l
LYvoPk8NwsthvI4WTR9lG2u1b7+rUKEVjiWZBxtiOI5suTl3GOjowgKyI1+VV4LOv8Rr6j56gzrW
O/mIL7pHzQlvGJLDfm9HZjH014G2ii6RMJYa5CpEN97Um1pL+yxheFhCLAAyXtNdwTiVgZc4Lj3p
ZZ5Ie9HSiPxjXOTL8jICv4tajvb0EJ52ScVjDtd+x18fzJCffx5N8RYl8nkBXb17IioN7yddT4gV
kxKnFCGaBPBclDVLxmL5340r6yYYMPYTS/C8V9Qgv6kfQqU323hV0MeaQtsCkAuHNVF4kvG46T5N
z9jrRU4RbMlpXdnI4VdSNVZqoS8Q8nUK0SSQ3uCGgetT6E51n9Op0SGm4dHUf5BzHNgDmQC9VIrm
YqeFwP5uRdc46QRU+mc5tj8phhVXDEA2tA3BvYvMeNAswlMwftfEgePr9YQ2GfYDT1cejM3j3kMi
TJe6TBPeC5BsS6oqKd5nCGXjU1oqpUkwAOD5ure+LDkI9B4CbwvbQ8F5F90fLxDMoCWCZznA2bl9
SPdsC3U0FRJco57ATFMpOrJvSN+j0/a8ivc4RHCzZuvc3inhT+7l1feJcBTOPBehmrRut/9SqLPY
bL2s0P3EnSMBqJQD8ysIh+ViRxDs0Sh4ATLkTxptZ8SkQMMiGirVwuO/B2Cu1aIrh7fakrZobaoB
1NZ48tO69rx4aP09h1/SYmETqbEdSXZI2N3P3umD09Af8SVl75rdsXiOf9S+HZnT1PBaGBi6vgE0
rJbSBcsYcBUjIDBRDes11xnVxI0NfWoH8XtbzJcWyT8v2/2AUu+ZhLAewWXxYt0cM1KVHknCyrqt
lx0OsWITiuIx9Cnwvpxot3zUsxJmpAYH+TivZUE4rEDUKkOx7Kkc7rYhs1GCarpEKt4h1bpHrqPe
3/UE6fKKonAOcNTgT2b/F/VBlVan5VQV/RAJVHvxXIBv/wYyBzV04h/bwSL1HGwdwoA17+l5klF+
sZjhS43TNyF8juVm3JGyoigdfNQPb5FkSeN8PD9qd5bHH2KcYUVKoirgdGPABdP55jKdUI9ZfWek
q3DkU7nWvEYgkOzQc90Y3v6Hk4GgEv4zeEeBWE94ywY9jueTSkLALHmzeIhDrXnaa124adH5a4z/
zztIJBuFJMd4szvcLYotM7zLz4obnsg/qvRUvbzcgNlVjxFtUWeGPIPNMMmE3qYIuXq5wuv8perO
oicTYfoio+1xg3AqGm9jHcLIyKITU+dfSQyf9Ic9ir0LYWS1BVTlNiAvCA4BTzqLHIBHAKHq01O6
2kfSYCylV0GtHk3YST/sGH7YRo/Jc6TMHLUxbR6la91D6iDctLpdD4x7Kp5ZIICndxEXxaPvr6yd
6fhz1odeWDq6usOTt/jXT+qO60ZWUPASCzOSujEOOCWh7BUUI8n3lICGW9IfOd3lSORKpKA1qtZp
mpix6QfS6bKyQtwogbkxu0j3aQm77v7u/6dagmeE6TPd8/P7dJMRCQnuRWHnhwQv302vbZ/wbt2R
8RWFi/LCzqiWZmhc8X7YH4hJQQHpWh07zQQoMSBOMQWEgnfjGtdc/Sa2XucS/ZsMwZX3uCq1nPJx
ZeYIu9SP6KOCUdMubHTN+uosjI9FZ8i0MfM7oooYJQ3x/F1nxX3zsImBbIVU3lwMaUm7YRWysJmP
zrB6DFKRrgKfRg1ivrOhpxBRbzVYJwQE3A7V4y66gyYWueubgCXSP3D6FTni+e9fUPleW8935JUs
7pxekAKY011zBuunhesPpdLmLK7fUsi7E/ti/7NXEn/YXMa14atZRcOxwqaiKnUTqwdcnkOGG7CE
Dr4xMB8mciLH+rn4X7fjiPEjVnAvOHKpNTeFhAbKsDLsVv5XtCfqnwIVNgHzjuP1z2N7MYNr48ah
W3O3oIPuimBtaceaRK+gyj07P8wquy/spqeyZGLcAUs42W/SvxxRXmx0l7Xmd9m9CJgoxR7W1cc4
pxxgR+RGDOVZ0838t1lRyCcUtMcAhpp8qG3Auro53Vegnk+s46f/IUtT+py6Ls6xv9b8fWxP7XLU
b+mGa+Tr3NVNoUo7dpZ/x7w4gwEghH9dN9rA8jpxYvpl4DwDqE7dIPVHJCliG4G5kMjr5JBJhP72
mDkXOaaXQppCqwKpcZLbFnN70yrcYwj3forT4hnEe1thHVDcjcCzAvq+as3ZrUBE/TDHv2/wIpjn
imTH4mGTsjywH4fezLBfyOz0GYj+U1HfJg4Zjd7rQioiryVVjcn2NwdZ8L26po2zGdyIGjw9sy1j
APP+cy6qpApuLYIr2cJSBHOmzDrKXt0maKGzBxTVe1G1I9frP0t10rfztJr4QxXCaJpudE6hIJ73
IQsNAEi+3o0jgXXMW6tEfD+/Bawf/u+Qd6OAYF6ETgdizfMnrnDA6v9Ye0WkgMudrLssUfcCUc6P
Y53hcXfKSG7eI5ijnqBM8FjGzAaLuZ7yvtdcI5ouiLPTKXHV79RmqnvCjK8PXrfuqCLb7ZmJQwHb
2RXHiQqN7cAIkGESKyAa1aqKnIrSYTnmN6FnzsinGykEqNVxexrO/dt946/FEjo2yzGelQ3kFuUx
FdRxygCcBIZXT8xcXDbVy1pNRvoj34+pwo/PIK5LDkkcPAWwh2Q38TD8f97cK5h/r7+7qDtUgg8P
r/dGsnEKeHZYrYiGG3Bi3Ta1imbDAggXdgUbOhi8jCLJpqBTXOPne+l0Gjg9GqF3CfklLMrXx87P
bUMzyqZxkPx6GRyOlvfKQemkXJxxCWgpVVsTMI+x0GLW4aNlupx2mfjTNP+zi/ILgGrvzON/N1nF
mCCj5M6g0cEckzCa2TEZTp5nlmym1f59so5onl0eMIiMwOE3su/xX41VapnUza6lzjy+RfQd76L8
JTdcVpkM+TfgETOseTwIthyo5X9FXGb85W5UUZX40fwTCyasKIwsARzWXFY5E+IlVXq82mGy2Ihh
xtNfJWy0MI/SDp572O4gvHzJ2pqT6HqLYlCegz/SqwFzKL0CuuKjFc+I1gcGGs5B/VbMh/KdZMOU
lTbG/zEJ4p1l5SO1RxpyBwVjsD6MTcxrfwMLVGHAOrx9KNRrIdzykDF5XL6Xbn3g3+gvU3h51Rh/
8qIzKvwAar/qjeQsXK51FpErLNVyEBFRg1IG6B4Ca7DMGI08uC0eKqZdXWKDERzHNy0AtSKZrYy5
WTTJjKCzpLGFQK+3TpZq7FNBQs/kmRAj6jJFMnuheWVQjqZmggBHawJr4498AYT8hNvx5dEIKWO2
2gVndQt3GdiXsQXhXkrkP37rjd1GVE5/BZ3TqyxGqWKvFNxfm7OixuPjAs1ZEEmxSOBZCDEgqA79
1FnHVUM8k3WSTB963HCjYxfYjOskHM5Tafb9UNan2TZcNH0Mp3XMO1iTvS9cu+KLjxGEukNGeSvv
lJ9YWIY4Nzn3FnNxIyHIhbcLIxTfNFrGTRhxsX0vsLB08UE7aDyAPYZqfQY0mcL/VYfgK5w5Eib8
L7ulex/NjK257blF0lULOPmMkC6Ej3Vu/imXWN5pWMqfrE2AbzPdohXNWhcFMoAagW4sxOxEP6iE
bWsdYs1bBhok3TMPPOt/ug8CWfEqEiEtcqGCCOPMG5zxQWGOR3sLPeEM6lfLsZBR/ckxEdjGVRqW
eFgnJLkxCI3AsWuyfEp45oLZkx5PbBItSv/3zjn7XcNckFhhJqhSFCKIlvOxhR16auHQLVEH1+r4
c5AQfNIbB2e321HwgqGMa+J/ykZPiPm8MqTRi5KaNB9MWKb6N2sDPDZGtTPSq0FeNqw2ZZ1XSUG5
rbfWCCKEn7HclVeTRaq13Ii/+hqiB08mnqCMoyn35/RJubWezlgb04uOgcMsQbzl7kYPgVkngroB
vuYowRY7/EBwNd9O6ms34YsEaz+qS2cKSiFxM38H4bUyKUFyXVl3lx82aYxCnpkcBQ7qAYkDg0r6
pdqrJrgQRRYTwI34JSs9tTtei/SoE0y8jwBmmJjR9duNNabwYvNHC7kKmv6UTH3hVkxKgiLtyAXN
yE7970gdZ/9d9ppnUNcHL8bDQlKe6UgQiaVi0U5rWjPFd0LyxI63sFIZey+ZRCR32BhlRj2CpRjh
gqPECfc+JfVUx26MWZKAUj6IZbzxpotxeBbRPfbXPc9mrGuqJ9cBItSGeFdvPxm1dA/F4uDZRYff
hebBDRdsk5sh8MlxklqBm0los2G3sBzisRNLw3B+cxgM5x/Z4k2+UN8T1s27EzQD6uWfiPqt3ML4
jdphWeSVcsmr4Ao36Kix46xZnGcM5u/uVSLJtY/ch9mzR+9QenjEDxJIJ34ERIG0oL9GGSF7q3YD
XixEjcjiVWwDMf2JDP2tBOvclQx+NxenhlJc8ju/IP4ExWE1a2d1IeNkDNixWCMMApIX7q4ktTrA
+N/SNYV+4/pzpG4NOXz7CeIEI5DMwoWsOnBzrEtkcH7U4xKpabTNuHywrADXNOXfALiv/ChQ6yiA
NVA72DMWdQ1rbRDVPy+Akro80rAswvcyqKk6h22P1RDm4ZTDQKyPvRzVks4RxZqOR8xgr4fsazwg
M2W/gLY33K2Hrs5/7C6aeD5pw5b8eVWzcgW0VAklerQZq2gJTrthjiNLf7OwB90bcXwM9qJWVviU
aV+yfIcqGe2cH4a+Sm24hIHOR3Uo85/Hk2+7jwCrsJrNVKr0mQPpPtwJwjMn7Rx9yG0xTjEuYB9M
UxKr8Pxlw/iCxd/hqt0EjaS4oL0wpMEBxbuaBWutUWAsGug9TnV3skUtL+QhhKllYqh8oGJ9uRbU
jC5CGjNUO9EWwxeldmixRpQLyAv1yvBHdzKbHAsR1IRQ1Ru9uLw7JgzqaAh3tGKjmUSw6jHJ+IFg
27qbvPmHG0vgFoQfEu/LtXA5fCN4VSDFbeW2YggMNqlU/J0CZ/ysJMjGdNBCGpSp3WzEXGkakPcd
QYwlT0OueZG5arxfEJ1NTLMlA6OoS5mCXEnzLTbqFjrExeRHRChqYySl7yds4AqemU+VeW4WVWrC
kuN98sLFJo/aOkGbJsqQJBQIb2ecd9Ubu3s0ME2a2QCYOrdaoRMjCZOI6zCY/D5/+67ahJPfj/aN
Q5NTfjqCtsA/3hxmevDMw6hz3iXbIsceJL3zYyA/6mb7HgVaPNshTz8jvC0/85Fl3MWm40cXbu15
Oeb8MVgmgzEyH8DRuePdMG+rO1rTzDLKd1aOXIoumt+ZJ1IRP1VPgzWTOjYOgDmaMmLaVVY16oSW
K8Wo7SRWHxko0Y1FmNfCU7qqMulKNUiw9L8eG6SuREoRs+uv1CEe+50XddD2qWvK+lTieJxG2JGj
zDeGftIHljpvywllw5grOgaGDvrPuoSB3OS8aPQGBQ6Cv3K47sI+nOM9Z779xWr3srV4UcZTIlXD
ZRcic4OLiWXd/xzUOxLg02UctZuVN4BFL4od2MZH4hAlEq6dkBom1jAiaNpi8DkpjJhuj/PNhzsg
PjtgCkQYh2UQqH1jqGR/fcY/5h22CbMu4PUQaTwnlGwA4E5N4PHB3dfLaCSjUrNdXPzbKAF/2AZU
OzSBptXODhoHsTgmSN4Yh0sotytDYg5fDQsvmCBEwXAJ+C3r0fAr9pFSkpoXQu75QmSCe9jTBdaD
EJlzpOswNiyORBH/SEIoRaYBXomT+EVK4Edrt9AHqKPwp6yMR6+26klJv0pWSf6bCJ0cjTUdjZuu
JruyA/774B0zjU0cT+Xw2oI78M53qcisafuulqeByM+6zMamcxyXBp0wl/iyB8JeLwCSgVT70wGr
3Ai5vEk9zfj0Fjh0Px+PZsu1A+Pap71Nj/zBAW9BpVC2iB5Vg+NP80VhMMY8LaoOb3xN8Eke1IH1
aKr2wQFgDniq1nvgP46VZ/6+ax2wYMTTODFgA5VJc3FKiBP8sc9A3zkaPeLUYYbIeqIlhhkxA/ol
QoM/Lzaw1Rsli3PHQuCfijf5KBhgRkViLBrUhwJilLYOrET6D5pTgryzuNaDMgOQd33cp06VnSYB
+O5WeEx0IJfYIxq6ilLRhOoVyatBQm97lt2tywrwwhkp4eQKhlol8SgOtRLqvzpHN8YKMJiNwgcl
uJnwpHqwlf15Q8DyNjBpBuswBzj4VyT0Oat9RB1NccxfI/n5inP1PIiRTfCOtmsZPxzvgFltwVdc
OspJ9I+mpRX2hDIXWB/6Ryh78p6/G0yeP4EpB3LhTZ7fWVxcOPgpkufoD/v1B0bV6XVez0MhdkAQ
eFk9kTKdQ28kU6m610mzsNL6wot7e7YtEGa3AtajRTibucv03fXyc2/eOsrIoYf1LxRQ6zDA3g52
NgTKHMJK8uRvc9L7IkpWLY/5JtbOwLne26pzLOpwZCuHH2SPnqjvoAUDt4/nwtcKpYUR0F51ktIE
OLHQ7hHw74NvcJIuwd10GCeN7UMn2uKzuScpcIjTbxlPuaeTlSQ0iQd9dGcRVyD+y43X6hGCx/yq
liWLnos9H8B8rrqgn2+cu77Ku3sMUvMAKE3y+P79XF2fEUB0Y1WiV06U/KxM+V18zpDWZDiDqqpx
GZj9sDlF/P7h0GjQRDuEHXzKZHBssDjQJlEqy1Ja3G7lPEQ4QCRF5l7e3rin/BVeGU9t5qL8UDLv
bKVqrklomiEBAPNzKnxLu0ovbQpKNc4GXxKJ0ExfxtuurI0NYn8h14todvmiW4ZGQeJX050OwcUQ
WXb4JK9N6Ay3F6NXoeCe4lWWB6vkUJc4LMZgQ1TPKXyY36O0aalhS7pGhwF034qYBWCOC5LSpdUF
BHUqZir3qHhEO90FPKa1ekhpq4wzDoKUtvdtUgmEMAREQAv1UOj3PrRw9PiI4QFW9cXMSylQwYum
YyY6Rd05kBDwV7J+R3RoNY79geOJqbS5i0D3qi1uuO72hNOaG8/5oBTq9PQOugpI7Nc9zQS5o/Os
wlBagoyWdYmVux47g/aNJfBFn8su2WlAHLaVKxDFyQTR7TsVuEDNDD0bYgpcAlfVqWAOGtCbCC6H
rNPoT+jE4xZ7dtVrl+Rr2+UQ1sQRHvJgAH4lQ+QXVvgO6sNUU1CfKlFJZ34C8qwrYCHGpPL64bsL
Xn6w+bB1bkOuzD+l2SMYQBfsSMhNhzCs+uReEsZmTTMASolm7G/KIbQ00UvM6u/QQ5gfdEGdaQ58
ODJ5ijK0Fbo0P19T8RAuiTwJ2oxdLbRzVB6oxpzbrdIytKvPagyw+goqAzGYpIs6aLVmi7L0y18r
0HUdplOo623PeY6P1gC3HYmlOhlVwuZGpObxU9ffQxUYhINyyxHp4EvUS2Lqsra+fW1TcBZ8nXVi
nj6D8HNN7oyBOO2dMeJmMg/ij66dygagj2sXGr7L9HeARYgebP7jb4Emxm2Qgd6I4eOWHSWx698m
nUiw3yU4d2iw/oRgezuW1m1nytymcNmumpOU5scDJtIOB/NUU6n8ZrKTdCxIKWc6Q55MnYk+Ifab
am5c99AVT2/3WtpsRR9R7ZlXQhIv10aJ6hFpF8WzJid1k3sGg30OSwN48oQmSFtabI9QdCRp32XJ
F7/OoTvxdaJHeUfc4YkJWfmDDc9DvSQYvT+2qLkkTisbSzJtzqUVcqrQAjtiDNIpd85blaYji/On
2J+UgorW8mSq4Rg9fPXFIrQO3MgrpKMkA3+aU7HCAHeJdAPEm8ukYH9verwZTty/3vwpB1y6/Ddd
OgiuNt0/USZOTelklud6haehtgoa8adD9K1WhhQrCCwvcyktGe5jM49tJNemVuMaKlX/S9gUHfe5
F9BJAC78PYOEK07siou89/44DR4VmgMi8ecApX7DspICRU3moGCuQx55G3AE2ptd/AQaLJX8UQt8
W/RfRY1wGzy79wFKY/AE4UIQ5c3RWGiyOQUpJpqu/C8F562NZQidc8/lTGB8Sr9WH2mmz47HhXkZ
Fh/dhtu3zYyz6rZqH+qLFVkJx3pNy7j8Eds4fGoYMTx5gIywiEK0abart4viW8m+SjgVobqFM5Hw
K7fe99oxpuRsLvHIce7k2kNA4e+5pyZqSa028Zax18k50epOjb33fwQr2nENgtN0bvL4oHkC9zVy
A4FrHo86DEIWOtd5YOhDBpLnnHOmXvePeOU45HQVGnEH55IHt2tvm2SZsX8/ODotV1273lKAWDJn
3U6jy5bqg5C7LYB8vNIcawlt6CBfz3Vcm/P6EYIr44FGOpNPadq78/CmJIxE4h9uGW8fnS0H7UTi
3lESSSQ0bIZDtqjd9gpGGtI1/L5U6vZJz5x+QyWAzI5i1ls3BJhXH5iAMnO4ez1vDJliG+wmROh8
T2zWNkhKEGp7WHCZ0dM4IkFqKRtYkLiXmwaXBem2QHrbEJunmSyI2Oba0MKMg48UAq34rapSvI2T
bEyhk4sxB1Kh96RgkGKgCC+0mwxb7RaeWhvCPlCQpMB6dg3jNGbRqBxFS3uCv2Y3Cxc//s9pfvd5
QbGof9QZcJSdHPcRm+DheZpz5OFFno5XZ6SYG/4WJMeLKa0h7sWi2kcpfWg2btbOP+egOoZ2h0p0
gOJCpMSjtjgPAyAJnV2Xcwrd7gsVYsmCX6y68z6gZJ+acjpzKELVgpoXOgQeDdbrpVMPzjucLw45
GhWfjPjev4VMbVsCyHy7fQU6cXud0ezNVpk79cnIgfvohIqJ875PMe3iZlY8S1ySFgVpQYah2uz1
STeu4saevybSi9i7NsDn2WuIlzf1P47YMLSYmmF/LqFZChoCGYHoVzklQhslKRU7fg3qNpk+8Add
4rVKASIT8x9lFltc+b9Pb9hQqCowBlSe2cwX+ffNlAwDIAhclR4XwccjxVZ967/hBVK8NByLIe0N
ds1YOqTAQL6LqV0JVPoXyH9MOxkVWohi3oQIqFvfHWvAkk/Y7tRklmDmRKEHHe/o4MRTrrdPAOdN
7oXyy+ObNMumLTuk0sYscTfWTOkd+2RSRNKuxwfSROhLdOrrkWqqzrSPugNwSJ8u8l/+NaZPpLrZ
GlX0IChxY6sXMK1jEo/O8gvlrE9rYIjZ9/gaIaw8z5NeKsKROlm8mXXVpn6oVIRDhViipfVIybqj
3mtsffx41WWDIO0SjYX6E6brXEzh1Jhi3hCJ4j4qjw03mxuvfkkD5wYS3//kqxWunqISzRXviuHL
WERXCLEtSqy1n6rWsuGTtFtjFnIPifHp2Iip0BiIjbRqmPPGvSGjrXSvLEhyLctZvgMU8P/aAT3W
EYfYwYiFoAtSocjlcKUDV5Uptc596AsWiiVekZtLRN0WKqVTrEVFRnqvFiN1I/auuvLqwsuCpzmT
PsKhCyIbThKXcbFV/3+7ZUR8yol9f/USAccxXUKgSMMQiwU57YDTv0VXsfl3IrSCBzLSxLbBQiqX
73akUtMD1J98BMMfb17pGnZaQLwyIyXROy9W8pndkiRsYTM94fn5n0YMJQ6xbSBc4dBFr0TBd2bj
h5UkEzem9reZdPPpxVBdnLP5WVOceh+YnxoeKLkRtn+9L8JLpuPXAd1g2WOW9ra/uCkiKFHuzSRM
odaWTBfjZaCjMntyyeJrEFMbRlfpLgvAxTPjEjXzXm2WDtc8P8YLMSsJDYKrz2CX8rPA6miAR/f9
nb6YVumkEQ/6K4vE1lw0VmAOE04RIDGpcyD4nmQHr/4bkeR8cfLHFiixInsehIRxdtqYN0yXb7Xk
2Zgi/XhEdcdfMmtWpN+kkYmda8sv2dAsmj8imtWMaerQ5lQp+B1g2csaKay5j0HTF46KR+7HQb1I
UA1avNbzQ9gQmvPIKrgYgzp+ryFH0ZySYCRHI+EcE01GfPt1mcMHr+PLg9ckxr3QKJvRshwTNqvS
wCftGGM1uJrWfqTJwlyAdp8RAZcE/RWE+wAokc3Jcqk2fCdMo9iAhzdUm+Y+u0rONgoqAmXNjbM4
/dhabyvBnlC2ufq5/JNE30R/EML+s/ruFJYudE1uFwwBL5VeGu37CneSrzV4aUAFaI2nF4lqwe/n
qcSNHb1YYttb5OKEqHtwKYtrS3e78mZlxfs04ATmOLKcjOPwoLrURVzwyWqKw3bmLuisIUEuQUi8
1hi7wPD1XvIK7GxQauDG8wXKoQCFhTlTBjdhmk8UvnXOfgzApjsynt7pIB0re+ybmxy5CZwDPC2U
TdUzVEPsDUn1TUIJZfYV9tK5mbfwNLhHPFjNKT7OnLi/OzKXm+X8MHtawlGyUtFVQtvuTiHmMdVZ
2oVVGBAjJd7VSvlS+CkFlx55e6AT4AtVvVnzd7jXoPITtUd8OZXAP8ELefnRMA1IHQ6AG5Ee2BZV
W6qhmNwzE2R1lQQy1bG/dfRO2w/VXTYKZwAzJChvz1GC1rQfNw001ujMAqGXwiLwqNySvIrQnGSt
aAesa7L3NIydrNCohCfKhSMFstAlcBeZPIQXfs71ODlA2SfZG8vTVfsJScN+pauaEAmcpa1PNbxT
vL2s+qPSFzNrmOXjPZJRvV8NCai6ivCH/XkdN+Di+ghR957YyYA//jQeMiV9YEGltNOH/xOiP+fA
MdHdY143+QiYBxZyE4Fc3HAtSb622SJ1dmVeFM/jULtxS39b7iZMxkEeJDmcAIwMYq/d2MXTUr9K
0GMRcCDF+M9j4J6QLLyCDimT+ewA1263rtmdbDFzeGMsOoJLiK+Fpm1TFuw1kOZZHVwopY/MkSDA
I7rhRaWPOrgLOM53K1vUdPKtDBLc3Wg5Wm/wUSDLInpPPkX+4j3tQydYxoAKDJVdzvgvQe/dlVtC
fMlFOkrrtchvM0oWgkMSS2XVFy3rC08BDeohvQU3FN6DgByKS4mbaP/AY0cy3ADJd7pyq6HBbHUG
/CxOawLhnXFJLcYBOMLbMTkq/sb4ubK1cvZ/5ZJtPYakgCYNYIWrQp7hN6/wwXSP3hX171fbRwfL
Ap2fKZhOukT6FdcZMi1Q0Ksuujq/IXj/vxdSIcLabTelVvUDqOMoZXlZtCxdD53tXUeWemu1advv
UKN+mRSXOSW6ybok8+WyDZmv5KsE59FKa8Xy70kTz8XYUJE/dTCoqkKy5FODlp/dRFHmv6HRR80E
SWbGcLlhZtPoy5vR+4oqqZxGQJ/6kelpr2kTPnGXpLPBwZ29Mjim0FUwM5K2T1pl8Po9LyphCTi0
DQDqniEjlRqhWJSR5Y3eXX+X+Pt+ryHOXY2NrK5F/7j0tx6Qhm39K0iiJAVnF+1cOl2q11AA0c4q
b322cKZzX+rof5vi68RpJUL6WeDmmvQT1qmIqwamou7BdnlawIfdJYym5SJHBi7UXI1UBTXqh56+
yVPviFdPrgDi9eKN6whASnARlCId9ZKpzgdLjNsIiBvakO6y7baNZ9GdgQcNniDo8tOjqLZgtCw4
PuEWgDzYXHWvqM2ny8xGiKUFIMSqwCAac9QL3Xzeitpm1mfDTdACC6zVASU369ZoRHfjlMjt8kds
hoeJn1hIm2arXrCXvU9DmIklt9mr1cG5An9bTkMtG5/9u6ziSHxk5/xadvjSGq7uqXBDlmNGBPcd
MslPeYeUSsHgegzW+n4LA34e1nfF8GvTKUZOj85LLEzdSZKXqPeB9P7rXxdHG8Y9qN0Krbya3W0o
TiCZk4kFJ3cZIYHGjEroENPXo5r16hyWJlIJb3kREyzjjpwITcDFvT2FdrHR29bL0DhHvWyU25wh
XT1EbaM636cpvzShaPHFByOFfnSHN1RDVtfQmF4hG8yJv2E7w5ov7FG8CHds1EunrbiIWwTLkvT2
ShlVz/mfUoGRVXt/Bx5jqPCRoYoBxqnvfOZGsMz6niPAea8egEJnkUce6uhJO1PmxHwWQskW7KCD
eI6PN/Rh9LS28hfcyF8jjBp+2GhXcM7T2mf6f4Cd7heU3T6gBcoh9rdsmCV9vw+RkDk7PitJ8qXF
82XO4u5xl83Seqv+5IGButKXnb7k8Fv+DgzvYDhrbcw9A/7C0u8nEgA6aDDNgCa5H/wYbmT/MHDO
Mgn9zJbNzH6UZT+lJi9FYX+otLr0pVTMtZBMJwBDnNdCnCV6Ao5P6wb613XTvFi761bmJ2YfXIJg
5p5qWdHC5zu/CF2e1yGzxsH1woBCg8VrGiyZZ4MxMSx7H/Sh9aviTh9JZQvd4l3lVtwZDo51v3aR
ici/NkY0wX2andHpBuv0WSJEyCIjFXpNeDyfu1z/DcT5E4cw1aqTWDUqN7J+i/qcrFdj5V7MBOkG
g1KNUQzGIkAOOPepiI6VaRW+WTAuLvup4t1m18RBfXhiZRazRQlHb0xO3dtepKlclgNvjXWcKIKp
izAKQgyxCwajzNsGqmk8PRHA/BVLXzJx9HpgAGTaXMM48UnR0vaS1+YmRMRqC4xsFLUXfSZWsDPE
0EkUAOQpa76IcNYvU2ij22+jztQUx8ASjkpzzy3iUQmiXOrHpmRqJgJxpP1nLQqYuUATBnZEmgU6
bq7E3ZqiFmkGrfcAuky7tmoD6JGjRXziM21nNMaM5R7UIXPmxYSnMqSVsdIphuQy5h5clcKb74w3
g+qpXZPdkkw+yGdoFHOGIh/kzBNtifl+OIZFxOufjb4BcwPrf320a/rv3YyOf6/F/2JkZHDiSR/G
lVGPfUGKIkc05L/aiEhX7pLGCQjfMcizhaboxvfkyAOMzGFSstKFyVMSsIrFaZ2YhFueyrvaQ8eo
2Z/XDrcZ6gpTtA1YZ/1rZZTxMC0l9d6UPnPeswfn7s/FgIGTZ9EqVSS5ZTd0NrQyeY/lFfn6ISwB
EqgveRmI/A7KcrjEquYutqFCktLtZDKNUPH8GpmMQkyeS4Wf1lQAJ6VY6CJWdzO/R1of74pvJlse
v0RbwtqOHaTz7tlmG5UM00Ryk5HV4uWn5UVtfFq/AiGmfwJJ4ijMWYxy86D6fGQE8andbY9xag19
YT7zeEvdiHWWPEyXKf1OakyQRhKqdg4AxZpgUpOY1fLM3jbLcwtky/4CiUg9OgQOKbQJXRfqT6jn
jmzas8Otn8OucNg5Rjda4s+gMdeUCZE3bTz2mrl76J5AuDLBOthulUJwBqZ+Y4Gc+hOG1wIWzvgh
k3WtW69S4s8QlvbOjx3m63pEl4JfudDpz1IAMFDf41S0zdgpEHzFtuy2AAeWhcKqsg7Qk1vbE6q9
acrgQzK/9gl4UwWfjUdmbsAilTPhmADQ9iM+0KpT78lKQZqGUAiVH6n8WLGUoAiiBXNPVrgjfLkK
As2kRnSyFVV/Aru1dD6xmWX4/5yiPo40+GMZkGab0OKxokV80qmfpWOxlBXdYge9i+FeGDJYIxmU
ZMiXd9k1/xIwwZk3xL/pTnsjCckFKelQxdpRmDdZJXmg67BZt6sEmaH92PriCoiq7x8JHL9hrEQx
S2rKZA9Z3+mCdY0Ne5M0cRetKQOSwed9Dwl8ul6HIaB0IYUA9On6ymAWcGSes8S0yy8LBy34UHwD
jzUWmZCng8tcTRCWpoZmhzTgkTpXXNxXHrAr4sD0gy63Hm74dBnSZkxQtsg4QoCI+O2vy4fqx0nm
m1XypPHCbfzrfKhIC0uo8Q1eJOr5NIYGPFT0i54QJ9Zzo0nwaP/0MSJYPYIYUAa1yca9oufWgJHB
eapzU4/x8W+gKRprBDHpwLlPY/2DMxwdsw2whPwCs6MekTjvcYjAUGEhRmVbyO3AozjvoCTEVsPd
PBoK+5GpV0d5ZDPNwxngBn0XEO1rGZybHJCC/onSfMvnb8Q9Q3xA9h8cGEE0amtF/hYLjAqa3QSW
YzmThTO/KEL6qXaTE08IdHcPpsbZURWgTclvRkgHeytvBB9fu1L2pC5aP+VQt1sfavVxJ+uiTKS2
SxyUwH+Co4D6m7U/TK6OfjBOcee0AdXLwatBk2Lxk3YNAj8F3KnBHZNYbWY6We4P8/QmbSKfKrgP
01SfsqcYfKTvSRjuosp3uu6ZL5lJspOGbkYZ4FdUpS+1JMbVGcpJI8GBuBgadq62N+hYVcSp7zrA
bAMXc3vYqBrGa6d33vgpHFmqADQ9tlvYqzSxxYFV14Fzd5ZSR6Cf0D+7Z+EOwpN4/sT6Zl8WE3b9
XqsvVgdqOvWMBQqZjF6wh/yWH/mjjLVClWlsRFTZuE/wmHn0SuBwdsCC2hOo/ZqH176rI+fXq0XT
K/3LQJiTPbUHwwcMct8QZSF87sfLeJK2QZWCSXAJIrMtwZEA2iw3c+L3jYq4Q+bmmn6l8qcdJWMN
yiTq7qnbr0FVLFZsOr8qb2ZKlNvkMZyXipq5ZSAyFROesIML3QWYoBXAhd8Aa7L2acgIRitxryt9
Snwqz+klkrsFXGSaVtK6LHKUEOMi9aZxU+3a1msmJIh+gu2KJTufc1lZkrXvFDv6q3IskDUs30vc
HIhHdGo944tbC55WYpqDyKd84xfigmjqOIqTTfYU7i4xPIL3XnZIB+Te3REaMXZdMQWYnm9tSXSF
pXXHjf9SmWIT8hzxpVjXiSat5x6fm9UJaD92+lkCtbyEHuscVNLUKcflEVK5X6HkOTDCOWEmL5ap
QIywxLPnqSicN5xYKZ+scH/QV2sEsKhsPWwNLrAkys7gTnLTgw3KLQkEWEO+LtXdtVb6IgvBvq7O
UCpmW9Bkd7H+QsxPLmclWiRNh75VuP6L6gjPWGAtaFIVe5OHaz9vnh3e96bApbi6vqq+maAfndxE
D3PGCGqXpnBfHFamf5e5yGZsFplJmy3SZTtMmhP/gJnzaVsBrpAwXsLt4W3T2x8btEhR6PJkl3vb
o12wj06ldQUu3YgtW2B1YPs2Ip+3aYcihERJ9lfc7I+QO9WNNGF/U5+Hh8NJIJqMJ476WL1nz4qk
aActFjsW3ObXJZtsHamdGq4dDZkUDsFcEninMPlpJkjhZcie5ykUKNtYmvB20kEcPlTYG6Vk/6+4
eAuWVTWEJHcDlhqY3PxcgOke0bvAf8GqQxuR94yvQnkynuqsP8hTG6KDUDPzYsA/l8kQ5yqt2mF8
c6dPoAy4SI/bhyFGFjwZk9Nz0pnWCRJqOS33i9XqWsqRPJpMbl9lsfrLROPF8c4U9WhWlQSLkUcw
W6oIhiuRyKwREPcYeCwkSAWigj+sWB0QMduS+c8M4jkDDfD+wIhyq5JEdjLJQHWKS2wFaqiN/enn
1BZXCv8X4DaQHXAHGOS2ueGsw7kOWlpzvMIQ2YC3UKJ9zuSoS4s+F9qloGD78q+S5q7Ms6DmTdNi
Ayu76Ur9D8DmVQsKT0vVamZ27XoRYV5BUM69YwRddG+e2apC+Y7B9wmuczOcM9vHHb8e3XmURkdW
EX2PJXeASWBPZdQyu64oOfN4DGPOJST7S1DjCB2PzOJn5WmNaM6oRyA7olyuAj4f62D6WjgzoZYo
KyEkaxy3s8eCInh4/VokeHpTfcbLOaQTb04swCobP2bMRQyyH7U5AtTzqV4I5KqGF5p98fibmBBv
GOrglxZ7rFuV4ibXIa2TBk/+lsqouNMLzw0kZXL/Dzdrs8ZurUiHDy9a/v04rjy0k6Q824eabDHT
GmBRC1R0zO+W2QdDJuHuwkMDY98RCDC04JCgfAWasFAIPOaXuh6TZpHyXVnsuO4nF3JqyyhL45oF
spWNxCum879/hl/A/+9iTfKi6mEq2VxfkLbz9sDMMWySbr6scxynfOPZcZUtqjhRCgWVA8azqUaU
iyx0gR0ayEbPbw7L/gEOXJk4XS0LEcvCycZvEk/wfdL4xZ+WHDsfXxMDLpiz5YhZnEGBvC4uNcwo
XTi8Atg6vx6IY5ZkG8yp6AxqqGP5/Qgq2p1de9le08RWZnvQ6wLi7WzxlXnguJ83kpcEbjPBcOAK
Xp4amVOuv9HbAVU+cKE5TUr1yauhcMA938NVFAKba9Z6RLS2RjKBi8O7j8pmTxETVRuiojtN1L43
MmCUIIhq8laTYXiL2lubIST/u21eV9xCi3Rzc7G62viy16ovLryP3acCOtYjAdo6r5JO1x1om7S3
BbTh1xy9dd8zoad3Q+JLpCS0A8zUmNgj6LdkC2hacvhvC4v/0aG/OP8dlr7EpVjQakn+SJACDp8j
r2h8qGXkZSZIRfZPjA4lU9lF+7BSJ3AVftXSdMKw5v1lygo7ebj3ZtRoWgsEIllhfjSkgruBmr0R
iUbfVN2x+HN8uOcIllLYxNsADfETU+4GU1Fgzjwj6BkCkgmAsZv4t+u2IQhbn3t5pBR44UKh0G79
kpVkMImb3On4KxmxqpOvsrIG78AP20JkSQjvnu4RklENyUXlF6fbvdF4X0ASquY1X/3/JCi5M26a
EIelN09p6YYSt47nb1i1c2LWlOpE8sLsejjSCwstPErlYFVw6iEn9NDsUpaOB2QG0vSAyH31CsCZ
Yj01beqOlCMkV9A/EoHbk9ckCILJEa1DIanguwVpJVU7fwkYM7AAjK236eiEXTsSaR63T+ywsv5q
k34e6v1panRL4Vo5wwGN9z3+8cVI0pXGpD3Jm7TBfBp8Oi8imNVAd5rMoYycG39muNUWjGAnMPz3
8xutakg7w0irhbyNCcrK3MpG+WJ3qKEBG3pNDiiVIFZuVgKi7OsNos/hAZHVBdFcaWMW+xJzrIDl
7X0X86K/rFmKOf+Mgz5XO1kuIGPdu1NXFMwTkQwQ08rGtjSh4u8EtowioOocFo7G1J+cpjk8KjCY
5JltfSHgNx7HFNdP1ejEabXxd8WklYjQVCi3lyPKueqVfgonyx7/hST9WP/tEOhtqlmfyE6A9pHf
PHbCqdtWSSJNpbQ/aVx6J/y8kCE1/tepS/sxQzmiLfeRDmCCQYT9RikvlFEhuH1V4HW1q/qncgW9
5fN/FnPA7NjYJrtbAvoUcFLpW7qlgSLKA3cTiakY3NAgXNMQRW7nrP4kxn6ORfI7sogYURAjPhii
MYV4QHqW0yxukviQsfbv3TEUQvnLoXSp+Bv6L2TuK0sn18NHtLV5XI0YkevS1YyxGse6FD8S2rVx
PliUUZJm2AcYZS9LEJedxF4ds+rxUvuaBgFlXC9NfilMwgf8+/znY3zmgjGAfriwaAoYnycwkvRq
QnYLpQw3NLPhXq6mHdt6Ocfe3kMYAsOTY2OQn5HvC1/XemKuCivBmF6G6hL73sD3ponkBTZJT8s8
u8oGp57p5DU3dI0ARzXDP7JWqKLlRnhXC1kJPeYfqE1DbScLjpray6vhvpg2n/R7hwQaRBuBGIMR
EtRXrQmrHv/xAPMaPkmMFzi74twuO7lFHhCyUsrGGZQ2FL3uKPP0aCTiBj3BIw0IuIVxbgVetibI
rAnrlufdWRcdPklAQFa+olnDNSN7gSaa6RexnU8/imKVnvkHiJIY2Je7pYoB0T2f980Eqlf2ZgDd
nSg60ALZ8ymFYhENpxchAgcYsDcSjVDdrYWkEnykuoRBBsNPwxtUQBGK7Rr1dTrZdWLB/KATz+EV
KaeouFtPg2Q/aKWoEWL0TqKwEnhjz39NXPENovijd6Viu6Ozg1UccNUOQlePO1TPaSk2LEf8c3vC
QUezjbdp+hMUkQE5Lj2D1ZB47YMzffH++W0w59JzhhGQvUPSgrUt1pgu90wvIOsbBqyUx7RK+wfG
OvzMXZGhzKlLoeqNdEWI7CMNHrVJFpEMqdB/FkKUIr3yLWEEfq+408cokLpUbgc+g9MkEpYXHl2J
aLngJBNGlbMmEM+qARCYmCfWJPBCrn9PsRBkVcEBEj6oBqQuNUN3vVU2XNCjIFpJ6af39wvp9K+7
SdFoytXbQiujlZtiq7DUcXNqZeFfYUeNSo1RtlTbzlBNiWMcbihKP/6q7j4CNNfsZlIV45CibHEn
SK9XE643DpecJqwSkdA2kUWgPMrA5f+HhPl+61UMx022hrmtLb3PefBU9bu6SSuucwRFegUb+xvm
ZdCaKF5WHwhfrNC7SKCihf111LUwBwnz4eWZDiDHLPta8bnF66U8doVIWSVwuWfpZUy4pSSO+1nT
2GQTiUHpY4FjlZsLABRbLyqx2plcCxGKG9GyF1kjxalk7M6524XmBlMYPyRnTD3n6peMlkcFsM2W
oGLO+nuKaS9wnyK4GpdgLUUSo548ygX6AyNW5bhQzYQQRdd1de8RZcJaQ8Pl8noSWC0fMM5im04s
SZlSbwQja+HQrjfrEzzRVpV4Fpkim3CFm8wDXXGoYd16Wn5n1ZCc6ylLu1kEKeWSAiQL+s9qGwQs
loGKPy/SH6m67ADqn7w2bQCz6yI/LY49+xk0DHO+FJ76N+TwCEINud8luUl5aMdUzL7EC5QAvkmc
d5SADH2rQGmZRcvrO6Mw++tOhDYC6VVD65JdoRw8h8wkb/fJjdKhwPmYQZejfrj1cm2XfO3DV73V
BVb1HY3WcTsmOlfX2qjitipvHmeN8/oLirxKQKgSsmEaxcJzYD+G6qlQFqZFqm7h0aqepR0WxEnp
jVZUUS9rX2coClvknRPWffjQhKnc9B81SVKGhZL+qd4B02uN8Njl9iN6BoblTluwVuH9JmRvSixv
KhEMzXJ/D+wPB2PFNxgvR/kQl6dv5s011DcoN0LSCZoprDrN+zRkvKegr5ZvPEev+4SS9i6mucN+
UmMfC3UCBXrQFKq/Ns+M4L25KgAOA2BH40cz6GZOuYYps052ynfQU9MzAA+71NG2389fIwuw8r6d
4WFp1/yy6fwfpJoq0kSZ2ix1Q4EKUPvjei3i7hBN7c4umaP2Zhg1ZvpMO69w9Peji18uTEsdaHVF
1NId937JDcVd9wkcHdSLM7MvwzXZ+Fgc5tvpWP5RlNNunowjP0fKXA+1lIl6OkJWyPt60Xbpc0Zb
oWVXOBYvxa3HqBRSoMUQMB7mXH6yc2qTQ/G/N6OmXJqCqltLLRhX4Aa1onRvk8wiifS6JQ3k9dmu
wjGYU30Fhjo4KmD3xltK4nKqN91WB+Oo0CRtrMzt1w43SsUzDGAhN+KePd+sfc0FiPQ1kTDlPZ72
epif+jokFE/2dQu8gJKq+KH7avJeGr5RMAKMBub422Kp7Qj5wmbrv6HKzpP+14q8xrTXsMRTfyQ/
Z4u30cv4/NR0MOy+b+/BODN6Zp6suCy5530sb5dPG4GSWx84z/zdp9ZvhRDGCKBvTw6RuPiR+9r0
aGXddJLgw75w3/QddV7X1Gmg7ffdTurWG5wfyG+r+cZ4aDW5prGnXF18n8CJ+dTe+XgoxHDDXSvM
PJb99IHB/TPK+F4IQrfYt1Ly/TcRgqAcCddZTjVDU+tbdfnYy5mRqn7zu6iIn6UgXbuPCQ0IevCb
Ht7k2pu48nNzwr5J8N/yh9nqLt1YtolgKrKX53YEIKre/qWuVANZTWIfar+ra+gkeEc3T4cr90k5
ztxCYZXH+JoRue42QfzOqWjn/WIWfEtdTtGvkF/wwUYXGPWWUX+mRssSxx02BM3+rZDFeQShxReg
waOtOzKmBIc7f1sVZMSwvX4XSTKD338vx046PtlOijdcnPndTF4eFXN92Hy8bgY/6ingliMDRgDE
xr1RMYuNh7Gwnl2Z7NH5I5wfg9MCSOUUVipdzOZy0BprOeumIIdxtdhJVW13kHwu/U121Xg6E6ZW
dm2pU/NhmraeqyveNCVtaAuGr8aYOV9FJdnpTMCrljiGksWTkgdhW/RFm25u48QwqlTTkHFkxEIB
yubWLYpvPzSTNptaX88xNk2vbBTwZcdLhmlvfg7u4NY2ANxSZdjbno+TCT1DSF2XSWyw7hpaFe4l
DMlAAK7BbgmzbtxRxJUjq8drXqWdgoFWiY1y8My2OzNW/hX5xu7Q8gieReRd3yPIQXRgj6AmT3id
9OurcjDr8p/nU9AlpZ5sOUTje3+JmhhoPU+QXv1QMyOa71HeH+EQLfBpbhw9nQ0JV5C0LdXLCxeS
DhYH2VgYxm9SSAIjT7M+h6MMJ+eQiEut+o2Qx2hbW7g61TMuRgv5MdKGA99XQh5KUpxeKmiECACG
PPayyN0BDWIJQTUu2Y2y8EpS3I6lEz8btHTlxY9hP97fCRTdMsvDXnS6HSic3Dhtvoz3QOjuXpbO
XfIacT6fklcIkKYLzfqJKyrU2F5ZWOrad0NNrosw+jocItXt+UDrsLnf3kQ6GZXie6YLU2CjSS9v
0+9LXciWqIIX0dibGHbGmdW083MLUheJmnLMz1XgD0+3rpSDrGD+/RvFTyOnTsz9tAzgva0lQvbs
E+LDzr8qGcGNRQiVATrytmSgRnEY1wXIZPlCKrzpw06F2pffpoHsSEZIPCyxmiSN2jtXil/FJ2kB
ub9rOxeX5XUz7txw6Gze49JM0aEgQiSYN6nb6jPDQdStr5kP1Hu4kGEYSWumkDJb+qFUWIMlZlnm
xjShdVc64gVaFm5Kl1bWG0GUp7j1ABWD/1iKqx4luzVD8H5jTaPsLk065bWE7tCTZVm2a3njuzdK
bXcVGoOlmnWEv+tGQj822lAYWLPiuTjYDJIFn4GIGhByLBT/01s0mpD1w9jgQM0BS7UMW2KWPLrw
i/b7dwVuG+uZzc/4PHgoLU/fi67U6kSNexzOBAmdnCc4vSLZ1QCECfJDFXi53nwUhEIILf5doBHZ
GAdiJycZ/KwGvLMKBaRJwInE5SPlKCrI+PcVoaAold5Q2g6dwtEOOYeouH+Uu5u9DIdpvKq9pnBR
TyyKzwKpo28NvTX/sG2SgDW2mxrg/Sok3/1rDfaUIPDNmeCo9XREXMdQ4jVLvnYCkhiueVoj2qL0
Y2Us8Mqe2eavomAGutlGwVOArxX+/ndnqkahlDmz3f4BPQE6mII4V0hlLlUIR+N59K+3KFOKge+k
pR3rW3FoYV3XeNly/e14zaOdQNNEqpovPeLWgVOJgHkpUS5AOVvEdo9DUCxIJK1dU5Rq45ajm/bn
50qZqcX8wREtZYeufoujhiGtpnYePCedmLfaapbpvJWTZDvk066nsQTXuem+nlEelbjn5MvIi4Jc
eOYoJHPrMnJ0Xp1kGzumDkBDQw9oNBwSmGZLMuvlHqFw3xo/tBCIsrRd9QMVdzLTy4nuj8h3QIYp
0EaAIjLO2IaxuutvhrwAoyVpGJouNcWTRHa0+8eg9xKwbjL8cBXMgdo9csZlURgIWe+uFNU/8V/C
QETfRKHVjxocniBDPoiKyxKGBaXSnX6GLP27JAUB5aZkvREop3ep3R+73WQYU7SGFAn3sYvK6HKe
pBnnShRFqlg8eWdYddCvA2zWFyXMorWpG0JPq3O8oakCpgSgJVbPsmPmb8aVmJHY9xuxjJLQmt3+
CgFBhg26ODbOs/m1GaDHasAriqTTBuYzWWjheD0cMNVQXd7BQfe2UC/zIuCFuqB2omZRlnFjFQLD
8pI4lsxEYtUKNZa2IjqNl47lrv4OpjmtNodr3KJ3SwfXlv60tmsgq4wWXZyP/l2Vt3YvayVmJmJZ
HiBAyRDqgGbvLkOWYz1DorKK8bSYr0vZz2/lzc/zZB8rsK8cu2QS1OlbHesPNkOsSbM+UR4afPwU
SWXEh5hrl7KPZkZOuqbUU6PI+k/kNZeOuOCOrRby+qx+4aAUZo0eME2VEYp6sViqMwUdVIpH98Rw
5OcQghjmwLPu5a5RIF/gKH1nk4DsXt5u17J+2L1nxqew1kgQpRL6DJzS2GIMjkt2oF4CXb6YhsE6
jQ5x8VZp9yeZlRvHVoJF/qkQ6OaxMyrbtezlNwRFhxqNJSiwyzC5TErOXs788cX8fb/N1upe37B1
4pYbbcmKITsbI0xqaoPIqwGJs5OLqsVfpySgtOUtBCLjKTCLBKF68LzQxms+ySuX3chYmCA+GOye
jUGOUtxGdjLL1O+q5S9Vcj6kHpvga3TMqteBa9yK7Y+yVheCAJ4hGFR3ayt/pHEVF6s879xrOhD+
unWgrIusNWIZZcDh2jT70XtmUZWcRX5aC0XkXIuLbhCYTED1wMrCPAYfTLXpuN4uRrpJAHnorVB7
APniRjH3SslMG2YeVEMVxGGQ/lCvSLPe930NjqMCT+dXKlQvYq+Oa1bJTtY403uADDQh+9+QqfSI
CdJi0Eh2mV1oHXVYNmden1rqNkqRgKTKorfixzBV00p+NaqRw+6Vqia+4dvwwq9yY1RI+5x8LMqn
c8YJzbqpUj/Txtht7ayr76up17QT7TYyIpf89+opO1GUgMjLcm7jpDoAOvarhjc3/HMkTVcHavP3
JeP/0ZyqWAHTAaXga0CdHQ1F0G3ieBYpiQq9B/+UPD5h8AjFNi2Xym1W0mOxtBryxHCPwjEV2T36
uRummM/aLHAyDNCWHmcBOV3Y7BBF72Q3eakIvhiwqsvzBDklRSmzG4Zfm0TcIcAk3xwr8gmvAeZJ
tNIWrbCfSft5/6pqR7V7/iLiNEeH2JRt1JCRYUpOcCD9M5qfTKTqSmRWVOs85ctgXYHaRuaedA2U
ZeT6LPmpFYPwUluhV4lCeT5vt+WjEyBDhdVYDchTfBo+RqrOvF5UbrHELH5BHfyH54u1PySthVKp
7Luc5sUysIf6AYmvURdyW0eQTK1zYf8vHzVd1M9zghN0SjT59txwTiydOVYqp764D/XXy0rGHHfO
d0SFZ9Xox3dtv/LPsHpndX/c4cxRT0fueZZ37VnGe2jGJur6aDotjjjBinAFOpp4TsSFXDTrWQlU
XBOz/dkauWVTNboh0Fa/I4dZwCMRPxJAi9qc5fM4AZOf+NyGCXsAT2QITdErtZGPKa6DCW5MuoEe
5LIOdTXeZ0nDRYA778DnobvrUC6OwsAEbP4A1saf+y9yMo5Jb5W4YKb50ogUItASca7pWwl8V96F
wtrGXVZ0tiDxQMakmTEBvk6yRHYqTK3YM142eRsXe2+4HjsYdpQdvQkTbvoNbi2wBgg17mhxaa/3
pP2+0Ocv78//INNbU47TpppcQ9J5c7isUVCV/JwAM3/gOrjecQNBaw53ZILXlo/NzxP0nN2ey6uA
YORk9DDOmBT5Q++cnwJ7Vssuse6vZLXpUNG3nVvYbzHgn1o+V11QqJq4hL5aYDuiWdZG2qljykKv
N7tDOyn4x4jz4nK2ysdvVlGIeYs7xuQcK7Q3PzvV/mLqr/YZ1PTCziKSxJYaVxHLWWix/CnxJFJq
q3n57xfOCDc9A3s6F+kd1MRIdRDw3dUL1CbcjHSL3F4B7sRgAwqad3DtH1+z3DfIsR0HgNV9kHRi
bP6HGtUIdhO8k3yMWHJgJrvq/GDZKpHHVbh1j2odOtMFgKb8H8r8FxTVPWGqWuVUwj9w/XsQNm90
YJxJy8/rBKNxVCVmagGzPhq5hzFRYsoV86LIFHxVVxUPbSmLCudg+/WaTCLQ5Nxl5vtJx+rxbyjb
KYeRtMi9L2h6XfiXj41SjiUmNE1HgXqtHCOj99w7B2kZMywHcwT4+WBkQxEVaHaHyA5+aj952Owl
BAq4B5yJAXEUFUUFi6FCVgrpTK1tZYfktZaI0PIMPsz4aMB/HMwnr/YuWDjhUI0MBjWLYJOFzRXa
6ICHiFLmn9Zer8pBPm1XiDQjxNbq7jmnRl4wxGeTS7HUkHNLRUkHt2S1yqZyq5HcoVPGxNNC1JCW
E+jwSCyDKGp+WxLNLJUm3HZl+91dEQ9bXts8pLR6FsyTF88pR2I6y+xju2sap5MBoLEmor8uGlSs
bpvRBj955GLXoPHBow/dNO6RPNF32sgxBjDTDlHjLBM1yJNm8687Hgyv9kxO5GzL2LOH6dgqiI25
g0XD/9XM8dxCsuGiFlr6y7O+xyCk2IAAYzCh5Au2GhHsmXF5W+2CW+zUX0fTWjS252rN21GVsr0u
WikhaFDBcWBsi3H2LJeFISid5KF1sa8KfCe/mAxo7jGRrktYLUE7LrPZ+ch30CtVew9cezdChSfn
7h2C3JA5Tnv00gSR+S+8uzG76vUep7N5hRBtFF3gFQoyMe6wt3sSDcPPIjl/TFqBijSiWFLwCBPy
cD4iRSdYk4CTi040Jo/CTujEHy6ALOSVrqE5nE8zbMjAcI5HHpBOz7W/3IvCG0tTddyoB2r6xpN4
xLD98zayLQZTVnGcKCyWd7ViEhnoTtUl0//TApL0/bfQIVvZqDb/3bMGuQfExr1FwkkxEtNCPxzJ
1kHD+EKrMn6yEyCLmWZITfjW4A9XAdkYDpZyiaEKikZI7IOJdbObZC7Ib8dhhGfPnzLe7AGdsgiE
4fnwP5/vzhWV1bUcRVymhGJ6Kw8t/+tsG1vyq6kWWwSMgWXuIs76UreXiorw6uwWeI2FtxJ1A9QH
2VlTO00keb65q+zxQYdG3AVh9OlVglMJP24p1J4+PsAQnegEObKTIwDmdh5lTVtSf9QYua0Fx/Lb
JPhgKtNpr/Ji+jz3hvyCYyjGGIuZ/ivxmlSzr2lf9rlDSZxHC/8v5htBVlVFHtqUGpcoYeZXWLJh
154VRcp6FcFlvvjSYDZPELgY327GUH4+ZYBQhxn24+CkUERLBI+P/yOah7TjB35SVBFlElDpcRKq
TQGLr3Y5oRToalI1RRn3b4ADpaGwTfRUTXc/JuKqxEwe/ofaAiD5kgKgXolSM6RgyeWFPQXkH54J
Zv8Ya27bOocCjjOWtoIeqjDf3M8fn3tH74Tyb6GCPbysMzvOCMgc1E2BJuBlYIdGr1I8RQt5buN+
kJtH4pEZvHzH7Yecltz5Qx998EYDlTM5wkw6QSvyTamhsSkRg7StbDX2Kn3Fir01sARkadJk/4YM
FZBRCOdysagWxO0ax9494KZXCDgLY/8whjUFtq26a7iQtrId9qk4c3adIf3iWwzbPMPX9oJfITUM
P5czT8t8N3H36gFARcFn+oqk6uUNAVRwh7QBzmWsmF/GwZoRm5i77Wb5YIcitdHTCQw485m2V1HI
RB8l74HVPpfpCVmyt7Z1ZzTaLYeS1qRBCrrVn45uKkw/kjZdUNkTEAAgaRoOt4hdu6dfu03TRPOn
eM6p7CAP27xr5m8ihE2BToAaRUW2sQK9zsKCSh9TTmeRxHw9kAKAMVqWAN45XDYx/gIU6kmNSbT6
zMTYcsUV2pNi+4MvFTP3KQjaHZx+SM8tltiJEdPY6lDMLdYxXjoqmHJ5+HTzrcMDBz+uuO/Sj/D0
KbkvAIbFhKC36Fz3o5mj69mSLJRU0DLQna2nGg9MiK6HulEWnlb++4/5kbx0wc7rROeoDGUpW3MR
/1PFT2WkRWlr9yBpEruUBF8CeW2GP1b1PCuzD+orsLNowUmvR0N/QIKUMv1L8yPg2LmvVuLZjhOc
ZGPub9EI7NLIJ1SKI8d3dHaElJxSQtefgZtf36rvVuPNO4PO07MSi12r90BU4AUa/Jh/LXsHzGFV
DbcqLXeTmf9xXphjllb5OuMuBstwf3toGjtcekeOCZyZ7dj/x//hharZ/XB8VStRP/KYS6ZNhmGq
UVt96V2DX6KaMKVYrz8/g0jp/fWLiamz70PcZ3PAEuHXA2blJvGTifcy27SYT2lIyeo9s6ydKLbe
M24ZNMSbtsH7cUZVFwKa9f/VaBEVsb0goFjH2JNVQN8u5FS7jALTy2uQ4SpojouXKN8dSyqcXcop
/ABMk8GHPvlDsctpuXi0T29wi1dyix7xTVpBKVYi93KMVf0gVcOmWqYhdgRETzWJe5cB0KtbVrK4
pRROfyuAL6224Edts5V393AQHWGHVfszX3Os93P9ZNzZedIEktoZ0YXuHHiyEIbCV2w9Nwq0zbqB
PHCa1Li8rJsJdZK74efOOskdS6J1KlumRMPimkMLreiGlMfs3YufQLbY8nWS0rYoe/Zvxo200MRX
/dyBKeqGNmMgwhssy5/trG8HPJVUD/I/V4ZI3pyU9WOCehbg8OLv2gnWBfVFQeenkTcjE+asTlWm
tiycK/XRg4Siw8LquV6XexdarEEog3KHsF3rH4OObyUtPeGsepHrdFrN5mOYCKshWT3d1Xm7IQ4l
QwHd9cSafAlFA+MF5gSJdk60zz6NcJ1CCUchRztqgAOe2YaB+W8crS+VSuDBjL6GoetxLYjCK2JY
Q3XNBSzYGfBO6AXBEVcP9IaOn8edpsjTTqp99BL8cPTlD1SNEPZXfj2rAlugtB5IoavaGOa0nfmQ
J2UpZBzR8UuEkEs4+dYXiGPX6Al/eiq0qeUD2kO1gAi+smH2sP+j3ARIwjxQpbI31ZjFn801EQpG
8P2eJJd6rhyLgsrIO3B5GsHrXuxJfuvAUIVx1yyvUsf9O24mnRRk7hWtXwLm5yWsEAr3B8Vv4eYv
e+/hEicL1svfpW4VVrS1iiRqlk+l0nJ+7dczSP7thWr8rPXAZEEhEGWBwrGrOEXwXsWZECd/+Vyo
2edufuZKgJr3lTL7SLFbEzK5eILMvkLzkb4HcIJnGXxIXZ3IcEPpLsApxzPRSZJepIq3BLf1o1Os
3ymdO/EuefiKRnxdL0ULC+Wm26i5XMZn8YKzb8TqUiJjKZHZzt2uTpsRObP8aKJXoDQLOa3alkKn
6KL4kwmE+cIzVjD4OB8cjqeuvv9qWAJDwF609PI1YTlDAtxhnOhz5NdogKTXrTNSf9UHSR8Zdsde
67M4l3ykBcXMLAGcMhIaJmtbhE4tE/ofpDVpysV3a4RkVyk9xO4A/VuLSfIzXPa/4cHYr9zaaOKi
2qKIZrChLcTJZZvxw9fNDJOZL/akHn6UBz+oTYGMIkk2eMahKbrktVpZ3EZwuUd1h0SehJwK3/ok
+301bGfuufWXsrYiyWyUqp0tcKG1EmbhiluHbDW22DpiT3arcZMo/rJpLr/o+RKmrDTjlqNYwQ78
tGCe9StapsqOv8Mq+Ose6N2ER8+NhIQRA1wDe+F8h4BkaAFoQj6FOanxpvbG8twro9/KjhiBZ79e
G1HQSKTLzEGdyz8Lo8eYKpHXEmgtjTtXc+RBKA6K83nW9sQ/Jumi4PX/P5Svlg5UVa1O4dWDlrk5
ssnwihwGsRLLBb2SIW7NGUwK+GObVESEv2IlP7dblOtdlKWe1H2EDtMj2s0EVI9+bp0KRloqWeQe
b5XM+YF2344a7KDT8G3cKrV3mVLeaTgl8vqmjhROLy61Qt0sBUnnxCS7SP4B+VoaTPOt8HNH+6y1
X1tny7adQ4PhCsL6m3upfADG286ZLQSGjdSO0xVggDgE2x7YnmuRjLp/ySotIjUsLr1lZw89YGSS
+uAHYGdljGNJoxNsBO16M41v+olTZhX/ZCFZyeuX2vNjsYB9VaeSv2+NnkUpYzgXAq4Hdbmo5bnq
Jx4lKEgK3Be5S+5UAE/gulJLWfkDTVMXxJjn0+w6rR30Ij3d9amZ4y448686p97sVE3YazEI1VDm
Dn0FhTfibpdRiN/LsXU+zUbDjQIGBzuBCMXtEAfDh/VKIjm7jGOosTqXB136UKrwnHyZpx5puUT7
4ALAln6lj146LTTTON3gnnhx3/g5hG9DoHkwqXuFAs3RfrEPZcraiXv3ZWK5IPpudlG+tcOWhowo
AmmVp+aR/pP/b0T6qGq4MSYWkTDIES1g919t+SaIwWgirkL5MxMMOOPqS1QKNjd8cPYJEraBFVJv
GlKvoAjEq1qpiyhlJUM9xOM9JLzNUZCxSEPMIFAUwR4grhd0ZYqR5cx9nGe6l/rYFskFrQbVskQs
hJ/tQyeCuGO4qosFIsjIZ9HejgL5hl3Vz8ZQSbICa2AegTce8/hKryyVtyBJZgW/5V3nVw5/lZcq
biM9Dh2M8ljC7Uqrsjwi6yqNvH0wMGTMVsiPrg5aS+jfjsnKOuTuu57Bn0hNXUHAcaov9LLT1ra/
Dt64fGdImxmOtxyH1/F6ZLzhd8PiN5EqGAn4fjIKHxhcb0zMs2XjXfKicsp0fzOX5q+GcGSOo7Wj
jNmZHNauT02WtYoC06celljxNncJZnsscxbvgHKiRMSi2kXgXvGYgBFE51CsN2ox4L92DONui1DB
bhoC6XuXGzpC1+utTYP4PXnTwtyX34b+RsiGBCBc+s4O6nYKRg/R7zNmKKlcg/cAWG11ffARi76Q
PAvCIOKX97U4LacNi2KYP6ZVxG7yipK4898+CX0IrwIqehpRUmWmi72uoF3Aeg4ZwZV5oaWCYtLn
72bmLxCWCzqlUB36FLxChn65XD/XTCqmMBnRSPep7QMWDjXd47OaGB4gJ3GTgaK/ir7EU+vAtERv
TxkjyWASFkL+Q8uTGLVAbE2YZ738iKl7fVBFN9bmCoQkw/gIaujnGa6kSB3/cZYSd/gd0HawNej9
sEK+7NQzlX6OMssFmkQbqbXdNO9j2opiWI3X05oKSoRz3uFQj6LYNxu8eeMcrYIKxPFVL/yW1i97
XtvOyBkZ9mRp6SzvASEFaDg7CUUs+FC8SJTLwmc4JRJWSXUEndrYAIVZ+PJbpB4BbY8B24r4mOvA
lNEwv9TusqPIfoGb2LX0aq+qfGfoF6cr/phn28+PrSInm/BehN8SweuZmjdgs6VYUrPYEF67qMYN
jFijaiwOyd4luFvxlTSYXA2/wNfUM1mJLrOx8mkc/jU/Szy4DEKjsydcb3zNn1WiwNi797/6kV5v
4M4CKEKvnT+MpPgf3pGN4x3zFGyqVKvnrlLxFeUXMANAWcy8dq3ox3mWG818IY+Ex/3DptvC1nr7
pMAY3/aNhPrEuI5rsgKetvYrHsf1gpQomVvWKJVMDqqk2PH1IDtefc35VZLHlk3ExygkuT7w5R70
nQ6ntU59XNp5MFCgn/IPam4O7n5IrE7Uc6EakqnpfuTRTwozO4aWdeWB+siG644ASYHlvsGtpkdm
as2+OMm+S4OexixePgixRc64tMrK5qSucOBKAfghw+VbQ59xbk8zuJlzN2LZJbMgQWqZakiHJ3xY
3s5fgqlhdeE2ZevhJ/0mG/aaUBKsG9QyENyqrY7Pxl1hLXna9NRFpzAOSjbLnXNghtQX9Cm+37fv
+AnuspMK+7SIPA4Z+CXulej3PA0eU+sx1bNozz0i5hyz3hMb9TQxIKLm8xDeWNdwylXaEftYHfol
/eQpxE4CYViAb967tuRubxtsOa23MWhZ0bSMe0dDFtN0MvIhAOqmBV4UR3KRFSWAe7kgthunimzK
ju6KQAUY4r4egV9hOZ7A7Xmmm6ek4N4rSLFFTeIpITPHSMGOeV2QsS+7ni97m9fwewY+gHmyRIOr
RDaegbAskVmmds687nHaLAOwR7F1ma23NqXbpESecbhFUxwx10Tkrkd8KnZMJr8SQxfyJSJx3YhC
V/KuDhxGN6KANZpaN2iMxLGAZvZO+9Re9CfXaSgslIwXIsvjkSBQv8QHBHc7lz2f1HA3tfWiMudL
mKW6qavXDr9TKfknaSxRRBhc6zuDrcazBFtWgmwsaQprLKobT9j/vAK30s+CKprT857WIVaEeoyF
rlBZdyhYYOufGaz9iv9/FsBOvd421C2+idYzKMAVvCvX2ZT3KLLmjhT9C0uIpY6kfOKZ08rigqrt
4Y8+8Xoga66sqscrLDeznww/mQBZFhyI/4C93aIRBa+H7MIZkW4xACal3DjCxJM8QAF1u9KB4Hhy
DaI4HC4sewDRcbOpbz1XnPcaZodt68J+oJ6s+Gi9aEWvYGhWYlTJVPXFWtUjH2A//9UjoD35xEd6
M4VVWtAf9dTIprZxCrYCzbFQNwGzTWg26v7EEhe0HrgAjWi4QN4MUVUmxOxrUGDd0ffEJidq2E/o
DrxPcb3v2UXts6LJW5Jf+g+el0oF/zlFlHHlvxpAl+HZcKW9gcOCya9a/NRH19LYVhjEq6zxmxaP
pW2s1KZWN9JOL59jI2PqcUPDpIpnl7SNPa8tsDFdDRHS3h4f99Kef2QyDArTn7rK0nJ52BB2Q2cC
YioeqBJ5EtnPGLjlPoFfvAVkahhbyjtEnm5QBxm+OAvZOWzwcueHqfjWbhCAbRDA5rzSjelPrvWi
+6rd0YHb3+S0PiSkeMqZfuAb4GeUqkCecFRy16Myw+MPNtM9AUjRHHZZVkNnCxURUmuKqWArpaFW
kXHMYxFiWObU1z2bClJ3tZxgFBpoudrnb6s2hvKflYyXUMGQWbrUatri6Nxmvd/GzS8oiM6XrPBe
iNHBzArMmRyteCCDXtKLmCvAIgEwWL4fqGHe1AOuLSwAylCmwYws6n/13KQsN3rt1SI2/RI+Z9pP
Bsp7AE5fvC8tOGFjwDXZbM/qS4a6ayG4v3Wy9eKqnCAdwALkNuPIHn1i9ZJngh6r0J4oI0LClHqT
FEmEBbatGbGK82Mubd8GA0tZZotMB5Z+dck413/vUC+ARqcEeOv/g9g+lHBgIwlOoLQTP100Cg3h
0tMBaw3lAX2vOe1HSLVmS+cZpLm+HtarJD04D3efNn/rHuYOeMaXwcxilWpbjPcg9jXVNr38/N7g
pfLDWvfUKe4bdVVGcjgX2sN7rgfQAwb3PAhpZGRCikwogFcuClfgdo82ObvjaNkW2Y+tKiervsj7
86X+YNVQuiq1NLJrAGTstM5W42K4gW8/nF05Y9yrzYR6tpMnrKJRzmIAnjJd0O2GLrKsSXkK/C86
VEwbX6kECz/dC2NHL6H5drQzHK0qYefE2xf70mkjtjNqV0k8/9OJ6ahzNOnZclz08skZKF8DBn4I
uOCvK8IzgXD03O0018csz+FPdUbqBT3APbOqg+XbIo8tnuXA53jbofTkHxSr32A56LU69fp9vYPJ
xFZkqlTUfeuO0bnYPPKveXAmDWd6gMAJx+c8jjibXiroJy++3Qq023vYcRkP45T8PKkUEdGw2viT
Y9szXFk4SBFNrlOtBkT6EpE2p/A2cI2MK7ERFdusTjmYANNVhUzRQ6ngRfKJ+ZflNpo53VidB1+F
nNirpxrAhBQodclLN2TPYe+m/T4aSLPg46QoLz/Vd8QK5QkI56gztUJYcvxLMSdCRikN1SOnbzEX
2ytKGDzrfATF+mrbE3psUN+iOMpWYIlAq6yIHZwcgZ/325odfkxedKZnMPAhRKoLJ3opp0X5VPaQ
mEMpntJKH2CJMNsSqN/UHh0iGjIpFLOuMISQsq6odl9aD8hoVJlCPgfRNeQf1I0fUDPGk55yqrMY
curXArGw+9tV+dwH0gPjiTxjM/W6smXJSYVTGJ42uh6On6zmPsOVisirZbcecvU6g3Fpr5iehQzn
Z67EyQwONFG6rltGUZekECcNYOFMl2XzNpVarj/Dewm4HIk56FKW45H5quIrgWkoq3+KvvGh4+LH
I2tbJyl1cXSi7q8UFnYhR04g3px9+oy3t6/zLrl6YoP+eIO7EeY6pYxfsEo6SHhSIWcVx1fx2Lbl
Uqxk6m/cSSuMjWRgFsGdBHg6j6Dg1Vmq4Tpi0m4vOmJaC6DxRu9CjOwXA0R5p/gf3GlfHOPjG24a
jCOAx/n0h28KzQOKydBzBLOizZ7Op6UpiWhn9bCe2r897maNoiavF5mAdkG8NKRkhY/iISJTrLZ7
LuS/cyjlCjT8bmcFlfyaKduqROMl1moLseb/qS6yxE1SBuSWF4S9i5EBKCivP9FstbRRP0Jqy659
hkAJrRXIFPEaxzLZvL+t8ZhuEcYnhJ3ugZzjtdMGRqCh2EZ1BL+vzfV4dedUzAoSWGJ5ebwVEN8M
67vE5y1aOhQHliNrndV4XyYyr6Ha6rt6cCGDp3cVLUxP5vXRdoO4nXPbP/aAqHAduATrj72FakiF
qsaX1OcG+0D4OZHIJcgdSymIOipWFEmosBz1G05G2FX21g5FYTQ/VnNwQ57b74CRYz/Qd0A4DGBX
vD2GI08b4BkcNe1PcYd6or4r9hR7wW1uLOYqJ9iFyXN4YGohC47oLIIvgNd2cZS4+DCcHVlAUOP6
iZi6xhmBd/k/8T55otwfNjy8ius+P02Wl5tPEkZ1q7f2C2MM3b+unClchiR04t6VXc3Pu/nltEwB
2dXdDDSTIduTeBS5THJU7E3Jjk1A8pWha+oIcNrVxfzxXWYE64eiNujslRtHke+IQy8V3xJU7jo2
WSLWf3C+i9xVAlC/scZ1M+usvuXmDrHL5GOTbL4D2STHZkmn6psxfr2vV/IupPoqZPFAwxFP37G2
vCD5PzgZ1iNLKq2ZZuVv5zufPqPSOVDtBOieU2DqInVze0HuBH44Id9+UrMLdUGsOv/cP7EjZcGS
zePe/isSI9b1lOjLQIq7Tpop6R0AKxLGHY5yoaPbuba5a4W4x01Lywy7dj9w/RY/oTbVQFam3b25
E/tZfB8meiSgxOWGAP7/GwNwR7P4hzjXWHJD5vVf5B31N9ExnnIMMxfoiXrMwFh99Fw7ZsaiOamf
cNgobx6B/SHdHhm786L5FwW4AWInHFlEqVDY6FX6xGJDhXuRjaqDAeooyIgpTr2yTkgkiuFar0Mg
SrXPOzR1DOTHwUscm3+op5PgocKqLmPPapxEekISNyu7eZoPjPHSc5oG2p3hUXiFEzGQyUGvpwan
Amzmuv2xJ3XKgR1EwOvgQ6gumD//g47yOhd/vIpH8bz3w4plQMquNzLKcoSjNr/FBO35z5xI1C6P
cPo5rD6gCf3aVNiHFRGZqLfz0QYuMRQ7OVxfQVO+oPl9xTvqRI46GnSCVRNs9qRr46W2wI+fZSEo
RbwTRjUt1DyQHWp26OQq6QXzr2PWlmQFQx3dxO7Ca8jMqSplttEH8qD7oH4Wi7xEFC9UiFnSkRAh
rUNUyuBQPDu3f2Zy33kEupa7/hii0jH8wrYBLSP2OeOq50zu8MaqLZJaHzEeDZQXEcErcuQgEnYQ
ht4GHHE30E0jqXXwvBIfwXDKJTHk2ZRyIUkF0qKpTnB1k/8kbxUFPffnetP5Qj+sArT7RW0DZ3PM
ui4xXjEXfQ+7insyDYO6BRH4DAvo6IOZx8EXBR9Zn1LHkriWfueXY91vL9tGpyi/DprCy8klhEwg
v5RxXaV1++xJ02sBxrcAFmmPN+HGU9l8I4Y7A60YxHA/VHLImCfEy7jCq7pnLNSUx51wKixGIFx4
jULHtHF/rtxQ25E1ByYPlsMsTk5FMFEqNSw2oDcHcqfX7NI1dji8R0T7/hmr7QOvf/ZWTCQeAYcr
qojZibmY1PVoBVMG6al/9u2/YOEUqH/d5xZi76MlaSjEEoRtPsB3PJwyQSUApLBQcDhfgBu/NObP
+JxU2VoOE6Hw1xei8L8AVSGXq5WWh4Eb9tddnoPxhT0SJZrYPj/n1MsNQ2njxK18XxPlHv72bSRo
hDA97tm9bezeDIcxkDnPU7glIuDAbuA1sHdUDjffdrCDdXqK57F8U153vNR+kAXwe46MDRqycJOS
Ikv5naT0diRGcShLsecksJh4ykX6xUXOjHzPFt8O1FXGknlgTSCFidCqLaPuPNz2jAXCoWKtHrQM
/CRlkqYeTGGe0/tq9wy4d+KKdRqCjFwXBtCMzqzmZDy2FRmopVkcDaaWoyOLV0zHwXgyfHUi6x4J
f82TnrfBychNEdng3cv+GE6908eX6LYK5iNxL1Ua6TCTFJfE3rBZ7oApQtlOrYE3PMsrtphGs+f5
dOM6Dqr7LVY5wQmbVwpGSN+ZQWGtMOYl0rkj3wa1wltqehw6q/okWCyBIQ0mgo0kVwf3LnvRHBKu
LRoBEuIYwEVRPF2JS8Dvv1C9waPsyF4Hmevhg+hi7VFRo3R8Q4Nq/GU0AuDnnLw7yWZrZrxiWvTm
ejkGWAQsPutL05iRHddznyn6fxx+48W3jIpan5r3zZeLskmscKYn7EDszaCrVRGo52hcjGyu6cMt
W1AMOYoJywSUY8g186/Lo+rYdUrgFmXbEdRmdgBqia6gEVVQXvpdn9BuXIG7uHD7lFuRy97hWpqe
bNS6rXMsJFOl11Gways8dnaT3tcsuer0IEuPZJwO3PmyHlMXmTWL9ozWUoV+weglpIejXYdXTx6J
TJ3fVTu89r++J32fhhGg46XjMeUEq5nmsIcvubm2ZYZChq3dv1bgvD66z1vA+JVpBfmjNrvi27Cx
69wKLX6Sf5I1xSGRA3xzdZ9lUiREMXEXnD4k80Wq8NQ9qYfIs3BBizkZfGPhWutoQ95kw+YqbFx5
zkoX9Om3H4K+lD5bNV11F55MeDtduDDL0JRN/bPkmshiUXAD3owIVVz6HZfcg5Gm0enC5eWLEIV3
bC1LYe4AAwI9PGMOMuc3tBkOyIs25+szP+O46z+zEs1tSqeSR96xV4U0/pRazsJLmjmo4EYgoREr
FzA5DcCVnooGk43DcBzoktiuN8b/Welu2pMR/ZgIlAKsy/HHYHHrav/5Hg3yV8HhMrqCis1LJQ+t
CaaIytaYCFVEUD6mJiHxwJPs/OArDSbonS7VfSfePYtcN9JdhQvZ8w9qrAD39COGN/OK8hyLShec
v4HcPfCTEEhkz4QwFRpNPEdFltirivf5K5IHUXsiXpYqf4/nXKbnKH9x1lKnT/MujxG49XjxjC5g
GSTywK2EsnFTh9f2dGaLz4QH8O1Wydm9hlLo6KrmBKiRbQwWlXmCwK2SP/SrkIYw4MNZitnddsUI
eors4HY/rLwaYpaBs5EIzeOFWLH8HrF2AsBf/RNBqwHFzMWSjYJRVx+InKKoh/RJZS+jU8Dlp+V0
kJjUoQhjA0fP0W4yqQ8UGISs1njZoBNusov/KIJfrvVVXtNy7Gm6esVir3n0hBDvUGNI654BIWL5
Np2tzgOp1s+JDSmOfDfl2/nJI5HPmqXodibg0VTR15XPXalIGn7o7E/bMfjOsaM4pyIGnc4xioin
2SyPJKA31wtu42jsbEcZCxEwxlLmlB7ffGKd7cjOz4iRNWq7L2AZ8xyirsEyxLxwOFLk7C5s3ULH
gI4m9OTcz66MW3Xz6TtSUXsbmE9gcE0KGCIgUKlgL4vTglPd8UeZXHXALO9AezD3oykwZevbxK6U
isOQGBtWSRwJDxef2/ABxdddd7LTyJp6aLuFsQYlwxjmaa7LQK5DO1Y8oy02fGEuQCHpo3pJsPVM
uGWxbsMpkzedcTUcszhQan50cXfVIDcrIzKMImwnJZYYIOOKolpL8KPdwIv0gzjofuGALJGK6Plk
fG1fOOZHI/pT50Y3XPQpJSp0dAc6TfFDJjUkqiJvD+Oz+JU/SWVohNP7c5zvXT8QDM+y/kUQt+gH
OSWs4Rjzp4oHiLhxaAQuLGPWLuhJci7+usJ3W/4dhV4pmmCnAsQdDbIRrQZpQnEkOwmyivFePDW6
xrhCnHn54IpeTz+aupjUh/z1YnZe7FKEyn5T0Pewd3CSqlhnkYCw/7Q+kaVcIzNXtvIKRA0j+Ud9
ydVeX4ql1gEdOLmsZacx6Fo0g7lY1R+VtkwLEdce6rVVp1YubPgDasYc05slyPuFozmEg5JfCeHg
iF2QKv5WmvGwGpbCBGVU2iA9kE9TvAZYkW7Qk9krTf62rDx4gKA5I6L2Nj7sqxj0f+jmH6DJEl58
yuNcs6Hsp6S5G8t4yMlyK8ML0FqkoIUdmxBR7+3wi1ZFb8ysT/PcDYSs3nnF8sp0ec2kT7Gdsn/t
0IjRwVAKlhHr8QbF+bY28jT5+qPL4KhqS+1KWq9ay38Qaf9NjHkVi7wMI3TtMtmrk/sKY1K9g1v0
zOvH/Dn+FkFY2nCTA6LxXzwzQxj35fBDzJ0ufV7X4r7x1+q2BnepnbUJlnpQkra44zL1aYK6duvT
0fj+jhEQJY7ZWAYOlaSMhz/bR7gCYQgzEqzfjXWTnjavKET6C5/k39FUrgXvgAUF08wqih2XMLNc
ctLyrAbxDWKNXLdVAVihmePiWFLwFnBsdQHEgUYzHgFhLptgz707gTqPcrooHIKFzfYpMuk+SqRK
LdWZy+tpIsuOAZWKmVwl6TuqonOfuYwYXf05+cPre3/Eh1x/8tYiH/oyjGKDhYIUwSFplZDaM+xq
TL65YiQsnlDyQfN9ibRyNBoa+yyFUWZqkHyEcLjj8GF7Zkq/Jh1NMyTw7b++Y7M3+DCFjFmCTZUp
IeVD8y4du5yWvOHcscCAVh0GzAje1oubwYjKVfZHVEds9xxXiG2S/swI2EJoYm9hKCGrZG3zGH85
ThNW7ACawjZgolLfv1VqWKudWxNVcprcvj+IBRkLuY1Ebp1TYzZ9gotUzwkJxfNAAMqMRIB1ogqz
/12M5GYaOEcY9D3pVh7PXQ4s7KKdyRLbWJixG8iUX16oGOtqnG7T4L0Q92aFRmOUXyiDqDqSr7et
l4F3zJLdoSOMcGAFHntwe51cO41ZY4cuc86vvBlCNw7OB0u01JKl7L7s57IqFhRdrbiG5bE9BZ4M
rnA1Nyn6fkS82m+3gnh7CIWFeGlsfzHlnU7Sq2aNVY469vW2iEA31U5hgZa+/+bn9FKjyJj+krSr
g0Ps/WIE40tPlZJzRB/+ercMJLSAdL5dMtwQHwODa2OVI226CjRaeTXCaOu7NwyWQD/GkO55jR8I
loJ3vGLEDB+orCtNoua9OF5hwQVPWfdvnRcKiSRBHDpClwiEUTUEgHHfrKsiMko27niPBXoR6Rgo
WTMEmxDI00cdB8DIrCu44HovfsSCxLZYcTU612GbImgKlNh22R946RfJLiVzObKz2Rf9Nm5LK0D/
lnXqJS+zOfjZO6hpk2RiEYwIQ+IG3V27m3lpCIMaVQe/Sq0N6rlsu11s5LM2PYE1tB5/B45trlaN
vX3/I0f2iexm3LxMqkOty7ehPkmbHSPoD2lnaSTC5timMU6yKrYPuRAUS6dzjftM/4mYL5+1MWRp
naMrL8+SwtgFVQII4WiExff0eQVpB135wSHM2SziVm/UNsPGaN4Jos1Vkx/t7c+EwXzUtcbJhCxl
Jqz53QUdcAy1fDDtELwyVb0Sg+pJeyWPErh3UyusJ9yiWFcSOtDGtMJk2T7ptqY/rOTJjKjC73L4
pr9KPSKR/eG59BpDqaSxemu9jijKcEzO6Ep4FOIKELqvlWBXhbKgq/9q0wRBbIsdKYnPuEkg4ohT
93zYumbmdLE4uB3ZcfHaX8uW+0aXImYIVJNx+Ed0qIAPjpmEWVn3Y35GTRy9naZo4hi3ejdWlXYy
6hOm9gFiPArAKXPxmC/7yY9yXft3vnMPAz7tfgV38zwRI6VNOKWTKvVwdhMTyLU1qZQezaevq/7+
D4ydtX3VwfSKpIbwGPamYROvr6aFKTZseJYnxI4fZ2P9xSav5WL1+3AYT2b3DsvngW2aW41meug6
8mgKYYBHUQplmCzKVwWsfWDayPGy4qsNRqP3spzie1vMj3GJ52Vz/eN6Q9xREA79bh5IJtb3wlDo
BrYFPeOZmhlWBM15Kv3b2C7nbeu2uB+LaccdXSLXBMrzCXWJKWlb7ThYVqgx61HBpeNVn8672Cle
EsywZDK26mtd7kwRESj7gX4lzPxSVJ9sw3+SIl4PdHNdZs6g5AdO9FQ6p1jRsQYwNdDRWhhCnuA2
ICmA+MRNJTRCh0Sbhr6kSRu323TimNZHbnyq3PnbhxB4EvijgZSzlzf4qXIotp47ht12opK2l695
zpTY7P13r/23DhWEjSFRIZj0okss7hZshdXbFIbMzELdeCXeCfYvvt2mlYw4HRGF06W00qwGpgt6
IZpiktczZipTiWKCEwcfr/Ip1jFuy9KqjIcHczB3Z6L3Ri13kk3oJfZL79SCpFvOpVzgKxny1vNx
SNVLyuGOgIdzjohhvqXez52KuALWepFAhecF2GGYUc40zLuKdvErZGQKoT5MUw2Dyj7yYyZavfjR
fdWIlmS5jc9sTcNjVRGQPPbGGZzJ5YshV+iWOVAqEkvyyuOM1pNi49qlkR0EADxUteKzIKQAPp4E
J0PDWt+604kUx8e1yFAfUT6CZJKe+i1HA1U1eR+cMovHlK/StLK4wdPB9QfzVwlvJ+vUQcH6hzmV
sOkuF7UwXaS9pPtKSjtHX5yse8FEHQYfhTQ5phQfId7MZcxHZJCgsGIUhg4cji+Epl6eM/Nnala5
AWWatNoIFp8tZIGv+aywujUwZEWw6Dbpb+xMiLJU3bQePRXhDj7XTvDA3wJmlNU71w04raAC5adR
FG1x/6i90Yu1k85G3+E4MpF+4OxfeXw4GLCR9ufhAKEBHed9tF65HtbkU6k/dLmWjD4YX07RxIW/
wDi0+06VOcNE1MXciRq7hpDlk3Yai0/CO9HesIhmcy3myLIjcvv1FT9VoFzgV63S0EkIQCSPMQEd
JpIA63q2t8r5CRakNFXZCwLlgemmQiKv3LESo1imv/7ssAkOrpxtWkar7W+cxIuOFTVczQf9zSs0
XqXYO84/Td97FhLhk3e9iciRlZzXxgJPnkxRMM+PstmiMqmb+oQITfPXPqgLnhDpboyCDI/cE8gZ
4wzdiMIVv0nuACBbdF7nHB0Ds6TOLfgWF35dXdGHrut98hx3Quoh2kYzlEytSQb+dK4yQ89W4lAF
jBNTWKp5gPCpIhsv29mHLJKIBMv1fL/X9Z9DTXczOBEf/BY/HenmaV1lJA6YNxKA0QMJwEU4fZKz
VBeXjpzDuXzcIrzhrgi8kBKH4LqM9vx2VEy4Fs5S/L3dqxYNa2h+3Nu1wXNykmq+GjMj3gn6qKrg
mS6ZQvW+1om/3rvbfaQngrGtV9vYDok0SZz9oF6SpCPy4p4McI8oy0GANqOAMxiIIUtY10qx3jw1
IYp5saovma+/NU7RDC1cyys5x4JK2K2whzOVAbD34lXVJ8BPO/s4MwMQwyX9vqCoYbL5rIKE1IuY
rQ5lE6KyHpFiESvYW/lE5KP9CW7ZFGXMxjxkwcg+RDpkeNnhg7XqMKbpWqHV61FzQUIhnua5fhSG
xZfIzZW4noHIlVeOItaDX8mMj9iE7YMSBmyrZhyduyz5HfvyrBMhptb1JFk5SOJ9igPmlYSnheIk
27Llv7NPZBumNHPXsqdDHFR4DH/JmfjqvzFHRET4tWYDbPJL08UKAVUUXtBYyuNJxJk+lQ0W8pN5
Rntu26XPw9O957aK7iC3rHNCwAt2IZIFbJgt6lwdAQr2phK5yGmGf83eYWlROepCUn/4pEkdTv5f
jbtIDYWuCBMISy1Cu+SqDrzDiyrRtogBBzZjgfDlHvILb3dfloAUNCm1Ep8XPIxotEL6w0S7jD83
LQ0++vGiRhMd1B/s4r5VbL4bazGodpKWZc7ksnXccakQNyX+VlSIGWd6BT7QUosKu4hwT4s6KUKd
b5bn9rm/beRvB5J2wRMQ6x0Hh2+Oh2aEC1C/K2vzF0p3NozV7fcGzhXf/Plu7X0JoE0Zqe8Rs6/v
3pPK9oTYAZa0U6Nh8DEMnJDewCer/squCexXXVA7DfIN2Mv2MfaVfMKmo/Uj2TywfG31NmODinxe
nkpRHY6Rz/hk0dPGW8mvF0sc0PBVDolXQTD/UPJdc2BbspZQnH9wYoxM2ux/TwZdvEGSNWoDijM5
MAZqewJwjvKpV/dGwx0KYIAzxr1ztL+IBCuFVYK2wzFWNn45VbWnaIbSuCAh8WXj6Cgn3TIKqLfe
UJf0e7qGUjRBMySxdnqzxcQIMIEl/KKSp6/MyMQlSRHT29inu/P1WY9kWlNKhC33FN1r44i3Umn8
Of28xkHvjaZHrS1Hc9MK8dz1qvSzXVPz1fKHUD7p2Qc+KDe5nK4goSYJvvswxLRiFkqRsAhUndHm
Ph9c3dIXSHHtt6nO6y5RsYq88QXb8CwPSWkQdUYu+9rTNDH1cWQOiKDhqFYiGgyPPBOGNow1VgEZ
ZxaMdubyRlLjIFOsFTnXfF8E2gKtwAiN+GyZ8+0dt2pzK8d0VW5Q6kj1VexcAOLNxv391UnKgZ3Y
bdxCbFmwinKvY0alO+srCV5EKuYDxkHynt0DX4xq12cHmEyERh3BtkEy1oMzE9yNN5H25lu+Kkz9
vyrk9qHdtMxwHk1PUaiCam6YNV7BNkcyIsXAQoBgGKMi8n3vB2Ia5cm5PFjgrW6kJYzPhlfy6gcI
5DguXdscdhfBLnixNVxBsUulKEySTfY7QdP15uSZ+1PCXeilHU0lRzqGPXoMzN1d9/O55sCraU1K
Nf29ew8sMg4s0BFfQKquNP/nsWPuMViz/Q9P+Pmt+eyEQGO9c5yD+FQJ08CLVjQY6tmnfa0I1T8L
D59KmNfJEiSyRgvDPNf56olt8H8tywn2w/wV8oMb8nrfekiJ3aa1C0GqNm5+j550tWKdHMLb2bRl
lga3xLfARXRWq7bm23SwZBxcq4IZQDnfVlLlpYsyNv/h0CFpKIfkmh6uvTvC5s5v0HnM9MxvMrZM
xo3ThIyEnTEI4TaKC611dINa7E69cnQ//EITtCj8hMzDZmt5XVx64BkPpourvCjkHylAMv4uE3aP
ZrXi7OJmzDcRfqOs18d+tXqa0yXVcwSLIw0tmadv84QqcKBVXKoqSHy2YM2tAlE0yyKMozvEd2oa
gpVDUeDmxtb8xdzcSFnCUEhEE308o92ZKfajXwKPC9PhO16UDx7oKejA1pHVwzX/Z88ap0/oOV8f
vBX+YSfOCX34erYKFsNy2RjJEqd5yahxiq8UCmwlTnoApuuPFq1+lHSexhxxp4MMNXbp91pUzNZ+
ZubuUml/T+20anD6nNZX62jpZKGROHVNI8CUKlacJVumi0yh4wKda4eiaWZ1bJoo9o7kfv391vSB
wJ3Am7MHDD2Wr1EhQizgxfmWT4DhOICyC9cjFDm5IdV7VS9iFEucYceMOOb2JADIQtjMi8ijlibH
f7ZpNgGIYXtKjdqfopkYgyNORU03nVIJ8cxWPHssokkypL1sJYKK3l5PKYWr8IISPd25Zviz0GCy
m98oSLE7BKYx5Q5yDPzNE7l/60QTLhhm2ZKvrhN46GaNgCRted7LEhuWPLLAduJhZ/WdnJRz9hST
2aVh6vqkm06kqDzvMAjqiQ5LZURorr0tUKRN9TC7eIhFms4ScwGpQxi8zi9gJJMKGUcrdrIeUlQq
W5TMAkrCm84wY9dtkrmlvLJy0W+kbzLirJ3KhPt2L9ihV3VmL2ptmdYulhYNiXFTY3QRdZgLJr4O
Agy8CWHlZ9SG7DPt/ES8bEvmUWkO8IyynoGk4Qd9rnJx7v+GF7p7kwPqg2cfsalHALMXWAhVUmhD
qIB9RxCtBXlRuVdmBHhjqReM2rk9jjguMJPSPoWX6zAbgnxfm5OCpvILOs2Ch09a08+ECbVTjd/z
aa18weG5ylFPAyPC038WC3LGBsQsR71pzTRjVrAov28QV9epqYIXbp9czFhlzXaWWgBp5TkkGYrU
PyI2Lr96fXvfMzxbzf5tbFu0kTas1tuAFmvEeQfMNTH2vCgssnq3ZTrTz4Mg5LkS7ijGWGjlWBYk
tb86CtgSugv+nlglCEpcSFAuI75hHWx2HaIuo1ZJ+seq6ParxTfKvLZEuXkUPcxTgqPFLYed3lmS
TI0GATNgdL4TKkB6eUiLcFBbLN9Q46qBbRZiesnd94joSepuTRW2jxBkzQk5KyRE+Z6nzw/0aCX5
k7GdBWw6+0GGUqaTiwVsI7aT2NkQJBJ/2b7vxCg7JrDyhXjZQ7zI+secp797XOt5EmpmOHkE2Dkt
iLkY0chcmbMV/hwYBJnbWKolKY1/rzHT0yB5yPy+BTKWi2DS0QSs9J+1xn1XcxVtb6E7LcupqyhG
/y9Zs56mKizuPzkpCHQcrBqYe5X0y1RWzGuwyDX2q92sQrFRtK8j5fNSc3JJUC7Q/fovoDKd2b0n
DGbHKvsm27R/2Gc4SLc/9+vKDtLmuar67kjFWGLrlDBfahDIxuiauBusay7RrGQa1YwaAY2rwT4J
3LbWU3Imv9QHv3TF3PKieADx3ZKWBEXUDDP3Or7gIsJdibmKlTUauyWfdUG2vUg2/ePNgZDI1Rds
hwDHM4Qs7yJp7YGUreFvllEkmqC1QQcq0yX25/Hns2HIW7hTAC2uIT7nj36fBoZu5iLi9WGQXuhO
khrDzhhMn7jYA8glbX6J/FU+rj6w90uQVO1iiQr93hEq3kZC2QqWvSTgU+pg3gj1ENywI0MsPTa9
6cRpMaK5ewXSP0pgAq2wNkh856zosVFRPa7A2ozVPUwn4qO5kbKs7k7yZzEfZKHtIZfMDzqt/G6J
IQr3krqy6PoXcerl8y/P+8cjAqmQFljIbTJku12uRVbORVMsXOwdxJYMNQWgEn7o8nBaS3f9+kby
nAlOLd6Mv4hX6S2d0SSbiqb8E5iCdXo/V1yaq2UFwftTZi4Z9ga0A9tTyPriDJTtnIIaLsJWSuQO
2lcHUGCwE1SyDbWETx0PVLsUoFeDdXZShetc5BOwynjqd5OJsEWz+/SMpBs/nV6DNWMsx+QXOqRK
eirbvIANz4UIoa9i6vn0lx1B2QMudJzTAXvBrneM94MerdDkUlDzzfJUlGFdg3Ljo/QgsApixG3v
TNJwsHj46vhz9NJSiPXEAR/WRraXX4Pi1jpq6ZsdoeVI8osMysc2JFFsUhGXMmHOwfVpPyFt3yVH
qMqL1ugUZDPYoDCPWNvy0WeFTSulKwsyFShYu7baQ6fGf6ICXzGlwllqpZ85doNGGtaxbjr7giyt
8jL0302NCrMqTMuwSh3nvUDxJnCo74Nxnm+XpO+l+ZOHQpYhCz3oPWAatMqCVpVRhXIMVaZxoXMU
ZLOaDyafRqdCoRcZ063vXFuUbEyYopM9eZAU5aHLe9iwgYxXQmK3wQtsoG7eBJwpTpO1bkftngD+
o4/3CQnZk7loCb/euvk+OPhN/GeN7j15JZC0EgOxWsctfFD2JfckXKuzcuTx2w32uq8uZPHYGaMp
VTigtQjhmLEzOwxpAGSbmn6ZTLWeCHLEmFzlNECkGA9dstwE3VylPnXDr87PlAvjNkNN03kcenuw
irpcU5H382nViFe7wHMorzDGSLD2IdkDfXXwBv/qjIHHVnbiOqhFONcCYaPNahZXO7cxW32/YELI
o1vQKtzlS4z3HEfZlml2B2q2qaASHraphvilUIiGiv66iAyHaYROOBE28ZAEtwwZAI29o620j5H3
vSNi67aLIZSUxbvr9F4BkDEBx21IcWNeMrofFnc4cXusgT6gHj5g9+e3r5OdCM0eKFF4Bnfkf4V8
tx4p/lXCImtVM9iyK/U7QCdyZiJYwNehEVOylOp2p3cRH38vOQX+Zpa5tPsodMLHoXU+aIZoSWnw
uV1T1MWYdIaXduk2DXkPnUM/ckKII4Lq25PJuxs6xFNnl1mSosHxC9Q2blIFfjhJnJqbIkDeKJbt
MqTf4HrSDIOoJUuUEW8GjagvpXwCK0GMfVGaHJTSc/CbTXMD1N46Qgq47XTP3q0AXxfDmOgtgeqW
lhzb8S/OldqKMGtaOwggSq2bjZjAphPIv64mcqIQ/7ugWnubVOWPjd1IWUkmWcrzkmBfDWUfs77m
uMv9V7H5fXISwgT+aZJnT0kg9WvVrTPQsQ/mlWRnyma8D+9yiEsjytbfD2sMN/6yn1mR+XmNxtAK
htuMlt9rOIAg0yuMRMuVvvr3+EcYoEyyOPZnUGxT1++YPndglWLLpu0WOIOBCKjemtCsVwNKaoaw
Ey3V3FT8uPgusaZ2T/INOs6Xp+4lQUa4pJ3KoYGfzqftbLq0aBqonT/WRaxqx9IubtlhDwe4mncW
Q6h/IMmdyscaXBXJOuWeNziDjzd9lekt+gMH5tjIHWxVuVgm+tK/ZnC3OjiscjG8FRxxHIaoNvXF
R38U13EHg8+U+xpPNsJ0tbScvfvGmi+7jTkgej5c/JmoUAopyFg8FFD//WBfmKRdC/e/LwNVq8kL
rWwg7FIrGwo2ACHIyoQ88EC9/t4OZ03/ByVAcgfEXKjlUpOHGB8eEViteauPlrzPDIfXUzIRjhx8
CUgIlktHzQYZfv76YdftZwLf0ElIMAhGBMJRQwQhP7UTSm+WPi3vt7ld+JVpvb6vJ5QgLVOcqjjH
XXx+7Fz53gp3afx3H7h0UuDG7U/WwcRrYxWuBchcHNNyn4De935GgY5QhCqeCtloZ4KhJdklVJn1
m2+7Q79K+fhTFq42CCydFMc5Wdrk6p8x2wH0elQkCrgNhKADZHGV1HreI/7ognc+gWIqucMagCYI
QLlvcR822YiWW3rPF98vj5rVrZjmRR3qSjzNotlL9ktsEAcynL2fIjsN+gCOJ1tKXdpoCjO22uVm
SzG2mHtEZOVhrO1tHd+somSQi3RedAuO2H/oUSvSIAhNKlxbpsucOmr4dJd4Z72tFUfUvrOGTeAl
I0duCVr9KMs055OW3yPxd5cWv4TzJ9itahQp5Ztf7ggnHUo0x0n4QzYPQn0+RvqjJeRIOWXIpE1m
UInyzj3CE3WUWOPtJkExSD/j14yMaHbauVVpXtVbqWCYZ1dYTpRCztQGe+4FkqYqaa6fJkHZYS2n
LQDu0Z079JQXNT+rHofWsr7ym9x1+brNK/uIOp0F68sijeG9pYC1UStn1uPt0aAujfXt+ydL7uZI
lfxjOwSREd4+MWhh3zdkr4Rd3fJOYEmFsrsm9cZU1KJsio+69FXF7WkyOZlcd/l/ijS3OpGxpD4/
FV77fKLOC7ij+zF2PojG7tl5NWV5UKnGltkUhO6iFRLcs0BYD9Wn9v6GOkC25Tk7P2gHfBhEMdfr
EYmgrs1spMvLg12o4fuGt8l9dW/hfem/2apicQ2djyn4mmWdQ6smjsJ70icacGjcw2YlrdIMzrd9
YDwsGPz6nFy8Tniy4nzL8sR9yO/p9ubrRE5sL3smxHADZtsH8zmNuwxo35+0pjZsir/k9iBKrBEQ
Vkni8P4SgDiK3zitEmP9SD7w0ZUyyf/48l5ygPXdzc0CduTINXL6RV/XZf7sM3oFA1oKIEjrv7aa
eR7TEkLymZD4b0b7IVVxQEUCTDO6SPFBjK0zMutFUfP1H+Y6r/n7nb2Q7WD5iSsWd39gtGND271k
rbCsMmVqX6eGGHxZW99YVRcl41khZvpowy6P4KR7PIyn7ki/7ua1zxRH+LJer0K2BBxjTNFje6ke
anUO3kyV8GN9UEjVfkfszYXzCb9TE2j3n8iJFV8eLTFNczgAjroPSKC20jE/nuq3kzNSE1OWrtpE
8FZoPWtR+0V4yBtn6ZOZ5nEovwzFEZ9RFW1/AOJsu6aij/P9X1Hly5uUt7oUVq9Shgo0KfRXqwAk
VZ4zXSKv8bjqU40cQGCqP7Y2LvuJpIQju/CcZRCku4gt7UemStuM25PeSMhL+NNQl9/LOCtRgZwN
b69hQs++3cpQiTS42SLT9air1cbkwFVX4MiAJJhN3HpMJFkwQcPJAjVbmkRL2ZGDzfnLrufqv+Kg
G3jssVL2g6UDPxawL6sS+SpT44wEbOMxCi5/7Q9Er8FM8Ipu131PA/6L9U8yCazEgxEQnBMPXERH
K42GDEAlUBKANutQwVkBS0XBoqpBl+PYtuJgb52tYZGx3SvlM4USL9Yb6LQ2d98Wmx1pyVyvEfKA
D94Ob6G5fvXdb228r5/4yJqQtZCtPqM+pvIuaO+9FN0lfAkJAQpl4rLrjpQEF6GuujaZb/TOiIaF
2yZM0NWLC2yODJf1pUSuv9sSgBFRPsx7YUt4MYKhJcNLBkTj+YtB2W6OEr4ar/cAJElUO9fQyHBl
zFWcyFRr75zdbvZHvEkglo5AeWisSh/3gUcvXErpt/U4hXCPGDT4MlHXqjHoJmyOlWNmPN/4p7WY
gV7RFw+FirZhnG1Rudonu22mPjeTh4drZOCaHKD1EKSQURCJFBmAAbJo+4C4vmXhYP8KIGHH2bx4
MjOXla7BcRRWDZodi7Fg6wX4oo1waPL7fE6hzLhXzpM33tOg6vCZa0n8psvd4+5EXUdP940YkOK7
jjS7JXuOQnOEhpk0cTvJz9ApeJcGMEVi2VZu1v+BMV1y/qRwl61GecRD4qahJNiowY3nfC9RasF1
neRhU+9ZSBmFWu47M0N7AqJM/gJSA/0TMaxhISIVdkwlAfkEhRqDsGOX3+Y6U4W8rZsDbCjBA+42
MstyjkMLVR/LMaX/RlyDpgEwn4qblhSP4VH3GW7kgZomr4+YQgTiFxs9QwiKPY292QJADk51Sdoc
N+l9YgQ+cAE7A2nKozwNy2Z7rmxF23yyuynLBgDe3qcjRzp9A5XALc4w1pGITg17rRSf8fBWnIAb
oyqbebSCCZO7sIe84eQ2/q6r0UR24hIssJGmNyiC1NqRgvZUEtXvo3YsA3OrHce9jr68KRzdAQ3I
/1BZsTgfWz87xcJ+L1vlOmLCGcMYgekbkZRBxm6ngYsEZL1N9XNSefwn/PWcaXqedHaAXM31hn6l
XP3AVActLPbiGOmwetai4CHESNPfXiIuSRTgLyl+36ZqL+eMTNt4DurysJ0RiNRfJHGSiS770MNU
GjkoaoMdzf/AmppUgDKZvcecPuQZ5VTQ7qHJNkC/8eO64OCYdosK+U4kxLtrjAFIDEj6/FViebnI
cmMFrC7TLYRnwAnvlZxzZskUCl/ZD+uTZuTJWgsShGd7dnhR0C5jv800FDMFPSOKraVbhM2Ymar5
PdFUeKCSOOOhz5/M+m1XW7FxH0TQCfAbtqnPMdsdwxKO61sPx5U5dTuWrAy0e8rKGO82ES1Tq7sf
YMonh15WnKXL3QSiZ40EOh706jZSIdDzsOKIzaFziSBLDMKPtQsFWs5hgBxeo6Dmv9seZ29rcW/V
EJMq6Ve+tN3XR8cjHiGN3X/rpooTQE8t6VYPysW+BV5Ew9HGetFJDcuJgSwzOj4IHItFG9jnXG/y
ZZwJSAt448TsWXH3lIGaTkr2joiMXFapdo1FpFgLSeCFz/MEGLSbhiN9ZDPGaF+Z2oNYoWppdifP
oLlFgH5x1b/Ya7edz0ZaXK7IaBnc2pDyP+OxGTcE7NyjilQxSqd+7iT5SPiqD42x+wJIYOtnECNY
zqBHylv+VzsawVMG3mnyvhERyaaSFRWcWPxvdNjfvznaHElSOomQdynpONW2ZBVfVc7tPH2CKqXv
cBTGNbfGgDa273mCDKb3vbMaRXGROEtcl/9P7aboNz1riFtKq8pV3yrgKdSuf8+Sb165G8GVJEGZ
98gzT6pmxQHvGRCGqOal6pVBF7wwfWz+czoZ5OAfiS02Om65iG0IEmicQZVtw5JdiCLueXPspNZu
MDvBbVrjJ7kKHusMcx10Notno4CSA2uXuX/0rZbAkCKgodPrecLUyAPrRn15cgf6cgV7qPX4FBTL
qZSbRYR2r3DpYkT4b2stAKhsiDrlKiAkwC2x8IUoaUtdH+rlIVLROcj0vBFQ2dH6sjMnMIMTF3mw
4HMo0yQtYjzdIVY38+jgCyj6BObOxZyvTU2B4yALnbCZlPFjpmsoGB2okXrI/gggxX6tZXJa7Ulw
K1NnG/4JO7lA6h73qsVKswieBA5huXJtGoP3N90XZPfuYwc0pXb1nCQV4AnU1NY69ugKz5cCy1a/
186D8RedEVwG2jwBzr7OXS+MwYBhZe/oMMOPCvrDF2x9HDALOCA4mPpjuKuvEYF+cSiUUJVtv4WB
IJWGPgwK72vbt87zt1Iv+lU9C1btQX5q9XlfFMz7A3sbkInG1pcNw8qd4EAIsAftsb05iizMZKSo
eXV+rXTgGF+bzurlcJysCII8s7sseHNyyqhfMpMufTwvcwmwKvZ1CETS4flhTeeTs/ATxpjWu9qq
Q6Brfl684i7INwxQ+qczFrj/PWND+ZD3xwNuBwWVlGrttLK+f7aytZddietqvFXchz2fIDDKJwax
G5jzlvwQyL+rjQFMkUuf/ZA+fZIgl3vOBJivmpVgBPMgVWblk9PpzfHexN4CVftwsMrXn16a20SO
y767xqCmrl78ag22sDwA0C7QHDY1bOJZ5rKMCBH1pIiZ765ioRHeyQnVYWDDtNOQnYUF4J00XsFo
CU8zs4p/B5Q2d6EjI9nPfpwpv+nTKpfmHHNdsN50iWSpAYkhW6K3dhUoCSsWjYXolLtsA4Vn5U/j
I0AgBIM+RGYjbzt3jxQHayhARdFuOoU2DgBckrvtCYZ0gYzoVrSo1rvSrZUbMBA8eHQK9pr5xmd+
Z0xpEfGLYRu3ocCZZY6dYfo+vCwRW0a/UqT4LQSzY48YijchAT3Yw7iAy0TSpnCotmqt49HoGwPr
9owSOX+431C0Ip31S/QAjNpqR9dajtWIE7GLFAYeTZZBVoG+rcDUGo/IVdK7E/dYHf/Wzj1jjEX8
skrIQWkeoWrMj15u6+GcPNEsyT184q9pu5ssfleU8CPvmb+MvEMtb73/6BTQ4Zz1I2kW/T/AozVi
Y+PhUrlsBrmFDmP3+2RBcOak9ZH69W6SWv47gsJXel4HqtuRrgfDdTuEqIKkNYWTIRDSGqmdXwKB
OkbKvIROchvXeftat/qp09gHo0MSuYowkMFlB3+FpW63uBwIDHc60kbUE1B3CUDUYgjK+mdApDNz
2oRZuyCI3hU/NG3v6TpbM/bqhsCoJwcej5Hgd4ZRGa2KivkdfODqQccwc7dehZplwdFCThjCjwg4
aj5gpfNlRqBrMWMSXA0zLmRRFMK/6cc7LnWK78aTYup1vDGb5S3kwibSvgNK+U16AUTtiPXT4uSM
LRBeAb7w1cf18hknmdPpMkiz0JTRBjlG6ICsBrpbfIBcgfSZP7QFfCXuUVIxV12iXoBIS7TqH0Vr
wpHLOPR657jJkSm0HL3F2NWohRlSDkRoh/De4oSuvH9rcYqx1vvou3Y+kCw23BAD7H3jzwxrN0JQ
E0HC3GndmdXTJrfKKhn46madI46pQC82ZTO5LC7nlKuLJmWYFxHkBzbfDg6Ve9m+sUBAzIo7fmXv
hEWrAtSYf539A4ERBgz0s/QXvPLhkIKG/w+k91iJ2+7Cj7XNXHUu1gR31NxIJqkVwPUZCL9C58cV
7rfaJf9w7bSdWbRJ8vHGKmzD4w75JGaP1nryMpVhUp/O9L6Rp3nbGT8aAcdwfs34CVwSTcYlMaYk
vsw0gDO5j6fbc6F1Lm26ZjTyyBK0yifHeTEstJSywKSBf36CRONpFQn5zbGjfk8HCGjFhPE6K/54
NPckg7MmFC9Wz6XvSAMat9+3AsW8w0YYwWONXpjm9GsMHNNXFI0KtqjkOayc8ZzIn+m+hUK5RLYK
PSVEYMF5AehMUUtmBuMrlYmuqXINse3wAcdRpj24sJPrFwFMkq9XXrAijrhia2NTIqArRqPnUrNk
hlpn8bYFYrJOA97yGPQGabrN593yG95GVAlO1vW5bmcxepxw7sQBqaA8VmipZKaBGn8c0P6VRSXW
5VNvrmBsnSeHNoAUxV6iPXZOy+5vtwfkVaDyDGU84Db1BiypmQH2673lHZYmR2ZfHsLbCNeGnoV2
LwMaSu4lYuMQl7OSJaFgvOTC8bJPRnaBSvMQanPI4o7LGM8pPOAeUBdiMMj1J50i0pEsfhLkG7FP
vBC+E3mf79Ec6pel6zdT2HB6QF6hRVaTZRdr0Xdz1K0C99c0LhJZjFKh7hZYmD/YyrYOiApLB65o
eHjoBIy0WKfNHx9go/0IwZbFne4D5P03aSqo5pi0pOOeAuIog51qb2tKLSd4aNhg5iX5Z1VrSuDm
M1CD28EOdTEa5AUVmM9mJL+br8XpTWCQ4WYxle5qSpiQqQ65qwY1hjLhWlgKsmjLVBCJ6w6Z7dju
kWzZHjS/klf/1ZfCLUsWZsV8DTnHA53SwIO7KAKxtS85srkfjphyku9NuxkbxcOXdcwAd6rOnFEb
7JxhWRuly/EWz4vU2TTFfQubVHfQilgK//5gDcFMk0ODrp2Ipd6+vzHQClMjaWX7hbTZtNrryPKe
V2CuoFgVGkBerNZAMIqTxJChTPoetrxD/H0NPWEGBUeSP5SVmzrMW6nJazOr3SCFW+5PxNoITpW6
D4hvR3pMDYbeT27TtxxQ689yWj4OMEr7mm2rVUzHZmuTL9BvXS/yGH5nZJuwEOnL82UTP4q/kE18
f0zeUR94V6HiXPXaaJb+p4RHnxkHdgkpIozaIhM6DzobaOkAsuiHeX6+OFqCZmRLJTznj0OKCWn1
HASdQJLnzzhdZp4aHvfSpj0j5vCJA0Z0TWm8YptGwSHCwtjknf/t/3JAgEAfJ+ktSCik+KOQsv10
QgqKTJrvLpeVofEDrjmKtMoEgiYxHwIcBQBZqhwOvG0eG9xmyn8x1hcJsjsMYAnhSMctdsSIRRpZ
/irwKkc9waBcYhs0JuEE2SWbZpGj9/KxM8vEw/WdMRM1P1XVF+gE9LDUnb/xyQoVBvEUjFgE7Vja
gbTLIAN2Ohtso0YOV1yk43g2gEq8fmXr1uVSGqVCQD0jNBNo0smgw8hGMQfNqAQ6AgDOUkXLmRhc
OdVvvGBenyqTn6VQ/8bXzYKX949z2ixKU0qWUklrvvpfpipPARWmTCYkShkhfMnHronu6uyMFmik
b2O+Etskc/ZYDI0e0DskNY/qvK1HcKdzI3rzbzw5pCLAIZYsAjqth4jPb/giSg1dSvCRsJiJfUx3
p1qDaDZ4k1lD8O+8dqon445TYX6rt4sBrjFp8X3PxYsCnBCSHgrahBSMbkw6IZF0udmytFfjjM8i
NjHQtLZnQ3g5M2BNNCrOwszsl+0SFunuCE1NNNpeUKpGpXUp/cqFqNE+yz/f5LslEzf2Qpw9wqL+
/3dS2VV2vV4aaBaZFYw4qpGaXxS5ORGixXQVtjHGBUOoMBxsiKmN+reBAa6kXr64Do0scFYStLh1
LTqF7UjzGP7W8Fq9te7/BEHrX7M8zfJiYgL7TmwvKxv0IfZccBI60p2+xF55GnYej2DAAQ0s8Wjb
jqqSS6TpBPAHN+BMOqsCFCeJvOS7lQDHqO2zaX+ZtQ6/wu+cMsctk4bIJ6F4ak3V9DqLkqeiuC78
rfg+7DEEP/w2J+jWuniEj/Mt4vKcK/9+6jIJ/Xyc2lIZKLe7YdTUoY2LKuCX71FtdNLFMhFkub6U
QSW+A/80jKvSnIr4xmXWkYdDaug90p8SRMI0/WQsYyQsaZaShMQiG28wL2kQfiiUKep8qzlnNfm7
+lFcwcKod6sGnreCog8Z0AWdf+Z21RyewyJVfkIgt5+UmlQO3IugTSpA++PFO+U007LMCALR3qjT
TewkZoSGdB61gSOpM9Ou4AFd+M+fsNBqOndTv8i0bUmUB66C6qW48+BW76+iDKLJuCOUiRX+mLRv
NT0s6zFUgRdL3AtYAsuEpKGz7vowsrrVQFfic/DyzxvwvLLtxfyQ7/XUxbotw7JdWvl3Uf4VhEU7
hw2mVwH5zGVqfXTZj3heX4whbWW66OY3hDkV23ZHzqSm117gZoD97DAdV2qVYMee0yVTIbQWINxQ
LYr5hFJGh1ClUj12VfRfeEchghARzO+P4/v9Jy6ILSWVv2YcaqimR2uC4c6v+jPmE5aAR9bbZe5x
Owg8bkqV9+LPCJ5xONyOjQQ36f/VY+9U/y7xnsiXGcDNtnjMY+1AZ0gpVh7YCjRWJi10wQNScuuq
UuCZcGKbrwNkGT8qWghZRKfFiBqnQCQGbB0eAnHxR0brufImJXNAIE7mZv6fHfEXtNYspVPH4KYd
2etA9d44Oh7BJTbycZb85B0TPzdxLE7YmW/AB7UEfZIQOXW9Rj5n5Nj5vz1tksX3Q6dG0sDmT57s
nKoWklDtiNBaCGeTGpzodL6JS5lLi7QtP7RDnVeymFhYRKCzs3/zNoULmi2MHki4bl2RdUGw0fxN
BIXNwRbxWbydwpC17Euz2qgh2Sfg75NkWt6jtoALITxZ5cieH2ESoVeI2bb0BtQVlD41Cer6ByoH
I+jjkC7NEVr2Y/oPbApj7JjEoehqeLiy1DhX9nWfyqDjRcUlpDxGpe/xSlJ9reZiAw1AyrCAhIFx
NRMeW7EeDUASx5qvhDQwjdHFRzpVbVt+CWXJy54YScw0hcgyeUnvjVAVFbK//aDv+DBbHtOIu37u
zoEPwJ1A9/L2whNso/8kXevVd/PvHiZ4xg+el3tDlEmJ9POqCn5Ak93YIIuflwySrdZlq/pdGRnd
+UvQzXjJxoVmwqggQ1vhAEsBSlGM5RSNCgeNtz9kTVQOZzQIR3cWpODUy8NN+DDsO7TfdDSOO+RR
cTBD4OhLhlepyP85aoMX8g7hH19N/Esskivth3tk0T3wYtCv/5D4NKL7LGjeHZOk57rRz+Yp+bg3
heynCxxQWzKw+YYCVSs3Jtiu7KFpitC+JYgfQVScGA35s3FTQTo/IlPI4+wDKZqoxGOGw8AxL97K
u/B0Gct/oa4JqAxKdpDykG6/6YctI4i2xLcY7K+rrYfdJ7I0yIOkkQPm9I/7/61OSk9A5FzoTjYv
gPCCClTqY/VW1ByWi7nrnNZ/JdRBq/Pyt0DVLjeYWhy3aFNlarIz5oSDJIKNJPQVjSh+IpRzgfO5
PFm11PU5qeTXJlefsgGV2ikYbGhY927fnnUNPwjiGJOmne6fd+jiN+cS/1RYSdhQ3sereiC/rmiR
nHT0Tg0VrxCLTYJjJdYW6+W6kO2+oZsfKRSwUmyYvQmB6TsHB9FKaJfrue3I5m9Q3cmGOYi8gAAL
rvXu4p2doS2Npqzz+BNt8zLWYy2MAkqvN7qxz6hUtm1hHkSuRgdaLZX49BKYjHs9jaoGsd6B8oXi
9MEHgSciF6FbW7AEAIhokrXUMUzc6WQjE/0JwIZ11zH9YPe4X0GmCHG2PIY094Jv3dpvfprfHK7L
pNY1mZ1VV11yhHCI5wCvpkGMHkwTd8BpEcPJPUpknCa5acrMLoQTmUkXXp2gAI/Kjo4BZ3vRozMN
h73JbSej2E0rsVWZ8ExZo9aXJtAR3atj3C2CuB/6pPc2ah/S3sHwE2GGZ/iw1llIavrXBNO97uiy
V9c8KfIj/JohIUreIShy5voEF3wgrQnS523D6k79UsczvZi6nJ/EFK7buQMt7A4y3tGuF+6EdNFt
+a/WaEdY6PTSVoXbTeQd9Jt9loZH+Tnolag8IwehF1SCIJgL1Ugr+oBptAPDCWN06cbzlPXpk5XK
EHJV9hRjXK5pPxqpaM4rwBNIG6ObIyXSyt7oG9MbUtSEKDFVOaoNfYmZ+Qa7mnXEXtaI5ltrGRRi
L3qbKL8kQkhundjhGEBChwX+oNcYOKjbiWYngBkNsYFdZ/01yK218Mt6Hi0rlx9AjW3y7iP/yhvi
shxZICX+zqwXCs+3cAfiEgUX0GsGeWo/jsxwYfnFJVmmP5j8gY8iMswF0sgPjjkrgQlYgRhWqYSI
T3auQyF5MeWMH3uUXofV473b7dzAM95e2Z0+GIFcGB0k63AlXMv3HExa8tjJch7SerVw9SsX2AKA
VKIT3A+R/PpNIvnw9+i8OLlGAmTxE5AewMV699xAxxkv2SAAT4OLs3h9lAciIZDq2i7Tz8rJJMja
tCcxP3nbOX+bFUncHXMbuiZrwtJHPtZNU1zenfMwzgknrWlBHDBF67Mw05MvPdxlsyJIvhtlIpUl
fWu9g+cRo6Wi//CsPz6E2AF4nsq5f0QBy2yza4nnxjLEAUhhH+kRzEVAanHQvGxNoFeqh6/cc0m+
WmncI2OHhTOdoIV9bBuWURVC4oL2FQ46jCurkYsVYabp+avv+tFj60ZcgR4oLI0/okiIJBn0/7+B
2JGTtDbv/JGK6cMtxlg5I4iT/ES0S46ojwutly3D4oMqJXZN57TrLostn0bbzkPTwiJ3k9eXVibf
P2lS8caZE6Q8v67ISUISrwAu4ThsczvsXwPjU4uUIJQ2Xdg/dv0cOWqiLDgH0TF376SSlQ3lpxGA
PtZ6nlAXvDgGzpXjljdFt8LG6KCCzWZFDNhb5ohx9AZ6rZiOs6Mfmt9/ZTeZIHCyZziGMD1fHBKC
5/4nHdUDCiCJNdRMHEzcBhDh3tD1osm3/dDuEVNMONANIL2JOVJHquOnh9Q7sTE07+UlCiAyMyLE
SpYI7duYHAKOGgtfJI+GasaM6dcBSk3ECB9JeM4iLy7zXpW+ZX2bOg4fJSKMHRCz7X4Uc7xUdqAj
OsutcKpdFUbNeXwMVlAQVYykxzpgqWMlLW1+5f92nasKETtTqwTJOe9k8tMiBpPUe11Lx29XZ9bV
0GXzxRg9msuHv7jC4TF57pcs2JOJ5/EaTW0I6Yt28FcPGkhUgVJ80DgZX5FgrPQUPE/i5mmUB02P
TAw/DTpQL3VfjLUB0shI/wZBUzoEUkOB9CYHuiCZezxUcaAG9BhTTXzAcDudIydYM7HhkduKJp5a
ScQNIyZD5Jks4fbLGjX9srgoU3Ichipv7U2qOCC745GmFfztpQ/CQ1ZjSypucf/hE/5a0eqHeuJ5
HzxMMNAGTKNgAccc9YjwNbonzYpyVVgBFu2W81ppLHjBpGieKSUsfNAULBQJxyYx+/efBDaOoF0K
igns0UVvA8B1Td6yRgSMCqkp4G2H/GAAMziwC6wZisF+QiXiYTLWwRiWcq0G3MOiP9IgwylyKtvE
7ngyIxRDjalUU2csHkjBFywQ7ID6mRK1734USmJZZ8ySt6vC2H6aOU7A7oSUJlFxg2SmhvO4JNFm
DZnAgkuET8KLXASjEadomLjD4KfopWgodpaGJYwZ+JjEN1YHKpH6v3S1D0rFVRiMzCHh4Qb8wi3O
7wlSVldXoi5Khzz5lP5Lt82y/YBI+Qx+A+MsgXiVxY6JgahGUF2ZoaEv74Cqy8xQrfNJ2Id69QwH
vDmdXaM8p9tgFyu3iV450x7VSmMBYSPDxFN51cgH1LgkFD08Yk3N52/56TuPBGh2gFKN1zHDCcU/
7KzNw3H1QwYaLuDDF9D7BQuZzRsdjARulf1wF1gqBbTLm90XkTS2g60RISb5/Zz0eGeqBeRpaWzK
y8kK8cC4Rq+2zZAkkmFJ1OMOkAwsIC/+g8swxVZ46j4JF82LPY+CriEdF+L8VLC3JvjQkbAx4HQc
SaPOeznrIFJR5a+fuiVfSL0oZ8B/eFJAmOTWK4OOFEGTy/zKaYOUzg/19szATc3xRFYSf2kObNMh
VeT+9phXCadP7NwHLk1A5xmuIbpV+M0B9w+aT6DkGi7QNYRSAD5uoecBEuPjcAnzcEVlr7OIumPW
ZvzyOFg2dR10LWBPHeaQAgWxtIwFL0AM7dsHhayURVel/Zg8NJ5XWiidrUJC75W4UsKi6S0A4nmy
JCGtryEmg3rAqx8Y9oKZpT8g2TGkmvGvndTBnOLgXmkR/VraajRfcSivk2CpS7FVTzthBx97vSa+
5wgb5htGbu3CarHRIGZHUCcnoer0d8+OOSa6ofIX/ReyXzfKY0HKp6dKjg7OjGyWZNeiPNUu52t2
ZPJiFy6AT+QCV39gOxlMcMbWx2o+dJoTJLyobaFVknuGwlTYq/hIZZp9k02SwktyViVA9kGHcjzT
Lj582uN5s+LjWeEJkCBNEF88rBjFQUHulrh/vcLPiTVHge/CuxOQm7Vl5lGMnDA+fk9xzjSvujJL
uWph9Mq4ej50QQwB0gIr6MQvR3CoS7Kuf+gZjFRNcP4ONDHHsrcovID4yrckILsY5WCkpEkxuUDA
Kvb4CifSWcYn6Wi3gMdIXbwZdnHKvPVm9voefF6zN6/E8rmTkX+45HcFZb8t5MUnOfMGhnLAAG3l
q62wN57/0+cbuSVtKdV+U5w639oHrddK2Cdq+FtkLtxYntXaOVHGDsrGmkNsHC2NF13U94Kwtpcn
zU9RS78tK5tsGUTYzt2vhyg9dnt46Q0WO7VLN4UAkLTM4guKF9dSmH8vsltHyha8nb8nckUubNXG
3d5v1hImhkGXKHDLKcro/xEj6/Qw6Dcfq0Vn5X+f5lmquX80s5HmQte9cm1vRPzFGeSy3SqOjXgX
CbmFZF/78cBMm9GZpHwHMcy2pq4L4qB9ZZcllulc83xUsdvmUrYdm+ADevsBmB3iLFDdWAH9e21w
X20kxTuP4jnonrc8aGCJS6Q6NjjRhNYBya0IzdhTv5aZvdEpWFHoLeKisZpFVYukk5BLW+/D8q1q
Zwuees/BgF4I3mGnqVz9q4IsGywTod21KB3GP8rtSJp7sK/YctkmKEdUFIcP10j7YN+raK5JWAj+
6HgaAOlZjEoyJHk5LJZWtW5cQD8oF2CcRH6iYhWtmaijbW++LxyBxESQZSHCDwyvt0EWZk75szEF
r/VcAR28myZZ2AYniNXMxfQt/rm8hf5DQNypR3K7Vug6UD41CexqplEUaNz4MdRI4aRXgoa3mGQN
9MCCanbKZqG6hLX7Raze3v18dWlQU8o5IbfreryyNKDmGaH8bfu1MunijDt2U+WcHLh5DZdPJFgZ
Iu08/92YyNoqYCVMRoBJZzLb0Fq/f2IokAio+ZX50xY5mhauhAn81vRYzsSmY7NG98B099yYIlHG
uO8yLPOgdIMvyU4WZxsJccswYVZUU4Apr2pK8yAIki+rXGPYXwSQI/2OO0o2Bs3djDPoFFu9ET4T
hIRkpKr9gAitBOFR/n1zMZnTN7+0jj4cEf5wXit2W8ojtVo94hjgg2UJJLzlXhwkiVJplVvwCaZ7
dz9744TeIIxk75dA7PqJEU4lqKadU2kmmds7GCuu01BBMqwhr+namtShm3/yEXs8UvnFLbJBFATq
qXVXm94seYlrMA8Zt8RRrOwcxx9m27OQjetqr74yODuS9ERsAWJqd+ADs65XUSoA2pi2/jpPEUDz
MG+RIN3/hPw4Sx/QoNGVo/iE0R3kxLnUMWSQtVj1+F1xM5bvAA7w1NWcfbQ73cl1zXKSmGhV77f8
2bNpdQ6m2UUeSX/MiCGL3J01SaDS2IJr/rGz4/U2mpE2CO7Lans0fzQMDUFoqUsxf6zUlCQ+dtmL
FepYYwdUl3ctsBPWsVyM5747U1v4lXA99XpRBdcSYDOcchxlXu8fDC2VN8rjxW8hcIilXxB3o2bm
IWm7dkYE8oz0xxX3tinf3to1tMpjc4mUDWI6jkHrxiUeiXJr+mA+21ZGcXYwzICp4ZMOSPVG0oZe
f0QkJRVXPi+d31Gt7X4Sa83efws7yZNnEm10GzRmOC6w5Z9xeJq6rl+nfnruFy/lE0x11MYMqhED
wbgUkIzOH+meyO42Gy+z/Ktm6NA8PdZt4eO6cWSyEvh5Gwgnddl4CkJSWQJuaPHbaclyiWe6IyAQ
QbXUWve7tcudrNdH3s8qi89t7Kky0fZ/bwBIln+TDtC8SrBjYylhHqkeVDOjyhbQQjmJvcykkdaI
Gz9DQ+NjUq4iSIFOELfsnzusEbGaQgZuEW19wBR0gsAQyvG3ClB0ulI/wku4ETrA1HcCxp3YDbk4
T/5BUBwvq9RvxYEgrFtdb5/246T7gPRBx6N9ijt8MmRjP6fAa34mQ5v2eOQtPrWQaDnCEWJTzhcK
yScD2J68VVLTl+kMVb4xaDbCZ2MzGhN/QcyoQyuoYtsQH8dNMEzqi/Iyy4mn9eoX9DmDgKvDAM/S
qwxcwjjxWV0+Phqb7Pn18Nmoi8aqfTAHYNcuCZGjGtW/zEKjaCT0S+Gpjnl65hjG0kWVL1GUy+PL
x2WKaOJLI1LiFVxDcTeaYwZTRVBUBSYhNGlG4+sHCqCU3JKiLzyfYMzg0KH/dSyuQnzwE841FuS9
OwjUqTR2DmAC5wo0G9cb1nF75LkpJT2Hy44bKmUbYjBwlwnUomHj7btyrLdl+UfqUuvvEVo7aIvt
AjY6iSFc5xqV9Z3qO39/CiKtiBXzlMWikVMwHb0+9i2SLjwkf/X323oS/2cyNPiqnj7JQGQO+LXg
8+Fl8j11SmdTl2os8czJXBsk37Ug7xW34pge1cpexmL1cuyEc1HJSHRqqtcLPOp5ghhbdZmFL1Xh
n3WIN+1YCag5gyFdJX+CGx+wr7kmoqiH+0lCkC3j8yyyCgiLLTceTsbNJ2r+DEuaaJQutnb/kCdk
forCllm1f1z4saToBddhybBisquhVXzLGdFRfcmXSYqqXwjlX7ibIjubYZ1cm2ku6bh9BpzPEdYW
GPH9/TZH8z7idOArcVbmYly52CUwA3Fj7A+Lj4rcJedtU7UIdC9TnqQ7Iw4uVH2siAy674a2FkW5
y9/g2+/ZWQhVtIr+go9ubDUvqawwOlcJGoINMGhJcQ4XEwcolCHg3DmtjPsT8Uq1sy8P1gh2sTRj
uCt10Tr4F/N9eziR2zKlDy2WtSxcVAFni/XOTVMlXix9C5GwDWWQhAqisd0zY43ri5jBN7wp2i2b
cpUY9GKJZMpdepYQzdSOCfztbImPd8ZCAdT52xu0FFGNo51UUQIVQpUGKFAlk7dlSrBKEmk/kJMC
iRcrwiLZoWQqDWHg0IA3Ptm/gBK98y16wejbCRYWXR8jVrP2e6NfE0+9SWKja/uYi7Fsr5OJeNCg
5H7BRf04FL5qoYysv776VxiUqCE3xMWKi94oE7RFqsTPb5JE0aYclDxIuuIWM2NmRzavYxQxU5HN
1jZLqrAg6opcosG4AVJYQlqkM7TvLrLgqmIda3ReDvR+Rka/D8U3u96qo+pFf+LIGdeos4QHGiNa
nbKWCt++5kj9WgBilMxt9hmi0yrzAz+oGdtaG3iJ0bb3Ad05h8qRN5Y8JKF/swqESyB6TPp+jBoM
a2NsQzKbfr8Nsjxk68udWwUznqoa59F9Bw15VbUK0KFoaqSxJ+G33vUvUHJyL39TYoetAL7PPDj5
oTnDug1ueTxYQ7IFCXLdqjkx42TO0jQn0+o2G82rS0ssE/mpZR3VEPBxrwph+zJJO0Oq6cG0fzVU
7mC/5AoclUGJVuUA5+x+l2QsrmQGBEGhXhjjyIfLRDM8vRFrCgjcNAMUl2P362L48fGoZBJI6cU/
fvniTtG3lglE5smv7G1YZ8ZTE44C4fZoVhrsz3Vv5nFR9qKTyENBBJg0zyun84RT7hvPHIQK2HJ0
5iB+kTF3cdJ0NOPiB9tbhMmrR4yWlaWRB4alFVax7RpblJhbW3BBkyKFrbvy3aHVMO/LJLUZPR1L
RdQWLLZZOsWK0MjmGfNo6wl1kTeC12AsMMs3bcYkHeBqHYmXErv9Q/uwaWRDKv9oazvOd0/qR4ve
IFaiaag3dX4OBB4EoFraPOjRV/38qE1U++iqnJTgp70qEazklIuz6PVG0gF3JPeh9kn2nNx77/FE
br1yxhz1KSrghYaWVUmoCEZD3ggdjolYevwGfgmD+roHP3K3EcnnrE4J7vOp95rCuY0U6O4XHB1U
jbqiNJ1VuvFVf/Te41job+jhlGxcAQ5RmTM9Plu/1UL8QIptotX8QoIAAuii7V8IfzfE7Kekukue
T5X8FguLJh6f+HsKPGZn2GjzVSzNUia8qbYi4aK5JT9+tHOl1J2noRLc8EJrNFxBO5XT6OAMQlyc
dcapxQI9w6UwcAQJnXRuk/e39ueMGU7IpJ3xxvYHe5ibuhUYwSkZ5uDoEHUJ7RGVflTjDz1+LsQ5
V5ujqDIUO5ZVCLpjRznqFo5v539q+9DtYX1kGAdg+Qb4SeCg3f9zvbT2Y13eLYB4XDW7K/TRj5sY
innY9Dy6YztnWC5zOqKxJW2cZxpoMmUsuRIayi4gPExMrEjeyUyx1tejUCEX1TZn1ibyGZ6HBGzf
JfDNuKVRMV0dbk9Ji4EeXCRJr77XSLfkIy36Rns/3UDFiY/L7C9zkEpjwrRVLsTEqKdsQXqCeFnP
/7Aj3gF2fn3ohXgftieHS8a/l1W0rs4yTm8IRD3tg5XALYLpTaNyRB1fc2adABjrL5whIBwTPkYs
iCpLBxL7dVmyKC+Q4tRfej1Xh594G006c6edYN4ugkfsvSw7eAzvapTTbB+e4hXwQvyFoZbrcR5x
L8ybvoXghKhJh7j1ZnKzPx9E+MiD6EnGKmLzF5ZKr0kQiYhpQezQVbUwKz4xnRLdHy+LINtBsiZe
103MOsDlXlbpxYEzLmrWzH17LdhDhYLJYHK6kuKvF+DFGAmylEIcyU9hoaNtbH/3Hk+gA/sC9rMp
W/+SaukpQL/yEeWcRi615lJT038Aqi5IEtpQxoMAK44vU2IhrCUKjdhoc6/XQJKoeoeXM1SFgSfh
FTY0SmhAFv66U4+P9qFSdYJG3ttT9tglqd4Q2l20f0L2LjDOd10OUNUVU39T9ePv7xJ9FaD5LICL
FtpqPOHY2fhP3+GZPAYldcLXHItj+QFCcShtOthh//q4CqFhwgGaw60zoA7zutxym3USETbW9gxo
ssVLWqJylmRZru5h/h23I8FmrhjzzR9LMt5ccTD+bMuXJrH90bC2SJj8jdQWyNyIb1Nfb2mkx1KO
VUv7TOdStgAw1t7nyLAe/S5uhoUbsQCJGTaBndIViDXcYOWkK9viJt2x+jgrtqXqUtvrSuXHCjre
Ge7Q2UESLuEGh1Hm2jfMd28bV8q/55fk9X2ki2ru+igeOWuDSNi9/PvwR0sfyUXwd8NI9RuiLjHa
+FbGwzvk/ogkyECSm0z+l0A5r7eI7lnqq835WsiNhLKYd3dqLiFz3IwNvCfVAXrPxaxZzE77Kaft
a8ugQHi+84GbIMqnBoETrWoL0XrM/vNt9tGhBxTl3/2/u1ypU6s3gsTGlEd+X1S2WqJdeCft6O0q
AEVYKi200m9uAYKcN4OxlfZXJJaj1lPVIGbImza9bClC0UyRbkBFwjQ2YpqdMhOppqZPkjNbUjaK
VHhRoVP0q9KXPp/tQVKTsstnDxC1QKlVZu+M6sYdQXSRFXVm6Ahu6g3/PcEu2fteWEU7AVLGKmiL
UVYiLLsb38mV2D9xH9DgvQiww4pIovdlG5iujPX4z6Yo8pBc4TvB2S6n7iTsZDJD9llQOZpUq7Hy
Ul354DgO5QEBdwypdWD6r17rS/2m7YHNtHXZoLTPO53KxLV2S8dcnT0KeAot5R6fE1vqdD/XHSCU
zcURMlwsq1H/hBqPbBw58sFSqm3lkal9ORwulz8zd15hkiKOLkBELZw39jmLRT95mcJoOef1T9+x
aCKa7PnN4XcwQFgogQk/S4I34oPuvH1yySI6uMyRdDyK9stPlwjodZ4z+qyg8JB7FhGVVfgqEbkT
1lu76iv7RVt3PkKHwIUAavDKdcXKtuT+fEwKdMBoMrLcWtnFontUTBe3UHFVsHDKD+XPRMnOzqoN
bQysZ3PWCY3Sl6dw75qaEfmiXSy53P//7Ny/NRVvjJBLJJxi6ZAhghCWjxqgfT93DfHi2WhX+yc1
HOtl6+l8/twJYvPsYoWBLhtMu8ZCYqQwIwmKcdol/ECXNNIHhVeCKmd68JH8ZKUQS2oLqFLSFBc+
iayo4FXSDhiCX0FWDkrnhcbA7IH1VuLn3npNh3klfF9iZ907qNboJnUAgboNaMIkvE7T6FuckCJQ
dQRNl87oRJOYsAQzTrawW8CGAt4A/1J+6+cpUboQ71dm9y4iwfhKQrmpl+mavVDgnK6IajKXvrBa
qNBTzxmMsBFFmqywKqGMZ4CMe/7AOdNggWwzw5oH5eFrhA+BRBFXMqOGj9avoRxafZThFjCEtDN7
Q/j4JApI7wv59shnhikQhBHpi6yOyodT5yCaznY/PPvQU8v1hIHa3Zfb6sGObRPh2J6XVHussWss
YWcw/K692C1XFf92tTCT9rz6BtL6z2uoy8QtEV8zlX+lkJ0tsj8A45P0YKc+PvSZxf87rNOiIANT
wIoxXUX4Rgc3imu3UDKdGnALWjU/ZZi5/pR7MsOnifJrw5KxSK/QSFOSznjHN6M5yIuOZp0Bc+4V
zbpomUD7GgU1FYUoINrj5cdydFftZYrxZLWoHwTW8oAfWobXtHWNrl4Xy5JWfsc+cOZrOCJYUA5/
UhD5eF8LTwD5rZRoA9iezWIZEEI/R7R8hc4oS6s9oNl8b41jVpqrdVbndoboyqmK8UPsPhsrzPW7
l6sSzYd2hhgFDp4Cscc8iV5UiYvd4xFqYUPezMNjONoYNvRWWzK+pv2PxnVcoMCxW1f88Fy+tszV
tVot1y1vpfJyqhH1i8vCNrK0OM6uNW4S++Wr+AhqnRQ/EuZhBbhWjhWqhNZkXrsl11XXe9qL03sR
YHM8DUAJbgG2/0/bzAPi/fzBO810paxq0AMV3n9QfVXbHWacYOq7qEOH+RPyI6oqzJU4A1FtI3z0
MeepGndw6RKQi5Y83det/MYO9yD1Ixu6+1aF42fJeZBIUymvdxBKFXN/fsDrQfPzygsvb9n+0Rr9
3Za7mVKcSWtN1EpCK17IocYvOsch7nYiFjR6T3fzcNnV9clI3Q7qafgL590cngbm60rDoP5Ub6Tg
v+CvF7ngjkayyJhGxrYlQVVzXb4oNTacbCX/Ydl6ku+dIFRewNuZgtt+IwyYgfwuxsE6Gpup53p8
3ayFaCljqMJo5dLbAcedUWhdgpdzHJf9UUdSwtlj6gPqCQgh4hB85vbBPi1rRo/0MhQuh3+L+o2T
d3mkyIQroRmeu0xJRkQhupAw4F4CuB5DaEg9GKjulJT3IsxgZrAbVH2fR5miB5zw69heGzI9HRMM
J5t92DF/pW8Nt0IArlk/rYLF/gEH5MjouVdvvQFSRCXvjaD80vPOqxX1t1nrw6XaeyoV+pgtSzEP
R3pfUDtTg56+7ITBhHpvEw3Mey35r5wHwiuwysaGE2wCUhuUDFV0IH/TC5KU4nCNHlQHdNVmtJ+z
I8Qc0B2pSsu7YIQDApUQFFpQu4trTdm+kSZbhbV35052ql2YzmCUyv9U1kf2NU29wUe9XjYS8k3f
PhwnBb2CxPcTI16ROxFTpD7xHAB0oHTNTx6YDTnHX7HuYsyeETigivSDwxf5yAMu9gTV7Cb6uxjC
GKdRYWUeAJEkGzpefD0BK/W1J5MyezmFIAAx5WRfRHzpJBx9mDjAGnnUFoG5AVqAdyvpcEsDMgGF
f8k+NVsH/dyI4E+M7Dfio0FJ4EvmV4uCZa7WzV6TjKMKwYVlfLW9hYd7a9pAjmoGf0tqs6z9lyMK
Pm4kuc57nfqTJ4A/OuPGOm2yN7Ol5OPUwVqMOpw4y0e8KS/HlIu/FrsCg+W0433phkpJRTGjUbyb
pLY5hhnRhxuBwYnWg9ZuMj//QznMDYolkd9bqdefA/Lbye7XDD+y6klUO/6KXcuk7vo6g+5LqN0O
oB5kv/M8nHxyYJDfEMrzPAdnQFBKUSC79i654Whmqkgl/Kjc0g0T3fxO1f8iiBI2BeDcO/ZdiW4H
U7AUkh3nd04E2V4jRa8vDooicFtwsTcr2hIN2aBItzSeDD3LW6pZMCuiSYVnT5bSIN4jF5i7QQZ9
un9FbcRJUhU3846Ysz19/kxuY+NgdCz2FXc+Ny0z+kVTMR9K43YwZPLpR+KOItViDKVXdf5cghEZ
ehFpibyT0uNpMU5FvZMDI0tQ8T8yVDxZK7H4hFPdEOvp4AamN1Ht6DTWLO8GAWzMX4pC6jbtJm3O
eqbxe3yiP0/EfN5m0qkZzc4Znw+krKMQJf+FgId6IxxkeUVnkgit2GtFpXZx/5h4Xrjeg3+8mln3
6k2JBLjWg5qvHfms+oTIXX/zopssROojUA2tonC0F2+paEgtEd1hC467BLFXK554n4EzhVE13FIK
G85O7dDtLJORSqiN+fy1QiKJvj7b8lgTK3NaYexuSbnRMPzKE1bshcKhGTmSEcRAQj8bUMLxqZJX
1+dFDVJplr4in0jYhFylf/QIjal3onlL9b6ECwqycmfnd+0QbsafgNol+T2nvxvCge2DSRciCgdb
M9Mex9hApoPMmTWYJH2YVxAd+btbEm32IkCBK6YcaoNH29SskOEG8eFPa6exeAio5AY89ojlFUKj
uB+BPHgGqCmDrtV3LQp9yU7LtKfmqF8UOmpHqeUaOrUYz4YBTh7hxnlN1oZN9CaQdnOQsbVI/aZv
ATJ5HQDfjbBhraB7n70eBWMTIcuxIcn5vApO4VP8PjgB4lPChnLTYQVqWMiORStfUKT0zuJgb5U8
JWwK3D7Y8Gx23EQHtHHZgJh6GK5kAkGUA2zlaniG930KtP+U8P6Vvr1HaD10RQbuJ8FS7gOsdTTG
jfvovsaqGcry5ZUxUfoTHs4zqWylwieKB2he1TlrpXWvVy3oo813QBNUwJT93kfOc93hWBnByzK7
eFDapayKBt7QFQgf89TgukGDOlBIEHtgDyi+UiNPQiLm+fmmMvMeS1g91nxdjz6Fy4bZildsh4uV
jJlKwpkh0OVNDj7xiYuVyw8IarSCucrZbiE/vIl8krRXVnwiXBrDQMFJ/hae3UcpMsknRIHjEZuC
oyDr6XCLXOxIq9e6CzcmHhSDy/R2sJo59eQJugWm565biLZ5hSsAINFQuMYPIlX7nfJi8Y/aiAAr
SiAc6du+AxjjQ7I1Iv0SvU/YmVk17GluflthIxXia2TErTk5koGA2we8N3CM1nitnI6KEa2R3tPN
IXyHSjJhNX5/EmVrXgsJflc1G4mB3FYKG4cwclUVo69/bw+QkxUIhMsMp6pYvtlA/Wj/1wCOkDYN
2tkEG6rnzOZjrhczWnfjc71tx7MvOOJp47Ny5J1dHAXIG3PnmLhd573/px+KOLNxRtWs7kJ7HpWC
zqH0yZDXi8sE/4OmlRsQRIbmDw6yex7dqHvA6SwcJjbbvvmH7lOnewaGJOjNR1Csd3Vz+psg583r
qN/N2ldt5qkiNeGniJ7kcUW8o3xB/K7OLpW7pmym+E4bv6fHxMGQ35AMLWZ7Az1UqsMq08ffBn73
QUrLF/k+Rz28zk/6mtxhxxWF36V/6Wiz896Xxt1ZlQ+cpbE/yNPiniDjhyEJvuyXsFjO05RvbktH
60fobDxGqXJ9z+bzFUuqqmikZDN9c95NQLoZb4wRE+lBy6xcKOTGPDb7UL59I75tpQ/vTi2j+eLH
AaYsFT5bQas27iHyi8F5dfOnIseKyyTrpr0iBHn4dwrJw0QTRjV2wV1RgyNWcJZO2K0TmWZt20BY
54fRkjymc7FhxXx20sdpGoDR7YBikR/Gu1MexV4c4ANQC5agI0unUiHGJ6RamymWI9CBXYAQ5p/L
IId12EimA9zQp7QcmtJIwMgYAH72rwkIADInHIFGDornURfdIEA55KXfOqiHd+4a3ChuWWI2ss7z
mUXZYtFmMEG+jDTh/h1lDkgQdt2Ji+4Mn9G/WnJXp+tQ50nFLMTbCKiO4gOIebhFJn4QiOGOIQNf
W7w0BHgD5FKnLD7xoFdJO3ugamQl/LUr7jl5g+m7J7kGxpLDJraVk/BwK0c9Es/QMo3/24Galp9J
EwwwW9BnD5Dmoho13DNbQEvxPYfovV24By5yVK2linqxCKdTSvsYnIrUpMy7TVJSNPDaYnim51xt
CGQG545eMPOxpmFLt02zL+6QIeeCtZQcX6pRoki1JAsdudvcuIeQET20az3q2z/xxQxF77OKfSIv
wvuwhqiTPCwJwMV+WVkeqSRocindWq4D7qIJqUKh22wMDIIovzZNo2rzjJU3TQYRCywVmbHwjcGH
cBHsi2tqugaKBxBoVI2QNzuy9M1EJFpS8rEg7jcpZu6AgqWc4WNfcd6UmTCb/oKf4kAeO+spoY8I
esep/z80AJlL1y/3uYwn9+YjCVDLrETOqsIrqspvDicF04qUWWKPoCHXr4OSIxCh46mn8mSsj/Po
F76piphmGUWsIz6scW+ybnZGG3X6iEeCvxaFxhwJoO+fgEivrJZ8KqVf8aGJd7dJk5LCEuniTLAV
2qq2xHFBnu+E97EiupqCVvZAuLVJAICC13TKKym+iLc5OSgrzoiDqqOuoCLBCAAKLP2I8i22rMVq
zfxC23jQOhWT+UgKWNIoX4N95KXJFinCVYJ5Z76Eaj0UBqf2HJvUIPzzRleNZlqBe1gMyI7bxqdr
U40GstEVYw1ZIT7eSjLSx05/JbrHVRkgztOG4Se7/bB3WozuTKvjNrNYw7Yz3MlG5SCAbjC+sGyU
brcwlnwzaAI+pC9yKsdFp+qWCwUT1hfT689axuBNP7k+We4XdLPxbNI/nTqvMDYuemRl4MSGffGW
1oQXQHPsQxYNb20ZsZjTtibwd+9QoeSSffedgx5QAfk1Cu3WUCUdv0i3xjQjhhT7BQyCz2yLvKbs
LDLdSly2wkVN7LBW0vt1Tm1wUm+X4o802hrWkvK9dc9khIVbPVDz+bSYk8+foev5D0H6fllGhqYW
R9/2S3zD7Iuyoo0+i8tJJwg/GAXujXqgG1d4EZvSTNhcpa84w5YOi6tu2D2eEwEc81RiE59SyS4V
ClijCf1h1ty2S50SpVyWaJ5D+YLYZDfGz+nJ46anW9/aLLW/+mXSFbb7FR8YzPNXf/XYlot+ml9l
TIroM6PdyzpLNj+AinQIuyP6MQ25Tq+bWdnC6Z+XiCg1E3Pyad1dCSPeeoP/42WYam7LXpzk6dAT
XCWM/EJGKMb6StN7X3YHapwYGizd7bIQTR+08GoMS83csp6yB7UtdLbeWbNiw0J76jfq38tCbU9m
2h3neWCul4qvDvxapJNcZhubYc6GtkEJWpUCGNxGphcvZrU8OcWc1X3TgwOuUcAdIkjFIhEzKfso
OY+0oX7AoCybqub1hxDhZsHm5/ojl9NzyW7t+TR8BhXkn/bmmO2A/l95FhWN7frs+KUJBwwPk6dx
oTQWw5MqTMfeoH44YphyJBq4GAgX8g+fNIfvcB0x3QfvuawEJnCwpuL5bKYA2SxBm/8iuOthvz0k
aVvmqEOOR4ifhRfcl2wKayIFNsYvKa1H2NLFvbudarRbg/bNsByZJCkdA/NgSQi4pKgbnOiqURZ7
KYdk8gfGYsZV4gYKMRaotoRK/U6looE6VWRfYopzcBYsVcwqoSUPBpOUfg26kScvSk0NXVz0Tsyp
crrm++tu7knlfG0zSvaOXD1N6lvMov5fIcpMcb8UNWTl960wkQhVBQVxKJX8II6gze0+xHHrQJi2
74F/G/LL10sdby+ZewHB92bju4NZJNB2ZE4tsPG4a0x40BBdy/WwSNX78wtqmHNGAsL24dhbbTUw
pfvegFFcp4PzAeS7FwKyCIC8vJTi8ZMXGMYR3J8Vu8SSMtUil8wKhxPUd1OiJ0Jx6Uza4Kpj0K5j
h0stApLpxFh5+UMDdHYKq6GFQ9HUkkJB0ithRd6zKjLhCsj4V81kA3ir6Nx8d045kQODwMHrMEVC
2gzTN6D8z5gdCqKfdf7yiUbov/ipJldgjmsBI8IxOWv/4fOUioBkT1FXxiLDTTT+FAgC0/HeAFUK
neyy9PDA8bAy+fYpgKtTeMgEuNu6FI6eQbcZZYnUoyZF7/fJmiAucUMMIA2mp1wUt6V2o0XeeMZO
BLJIN2l9f6FciqZhGw+sSiiw3bs9ngM17KdtSM/ZNTA2kVguWFAanV/fBdxhKQRv70Rj7oYHV/vf
WEbbg7kPkaiXnWePiV4aS+j1+xF60EAhti2lvBmxWvCbg24HUSMR/WRmYCO4uzUdpabSNEkv/bu3
75EuR8CkIGnr+dY7KjKDO6B+GO6T5FtRXljZq2qEqzykvUGJeEXZSuTyOTNEak5qgqJXuSvMLwdA
fCdBJanFtInLswZoWpdpYixDsqOvrtltnCUq1/FI3EDPa0JQtLBB/LrL2EPWWfvhOI9sDteFUyhS
SzekSDP0KmoptLfXDpNNMvVBM7Ffl1JsNcSUk3NdWtObdvt+M9+afZCmmQtKHMGaC79dfZDY4bZ3
N3vs7lkNs86QOq+ao1Ula9jfO4ea3nmVrtAaopzuIc2cSO7R2fgf7gWIiNXYOXIkUP0ez8z6d/1V
krWFDYUAlDDiyEk54H556rjEZgcjqPmiuO4Y8Rv1teJBMLcmFFZVoMykdp/2uHqaIkep6PwQsrlH
l5xlyZvIf0q+kb43mXdXkyU8jSRSl0frdz/hzI36w5EllP7t+KepdFsGIsnPmszAaD2nlmHP0QyA
XOERWHy6NdzqvH8t6dNHC8JI9jOzTBxasx3gkdqtC0zsrnsvESXiZgpazhe1bYrTUxSNiOh5ebGr
iPdzPSTiWwiy1V6LTfYMBsPqfN2JqAz71CdA2M3zOhOWFiHNT1pM8SdEVjMvOaXqKr3kJmh5WDgS
+sQCCwp/4IIeLW6iuX4vh7SfIg0YIJ3F+qxQv3BqqF+BWszLaTEygybgW184tjlBydIazxXZLLPH
SrjOIhvK5C9EJ7IQGdqn9aavJYR8xlblVUtW6/D5L6JBLQpmcOu1yKWC5Ga5cw/n5Nxd9OwjFGGm
kfDbzSi0gQZ7jUiqDmIDwQ/h/n2aqzy7B84vbEo7TwupotoCDjYgsx24d2fAe5QO1zdMJHWvhZsl
vsAtxM7MyJnZJjQwdAqyaNNjjOmFh8lYWc3vgcxKE4MBErC7nZtkrM0Wn63T+zhB+Y7ICXKnivgQ
IqaXKHEDX2ThrrlyWH5cU9RBcQEipAR62g0VJ5Sx4dlciRhFpgw+9u99NYySovByAVeDmT7QtmFy
yMXMzxcLxJy54gKGNgPWPF3MAoKfpm+uQHJ+aBrveo6brSsuGK0qzdjVhVQZTYwtABgi22rE7n1i
zx2RiKPTZrWvG5CR+iOKMbVRUR3/JQNOSDV9eehyTNM/WlDYXACohP48cjeHNNXz8v/KTa2Briup
8wTbZYssGT6h0i6MpJuUwmWDLBbnxDt3U+YOkF25BYLYUTlqk4tHuWaGlh0Ox64F7fEfg46rVCkr
LO/tV9dbHH3D86lluucca6ArXQZ+ZTnppC9M6LdCZSqDwGxtRNCbThPWVTsn/iWsQOI20A3fLO4d
saUWQ+mi6YpK8fmh6Ts7j+T/Vvauq0wKd2WjKa6vQtpKn3E4fSsfyyUxlraKTt0CCJU6Oi1lCOp7
fXdoLkXQMlxBKOwnZEX8DVHKTG0w5dS8A1AcukExPEsLeAIbiUD/Iq3Eg6wUq2i12+CLEp/frsPO
cDxGp9fOZNL3SSJdwcouwKCbMRq7ctPk//YSiYOvKQJt78vcGqyBs413Xoo19bToW4hhYrXAhvYW
z83tJRE3g2abCtI5ewnDxRkuorGvQCE7/UOf8aRlCIUsydO8+OYNH2MSspJCmt7A/2/B5M4sZMSO
bINiAyNiSl17d09SpxKnMHDrr6WyYA/5vCvLLfiv6UgwjirigXLfuPoh3e1qgujvxKT3ZIqDPNmq
JoHHQ6eHOZ92b0B1wpTgbSKTvJ/6x93c06WZp4Ljh/bAifOYF1p9vWegOkgW7Skv6p2Elemlh0rS
L1grR9Vzcz5zjc4i/Q1IRKhdQ57oYw8BaZQnnVhTIhzA1NPvIE+8PRBDwbgNBb+Yk9S6KP1gIYWB
niTDOlgq1jPPXaLkMS3bjzXAuo1/CuNA3rXMWoUNbOL3M2qNWRg0uqlh9RxDFDYvOx7AA9W9YRMG
3OdVLs72M43eJ43fsV6IHEsUG2hbHtsf/yxcffPYEIfAQiLJuLdSJDYZbteGBIVSrsMt/k+cQS4Z
uFafVMXCnO7ltIGZl0YrBXl0DaU2AHpV69dODi37NCn0QysV7Z1Y+MFKyAULQHdPXFdzXj+yQ60f
wELTtcPfT3imoolxfEfyoV1C8mhV8gNeQwBjQDuV9ZYYsCfgD0SDNJeTPCHUPugilRUgdIzPuXOn
X3pi0VlUw3i1zDdSSZO944miSk86rFN4XCA7OnaNBNbspPzRMilI6qSboZ7JQvkfD1LPXJ9SUI46
fjdjEAyc86TPgyymYUQks/e/G7hifttNJh5j1GPy1Ra9vHYcay20eoUFsbEBsQtcvJdAyFEug+f6
f3EQmQNjWjMlnj7KamxJrbezCywfI2YXGLHp/IkWrRGFe2/KVP33e7mvrxhDLQhGZpxguNeHkn9R
QJdUbHYuLylEE/N/TR5l4v5/dwCEoLzk0gAmxbrJEDs8HJPS0EClklz1AR88HCk6Nzha0AQJhb0D
nLk/ObjwlKUxn6W7mnb9TUfPU2R37rIU2dXCvZP0oP834ShjQFq1dULI80x+OQ2D8AlIh3z+MPea
EV3qkve0TZbJhj8XlONXT41sdRbf2FJPaM+0tbFUIaTcofqLGkj5kCZVNVxCAQZBKBgIJSoVAJlx
H5tr7QdH4+u9IcUhVYFywHJn3kGgdz8lTYeY+gmLiSlQSwysmuWs+UpQJPv/X2z3BXX0HT6U6ahK
1uu6KNRlI6KBfJCycp81MF+cZhU6k9hJPoijTyTcfdMsw3w+iN4GRjkwZZBHnhDCDJXrgE4Wp78/
9j40Ok/RY0IyxdcAjTFSqVSuUYrc5BLrhG57mkODOcXZ0b4AMQy06MkdvT364xmeL7fAT/BvCB2G
hf2/Lki+CXd8V8oFHlUFhqWJOi4W5bU1CfH3J0EjLuBCVNaNZVrMMzlJZ2mGvcekJSMcSVHd9kdK
X99X7dytLD/IQ3Ue0YNK/gcurk6M6MLeTbseYUdRnvzu42GMijuyw2cN42g0SYF9GFO5rMWIwCBn
QejSRVjBWmP9XWqetcd0eitBD47T3BSkr34carBKs1yYejm95C9P/E2jV4ZZfqry+761PwfViiJH
BH8P5/fynHfN4HGdPTxCPMO06wBqFCwBmo9k5AcQK+WFY/VrmvNrZsnKC3JNLLN3U/RKxqrdCxWA
eUPB5FRUIRP7P1BEtX1GjhbKbMIuOsT2v6KV5wK2ayy4bJjJwf0Q7HtgwuqI9gmQ/pKwTZmpdG0h
9RvRIooLN57ROubhIHsTUT8kkKRTmWRFMAMYU1Vb4HXeBcI/RSueYYqMcktVxim5qnypLpOuJ90H
IE3XFMPQk1nVDNfJOgDV6ofEVj/It8QnmIngcsYlV3wf2easlc7Q+ir2pcucQDIIB9+r/JLmmnAl
KLiFGxCS7QQ6ZmaEauxyaYKPshK3QuVyMwO0pVCVmKY3albBo8J2qzoz3WyvJ4gx2dsd5uaczOq8
DqR42EFRsYED7dNq8jifSk11bZTn8J8JJL5/WYl7aKHDm7KunAy8kCDercRnYMdtpO0dPUc8L+V9
FNvA9/mGsSYmTrRQs9/HxFHt58EG4cGuPUaPayjtlBJJNjWupHXIUEywX9USO3KCG8uq2rqBB9+v
ENIHMrSo1xSq0gSzWXCG+lYRqL+uVwxRvt+g0eIXFSnitpTqnHUr/cg79vWBzWQJWEqOP3aojP/M
mLZzfK9e/B4liSvrXve3V30oY4hE5PhqapaVydvBmaUSI0jeXZ5zTK4mfywvJoQUHQczw398GL3j
OfjheOFHGzQ+oeDempKAc+LUj57H6ycmCPAasPlVrANecjYetSys4PAcTGUPW74iYc56WRgGwg13
ZwQtkQnN+1J289TLDQ6cp3ibNdreZO9ndoDquMYSmeUaJu0HfG5hFXXWf8z93QwH3EDSEth+QVIp
oGb0p2Ut4ZcfQNz1qR4qk+I9JOwu584Ys+bNwot5lOzqQmrBpIRdCkPyVC50b/iu4ySaZLrkPaRE
UOpKuI2MwNoCYcTyTzSkl2ps6FM1SZ3p//i721CH1JUnu6I6Gb3dVsYWigGQ2pq0VHDLWPZ18nQS
ezZ1LJPVa1jZ+5PEzHE7lB6zcdjMmnC3Q3JX6E2d97pJv0Uh9LwosrwQGGndngOR9A47futSwQiy
pY26goakIUR57Ib75ydqZCOxITGYtVzsVojsdWK4Fp0RHtgcWV8z/Z83P54F5nyswA0Hweed1UPf
R0dYzshOnrZTZJvsLGyQj9cBmJvJUSzoaNNY1asQVhDAOhHl1aW/r0GeQZRsESYPw6UZvsTlR4sJ
+fvAkqVsHFvc6wp1u4gCkISR2ZCi018AwMsj01qXOozTWXjXX8CrdY3IRixAiQ609NmMNE9bKowi
4rgD8P5Nypk5mrkc1PTtDhWaGWMezT0ijckiSSo+XmU8+LfWUifY7Jr0Xz+pcdGkIHMTx/z8AyXA
O+jDt/X4rIa2zJfkB5K2u8M7S5g+fUORMs7CJuqRKK0kZYgvgOcZ2/kFTkY+7Hxy8YNCUPLAmreG
PiyloDqsCc4//ER92RjM61nHxb6ddQqfOJY+nQAWii5mw3UiDZuMX0N4CNEyes5yie6xr2jXgYGu
KthlfJPWMB3qdT5b6Xy7fzW+ryeqotLhkhZayOX5eZn9JCHXC70jmGQo4fUjzPGJl/0ovUe0CO/n
eT64p4QmmZdw6lZPgwLnutnqgsCG//1BqAWgHOZeOgQULcqSPerKShvnDspVfGZIp+D64JG5AVhf
qQ7YgZe7rGoB5hIP2Alz0J1HUi3PeY7ATCiIVuV6OE96483ubzDJZa9L90D3SG4k5EC9KWBUFc3x
Tc3SZiZWKwur2D3Ap2eX8zvbl5zUvpA1n8EkKYJcBe3bvI6Q9Pq7qpCNHmlK0pW2RTdMszHVMVVc
t0F2IEVxjDFfs98gMkq8MX7339ZwDkCdPpqYF9GrZJEtBwiOGx9wiksWOwK3+FobiFfeU7CK8Zws
nEuh2a8lORXhDFMmnduYUCdDemi0zsrPAhSQi1yI3c6qh/9C/D0xBznEpBzTWi3f040OPwyH3yIN
PfEJZnwEJyROC6U6AkbMHxJ2r8xQ3AdGdj0XEud/vXMtGG2iX3rPJXCh/MtGDYwAoNfinES+Rl21
gloXWv7aRrgFUe8EYFro1JXASM91kvlTyaL7M9URECFgjJXJwMUJvK91nliX7DxCtbX4gZKu9XRw
fh2I7TXiF97MkjziDPMG9RpW4FZ+seSDXipGwnMiHMkaAjKFWp3UIHdevuboOEZAbcvN355amzMz
XAqZfdDpmC9T+jhsf+iLbm6WKlgiF+s9f42/vRxKyeXoiatl2thRmZA9TWs27h0VQIwgOJZwZv54
s0VveznjF/1RLtNbb/BQdHKhEP2/+nKR5QEbd8p0wg4+1GN1urEJqr1vJDClE6+A2qp2kugZNlE8
4cDZG85anJrssufpVMHm1KkJpx6zAnScyo+1AzvszL00jfZRFL+7y1GZO0jtCNckS+C2XHDYmST5
mxdUgJE4sZ1e821GmObwPDr1yUjAvtuAohv6hBsHiXGwZWAegqhuYxJbutEptfVXZyx656bT61HY
PMOnDiZTKT0NYfKGmelKm0GL7bca74BuqvwKr/arGSPUwFa+qjx4zFfS9b7+nQi05sONK356i9i2
9WbxOWTD2htkntpyP/OtfeE0+JxtoPeTmm7pwkjlf223f5zsb6tBSVOjwDS1p8J7i3psfGDsOXfv
nydtRS69k0O7WUrpdXK5g5BYLZ0DQwBjSjrJKyxYkSJlwjGEniFTfLFQ+6qALMzyGGWi3rtHQtvu
6MLEGg8uqS0Z6CWYKrV2Q4mxdhVuTS6S/uq+JhBlrqJdGv7Rt5x0NspYrjhjCxYbZJQoNrst2imv
E9q8aPx4snpxybFlHRxPTohumHa2kQ6H6u6JQjUjbxjYA72BgDV151+7NC3mpRmbXR4+QB2KEYZ6
RXvOxR0r5Atb4vJcKZyx4cX7ybMMp0ocaZ7ZdLCkN625NfMFGtUEkxxIQA79BenU4yx3WWJEOHir
M7LaBDFxiR2rk9jKK/1roc5AYXPL3I3opLDeGwZo54nY3Eb4DCiZUqh1fNODkRfXxi+04/QICyed
8OcA/0LTUoiXZS9sWu+ZUrdHUWzlcAtHZ4Djcig+exnZ9apZkmEMbGsHXPlSX13QxW7WDyU+5M08
sUwrpsXFNv8cYZs7zb98FoU/abFNixiBRC6HN5jQ1/Fglrn1Fwh5eZoY0zM5LIFFKY6rVKHlPAk6
9dzzqpa2HxTRQf50cmI31aB8BLpyt4WwTM8+SNCZtUDN55bPywVPXZk48zXz775gaIFejA2sGmIz
O2snGWRy/EwbWbjwydsfecG+kx+mi/FwJTstQ2fWDq2vtavWwjHWZLILhQtRxLvssntazpL2ytTa
YVtncStFl63phOTN2xrWki0w+fw9jDPTzq6h6AQJgIayt5D00626LSMS7PokMsixmRdtYtoQ1afK
bsVJc37KtPrBAfET2S+RlfWAs8DRQsho/+N7BepGq2p5PQnYgxnPDVWgHuOzRyFElnKtbPw0Rj0e
LVELwYLHB9QmOssM0pLKMvmvqolyS/hXFOevifBW+OL2b/VWwUcf8IZRqppmgt9qy8rGclEOXian
tiFOrf9Vti6n/W9tKBOlY+PrDiwpmJDkQEWEjj0SAZxliE2hEOV15kym0QcEkyxcD1HIIyVaZ/ur
p+6MfINTDImIvW2Xu21nIPOcbUeFdEsc0Yr7S72N/sDGtEW015EwYBSTOOhGYlrnRL9fCRMVwjbi
FkpEuXTJx7RnZwKNGbBJkUoDBZKtIps/QdbpjG07kpPp/+6n1UqTCNm4SDcX/gp8zgVd5x2srenl
w7RK8JKdZwy2jPZrC5zG9ofMaJ5cJ7ax0+UJ0xmk5kO9UiSuCIlrZ/zqxsfvaDZCXIBBVrFYnZz1
ClvTALrkcJSjnjXU0+Zl2jOW9pbrwiqfmv3F8QbvjxIDN0CwAguoeRXvLr41ZKPtiErTzrB9O72D
zwKkXEBlpaaJI6h3knKInh7Fl/KOUCN687ti63QC5RM/3lhafPU/g75KLGPAfhEM+Zddukk8WA1z
uRYnWmGPPCoVm229DL1hswWmnSQW8WmMjtEH2jWfVZEV0i2vltxkxvq4vkYNniLLbinWkv3J/cFU
1cWuWEmXUJZxPw1OGofkGZrhZhYjQOAhODiBLrnTw6LZORPklj++YCMIGdqDoBZxeKLenKmCpgT2
4KwbOpx7fvuIt7GLBAnvngbRTBBJo7MxLL9xk+gVyyd/I0x4SAe0Qa8iiu182O+cErfcGiMXsBzc
n3IxtylzxuGSg4Ch/3tp1TSQww1/6OEiMRwecG7bvzr4L/OLh0gjRjg9ftNRUz2ghhZOAY4cHHWv
Wv2I0u0/5AlYZbI5TO5ZDtYFPYWeytmsVJyx9cLBzAarosMYPxyg3DJODshts00iC4HlkQHiixw6
i5hM4fXniKgYzW5uRMIjVQIDoBqzj7+wAxi/xje5T52fn7wLWULb8aIpDJn2Pz1bbRxUz83pejBc
GMK54rNtkskHXClXrbmRYtFFQzEAoi8dZQAhXyxPSgVRdEtYRfJB9R5EbYjELDrUvBbDBQ/f1JX8
ZfuZqvpRXjAVIuzzKCvNmqeqBm3QXiu2LiLVnS/B1i7Pvd+hyd6nDb1ME+UO4semnOvY0fOWM/RW
7QoVGPyZEQuHc6poEZgjhX+lL6+tBEf8ETdbULBCOwX4clpqyga23Df57JWgR2TIcmPFRIJOMcAD
v17fXlPmApWeAV+9p3VUCvCzq0Fii+EwEDApTsiULdz4WWB8HSq4TZ8ta5l6URzK5nfH6SbYdE6z
L+WeJma//KgNVMb7+xU1jEdb/wR4sYUqq6j9o8A/WMsVOWqNe/pI7DUSWyvHfg3Jf5BilUscJMU0
wjFf+kLZxAUL3zwuDrkXbJclcqdOeaFTg3oNI9gagCLIUm+Q8bABJI9yJqK+WX9fXfF5ZAvJ6/aB
C9rj4JOfZ0ughJoJhuhTYeRowUJMjUFj4lsOLMCX1LUpZ9a3CLBouaC49nZHwaYAue26JD+KNN8p
qu/38cjGABnQqGdGT7b7IkzkRzoUTZbccM+8rplYRP1KSYd0GnjyGBw6wBPaLpS1Hsozl6jfqkB0
czuXcNMy67J3xgYNrAAEnkGS4U7tTMfTniVMewxax6namFNt2nA+BRko+k2Iaj97JPZSUwFgk1L4
AIOACTeOuxSKXGPK5XQVErTIclSAwRWjkblDSkyfuthegdS8ghQdG7Rxhqn2lF28AGQ9AXXzF6A9
eFYWw5EgUoygBUFz+BZT+aiG7iaCcqktlcAuohK5CD8f2AXElctgZWeVAJu3FhCYyB07SiC8atUh
cnI9BmUnGTHGTUhJc5bZAnKMrgkGdJbXPoSOZFdaEGMwcLo6WfUymxHk94eU33izJwoRbO/1bOei
rx8gZxWEiwXCsgKySqM5xU2mv7S44trjy6GZdZUTmDRf9e1BhxVOxJZ2WboAKhNqSpvy0Uw9APw1
oGPudJnPC0A9YjDEb8zfHvL0OZfDHs5ZCT8nwZxJLNQZHcJ1R7jyujsS3RZkHXZu21Fqeh0WYsbr
dmih3wZpkCI3P2L7P7VtsrMOyZHxUdrh1/DraO34rQBS06bv3HTHXKcoYWPm8lXVyWVh5NHnLUso
HFMShUnLWlspQFMaWyPFoSHfBygCrFOAm5l7GLC2n3BFoSdJ0sL8so2eQbDT9mhtDg5bPLNM/aXw
jKG+z5R2H+OXIIrMtaIGkIHPnKIvbcRghVrvSZgp26Dh85MXVCcq/eOokqussiVC5WV4ka90daGZ
QEuhn/x1HyAqSetcYK696QDxkLluO8LwlYvVA5jkgh/3N4e+58w47dqMRrmRpvSKHO4FxD4EemBW
k8gZPSoH9hbGoGO0EW+ip51RzcxdDCD6Vo+KSKvCMCz6c5cGrshm0DK1Yf31euoLJN9xReprBf/p
lVmK1EdTXZd1VWz6UywhHe8OdEn2Nh/RR+NlStKTDjPUAeTo6vcznOG8AFwwIKW8tjPkWqXuG/AP
ZXyH12fJVYgVpPJfjkRhcz/WPyq8mer0WZFJPR2XUkSz4qImJ6wxx/4XzkfnusTBJ2Nbiu4Y4Jkx
Nyf/jr5Zxzn5rxZjItJ3PiO5EDxQQZ5mXetMGnKX0aLdphCX4oU5zmLXzGS6CavvWKoUVdA/FLu8
9xCa2SA/9fDUzjMLxH1/God+/7/eVN90SHoLkqHSoCLjz+NmIzOchZt48Iype/aSCmrrAGcS0POO
7pNKH/qWtizaQ4fxHv3wvnhc3GW+5qCHAerbDWJN2P+obNq1Tn00l/rHtoZ3wK4zGVLxTfXQXvER
7rRrCR4WQyUeXKtgFr5QdGAKU77GVVla61A1jjL5922rN5yoIROATbCklx6P1Fhkcgd3/bqNlKFb
IN5fD/VDuMJGuK/BqmSlBy8FCpb34T3hhvQSIlrE+uH+I/Ss6SYJIJGKyE2EgKWIIKnUQSRAo8ls
S14/J9n+fmMo7W0GYwGC4bwlh4K81s5sUgYNg7CQpnYt0RPRIiWucnEgc3Fnmy+n0Km2aV4HABDL
ifh6tzp61qPXEtMWf/EOJm+WfwcYUm/dk1Ik2JWIx4juIIV/7WxBmZCMiRyxgO3ehqyor/dHg38C
B5L7/nksp8s2LoggDTYixs5JsknH9obXdWH8zLElnJGrM94YlUjkoDToZKyjftev/rbKyXjIvlrt
h6YXApgWHsNK0f2fzMdQLSpcCHuREpfTFtAqwwNTyLD90lmlr426JJJRKtwA3jPB8hiZcaO1590K
5LVtIDTGO0n/2fCrC+XPhcYaTg6ZyaRNX7IFaptvq8S9JyLATRto5ZRxJn/83EILi09J7uCKYye+
d6oQIc/zZhZ4vUb9voXkGi+NSjZzF0eVBdbLgaT+bDfvWopA6xSvog7G/J+qVUFZjn26eqGUkj5W
WWABQFE63YYJpL82xFMgy28lmsZq7yGvapl/EXrJvX0lP3MwSCZW0n+HF84pMQolf+M/nOxQPWEo
JIXNRTtE/WqGcXsGT00aHKC3DgBhgHqjL7XnHTybyhU+FIWgWmAQPtzmPxO+bDO8lL7pVLiavdtw
cFhWuo6hfmTLZIkNGho8lk2RZPr9grAL0RA7gPQp0CJvuci2Kbs+7oJtsDjSRr2l/2/KjcnAtmSh
iGa92QFdBl+Z0SKZOBbAO8WZYSZbDegxb73WM7yxp/4k8ksvtfw7LZWVAmPzSz++EWVKisSAnAPV
UOFENK4ZomFrpOOK7n3rjia+tXWJ9h2sBUe//YlgCO7V+MVYXjteCuNz9z9nCe2KiVM/y8US6dJz
OzH7RhF+6xDepZdUn/28daejEOC6JuaQa1aQ4M5AopEy/UQUT+mCEALaSW6FIBaP8WovJvorvYue
US936r2iodMvnggvIluIxhHzGZ8IOsdNZ32jjv5DIagqopbygrTBhMeZoitXChsfeDlUzFQDByDy
SShn1jiU4jGTE5T0Q8TwCgLOlZY0hZixFHHtVcr0RBAnl5Cn3ra+kcceP2ixW0Nc5zqegD1ivX/5
8jImck0nyRzACYk1T1TPWFfiTYLBY+lsTyFyqmKW3UGJqupCRZXLSZCx2dG7Yp1LDbhb89Un9Ssf
YCLF1LluTYJwvoQNZv3DuZInkC7kvKwLEHuext9GTIqRHafNzTFJXaLZ6Z5GO4/LCkAlWHXABr6v
feV/+WFHP+d5tO8uzPf/4Ae8W4jOLb4Qs2Q25vQZ4rbfS0AvsIZkMcMUVVyJ8Ze3IAU1iMlzpheZ
VjcerJvSmbBGv7NA/+7XVWnklHlYUAaRhw4nh+uS8VPE+oq2NWs4NnQLDjTDNsf2GhuI48X+VefR
KSCbuvfty6vItBAP1bOpMfiRIhZTJIqAk8AWla0X0FM/t+snwCVrAotqSLBmDXpG6W0MIOfK2/os
XwTJRuQhPxLwvEO5lAVk63CLQag9ACZnXsbJ5MbpY02xHIljtKhN1ASe0Uyp4WpE1+7/s8n4lDF4
i3utyrFwV/HexM7zNP6XCfoC2rfABhQxHfIW3DuLU5DPU47vs2aRIGQI1pN+mVoj2yMwSgLPBDp7
fujK4JehFg6wWtsPZ7u7aEuF+jRbsTZwudqEfbKJ5y9jiJKBk+g2lFZiMDGo+l2rgxhV9rgDQabC
J7SGsXxp3prFyc9YTikbWakSJcF5PpNQ2bDjsgpREFltg/uCuaQT2d9rViXoJnThmHI2YIIWnCqO
yrL++vIeFM4zHcheR+fP+Ir7v/nnq8xqeSWMuooYvHq9GigXjGoWUSPinuZZXAI0tpLhHj5VOMVo
+FtZNwv4tqbcHwmUi5kLvDkKiO/0utEGChJjiA1vp7iyRP1zNAnLw7tMJtz9Yp8a3+J//aRCaUwO
Kza2UloBbx8VYAMPuAf647XhnHNapnjxzxqpxldiSHi6iQ/+zl4uFdaZB4ZNIAyW7JWeIe1NM6IV
MKG7E7IL9A0MvG3aXxaDq3sUXOwU+31b1fywSdkDK/7PRrZzi+2PsLYUxaj4/dkEdpOxjUYLoifd
L76qKZwQrNlY+7LHKYHDzqmUovtj6AbDS5JPu06/PnUN3e7VykDhzqBd38KfbFbvYyTzelNhqQRa
z0u8ssG50j30VMBAGAs+EOg7+eoMAXGViQUzcdpnxuAtwmlwkC/Q4e/JjFC/kx0kaZ8hcV81DOQ6
D6Ky76T3xwCiIByS8fC/Ga88drq1IL9mz9S6r39JKWlV48nSPpKLv8Z13byOq8Q68OfPNH5SFiDX
6NKhGd65vBN4p80HT6pu2cC6ondNih8fHqlJXXoOCw1TLk7LOaawi+fh5fZ87vs4EThV23K87OfT
nS8gOd1nmvzTypT2KyxPCCAYZ80OFO8BUvKjfQG6Nzqz+u8Wt2ntaWwS4bqpDN/AC9T+N1CqEf+x
Im71bYauR5tPh2HxkW33rkkribD8iLTiZuGnOOqt/s9PV7wMZt7Ax2n+3XeaGABo8JZ3nz+Nj7op
UzyG/myUDb0evUNBZHMBSzQ7EGZEze7x8HjECvm0gDFfJDfwR5YspORqWGpH9UNpM/ZpfqKJOu4y
z6X+oJB4jlpGlsyUcmxtbMp1sPNT/bqiV6bEYn+PlseknEeiOVKiPWbgdLvmwOBOdX/rb0WM1/YZ
jJqEnLTV7XApxTB1DkJZ81Kot8LxVhOS7YulXxa5syWOi8bQDMUm0LGjkf0JD7LrSbR1cPDSKvmM
Ayge9PZX/xpnwcSePyMvdiG7Cy1yUxj8W51lPmN4Wi5AVqfgs4lixhBZRRiM7aDcZT/oFzK7MxyE
0RDt9Wy9Eytx9LbrQG6RKRS/xeuB2HtWUac6DFyZBxk0AZUaoJM7V3mb78LFGtZRXc8xCAPoSjvt
ZGnKLBvIQ95Nk1z6JE9OMuVHWd0RECe9oijBd3gXCUk15kuTlFQvEtuJbqs/przF+ILCf72RtKRx
4ZQmBrRod0euNlCXD+ESwZD/aK2RoL/WWyR+IPeUJw9DiMBKmip3PRLceJ30YjYwYgbtVWic7k1o
lX7+nc1MzqJSEGMrRCcjnf5yzAsKM9AAaA5mHfgdEfCrQxBuSXetqJ+cV82vrbnMj3dUiK1vvxf8
4wF0GvNNWdjVwG18A1iykZRJAXF+VWoVXfEKjroOvT0Pj0Xo6d1IxAPgW3fiqGzF2+0tl3BdNJxk
s1To0inVTfcxXjuxKIwUnPQfC7b/Nf6ve48UUFa6QEVAG+zqqKnxWur/E/4dZCdLeEWsmUrLEZL5
jyG04AcL982k5rQ0Ok30xMctctUU/jHBVfZQsWEfs3Il/c9sEw6uPkDV4IYy6TvCqM3LeNEI3IWw
Jo6ZnqzSm41pPt6GtBLTqGidEUTsvCLr7yRLoxXsr5BlIX9mqFuHiX+GhhcmoLlaTV6BgEX6f9M8
06daiAFd2Hjpsfh5T7V7rRk4XFNOEsNY6j5LUrFnH73jO48xLCbPQITzNElU+is050jb0cpZxvFv
wotIWKY5NWRbdJcmL3MvBKOZwfxdqEuNSwrpw2CWrVgBcTvgP0yISeV1uvFZTW/ZTHh2dxm+sWkR
FHdMMSJ28Iu+AC3G3JO1HavzgNN1+NftRR6iLzdSASleVTR4FczLYjRZZ9P77sZ/eydS8U/BtMBt
892CBpkhDzKDYFloSi2JE9wcTipj/02vGowjTXGLaj9YmX+zBtTQz1G3MIyP9q7EZiE8khLPcrqJ
sYNayYu2Xb2DiPuYQMaN7mM8tTByyu0v/czuGZVKsrt/CYWwpHFgLM3rjwJnUjYsndZDCFxyppJb
1191zAOi+x4FiQY24gaNx6eB3BKYCNYjJPkvWB/yIu4hNlL4DPS7o3yy+ozwvxD7w0ZZ2cSnyXOp
R+021KUR9LoYCmB8zp3HL9ztX61cMwFO9gYlcK3zlQOLBv/swshV1u0A0ETo0ItNxXQS+Hgt8Hnf
mQQXUkT4h4PRY8Hy3aO/EEV1di1lAiypshVO3cLUgcKhiRdqSreAEthGU6o8t48Px7LAGUGvG5Ec
K1DIITaHSwQi+ophfYlQ/Gl0r8DPIcNDtydkdQ6QSpevAn4W2iSVkOqKIx074td+K3srWsSnt81w
7tx3HKxXHIPcLRUZH/Ic8G/zUNAlUp/n0UeILXjFWrrjdP8k64P/wUSel/lC5tROkVH8UC2RszIn
MTndc06951ICNtPgayNPaDe07w7EVOhGBUiRrU+VP0gRwbqja8EMC97Y7dzSgS0QhKYunqoANeEU
+6hMN43+wF8xLjzLACt8VmMTjszZzaLiHTGpJU/LGBvWhQUKACN6jIHYUZzakvpJ/79Ry5tTkRHZ
pH5eA95HC2ksyzZdRjjsbxeoSKl7lxIpzzVD/dd8n4jm5Y6J90AgO27oLVTmMrT5JM8aALnSC3qH
lx2jIszF4RH+cRjv83gLWRyYpzr8Jc2ix3wYNFoSRyCjooDIenhpdEKzpfgGpY6AI5IhBxun3C0s
qsQc8J4hAHjoZAfTJYCNSszL1o9G+zpiv3A63i6yrrHTxTrTAcUPjMgGlKdmxSoltTM2zZk+ZpjF
KkF+lZ/Sb/CDN+G6g/bW/sA8Sa/2eVk1AnX7wstYGNVylFZMLAW9P9tpAf/7wH/6ngEzKDxP2dNh
JbV4tTQl00jbelRfmjuLRN7QFNu7a95yGjLuiWSLHOPD14Y9Fwcped2NCQuzQmpi6wweAt6aEIV2
YPEKzu/wmFMjDcY/bURTorz0rGTTFXceectwj77kZpBrX4uxi+iB431RpFNqJ40mjckg5q/saJdh
we5kcKohFvbIq++/AlVNOYn65vM1URrujetVotVD8pG0a2iFmu8InvJx6iIKmS7ryLp8icpcX0Zf
G82ylCz4IrjiCnRzHti+WImuZjMr+jawW+fJx8wbDPwzSJKvlZeDfYERv/J1j3vv9+4kkNFcq8Cw
J/ouNLBFCh9lPPGSMUZvC+FvKoVEcFwliUQHA9s/wwvrH8qnSPHk7ka8qbE3gohc/boaNv+0BxZ1
aynvJkOn12R4m/hmpbnM8XF1FikZ7Ast7TITOUEBDr3Q6uvl6+MFSMCwMDjPWD+/TcWqYNf1N8xk
zde8aUUqN/dq234C+YKMHIELYnXzhwgOmAeLC6PdtnqSatlTy4hT0hYCIabpVUraISHdo/vNDj5p
GBwpMteXtBVvC3xd6/tV9PKNmk+6uY67lsqV0XKnM3bWgOX/QPYHE1RBulJ4YaC+ZJKk5R/aaqCf
YmB1BV9GIxfebCuO9lNm3R+lqCJijbTWqrdVuXyWSwjtyCh16mgmMC0vbLGBwiiQ78bbfx74MLa7
9cZQRgRrBXz3GTM2lRh/ZMwFjCRVbofMTkgQSU+e4+mk+UYxZ3r5y4u0P0rJIMCUa4nyCKLNy4LM
5FPSkR7u1EoSkpfcSNXdt+knEtkhFXpMGVVRFap2m9tHw3SMDc2MsZmXzaEXENB0WSrsyRu3Rc/q
X+hO54IAn8DOn+rXxTipbwWRdfryd4bR/b4LtV5KPM4XLc/6H6GSWqY40JtJYKSbO+W+zNr9ji5W
PsuK/e8/betO3+8HyHAIrv8WHxShkHJU3z4kRbEBNpWa/VYJeYtXKXqzBDDUg0aLfWgl3FnNYvI4
dnAysAoP1dPDwkDwORS3I7IlAH+9hnZkMKqr01A+rpcv2yTTgT2LEuHySZ+k4wXV83AVIrlMRIIu
OYrdbwn3ulRq+Is+kl6Zx8ULUFxrmjQ7/P8dc4zPVE/wWilF5nZ0wlIJMZHY3V1o2LuvOeRsRqRt
IaCjy5x3HUoO1Z/UAkAER3jf8q4qvXR5In6LUwlnpq9zfz7v/ek+ZwZc8RJfVAKiJyq1POYpKRAz
Tah8ty4iwzrhX5JpExkkSoPvP3PRSLo8Ms5p76pnOmGhafYlNTYBcC33ZMZaLC257sea5B/sWLz7
+VLjc63/UxkqnCRF5UhRDQEO0hUaA/yC3TsFcbKltwhqGDkiQqpFo+SXkoARg6bVhUlEbseM7DIW
B8rLi2JBMS/kMIFg2IsvqAQAqxCZqTWckkpygZhAqtZw7uuIvE/7TmDkj7KROVlTEGqnyisHjqra
jULr4Ga6Omy9XtFIgQPSsY9wddmfapluLAtC4g84GJq64oJpZcXtixlxrUBvSp/91NloWWFQCpOT
X/0B25prKeP3b9Z7kl4fXwSakpkmsclyJ3Ucu63s1I07JIIdTD76VM1Rl1tjKXIxQWtzzZfd6i5T
8hzgCpkAqMxfIUDl+Q7lPCbhipX0fmeLPoxbAufWCNM23i6RcaVsc0z6qZtzd48P0s+Aa2Ef2+60
7UO+jxoSLfXHuIrW35PRdBt66f5moZVLh4TMXmmqb6uoR9SrDXtLqpxV1nWKLtEhKvmjf9VIOmt+
nLxPuw6SNNes4eCy9XzxVSjvlZeDQ6CgnvQh1MQatnduu71Ce2xSy0z/qKtcFFdXU5wL7dx3QV+v
fFTNTOPbqVPN7RxDIYKoOwCl99HaVyeZyGGTUw+z3IyLKeKgZVfx8Lz1fHJxLCtpwPa8T+Jq/D7l
TwmmG1Bv9+FKURQ3QbMP10StX55lBTVJDgoE9iMT2WjOmiWxlo3fllQtFKLNDkRpxERf0s5bkuCC
miMsBA/8BKbuOr3qsDE08GDnjd0LxY5sGaxl1PyjqOcdxCHzFoJsLC73qopeR91XlBFe8we8DNMG
DPcEyaHbuxosNzm9c8cJaa1p9/ddyNMEZHdRg4YJszn9GTXgrXBPb5KFSlqSK7egD8VziLVOfF+Q
8YnDMhDZvVpXweLmVRYKdq0HGO1ms2WRIEUPDkwqnJmVcwsGF4gqObP4a5qIAV8RVlIiZ78icxhs
hnwis24xvDz5HOD2dDLlwaZUK5hnnygV2TAwZmN7zcGNmo9RnabF0GdWhQaj6LEFceItDDLxcgzD
RtkuIFaAbYCYxWb13X5qJh52pPujp+O7B4FGLMBI778nZhKozGC/gfJxo5ozDAX4P9x8wrX0GDwa
4sBZoVHnYrQjkQ0ga61rLop4QHdhvNU1Uv76pdFSgBzvAWlKLrG/ITI5MwqxGMdALXTmlhgl9kxX
//sT/Yrvf0tnJhFipQeGk20Ff1XaRl4R/QV+U0EBRNgfCyENYeMZn5A/e1fP/aJWKlt3bAmYxhKl
UcIBoJEQ4tYGFbEgHf5FHGYgkiBXXCdR/zXjkh9p629nMFHqyxmqDq1fitDUOKk8Yzv1n4jpKdSc
0XiwvaVM+fDe8hrfeeKjhbtOZ7ygz4pMjjUVLjdOE7MKDSqNvo3WN1/DG3Q7a7c6eY74vLjaPz/r
FVfQbtZRkZeVvHzna/cXruLh7y0TUEzn/673uoXysFa+NdIMzusN5lzMifQWFq5HxYKmeu/20fVS
kLkAcOmuYUE+WOTcScTZKobwx/XDfjTg8QION3FPzEKJ4qhyPLQ7pzsUPpaRwhP2O31IzJwDMXJN
sgjS3ZW1mmjJ7HVHtkIOptFo26U2hmc2WZUky+tpaGXjaVgpu0fcUHr5Nx7bzju15KWcj1gYN38F
vioIuEq3T/0zRJC78KwwUdh9U7YfGcGlrquDKwwkJ6dgb7DoKnBP1WX3nC9aF0N9irgqiyWyuL8l
9KqptX2b3Gzve7PdXpQxfJJgkbuxbRGDRE7eistsurJB7zQA2DACnvipEv/IXEhLn6GoNttyGH4c
+Wl/H+R7AZR+h9BqHpy67SArR3Hsk2/ms5+/lxTZ0hD7enjP/Z1rzcfFLUnuHZvytJM4vVc1FOYY
5wpepkaJ0ZdUMDbRlc2JKkr7tRCeZTcJFWAwrOME77uUXvtYBBz8H9lQfRyweocj9q0UOiMg33jw
pifczN60qRxxaS3x/uZ8CUql499D4hq5GnCX8/BFcTdjzTkR4rTatCQnQLCD36iHaSHUtlKBZzU0
jFnSYyGFI3N5rB7Lsbq8xv2ej11Zp6bW3iWUALBfkm4V20dQ0ntxME3uKoCu3tWxx/KbGBt3bHXS
6jHmF3muxAAPKkEzJwbZTdYkQN4Uiu6jOTB5YwZONUwgWY7axiCeYUzlDEsvLRD5q0KaGrMpP6Sb
QukGxU2sox8znOQc3LkD2FzBYb88C8o9YUMXAKMMoswCIP//dtZbk7Ca2hNZxBBBf0aIz6inizon
oMzZV169ejriaRwBjCtXAFRedZ/ElaR20ppGWBBDuyluFKJXElR+iWO7TO7X/L/otpfa6RtrqRyq
/7CAGnxOfiWC+cUEPQi1XWy2ZZqq6a9rgpZwJLartmgfysFxNWJdOyeRDcnx3T1HjIAqTX95jS/o
8Dh1KlHiTpPpVeBWpdLUGHdt3L3Au+HCNdhq8dP6ZDC/tNFLqXIVPsq/Rl8hoKeG21FtNAS1TQbO
MChEVNDsGuMUo1LRVGVlsUVtWNKNpCDyRdm9GcUsSUEUjv4HiYaX+4K2FrwRbQkdqqzHjDE524QC
R1YikfU4Wg5MGLQbvp/2wVFed2t4CwOwxuvqjJaSMh51IIkYnC2dSZ6mcO4UZIeNyZLdtK38ZEec
QLbx6nII39i2dM9VqCiyT0cWy6WQQ2nuPW4vkfqrOG+3h7WEi5fYy9DrF1XWfvArbtFGQ+2dbh2f
N2mp904BpHj59NAgLC+GaaHU4e7hlAhYcv4PeDHTCE5Ug0XxcoWL6h7TefouGDoow4h0OcZmTA4T
qqqtA4gau9OtXmsTPqyLgHYJAaMQU6MLzvh30+nBGSLNM2zJbPY5UDIXfGhwSlhrGZkCp07ayM4q
WHOyIIXZEx+vMQ3tFt/SqxWHxEvlTxLg0t80k+8g/Ew3MqQcP7UUl7WYAdPn22UOL5bCFCo8VcOZ
BghLXjXTcgYKO/suT8gMGKh/B1tSyETr0mL6hPIYwcPzFv8cji3CCLD+s/idolUtcgbpCGyAqN3N
a6jWcLeNp592jjeKH29pOmnQ/x9XTZjGRkD0p2XOM+Gjv5nhT7GwDzFq0I9KasWyiNFpeWdo4u8K
gpe6bj4QWX7Y+eOmgIO2Zh/T5E3K6jO/bgZvXUFlGSfpTv1S1t1YJuTXeE1GymQ7GpkugrKP7zNK
BVatlbyFP3C5MSTV3x6fDQGebNzG3lCMju8sIsmzwLNrFg5q6Zp0gUTSgw10ONaqdFkqbgaiezfV
pcuZxBDfOcQGOfMONk10SyvQ4OXFcaSA40fpPXB/fy12JUw+NQ5hbRkqtgzwdi2Bv551n+C5ay87
J4CFa+wsnOhJE8f8P0YoUDEhsH7/2ESQALWrvCgJLokXHZxfbWw0TVXntENiVfMu/97Kzh/Q7j0j
ire81esqscPbcozW+whKqzKtpPeAUwP4x+oBHtjrjUlqNnEJGhlWUofD9rjkSDZWQL88lVYTE5wg
FCEWv+mw8x4Q8yK9pCE/HDtEijJBmXNlAQqUtHZx/iPlPy2DzNikuCUh4IWt8k+O/ZgrEJ1FQvOU
IWlkTbbu0Hpe1xWBPY12lM4Ggrp8PCBCscvMUYmzRptbeCiNG3u3sFbZebkgtbJ4vuoSbOe+TpMC
1aK/Od0ml5VZyJs2i0Z7sRJJ2D+mgqUyWiAhmzdqEFb2W55AoJj7vec9laW1oC+8dWEVpV2ohlDX
nf5IeH0P08AEb/3NKZv/eAgYWRrnSow1IIJiSZj7BjoUcdvbJqvPNEoDzCT0TukVvd1vj+DBkyiY
8sv1wotS0cXV+tFHp/RcxNKBfarr+TpYk7linwSpqFct9pID7x8Q3QcAAtQr+psHmgyTHzlKHQ2n
6v2hZBm1DvnPX0ew4KCTxN5Dir15exSdIPOr1d+0brGv72An1JzMEO2SbRKZT5CKa/OwA6QBNarE
mI+k8o2cpvJKcNC9AuW91a/Wo7U02gyN8cpD57/HI9xTK8dvxd4yBF2gObjohjBCcZy81a26w2Ez
8idhfyKnOP173b22dQFCNvrPdBlRfj1qWknfVVjfv0SfJnzMzjmlTqoJDwcLkkte9pJfp79Jv1Xg
zfVs/hycw3Ei3zdZDAmBPV2u6Ak+DVKpmdw77sZGV99FdCAbUnbU50iZDJogd+QtYDMvVdOUuDHK
D3iNd47rud6pQ/GRS0CU+mfX0zAwrVxdZL2M5XWkLJcQoFitvHCxNH4idQaQZ7D5uTODdwckOgST
CHaMvUnIBQXGiLTWftejxgnHcST6w7eX3ReCC8TCymcOwPx7CD1alIazjXzfNnfcxqxO0k/kA7L3
kmZbFxOsNTWxEzZQwTVNzQNGFYfiQA8j+ttcotOjZLfeCN3Hdsqwn0n/AC+N6AIHMIr8c/+H/4AL
G0D8ABpgNpxBFmWP5e4Km60cMEao5r2ookYTewkIgmv3mj9NRPNVTUkO+2V3ZTUR2nYokl5NKzTT
iFNQpKD71W+igAOtwYEq30wxbZP/zc4lVgijWQ47ab7dClkVqXzag/pI8LrhblXM04q0eXfuyVJQ
LANwpQttXDWaIkmnfTbYky+kGraUgXeh3jWW1Zpq8tVNOgp15uW8R316rHJPgDMVC20wfDchvoXI
p1+9ybgjYXdh0nJ1HbRm3tUK0eKa77uENySJmAIqWoYowJFY4boibBiUPF+0Yw4KudXFtvky5sep
THmdBlI8J9WF8l7hhawbWt5Ya8AuRJqtzDgfXRzrpLjunOCvNDZ8SNlZLO54DaKcpkvFemLtKFQx
bfpW6kJfe+FPx49zJw5EPmeXTWwKzSSTsKj631BrFeN5BSDekWnoVwh0BfAXV7v6vv2apSVGLcg0
GwFV/Givr/mvZtcdq7D9c2TczG/QOwprLJOwOKjuxSBS5j541pclHWkpa92PtkUwCXIyZtoVFO4J
khXgEo1IvI+QDTSALj211eSGSzNspEFVQnCpss22wdwcyqL/T3pZ+smL3lyp4Xr4sf/pP073Ca4z
insTGbFacs8/qMjj30feNVsd/26pyd7acBJAuVQ3SnYSuarYOVegX8PE2/erGdmQOUNCgygPx2MV
WwMQy3w9mcfHx3oDrc7uRRXBE2q/jVkEfBhBJ/rP9O92DvQ3duIwUJ31WhCPKuvHmiD6GDZhA997
t4rjUbEbcVqYV8QafHdNmdf+Rb2Zsn2CKNSBQEz/OPq1hWXx7U6lwpx4oOl0I5ecEqWIXCiJDRH0
dqWXeX09tWlqIJaLST5DQZ5wqvERE6mafW1PqJgnnsd757b1JLm0kYmQfukhuBI6FeWpaNF+SH4x
rhvpohVK1RIT707woSvVBDRqYusXvAihn7jGtmklE0Va8TKwheC2ZMZfa2caxxh3ILkU1899DfSl
oaKDoHDhWLAdPgJYFpTK6PjU8Np2Sb4A8tNKQcmFq/bFjsSC5wgfyfJE9CoIuJkINgBMCd+GCT07
YzeNOjKoycO6AyboddLNgbEBXI288gAdxMsVZC88Ajzn108bAwYdfBq/CRXHWzmPmCM7tfbwszVI
EUOvsYNfdxQW+zvN1sm2S5Ke5MlQ0+78oQc8MqRrA5yBo6p8y0xfrGUrsCM+bUt7+en6OJeBEKTb
xeOovOf2aZP54ebwFMqWRfSbF8mZWC7QvGrjKiTDztXZh+ziLPQi5MVoTroyxA3FksGL8jfF80Pc
XhYpXr1U8KrxL8proIt6JX75WaTnoB2EqyESnsqAmkRoJa/nU1hFfdak4QubDtzW9Et4X+EylNf5
JrckgP3cpH7FzJdHBRii648SulqbVfMmYnlMT8mlvw5aIE28L0p0KaGe487VADB2rpgTvJt7U7D+
+UHIWl34Ma2GoiEKJ19v8seWsuCwuVWgMMadAzBFd2qpGM9jwTC1E5EnCOkwc+V2DGSY2ihemOdD
RFPyZpaURQmi7Ccyy3OHyK5aVR/LA+8wo2H0wLxQVvVcB9geYXvSe0foL60e339u2ZddRe67eAPl
Axooy7wnvDZyIcyBK8Oa5Yp1jqK/4eGKeRyhpcnajhe9s2JgySqFb5UcyxKyXyIxS+FFxmOhcJGk
hBHRsCVM44X/6/YyTB0riQwb81TNRgabndoOKL7p9xL+wlRAOqrqyJq2/Y0V8xt48tAlHn1R0dci
v+PxSAfcGP5hNLDPhZ88gR7F2S9F587QjFBb6u63aAt9znKqfyNHEGvgj8N8jGvmO+62mHBbvQ2G
3hbtmysr2Gg9XKUh8KPKosE8RMp+9TB5uT/bMmMU6PZV8ti/35Wob0Zt++5A0xpENepeT04mlql5
+PImUk5T53CYIHvNGoU8NYOwRdliouS+YlAE+7zBiyEJok6twkUPcflWyalwC+tesvR3Sk64bZ03
3aSZ9TLdwMiUe8PmIG6vIwvhNwZkYHzsnzt3HtKE1EZCRMta/kE0vFh783U0F1VFTW4dCqBQa8JS
jr98xeN5sD9AfjUeWxcm9GjFXMXr0DTbnBeFZFuULaFiNt0Qv6MkK/heN+WUb5497HKf6cYe4h2c
3W3LOGr/k9O/H+4afIsYGyMEojiIYr/NdNU57T27BYZMALfjAa9HCM2jhYs3OjT5tcqbkIPZk65P
WPVOFSkABOX4nMwXGFYdKf9NNbgpY7EC+k+GZZpvzWl+XF7DCiPSYIhxFKM0CokGnrBY04hG/t6r
kAUxyCnAfTJhzOBO7/0k7HmnHvcs0LX/JdydQ8WukBNMMWKAdJsxXHABp+gZlU2YShhXHleferbg
ZnwFCO7tu6AwkJ5COKVlJkd689ZMNQ+0ft/hfKYcDVwpJxwEJHg6G/tpoMsFcjAVpSkeaKdbJTch
McYfgmLsK1Uolo0Y/s5TT13B20SgYLHwaPOs1aI9VMIkQ9hpuxVnxIZaH0Ua0j5Ch3w0EBITE61S
EAgOpxmz99oNyjwXsqKJ4uUw/9XKJjwySzC7PTIZWid2qyXSFatMxW7S47Z6HaW1l8OIQLHoReYA
HguhT3qqw3tEPgt8AlhbNR5YakVeMdPxdUrzpq03Sf1WQE9BiLMyZOO4UqujStYyKdfegJyV2WfL
vS+xOpIHFEnKa/cwBQBCrZSynQD4U21cgSUJ6HvJW7i9zkf8x4Ff2wYn0JcD6e8wmfHduE9yB0IX
W0D88grsvdQeqghzTj2+XyyurfasyOq/lhr0cExLmpbwzRrUnJhlShXFrpBRVv7r0NRrzlCYnETQ
tMAQeg8+tF00JrniP8LQ2ByIiZfCK28zkpG9zMWsBRpA2pLN2//F7Q7N1PbwMFIQk9S0LPIzWj+A
ldMxrhw2nprHzy1p+EOrc+gz2KBhPnHLzMtqQccr5pJmXh4Tx+Dtzvwfkpn5jqwVJxFD2X8poUDU
iixZ3pSbIdQamGHgUKMVD5HLzI7XrS2gSBqrVMAP+jB3bvn1LZMq1tBHUzmL7m1sFl+tbNM0e48y
NFYvyToKU5A5LWvDuU4Zpxa8/PX2ZJfHb38NcGp4TILCmaffgw5DFEIYZWkTzIXbDs6/cSqeU4sU
9whX+HsCf/jnvTkH0P2M43zAbw4jJAHrq8XU23vrlSrg4j96shhAxqpPEerFieMws7WatdObDQTc
IuVHf4/yxkOhXtKe+loVkUEbplS3h/qM74/+A7jpiXkdVRl3dxcl9VZe5xggUzJUTvJjMqumKeEF
HnopC6LK4dk9If3S2GQ7x/8IMLPXzdlK6mMTfCg7Z42R89ya+hJAavE33/W4TzILfHmfLaplnzwM
20qtz4lLtLpLpTDbikqlbH5356n9OPs19nE4ZBbbhJhbm1kZaB/irBLgaBl+iYFcd38OhFZB8c4F
Bu8mjC9tcI3ycMHjL7LRJWKuavwPWK1u48ueMN/n325nFtbxDlg4B2YMhlUzqQyMF0W9+uoPLv1s
Mvh4M8T19WCQvI0pC6V+8mrBgPyn5Sgtdl0R2JVIkdPj77Gl7oYAJ3h/4v922UzoshiHm1PUgL5Q
1uNd8T38R/4SwtEs0qOZRPT3TWSYYERqoaOqi4sBtElwF11siJ2zg1oQZdNcG7Un/X7o0rHi2Xft
36yK9VweIH7w1GOKCqOZzyj7qvKfX/U46hPP69aaUsPRV2Uih3I0MBHh+EfU1damhKqsHTN71yJ1
Xc+ul+fu0wFNF9RbhyNHZTCEzd+Jb110mLbk6heeGfxgMpIdYLBG7NSOs25RtTl5IU0VHJosZeCK
U3lvodfUDNPBSXO6Qd1+iNPMZOvOxjmmL2JWzz5Co28FOoliKpkOYPhYBrNnClSrzJv0gW3xNmnw
dbN8YOmmDu832nAvPEzxDlKDJKm9erFX+7O0VEI4ai/otPGaPb7nDc0WfLTjgVp76mskgXIpgIwY
ZBjD12BIgTrtMpIoAbGtbDyznEq0d/9vyz9z9XKWv/IbMseKlqEO3DZ0GNiqqL71XK614mAmH0c6
rSqkUzSYfA6mAP+UGjH9sO7EQCSLKUer890tDm6m6JGB/Nmhcb0Mo9O+Ndpf2GyORYF7jp3DD/Pg
nafWLEsLs4m4qsBHwBXGZaLAl533kvRN5ahKeIG04zHty/liqWG5AjfxM8RkwlYIhuJOVc6tugGl
zo6dEmvc4v0wEN/+jM6plEUPFbMd52MYoSQHkLhnNVwRid9sKpElbBe8VjAQ0efKRwwzdkVyQe2d
yZV5LDc1ptzo8F/WHFHnP5y4lCq5zpIo7lUdyPGgmmB8jD3uBS0xrCMifSKeuSQvRor3t6zCBYmz
Wid7LcDmv06peE8tsH2LCIQi6xT13mehmdIXDHQM0iU+r7qylFQxQotXYV6W6ELQqQiA6Ly7i1lo
z7HcNIjqD15ygD56GydqC7yb0BGosUYFYPAbpg2vReGeq1dEupkfB/dZQv/NhNwvRk7C+Zficlgl
g5kIAXHOoJAZgRegOH+wNiwybh8XywMMaazuXXLTTGGS9tJPYGTXM2JCVsZ1xkOvYQqGvbG0e+Ar
rQJOJtV/CbHZpYRyn3T+uRj4U7dOpX8dNGDjiwn9zWNQZ355iWtEJ5dyWqP7xcPsyvCAErRIkA8h
XaIZ7PovsIkf8bmulgXff+O3kUrrK7aQFzFypB8ha0I2hQ/qgIkmaE0xZQqEsKg3QDVtw3vfnyD/
iLwZ0IiMMXYkWzwE7H7irnq2TIfquawS9N/ORqkwP5ZxKpd2BnsNihNvDIeVrr8vqb1Exj8VTzc+
oNtLnBWipkGtnAlFIfnrS4kSvhuPmRqxT9XPxuC9zs/lTislpgj5ylTQdCIkIjkm15aTTDibSig+
7TSgysTSez+XjPS2pYxRI8lHBpA3Kxlg/yaNBxKvIN/2J1WFkprBpSniwI0oszS+lr1PEBcPdL5R
TzCwppmbROCL9YN5etR6ifhEbSaWcQ8EdYDe7RY/Bqgx0U7g1MPhSkBWrnTHvBW2AIZml5YjC/Ed
Thdx64R2dYCDxJlszBqmjvCJ92MnhSPDTVdvV3+3W/Eg5WYXxQbOivvhKzXEUG6KAofKzRZaw7Mw
ja6GO3x5L/sfTT1Fh1jHbAHgVLOd9J7IdoRlNJx2B0JxJ+5NWLtnViXdHAZ9CsG9/BbMtTSpp8Z8
9ma71H8xBaz5VR/LjcrOntAsdyLnlE0WYIgY1+6vEDlxUNauFVefcy4JaSMLVIP4t0hSEs70xenw
aWjTvGhlhdJlJaOBOS/lar17dX5F1uyrbzeIsTmHjJMxsQhXWifF3SldaeesiLou9h5A0khumySP
YnxQD1mGoWvEkK1P1ap7V8D9Uq/5c4benrLpeVTaNuwN5gCo+8+Hw9mPxA/defSz42/wxhSNYAQX
ze5DYsGWNEA7K0FJE78KzD533zUULM4GJ+cqQHlgWPPF8ZVjZhGINt2+INqQE/9O0UH7kfvCM5Rb
H4r3OU1acfmJ595sbJMiRqHGno722NAEwmNqHe4kTMm9xTFyFZSO6OJxQUPTcBhfx0PbO5boQ+0Q
pfx1TEf2wgcptdlk6SsikgfBeS+31bnJc5Fh2LmuIl+JdRYzKlETqyhbB3AKewmCD3nQvAVmwgu2
z0Pc5YkXv8pAYG5g8B95FfxJQuiphAMx6kbR3vzq9hrlj136+pfk7eTYSS3JfrfochIsx9BB5LQ2
OxFjs6zhDG9hsmpiuGw0LpZ/N9YbhdNij7QwnyqZ1NiVvvdT+hohkUU84gJ+BjhkJ9zVZ4FiKKCl
bIZvxQ2qu6njo5YIJfJASLRtv7pFwUGzFfFyw2fRJU8ZQaBzO3Fnan0Iq2n+gTC8SVOrzwIC9tWN
1+1bs5pwIJ5G/hD4cvp/Y01x9jNUjcHir0AgTJ2o2jsJmzrkNK4l+eehCV6JGP/CW+i2dAHm3A7r
+RYCTw/qesNquB15q5XPE7Xy/rsSAr1vX8eLCG02Ubr7V9dAlwo4sY7Ijvjp55WK2gTRDVxNA7PZ
JpTasYIgqR1vLHZLG2Q3TUj51DE0oYeRDM7TP6c2yLcy26mr8KIO26UA41B+/mFOJ3eYewEMPnJk
juHb59cLkmELO4xRSs9Pqv9PUKJtb0nu2D3pV6g+sWpNDw4ZcYmBbNSIZooCbltCgjzRZn+yV4kj
+J749G9zXatw/IcBqNyClcWMOmyxMDxw8GVztNkMkiNiFrfzCcO1zlQEkeVtMDXWUOzUY6ywNCSR
IDuzfnEyQ1XeEuoNp7Ev4IfRTdR7EQUJTnFZ/5XhtjPwEI0ow8kohBZdnlp6te6u2V2cRFc34QIb
kWcAtFxQnjeImUbINxm8Dg6xue2hs6zU76Qil8J0QKN0/QWz29tj+VfUXgaU9+iVJp6tV/HYdGXd
CkPDf0ypmy8YWGdn0k4UMI71Iyk6mvBhMB2uZwjfssX9/8bQLMsKdY8stVESkgxEsuYGiW7F67G2
7RyPstfnUvi31i6Utz9Y3we3IjM9yw6+/Mta0hWV4mSAgcRtzqQ9tVloadUCZ3LKAwArsLZUaF3R
Hm3PjrF8xWAWaEPKzgntV77WOkszzXiEN8k2X9QAQo0hKvhqja3/r0BlyXuKD2DfLenoCQb05hvu
aAs78f83NuA8lP8KFYk5L3ztyRBOqALe4p7LPmueIwsggVQ52W1kzpcTPw2TyhFsTxyeWqCrRYTE
gbgjboy6CZo4pnm3i3CB6LiiCET97SkIYzhSOrjrDo0HAqRFHRLf0i5KwxrktJMQdYqqlvH9QqNR
82DMhpdyD/mEJIdGCDH51eWFC6VvSeALZleQhLm5Q+1RiGVSgFOKIjdJ4IHsEFwmfpr2Z+/4vF3+
b/PiLet/B3Nh45CbsULMJ2cCQV55tXSWvu/t4NPC7vLrbM9t+UybeWj9OKVPD850iywfKZGifQ8+
nZ6/lu389cUFk+jmL/K6tTMYm3Q509oKVa1sWCKIDlHudatzouqzWqscNENlcrFm01SA0IhO63cp
oOGeyMOpzgB2RgsHTB53MCFVDCChK4C5ESKR+LqeAhZtkjv8zo0hkMfMDHC7451ZGzLzjy4dgN79
tpfa8cgs66mxJqxM8x78Ojj7ZzD8ej9toxvfie1Y8ihalGCb5RgYfg/BRhuP9UxcvbTtMQsV4Js0
C35ua67xRzTgWFpwhgj4DMkhE9kJzeOxNNPfUcyyknuinWpW819GqdmiVpMJ7NsU5hDBSA+TzHxv
5NrJGjyOOfBpFUfPxMUBUUj99iNrYxw+3KXT9cTG73KiYkfWQV1FqLqXFrFXxodIor9rkRXXXstP
6BAOghjP0MIhThWglsu/ST4MsBFIAQeqrMAOJgkb3H06BFjCoX4PRY43YWs1DKl9kDSzASbFu7/8
jzC3OiZ7kHcBDurSsu0Vkk0Pxf11bkBy3eJzt7R19UyeuTZfRPiMdBIbibYcHl11+1qlqh8U4TCH
XbrfZlNapcoA7ylEfZz6r4p5je6RKpmEBn01gNrM2jz3QjrgVqMqX79TxB6lTf2QFGmKzgbmCzUm
58kipWaBqHbd1DDO7nkcnFlwd+i9FryHp4Gr9mvwidqc3MTg6wt5DcHpaKeJZ8g6Gqk2lt+eHMkm
Eng9CFMMHQKIAMVnp6nsDliiQY0y7be4CwxJGXT32GPAhwp24kqbYvT1/F8FX5xerjyUoOV1MR8Y
EqsmhaleChLyBA+tieM3TH4mbjDrHx73E7aEqkhjF+lyPZBYLzEdyHX21xsEXir+6xtSpJhydMEH
sjnEpkFxS8jrguJecTfCfoswKt1YIjN0tL9NmdK4FiM0YSPPj4q3B49oskK3hUMtrz8uWNL6gMnJ
JQWH03s8q62PnZVpdHnl9JBlYx00lYIcP1Uw/nprw6n1DnUnDZqmAD70W9DggMyDHnS6ZN1bV/ot
7MY+F0WY9WRKVV/cbFiHxxaAL6le6ti61tXsSfxbIwc8GvjoAzQv1IWtmhlBoh3LX2Rl7rRm4MbW
KtigIRZCZAvNwPe/LvW0P2u1pKNos82yzq2NSfkeIzYiXVpaBwR4zA8rbNLIAwDa7/MF5o5tbHKs
lyzGo+CqJan7cYTNQKNmoMVlcVfPoDGRJIeAXAifHSl1Rcm25QZJ3bXNithBnCuD/77VY45qJroy
wk2smYO/ZNPJhsBts1GSKWCO9DeJLiLZ+4zjc/53DFyJP3JYyeVpmbq4gTr4TdLy55wf21rI6dci
nCPu6LRy12PgoYKfZ3JrtiYdlBE3K4Rm9JNbed9G8sbhw6O3ZX3KU3HDua6vqVNylQBF0G77S07+
dnms1NZoORABEPliL7bY4CDtefqZN5EBLY+0nVME07MAsB3KdK9XM0uA0Q7CgMtD37URmjapinME
88JOeuVY4ozqFyFe5wHr6ZMN5A5wMxzlhFtoHXICpjr2fJWpR6N5Zg+aiqlSKO1E36YpR85kI326
/Tow0PgwP2bq79RebVbI6SZiUGHrF0XJC84aINYUM0ADtPXkU9Ot/jm58yX98KMCkkKQhjMKgvnG
MHl2TEKHRpo61EwY4EPQmVsffsWYbmfOXe7sx2z2dpls3tw8iIUPhA9EIL1s6HT6s0+/HWWxlTQQ
psOIYr6HyiM2oS76twhVrxPaou2oZEgqJIgFSkjgBnR4csC1V++M3Rj7KfV6Qw5IW5F7UGeE1i88
t0824sy+Y5dHdXobItXSG+K534HkVqY66swe7itrnhT81+wYFM37zTYXfs7Pe2C8HWYy54VTdF3r
70rCTtvRDfBmXsnoUdP7p7769R0ns0FWM1wEIyo0YKFPyE7M/32SDiBTHvq00yUioKG9rcnaiHX9
/TqdGHyfRE0KOuj84EZLlGBi9vwY2Y/cojpdcsluobeQQGGRjIZ7YXBGFR9rQD/na/cRHC10Gf5j
72G4BtK6uEEYkA+uuXMk249WWkR1eFL/saDBM/kYIOTgYVtY4tfYJ9gOGz4qZ3qxJMYs0qy6IJWz
4UfVhRuA0n/Im0Pb86Ke6diwZvy4rhWhIE1CxB702B37h2bUPeuZtKAB9Ai/iSO2k63lGmL38vwU
5B+k2SRUDLWzPZ30qnAq2QgrwJYfcEaLSoj65rNM/WHHtovHeWEWfEWuIgQGqiZBMnyiIfyoe/jJ
Pw+iKRvLAcIxYC/aa2YQQ7Qq9b6fBnixK9TaThz32BO08L1Lkcakx23EsVB/tunFb1dCR2nAdQa1
Ka07p3jrez1A/vJ8wUpqCmme4k5IAhEG+a3qpodZRweL+5ktV5iLdy0WaIAPKZjPndfuL20Macd/
kSDWUZTTYCE4xDW86+NJMhVs+HqnfsiL5JqDmrHvswV6ensE04ZUEZ5Mt0wgElqXRDzJeKwS1uAm
PcrlzObKSKjudsE2rxi0J6GcGxJrK2xaGvdHC9kNTPUAg+odLwu0d4zJAWy98Z5AwjqTWVU32u7n
NH+0A7OLx8tQf/bBQKE7OYu4xCurni8Wq5Lo92OYjKNQFIMhWsNlE//TMQzFDIUEerexT6fjcjji
kG0hmI/gHA/Yloa4+YiqfzeoeX090RdryIN4DAKHt9zEF1I7QrwG7sGcxx8kjDWnTSkmdHuY8NPK
71yBwHclG41nVAu71s5q/wceYCxpfuWHJxpEV9bXkbubxEVJ9JH3/i19So0ktnZ3hdr7RjHzache
bqYI2EO04p4QwP7D/2hV5urGi7XlR5LXOZWjFHPjYC0Pyb1T3+QUPWNBgHb2UlT3hKcd+Zx+fY06
3k648lCmOK+x4YxXvVxrq1hlb3BL0ygbnDWG3uJUj9K+DlMsA1KjWWIhGNGszPL4oQrbK3oaob5S
k+Eq7HHxfPQCP3WbxewIHBV7zYTjRGup9Nrr3uhHJlDJ0QX45/i/gknrnaBd8unCRIRJy/tKn2xL
ndCHr5Ml0b5Cm8ob231qXkXfa1Trh1GWG7++l9YXA+NMTYNWNq9Vxik+aNRfG+7KCJ5MNNKqE7jz
ONwkMpNU7vk87skOA8CWQJUeCXPkBYdJ5Uye2H6bZeQ206uTa8Q5fe8JdeNrq5JIEVwIU36VdoJa
ukUWC7QL4dlb4YcYRpjCDupafToDH5YIPz6VQC+Y9ftDgKSBFuOs61qfUmOk7Y7ODmdetHy/cG5+
nmDT7X46jSc/0Xmiyoz0qtFpmxXbKQHF8DG0KmSXZRlnDKN0vBL5DMB4jMatf+Ekv7saaO1pHzNE
P04vDGiJ6feqSRfrGQz/kwPeYlQornB6epx6Z45TYHSV/qhJ8LW+DQnbfC5Y5o+YErfsQrKDaOCc
tRnQSgIqEcTN2kl0Foy2XFWmJJhfa2EVPE5FMhh5Avw/cr0FwWX+pfCvNdgjVx2VFcvQBqXheh+6
CKXfE8YXE8lR5mAinMJras192dmx2hTjUwjr+TjPG/HeJYEdlDWObq/+Z14nWeGtMYaXlMqgkILn
sc5yl3sePMJM5Z+RrIOARuhbm3dWVTSRSirXeIWVuhxSHsK3sFbLDf/6t2ZLhvqtSxRD7F6N1FKC
jdOItx1Im17+isB4IS6XLVxjXAgoqZUzgA8OAksjYZjzaBsuxDMahH1sgPOicXXjiecAsLhtOv/V
CxDTEKYtMPoaozfv9x/XG+k3hLKDmSo1api/GdTkhquGBeveuqDartJWKlx9ds4fWcymhpWb0W/M
p8A3hzg2ZVqFHGB9EUyj9meHIUZhoiUI8BdwSrFo2E+po3NH73SadtnaXohcpdjlwle0pIf7J8s7
no8gndE2f/JOuX0zOc7m5erqMpe2oXnzSaiqib6g/Wl+z8UXbuhwlcJ8vLsHid1aIAaTSPRFzNQz
AYkY00gePfjOakpYJ+N0kD+7a8kaQfFRwEGYoofEla1SkgnXq6HHolFFBibNe4309NRraIJ2WDPH
U9246EAGuQLC6T13VC/EbasAO3L6Ccai3uUlPOcHwUbYXmp2tcvERHx4CBvgcGOSeAQbxOXGPwFH
xek71bQOf8Ogwzacn3/MRtZkb9YZspdv8pg6j2WJ4+v8wxPXlNOrqLudKa4GTupl8jxUQ9YHMbca
RG86BRPD3qjxOjcLhF8gjTx+wV32ncL2lJawawSv7WwGx50cTlOZd2aEdXOR9jgBmAxPY3p+vvYL
EJwexPAQfyw5JAPFUp7vFgyRf1Qg0CV0c2DUaw+Ku8kMcp5Npu7nABeqGRi9ad1kxppgike7NWC7
Lk8UT9npfnVpG3lMWr0glx5flWp3pmvfM5IYOItB45OKMndMA7voi/T26dvmwkRpDIv6pz8NSmgd
UletNFRKMWFkNu02SRN0vj0lT847MobxM+nX7Wb2ZQKP26ehDTPOaWhw1JZqhHeDIk1gIRsXr4e/
1BP54UkhUDWlSML/L6KUbQNk6r6fXyjFKCU30WYbBdJYiweK+zKf3kvlpLu0WDG0yGb7tLGBf87X
wV3JvRmEq/8k6uugVGBpNXN+AZrRdMSWudqe1U77YF72UDmVnp8JV2nMqlm9aSMuSYQwaA5STxWi
VS4Um7XHbwTT9bI/GLcFBrAEZAPUcL7FvuB80hzba2RzCDJnxzH6jixLRENahJB0hMtZPlbQ9lEZ
ZMCuULzboDoNS79NeSkihTp+ibZ7ODQCKxmjlXhbn2wfDnnGm63kUNlihPthCzP+qEGtnngkW+l0
6iDo1bmxGEtpZwgkGyVr74Oq76zhD/Dal5Tpdps//N5JFq/HLdG3INkUgeHpTyzgEoG8JD7JkbpJ
sLQ0wd8r25AUsDwUnp1SCwwmiRYWPgwMifMQWwmDKlBcA1/nGl21LPKX57KJPRoPzqrJ37uRs3ur
Ew46pDw4uHNu3dS9ZI5ACiAMBN0V4fb412jkdp312h6b6HzHSCrKCNTxK40+Jl2KQov2NOxk1MCo
rHwJrRsa/58qjatXhhMNpgEDiFX0bMBVgJA4Anf7HvRzDWezBanJ8/eXA0IhBh5ihNyN0zG8grn7
3QCIy4SHv4l4pNUnmyUytkEORIjV8GQA92hdcATWXOLjIBh6DdYP89dyXCT8xdiZKiXDD7pDpkYG
cd5Tw8RwU3aZICl/eew2gKdY8kIW86RXLAjgF4PxdeVANHYXz6nNxbr2ZFrIL9bdhxM0Dcp4kUlW
vbQZ+9PoGTwJeG15jtaPIadXh6Hpv5z/vSGfIz0eFqZLt4Q3wz5MmFcOoMXLHbva1DUAbjc04teL
Dh942joMZySSkJm7UOMZN8AFL5OHdqjLk4onT6SHE/4sZRFdqpbtaKooU98mfBEcY1GxGXBlWlvI
eAldmi50nSta6qfCo8BJdZPPoontw+AO5o008npNA7YmOBfOe5ed59LgONQyaM9quhuWMx6fKul5
v1Pf3SAQ3Q2eKATLlt2Ee3oOtY/lS8iB6q8lLTWBt5RxTx3OGcXkbWOrisnvb1c+x7jO3Si/DESH
1yLUbswB7aKmMM0R9SV9dvt+Cr9bdVv2FdewJHPw0xGavEd5+cWH0wbz0t6Z0UVeEIbKsh5MP4K/
fMrPJrGV4dE9miY5smEifGfy/MdXW+DPVahVrjmJkmqyLTF8BHjaIRyzaW44kic+r4PHq3WOJ8PQ
GI/W9VXTijcaw5OzU5MDcVAkH7FLkX1C5znbW+LlQap24TOPkIITJTSwVhZaZvYrmptUqB/ESd8z
2/dYReLMwXwwOMCYRXRJOz8Q9EBsSwkuQYp8k4ZFsP1aI5q5JyZ4DHzJ4bKVukeD43EM36uClnDG
upVgcaPYmkT3ldB5+3N6wvjF6l0OXYbLRMN42qQp7Cy7VQkesfzAeVYo7Sk+7HBOmDHre7h+dKuB
hGa7i8dppC4KrpiLyM4nIybkUn5EesoGhnGhCqQG9pUnF+ZUMRWqCeI3rv3iVHfGt5m2GY5zgfz0
LWVnZn7peXCzsseuD1TuCgVlFte+Yfc7FV4hJc3fHD9XlyMeCPKywuHUSpIJSrQSfdiWsT1xAOvs
HG9CuXbf2dzfYfIlChhj8utTLx/XnvE83WS+EMlJrP/rqEXeME2xQpjnup+oc3DhAhz8YC40xMSB
1Gx9GCRBUnOdAPF7rLrD9T6aR7SYZRe2DBPeNKMyqdM+Rj8vL2vcq4SMITY+nI6P/CuPZSKCapUE
eic4/UdGGS4bQYz/u0xv+e/PiYpXpxUIW+dIDFAdPNcnYqzFbKCACxiTywMehSyfXS3fy6+N4VIs
TTjEpPJ/0AXozg5TqDySJINQHuUBVjwrM//QPvrPF/nnd50jFIjXcIgSihPC/F8n7ft5d+q07Ggp
+vsiKlU9T6qvPEsedPxd+0fNYai2InEgGQiRDoyaKkJnRlm3H9cjHaR0kznzRG3hcW/zTqa8TA3p
8RM09+vRP7gb4TF8Y3mhKKI6AFqEmZ6yJM+2pDLv9vlYVBhU6LF58l+ovlvikHEILRD/N/cmSGFB
XnY1BR2LsbCYBxife/6GarAPyP50Xp/nTLIVZQ3Y0c/d/Db/ZQT9We4yCFEscsC+WzmaPVycAPyI
bcWAvaobZyyapMW1Xvwe2dLvy5keU6s11BhyJEW+LSHK6woRqxGud4XFL/F0qacIjwL/ieNlOc8u
izhEQ2VmfeR7kmta9F7Go8g+MvQB6UYhfKTT2Rja5aRvdr15lO2OKXDZ9h585mPYffSXtw5IedOT
LbbBARo7kKM00t0h1cdOPhDTJJhqw0YJvUV7yqUp9hu557mtZDNDooBjV1v1U3w/cXCoZ+FUWTXk
aGdNrBFrXZFBZsz5WPcfTesiQ16g16RwVdH6LT8xC3UaB2cQtUI1ZBVJcpRyze2jXcGjAmfX5qTO
O2YMge9Cyy0QELhugMLKaQXsT/vln6/OwOUpOSuZ4ulBVVsYN3ziWjjobEhDZk2c6cB6Q2LAc2cW
rFnlTXe4JviO0INJrrQKE31flk+NDxXC0kfnJKnX6/nZcc4mI3+hGIRPi9yJSqyTdcpRtFtiJU12
+2WyLDD7HHTU3+fr/C5BsX07S4L4EMizKZdjcMGv+mPuH2FUDraLe5HnUXjmBG6aoyxMe05XNwBm
xg7y54CszcPGTl3k7uMH0mKaS1shT8kFcMO+thleAefnUFyvNobnc90LFokLAl5Uw1SygWIjFn9n
CiH+0Ntto33rgEubj177tsb908J1I3J626d29M78UV9mjMG5lqOcs4XLETTMEpvjT14Zke6kkv8D
QG4nzZXjIB27OiuU7cSAPFwxhXlra0qjaHPmbHW8c6jn9JjoJ0Ty1cAS8yjOEhge5dsOf/sQIY5V
HDlrfWBSxZx2kWPPNZq+97iXMhlx/OGiQTrqoUnYfyYvHE8NlY1YgmuYabV4lC5erdkyQ62bWLiH
lXTtwiq15DlNVE+V9wE9bnE5LR7swzfw5Y/y+o6Pt88h6Az61PEUEEdTkarcu9sd+cxA9wPE2gc7
Pl7X5z84ojqZD94VrJPElsXZWGoZIYIGb3I/f3sfd1B3eu36afnA63B3Ab4j/jFqzSt91DyDpZ3R
tt6YN8mZGqmVotxxZFGptNuIq81sOH1tVxo+bRec1+r6XYuLFousV/R1WOvW8GypYqqST1rOnLOy
wPqa22kOqpRFAvGfVaNee64BVxyyAicd/KfHXwSwzzNOK8ee7dTvxVI3GdJ5Cx1qj5FQvNnfiqNw
cJ8duYEXkgrxzTe1f7dCe2cf+x+I0jaZ2KwBe3zffK5UMV1ddkseYMx7/Ko6xg7kQzNr+8R1hq3c
CXL6KlciYLuzmJJBVqJ8lrhZExPyVY5/4bO9V0cNuXxgcSWPkoSiVmRCkSB4pIs4mx7RKr/MHFuh
p8SSVrod8IEWlJjcfyyDfhnkfHzOFIbP7i3y4Apm8vrAxujrLBEtzo7cj09fTrXfpdKeqJ0wXb0K
gzvX/I6KMcer0htIjWhwM8BZdtxtWM/UAL6HjVF5X0403/rKYh9lNZZnv3UiZ6/SzRDmybfu2FVl
V//+P14f/OnV2PmEVTd+BUQ+Dfy4dFGyBnoLsQ8Ad0pvvcKy3yMd9g97Y8kxq4ftPnHta5Q6ybWY
4HKA5kCTywffupaMr8GOiJY+54KdxuQEfddp5jpXVkhWyyNlo1N9cLvBELp4cDKNLkG+DSEV10no
DcbtPt9kAgKNt3ZY1fxNJBO5/KnAjgtBHJpzBhahtC1W/0DUuOMRlYlcUYIJ05ePpBcXY0zW42BC
oo4Reah5rUT+laflYDlIoMK+2Q/nZoTViDU7ciZ0a9G4Nn05nBp+5BEYwhYkL9VTz6jHYwY7lUji
VD9O+lfVhpEFJj0Znri0GvGTgUA0bpN0ZhVQ29e3TsGJ5LmepYhVX7rbEbd1lWHYptLD6ol+DuJD
CSglmEBa2fhR1zAJCEhk8DEXYOhNzvzEgmBFQ4+MRBIN4GWAsppJj7igZ9VeJdfRNaeadlgc8zNr
lIrDZJg80siyEZZYqkvh6sCRBy/fXRr6R0nXtLoQRpKXzdATqjIKq3BeKR3hFYmcUYqotx22Kb8D
GjC2tHGhbZQmKUKfX/7iOEEwxVNPpqiDbWEQTZIWNxL1R3j0aXbfZjVSFfzX+JFTB328MEmRSQpn
eMz08eXfuZceMgPcAoFd2YpjriYk3xtXKW8OCfFTujO9HtaCTkziQ6mNLywgQWJiTe4SpncRGk/d
LBUmk0MZnyakGDc2oQinU8RWtS5x2wmfj9qGsZJnR4u2yfESWGVXdUyhLwwV8W0+Q3RDpMh55lol
exdLAPufqzArV9ebappjngFWiwDeUZjZ8kYwDx0ziKbjSvmqWQ2k1tgsviueKEw2n5mp5KLt1sCw
wPJsHxwMH7T6A2viVkWD1EZLAEdSt7ZxpwlrmoknacfcX+xSqy/PF2gp9Me5v1psVvYNAA0SkWaI
Avuf7u9Hp+h+LZfi6SehaEhDshJiTY6EldhGxW4jWWUNrtqNoqy9gqBngmW/OiJOgfDGlyQ/Q7PF
GAK33lzaWcmUXRoXAR5rEXYImyiZ/DJ8DRE0ZclGpZoUaxuZTsxuRxG2YhnrN2IqSlKoEV+HHQo3
UF1IS3mON2+4EJlYzfkn38vv7KwyMeH86qCeR6nn15FxfR2VS0AIkA1c1ghReNE9z8DcMZMZzfG9
cITUL4QOH18fq3d7u80N0q/farda0AgB9NdbJPBcwhuNx4N40kQFsZq+E9UiGQNqPMM7XQeu0YIg
kGcBn0zkK6jZ320Lk8xfnsWVHztUeW2jFeZaPTx640rzPHCDxi8Ta3oQNF9DyHHxEymrQycfzJgB
LWl9ejO5CUwmtc5HCoQRUV3x2HoyPE2NrwO4DPci67hOMaZ5KtiiOC3yvFo6h3ZB7GnvAJrnHncX
oO/prLNGw2A/fotx/FrwzBKZFuOX6tB9gCP6yNPvAsnvjfEBp1+/L7gbSe2ts187+OmumRyH5QHi
sDRQvXW3ZLBqRlWuvcSyht8eolKY3Bq8CQ96sdh0/p0vLnG8b6oGekfyCxtQBxd7yoBmer1WxeFM
w6r6Rt+fUne9EIyXggk7X6ou7ZlTVGm7e2VicLUa03NnmZSEl3D9LJhvthnNFm/RKrz7R0e9U6f6
cxaCMluFVgcO51JTqMyChk9rn5g+p3VFJd/fegptqmYbRHGfcnPHsPLzJX2eT8+RSJPfH1DYJaFd
tiy5/ZWuA46mrE86uheXOK/Ai3RM8dXyhJDpAXYpRtTJBkGCItJoQvH6AAiii5Y9uaPszuK84HsR
t/NzR2KI91VfUmezG3D9byP55tJ+kLhfakEJG92jptXFsw641eNUvfhtx+SV46rBiGsM0853YdA6
oqAF/1+HaKoJC9WFAu0z6V4l3eheSlRT79AQsl5Ls6hu6u77eUu6Wh9EC3bNd6t6idz50Y5uB96s
NHGKQ/aBf8/Wsb7n+/0X0CDedN5l4wspDd09xvPkvoKMeqNJc3L1HZhl2EtOJmqqgXD/gAEmfYjp
xhI1g6ilDCSdYD8ou+VDsNvmSmi8ypw160XDc9Ia4/2UlGNcLgV8mYkZe6c+wZTwRr1ZMNemrf+j
cgV4vxN+AN2L2rwyZR411lnzyGD2zWCS57/oFo+4Az+oGMsRcqp79rbfxf8xVHn/i17FUFH4nCyM
9CHGwLucD8A2n9+zxfFk2NuTdbQAuBQFYHC7NwaHQbhmsL3xWHF9V/xEbM7Dyx4IK6JN62JwxEz1
eSWv226trNsBGOW+CdScjvj65nIBa1CwyM/7KensMBiHR96IVPrwh+qKKThTo7ymbo1ha0lyd+FY
vvfdKL6mf8NYgnaj9JhDrkOh5dy9+wSzDRLfakOzbMz+CmM+Cdzasejr3DDt5b2RJJk/j1DFmjsZ
PtRG+KCyK02/YpcXJwRD0yu0xPIhowu0X3otjrHZLT8mYJUArOihka1Y6pLMNByJQiFMVd4RCyYI
FS/SNULp6oFWFpRp3nZrLe5A5Bhsni/aisy4Ozd7n6uEYziOGswdhKvFUVfR4lpl8wFXnN4PMsxY
+X51D37DgASm1+yQc43IZR0prJ94qzH6J6/4O7eN8K08JsgmNMaUX9yUvXON40OePLlfwM8pNtXe
9aLMLzqaIl9mDLaA0d87pBx9P/hRRo0NxWta0iv9GaRQ06U0OamWskbW/O10NNCZpyKpc6lNSL2k
vRYa4ixYlYzqJzbCl/ctnIYwT0wGeWoQtm41zuYwY6qt8qccrCwvNExsX7I1pcwoIXVkJ2mBLOWL
POZ4g47YZYhkRe/4KlCPU3sOt6qdhjK72mx42czaV0p0PGFrcGKQMnfP0cIUYWzLyqU8kbfDpxfc
0Nh4GIszPj6U+OsIVEbp5c+PHRxqCuy5hM9Y0JhGZv2+LwDFDetrcUZleldiFY7GebT/faYM6opT
bAuGSRcyWMQX1dWMIx9k1lhoyllThihhQ216/H0sndcjdj3t/+iPqHVIPh1oNcjjvMX7uFU3hk7h
rkIJEhnQhNceoPzWbYKcg5ES+6h4ptQFyTis24qsNfGJ1OnBK4A8OuG3U/UxZVIoK4Wgl1SioDOD
1mM90XBkIL1xgDnYfM2/HPlI/NC70gQlgV1PLGmLR53Ta/ZtbCVFcixFT4bD4StUJomUo45gzUN1
X+wPgPYtya/AfWcCLfKWncluAKUpELfdqgmXrB1lWr/roYRHE4JUqCPlBYPXoTqIerazD1d92+w1
m+cZEdxThMj4OK+gjsgucohJ9046Yf8c1302YyKr/uaLVf5jMAcg8QbuTgMugH2Dh6rPJCoiM0Pn
GBS5wgvJqCAMTkXt5oXLFGmLniWOTPKw2+edp2F3L+vtmVIyE/GcsNIutkfNqVvlRFYqpQFPnOdo
mBolN2CS7oU7gQQS83xKij3muiRDy7XBX7hVCkkUuhcuDvuuu1auSYFscUhtHsEaSq08FIyKH91n
TigytgSsDF5/1wfypZCmrh1yh8018R1OhVVytcwIvWzrrE2+Guv+fTPt7O6+WrsVxmAByLMpW2zQ
NSPjwym88FQYJH2Re20Oo3zaT54Q/EoGuNok0dGGwsmLXbrWSHWeRISQdrY8QFFHP7aH6Gcw25Tw
Uf9uZpXUd83oQw4ViuwRO2gmVicX0nGZu0eJRDSo5fDyKM5XbjzEeXu2J0WNg1oUNVNypea6DUxx
gJP9sKTfcQNvMsNYNyCDTTvComBgCuhmRMjr2kLLWqXnSFrCjGDCcMN4WrR8v57rgUqU5y2AMEeE
ULrbC2Q73bzN7NE2ablJQ129Ct+zoejZon3u8RMMJn2LgxDjbGlIRhq7TWf6fnNV8RlbwyUSnyIX
Ok3ZNYaLhajQM4fW5Iw9GNeIlNsOZhdINPaL3R3pGWhANDPbhbUOrGwSVF8vTaynyhvOKfKQvz5j
MesVPuRQRv/riiDKg0JA4usT4PtBjY6FKvGlEO5m+kWzNdbSWOpEXuXsY7FC1Vzk1gfv/hzhZ978
OMROv3QDhy8iVfOvwsHMNYaIbhdL4Fh9eEsBH9ZiR8dJFk+k/m8oOAK7lXSgmQwgaRJ/ErLbaxNh
AYVzJNSnBa/eSeyam6VZUXiFtYE20CFx6+wKVW2z5R6q3jA+a3IBUf2XGwKqLxBdGDKSueW58mJ4
D0t2MLMJBVghqrFFkJ/gXJC79hOCj3ea52Jvb92LyRffg4CCBuzXEFgq3trIX3zHPGCAqD3XrhjR
OmmAboiBMIe4XEj7suGYK+VHka2g0RRdj2IDZUAsMTabwiHQuBnNyRKBvLm+fN7Wnk/YUlunBcMh
Uj6aezQiaHt2jNxLmDD9S6N8crpip3ZGpdtXOLVvsOkj6Cc8pZRvzF+sZJoPDateRE6FomKM+w8g
PYQCselQBtMrX3IzLTwSJj1Eq1lB+m0E668b6k1adymJ5JFCmiqj5Z3oJewKBM4x7DGq9w9e7yWI
kjfoewmUU5j7EsTdicoohkL/lFJi4MW7H4L4hucy8LNRYdvT/7kVKr0PBtLw+8zuZ1KtDFVRvgS1
WqxgFf6hhP5+FP3tttSLghz/tP17wxdxo11IdFradKtAer65/IMlkw5b/ET+DXlGnuHpgh62PYfr
PMzt8ylNLZtMhkP1YzTAGUo0KAHwROCo6UGbS6LHgYt/wH5MKF5/R40n9a5T8PkTBig+lPy6EVl5
+q6qURFooOHfQ6U94vzoalNYbM82akDiJeiASg3tWmj3gDzG2htlnEdPPoW8n0R2m2lePeYyoS0H
O0R2w+uOdLz2808gAYdX0r1PilbqOaPrYx6ivq9lZ2fv6O0XPgqzihqapVcDCn5HNQ9vMUOYPoRc
KUsBrkPFQOLodgV62uWxiPBinL81ACYlXA2nR2D09KZjZxzu6qjRWMbO0nUKNiRPMBkk2fsZ/X03
4kbMXOrXov15R7pNpVkcqfTCIRyNyzcFo3bDX15uvRJQyoMTahCyZR/Vjf/uFxszn8hUm8SreVCJ
k0V0j6WovQPd8GbOUr9WwPuU2tMwG2oYMbaXr5V0vdU2Htpbl7WRvQou1U61zUl9Sh9by5x7ddea
wY8LZi0QCHxtAbsRh2sAG6nmduwkNNl1WVxlhpTztik5iXaufa5RaSJgR1tUI6l/5l4Nw8xT5w71
IiPbkAFcs++z/DTrrALTmkm47qW1O3rKmE75EaLQ+cy4YcWx7SEiG3slvLQJnRVP1UKGGNf24aOA
ubajBmGswYzunJ4mF48gTw1uuMgmS/DsEX47soLGekWs2Jp08u+jI9PrAo/85ihaXNUGDkSm2PsM
kGRnJqOlXyUVT2rI8zJTTT/wSC6D6UZKEB+wjUO8VveuF6bYP81visuIB8Y99dcfI7EdSeMVd+Ye
x3WDK/WL1I675CNumM3voU1qyGyNnMKzP8uIRoKaEF96PloRG2ALMfy8dLlbmAQkkebw883zZiOC
VjCMLv5G3FmdG3OnOpGWITzsi0hkNK5NQeiG9Gi3n4d1Zqh1htIB/sZ3uR62wQQPsR4tc6uIZRZF
CAqk7xbHamvejOYxaMrCpzV/I97ZtbNmS80TwD9dBkWTIWdvYzfU0Zp96XBLyomlv6EiM6gcwRXy
qwMlMgtGK8SLI6PNPYcs7C1i1escxWh5ZP1KjrS3kh8xTtjqywl95okf2WzkZD7i841KQUV8QFl3
VGxCBF1eFp5EvtrRRJmOXZBOPuverI4u4sHS/QO0QpyKoIEgvzgl0pqLW/AEmOv1UGP37rObHgf3
WSn8O2mr/HveqYqXGJFjxKdUT6BEWeIpLiDzCa9tD8cvzCs/QEuF2oEmJwZJG6PsoQVoOtoM9SRY
HYt8adq0Hthu2sNitt5SNs0BGkMKWnNn1XeuuygqOLACZ75+j+Wyxv2r3AOQb7thTjbxXZdSbzGA
zRJh2CFkYMgnh3ZQ97i9O1joyb3JrxowxrgDyQPOPwExqoWN+NTBEHHOmR8HAx25xJcxD8QdPtDd
WIvoifnQ7+ewJBNiVQkAw+w3sBV7T3xJZztbjfzzAWTjHJc6NzNw7m80PVry5D0l9WBKR5ieuxvA
EwIIm/Qaul/WOSljQka/Uc4eOzjB7aJWdO9//+uQptXknNpUiMObKFbC+vjNORpXIVIUmDNFcvE6
wCtTskB5ls+6a31uDYidxK/Ezi2g4Hc2fqH1a3rgFHC2wIq/+UL/2/YwHJ46DdebUdgFkqBuZ8nS
FVSN08JBbyOxeAdJDTjrSL9epVuoELfoNPy3Kwzu3ATyUe/034aNKY7yXf+DK8PV7dGVr6Kq+TGA
X+ZJ0MfC2oLeBUht6ocOtt1Pcb6vLv6XaPYjGZffESr4AlJ8ZckZWwCV7Np4/gLRN9H21xQ3A2FT
Gkp9Oz8b7M/sAvyCHVNs2XpjEb481coAFoYB+FPt7Opx8jxi1XR1GXCzdpPRFaFuDvT7ubtM5RF9
7nUKy8Rey6qemY2UBL50eUak+iVmjTdKQaVfrQD8qjau9rKKjih0eH+5dFjzA0D9NfSjFaYiTCVK
+f+aj4PS/a8ZGLDiRtXNtqfow50KchOgT1v7JlGGfVu3N+Ailr9CrtJLt65MfddWYIviq3VA1qid
pTM5moB2b21VNqHH/c81ZfwUM78dIZQpqVdL1eS4SevSyfQrHqcnR74RG4wWhR69eUXKEgfhuKsR
K18OH6K2VYm4mHH/5Jmt0iLAf7ab8y+wJUOP13hqVG7bmucSlVIbSN4+lH6sh3OspQRwW0be/kbM
Tb7H+mTHbzyKQt3vOuXp55ZnOi7Z4B6UcEBJoxqT+nsTRlqb6muVlJJ5S6t95WbpsxzASDa4VQ8r
CYJH4ejAcVLMOnMQFbGoQTIsJLaWM+j7qja4agWuBCQBGzz3sCVd9vuSIoPqj0i2SqsWSn1/JgRg
Rc2c39rm7OX8AeNg89K9JagqLbZvNB/2LfDLU7cZZLCNTuwGFICQav8yAyE+HE8TL01+fK1Z+J2L
oDiEApAXPAh20hLM7TQw3RAp+NavDMie79rokiLnK5ZM2Q9uDXg799uj3JKH+jBBha8HG/iFJP0c
YcvI6PItk9POri4oqPtiag0WgBsl2kPD16TvAVz2paQHYopCR6VstMUJxFMvQi1Mz5DdKUtqeYAm
TPTRKr+ricz3/4Pjg+Qw6+RXMY8JOthpmh1+7tfbvUqBPdP9veqasjDe43UVHgtUL9G1d19efD14
1pOI3Td+BF5m2ZwjX51A2LJDtdRhuNUIBiAuGGtq5eUBxM6pxO5R5MEdVar83CbNjPHRkr8zhlpm
gnkQBxh7rqdznsfDhGPgYMwcrkd2sQZ5OqNKoes/quBADiGB02vLH7/dhJUWZkYJsxrK3JHvlEA0
B926OrYjlt2AKMU1QrZE+Nplb27p9QF7pMolQQ3DG83ANmmE87EL5FjoalZiLWDSeE92rd5CayoJ
TFAp0M7Hrgw6hf8egMPQTG4TgaOVwk7FGhkJxjBOBNBJlN4Iq/d3VEVfgdmpG1r+C38PnsH1btx1
icZ4cYM19UB2lCJu7tybgb/8dnR/HHUkL/0cO25+jp2FJcwXkm/6DO32B3PtWuZ9OI/Ma7O4NXes
kkWEmvX9zTnn9HmwOlAOY3j2Dp/xrhSuK23Qp+Io9nvfpCpsjQUk/chjo4/c7VYQGFC4xTIXkTsi
eAmzViJiLLhPDrBYZSv6wZLSbCQesiIl6gcHbS878CPAfCJiCy4sIs/mopKOQvg3wH8JIpbS47Cf
t2SrWidGhOS167bdXnXvuX9yIVvpSV+MaQGQInj1hf+ep6kLExxgtQVYGDSeyWmvwvQ4Wnp5+VwD
9gSHG+GuVbauHJFP/GiV/wCFXSTNqfG413rS9bN8MU+u6H66DJnjZxAi4JdbjXxoPKzbANh4WbuG
SIsZ1HPumLBegftsgNmjCH1fIBkXKU45naJqkEbxTy/gQwrwZK2AWBXFeibKru+5iGd2CMcATSk2
QH7c/rInCZ0WdDyp3arUSlw+96j+9MvsFEGf0/LWDdA9MYOA1Ow+6lCxy7i/7nzg1WvO0P56rx9A
GfQz/volA7+7UdYuG6LMz0corwm4HP2sqriCjz1GdhoT4SzSLfyP4nXk+NARMau3mKED8J+zG+dR
f+IDKfuwpqz7fOF/gGjDIqMPO1tSOBWcDwTrfivn5yegAXDR/TI74HBbejSnfaY3qZytfGlIPj/R
Uh3Zffdq2I6ZR8ZKGjZaxanjsQLZezREAAMMuN+SngqCAUNpX7qZbTEoVG5EkIJsL0o0sErvqVlH
yDsFSFgV7xUtLN+r8VtVfw8g7qpOa1LV7UlstSSm4QtiFPP2YwfZD6JUXUzi2wUh+xFiWkhYW27T
WFeHyGbzn/TdnBcBnP1NFOWEDjw8fUzMRwmhqkJagm+1eRbzwr8jKXDn5A3FFZN5bfaxkbl4H2FF
9EFXlqwqeR/4O7g/oguZYEtY2Fvuo2MKNQJEm0r3q9PcWBU8ra3mx2HFWwOcodPN0i9RVg7AYeDg
yAHFBt9RL+vm6foifnFlZNb2ijqoYusUDIsPscX4nNBuN6IU2DDRiyoFJGB1lrGHrh5rZY8biOZi
j/9dvrCRWUwpBmQb1zzNYywaXab+KjcSc0jdXAdPil7TJgT+KFUwfhlY4Ec0RPpo5TRAU+rUzDnS
C+tmgURAsRzFRLp/yD8Akd+P67CvZ7lC9l8slOAhTDCB6xFwNAw78ZR+kME4J6tyzGlcjhDgaPke
Yzlzyz6LyTZiLRojuRi8aJ2povc2ecX+pln+tn7QEQS3Hcj46GJ7VYcRJM5kqmOVr51r5LRmcHkf
Axd9s8BiiH8WEtMDzwk2dPqFjBc04h4pr3eYoX3tSH8LAyWgow3BhsG+I6nLnCAWQdumuwH3S4Tk
vL9qKZAerhKu5aAAZlvdDTIjtBaKkYvuF/3FYbgANp7mTpW16JC+EqkvQTmPJ5zvwu1jjXN2K3/w
7DB6NsuNKyFPZEX9QKZPhl5pHZc1UfSCVEZVrDqyYRiyHaxgrjlMGZT3oOUl1R/wJTFEmHeJbIvT
Q+f0Sg4Oxaodgzv+SV2Lnzn1RlrptWZL25WEpI6RzoDyRnlLSbJ1Ilq480C4iV2zu6cberT95yHn
VXunaHm9zerwvxiBL4T+X2yN6DRHHPhGr78xc6TDbeZ6QukLzBHTuXcfIlv58EkFwDubIwifMnVe
BYl51rFvKYL4Rf7eOz0c3E6/0jEOPOBOkfOo+wzAG84y0XTPjfqPSKwn0FP0AbB0Dte1Anb3eGKP
VlSB/N/AuB8xkTL/AdbpyklF3NHyb/l2w/ENJqFTzVdvoa9azS+iNJRQ2Rk08rzgsd96tI48vQhm
a5DB5mnB7NcnAvWpEyHHv5Fgj3+RMptL9swnaFvnpzD7c7cO8vwbhYFPNm6bEeQwLewqwm1EPBwY
nrKxpPCcV3TRXRtNJsL+8YLT+6qfxRTigaHXb1Y/nQ4MWktjPvx06ZhRz1+bJ9x4dXSzwtgTcK9K
o1Xzrj7cbCuFPK3ttoy2lnWm9cnzjyXl4yw25RErGCorlEwACVlWCdEuXyRhjQ+i6hSi0fotG6dW
7O2ow3DU+aVj7VbZ+LQcJdFqgCYke1nKVPOUCLl5+weZnnKQQwcLI1fhoHzw1E2GbZqxJ1RgiBB1
IriBFMxVXYzNiSmsSJHzqCLCW7xo30t8KMyjvIzQ00JRqC313aGBMYm7/2Uri0l+BD81ivNAnz5W
Sh6ib3ojJZRoaktnZFbKVGM6lK5+MOSU1LkfRM5LxbU/ceFRaBbn9RTehWw+/6fgqX/3V5o/Z+E4
uCCKfEnaNLy4jsoahtDERscALnV7ec8zSI9MIJvjhaYNtabAXG43wSIvn9TvRmxhF5ccVALctDdL
D7ZUvmfb24F3g/lAerZFy5ie2XMCHoxI6VRqvTvE5XHXEnzXSgfce0w+Jup/49fRBh6SXGdNIj7/
OwNFQKCG17BaOQzEKylrEfm0MnpASjtkaM6I1aep7N7ptsDcwMXhWlGanyZSUp61407VO6+IQuHX
z/oMvwtCCdF1rlRNEZMNLoeQTbBXP1KpgmzM5aNTUwQt6ENFlHPV3uGfK8zezmkb3ApEuB4thStF
i3Tr2aDrAADY9lY7ny8l0sWnEHBVKvnPsNynbz1B1qmJfvFdMLSEsnNrg+l5QO7nCurHa/jJQdU2
StIDDAgiT1/t/Resb04+7Abj8b5kH/4RTm/Dc1WJH7GWJHhEkq9M/aV8Kjlx1K+rpg2jJdRzAg+i
K209m3VnzwnbAX8rKDTuwhtT0H11oFD1SDk1oijkVzZL5D7uC8rpc1JFJDA7lPeJzM3spNikUsNP
EHhV2CscdRMIAPsmiExanxd4h0zCbIXW+05xT04eBeLfKFY5vVZZ7Cxz38LNx1miIfSE7BQQY2+g
cskc1PuVQDaYpwC5YTKn9QBCwWsVbyOgVNlJPnv/YsRzp1kJmcwglIoFAIL9e59PNFZynlrgaC89
INBhYYKop8JDddHQf6dXJB+tWH/TtY884Ag7DLbDZx+S/6GMcis0aNzVf6eXgEPl3RxV/+CxNSrD
BEAInj8RqLEoy9jGGMvMRVTZhgOkuqmBCii4AKFtoA+mxq1ru+C4l81tg29kFsXi96SZLILbXVaw
e3drAwCEow7PQEzpNm4nYAxsEEieQixdvgCSWO0om2fHlVmgRKdWGuWT3QRXKjMwM6ZD4lWk9Hve
yDGFVxbMLjfx/97//kDlL2mpCIpUEFAaIOCVtsoIIPS0wkVXgcqvMUWTdIhNtxdc/xB2cQwtuUnb
gSlWu9sd5jufRan1zfd0eg6r45tXIFa2d/jT8f+5d87I1b/vCGIw+pQXG20icJkoYOZQvs+DB5Ym
gnazS6PyA61YaOtH17n+JDhCcDMJjx/DxcrRTGZjCEjdVrJ3O+4xonCZ8Knu3++gdtcChEJtegkb
84jscVHvrUeaPLTM4udHmPFNTWt8cLHJVFjcwTsMOc9XPL9ZSfieCyxl5zlm85UbI1Llvq++1JqA
1ZWrVkzcTG/e2xqL/Kh8KQrG8FFHlV1oF+4H/wJ/IpOVJx8I4Aobn1ltJYhNOMZW181XMkE7nhNq
qEJyF6+Ij/oKnf6+RILp8IgNWp9bxkjXNuxsjF3DJ0MwdErRwXOZQbrr3zG9nGDRhvLHCxkYtQS4
QYXYG+eHCY6dyba04o3jieYVR0o924fiwnhWD4h0Cfjv1Q8HY8DNhtT2HAlo2YB48k0K3osAUueY
i00/+WC3s9e21Z/QntnBvv8M8hm27j7bQNM55Kh3qBBSv4IrDm8MIgJqTSoRImY4IHgxJjitTpqS
ZJgqoAmzSIr0QaaDHoc+AAkdUe0Z5FoR2+tvK/7p7WqsJwYtuY/Pxkhzqeiao+P0BYW/hMr+tskm
jMlNDrbtp2je/WD3ygQ3UGiIdW0313aYX+0pzgzrbEPggfYUWlqqrK2IIXFAX5GE3sdLLvdF2bmB
rghatggFR8nT7ijVPMUnnbjXz1C8w8WtWintR87pOXHVbdOuHAaye+hbY1kXJFrDCYYL+PO1RyB3
KfBBW9IocuqJ1MPSPXYh1n+k/S/ObMBXZIUcJ1vgomO+P4Hzr69QGvE7giZhgV9tIiqCkYWJn2tF
olMge7QMvorCeBHDSab7jkQZsqqL8GKUoEjb//GlJIjFfBBv/jMlOhvHs2O+Ll9wOocbj/DqBKdz
yTW4Ttm3qRAg1eh0rezwHz797Lm0Px6D560H6NcbXuNYyx1MDisEBhEchuLph7Fz39Pqi0dpTTSX
KYU3y4+Cpzw4m+DoSJuNGUWXMRPB1W33ajFgZuR6+JD7sGs5cRpty0/ys/N3zvh8xD7nMU8o7r5c
Gp+TqMHocgvXYjlmO6LeiMAyi9nHBnYRqHfG0yvKCm3SsHsdDlvJJ8Mc59j9q0ulwbu+4kB1HGNu
OeKXqpddYiP0UyqJ2VC49Dn8IgaogpVfmvpnYkY3MR6ZATiuz0H+bJvGQdlS9o6EgVoC4GVQJVjU
ht1wRBoZc5fWOVEJQTWXG5OQ3c3c5KLWnibhjJQqy6JBSXJZyJ6rb0mGtRR3pWHL/2kiArHFjrIK
G0pzjS1Y9UfsA0E4eiG0ljSYZTkLGppODkgrI4Wrmq6gV7kR8RS1mUdl0V4gA12daMAVzd7pLj8i
pBkAZ7wuB5aXIMdEZKdUv9Du6Ah6dUYTLcNubsqkzlNGs5V9CN3BIAwqruqx9juSNiiEHHbHH3Cm
dHIuLa0mds0a9tgkAx9ivsh7s14Q1dKVfJ0E+Vb7wnJ0OYwH++qX1yHY5ilaN4t10/lszZR7OA+i
GkOsfAd5kAGDlSBV12hfQfZlKlE3YR/Tx7+7uLpkkR+4EFnbJGAmL8ylcVkC6mofBnFxFT6lMB8N
sjJIO0VLu/Jui1InCDdbKSfOsZFEPO6/usKkgC3V2bU3X6bQpxwYHLlFSIv9dujtAsL0PQ/Gz5/D
1jAi8S+qYMdbSCQdOwHX+tIv0w7Q4K4P27nLg65ilvCQRylcEQwdTEH/mVey4tiNLYf5ZYTNkEYc
Kp7ezsglNRxOV1AJ4MCQvL0ZkgoLh0dvOV+tzvs+xsG5466fYOUIxyjx+226eLr4YpaR7Bgy0n59
VtRtMJyBHlFprVc2ZddbjVI5lnAoDP3tof4cjY64NYFAYWDhqeJmgn8Hw63CqcvaWVtQS9GyKBYf
W3DuI52lWKjFzJp4sKzO5KqOjLC0IaCV02KIybZd2rcoVLpPLh8x5z0nzh5cG4U1IcsaCRa547iG
PjfT/CPU20h9BL8n1ki6YOfdP4Uda/B7joAEII+iVJwe8OqS/IbP+dlA4herdH8NlAOS+J4Av/bX
7+Crs+bwCEjk8tM44ynXFsQ25quZTKLcWxWF3Gh7QJme3WKuAdr9zVFX54OiAbqjkTK5EowdeG19
00GknLUEsOQSHV2ROHPa+cb6Za4saGW7vym03iWd5MiS3j7caX/S098olyUwUQmplEzYhREQZ00I
Mct2dtX0dE1bXKCXOTh/zqKgY9rkFP5bhmCIZygC0B+XNJbtNaYCHvh9XixtcMUV1XjOa5ixyyzN
kk2YiyWKau/zu+HI4QxJoWNJ/HGi7RcAp0gOY3ip6haNpoSbf92Yy85B2IUAaGZD7avX6AArKS8i
m1JZY+QxVLV1wpDGaWmflD/014NzpxQRpNyWcBbX0TIF2/QVast7AWmPkQgNthoeblNOK6+BcJ7R
bnvQMFaFgn2IPlk8qnaMsVzW+pfCPCrb6L27Swb52DoFAxA8MO0u74fmXJwmD7gnXqOE8ysuzphm
6DOKED7kkDvEJi0WZOd9NJplDlHUt8bQ/CfHzigHskN2XvPtMYJxKBIcZSctR7zmUTHaDisxjFw+
LPSaAMOg2Jc0iYq3r5QbGoFyAqT/PFzx6rz0UT2u1cV1AC+fVVpyxxYBKtBcKG/Ij/xYwyifWWlY
uvtRnjxl6Cv7dRuXySvwWhItlg7GIK3WYL/OA5Y+sTR8fg+2ltxaJDEn3lSm0+UMMznrG5h1MZ5/
B7CdJetMtXDqX12JWGWAPvJf2LEqVcwRdmKytbbqUlsT2REkrq/nxS16g6V1qlAOPYrFq/+GxI6W
mtpM4iTBzuyNxHEKeuedOZyVRSIQrzNFh8SBS8VKf+K9YwE/WIOnFuKtQSqkbUzmb6zX6W6I6e5q
VSgHYW4uGu28/BD8PuTGP4JuQxlDHI6aTGb4+kLOYpcHj4jRigcDE4JsHPR8e3uHA9ESnuodPp12
9dbMvZBJKcLI8RS4l1+xuSqmuKOLqoV5kzTPoFkjQgln/BZCvoaSPL7zp2+vezmfThNu44saBqiN
+5v4+YZHFo7PxUbfdm3+QbCdhuXUyXDvOptP2r2dhLvAgA06kJei19CrHmfBrf+Hd0AixEvceTfr
OQFh/+620a85nUX5NsK3/fTLXOlLsbuCyGjLahbj7PiT1UHVa9ToiYncQptIwBLGnZg45nV8BW+J
jgU0BTghxmvwEk+t5zzHyM+V4xiiurubFyA0vI4Zu0csdtU5Ma8SBTNnzu7aGlhZTxVZ4W4cWP10
4j3+7m/WNxmx2xlNYvxTjoGYJlWm2iZKu9gN/TjQGefQKD8Aai484gVkviUzmpOMLvvsH3K5le1l
2ysw1etsOYvm+/BC9QEGaMohntYx2UogEv08rYVGLqKhOl/mQBEEb2a23skTgwnToIQwVNPfhoi7
BEeIZrbmS+MdYnswK3bJ3jOzV0QQvOcpJ16/23ihUPT4fFQkogo3/jhNKefQY0Ko9n7B83FcRUvG
Bn+w4JokFtgt4t6xXEdRu/SL8iaf8O8txIagACCBXdqVwHFQdb1ZwClJLshGWI+ozIepOPn4C20a
+JDCYX4jM8xNSAfilpe1deEQV6iG9LmqBvewBrEZw7JFy3GtL62MjtRg3QIyHwLcf8B3xuBw0YU7
PvRvbIZXbcVSMA89VL1KSXY+O1IMYuqkvv1eQeQ6OkECsGpJXohxEedRC6ekhDVvkECfjSKw18fT
r/JgE/UaJms8kpPPCPOF4XBQWz6/Z5QXuCYWvcV1bUz3DCEljdRWYuXRwa/XY29XIeQH6Hn2WIvo
lngRVnIn7rp/ZdzfpH16rpdDnk6F9GX3YIdfnZdQuIXS6SxUqP+yuJ8oY8nLucmWBRRm55p/KJg6
FQI3/eo9fn5Z6uPzwHFtXuy9mYLunyUWCFN4zTOjimFqWwUvuity4BprFascZJBftvTcqnuwsrkS
JcM+qmqZxzqNrHhDIPaUG+J05vK1NwqzsDQdLA8Jm+yjJi3x3ULkucO99SA4DrmkNkizzhEha6/m
L4vp2UkVZSDXN9mZiOESw4F/QYjkR0Kl+MZUYVSWQUjSQXinDngDuyr8qFniMMdBUuYYbvq5BY/H
xnvMhXMkRqjXLO/MFNrK7FwkLXDcivLJW+uQFc2d9rbTMMnTA4tLu0iFTUOJQ7QMPMKAfJYnLe6Y
nCMvFMxeGHJm4nLLy7xm5ktg2UUTspBGB1ZnlIkngv/WMFQOekWw/hDefkuWlbFFT+hCc02XcJZm
QwFbiX8yRqeQD4dfavBCIoQ77xb48UIkdBscljFoOLqRBlwl+aL4gTQH5q2sycKVLqcuecPkBNXh
Xhdfj0uRJEC5R3II5K36dHDopfqEtFUKeK6+D17Dwl1UoOJH7yj1+X+oq0Sd21e89b5ROBysUi0z
ofRX3kDTIk7VoGtrfRs4VEFd+OGN8ghAbC9Addiasf4IuxEJ273biJ3g3vLLBxW4BQmCnqYKQD5w
vJy+ml41RvXGDoRw2ISp8rq3osWN8hVgrHRyDftyOdEcSHFzOpNrCCVfa6OO/8PHHwxh5sOIQAus
fSIgjEnPcGg8iLtlY3ZWeIhAfHzcz9c43T4k6ca4Q3gt8RCn23T0ZujexzG+CDILFVflwhxy3Zui
ZvdTkK1zwH5mdpFjj/q/4BnuNcsRcGlsRbDbjGUNM/U5aYQwI4zt3afsqOdFovJEnoMFSxQVTzB6
HNuYkfGGQsb3PihZUKSkP0sNYX8+U6bRrNYzSsCG/xtJxWhJWEnu0Y1Vf0HavZ3vaiBhN9DpjhuO
yGAfeVZ2mk+SNQAg3wniA4S8dJLLSJ7yX4xsk/AP2/6sq6eY2pAJBxwyridmXiqqkXmC/YrwQRjR
o0BsKNF1cGR71k1AuzMyhH3bOBkwR/I57LEEJpy1/zdIh8a3ZYXHrajzZGZ+krnZdNdm30hLXI+2
/nezcAD3A1ElvKcv6HDCdgRYLvqFqob9FJdZFfPjTedeAak8Dy3qMljIeLEsL+daMOj/eB/8B/WR
8XhVWQkQPLFHDgo3N+oUcCOCENdxbV/QFTeXQatd9fmQellsTbBb2kU1mHORYq57zsy9Z4H9Gvb1
s5r0zcuotJqKW1/GX0QgDFrJSp/+eYPE8TjJSz2ko4kPtsK2mmsE0+G+OjMQPAAiWAUQDZwhA6h9
YMtKCnlCKZgvUUu6MSYcJ08aCySahaartgKZqVFe1g4FbGMNvXuI3pqs6fc3ViRaJcHROX+DsdzG
y7BwMI7YLuuW7qL3CpMn3lIKX/TNtf4zpjc/uSbjPDkZf3O+JVdfR6ze7c0bUBcNrkDZXUL1XI2G
v8dQr2z8hEo/Chla/HxeJcQ5AV7+3cOMOKOkz1p2XgAJZCJv5Ykc4HK+MQNaJpSU3KY7jSOcBMgl
y0lv6tADqxdPqVifyoE/d0RLgcwF4Ojwf5VrRzYm2LXkw6tV5AoTljXa7gnYE/2qxhZ0HZ7P5OjB
oobbCLLPfq3mk/02KPmeZ9BFGghIQ2frBgClCnhhVbs1oO6WuD4tdikBOtFQWBStyQ6qsseKmjMi
6x9OjP0EERdy94UJNKIPDQd/qB98cGLlmpjSKjIp/191uCyxVYkxsGX2SAAvhJmp3N1R720ORQlO
Z0/Kp9yXnSDNcJucfRvOUbL+yMxiUhQa8zjbfKtndXkAKVoyhUfou6gvsc1W7JNP25RYSV5JLrSW
yOLDAZdVfofO1CxyzBqkNM2kPLx2nbAayhhqsJPlw5oreBnMbPuKV3sV5cboalZ0XxY56mAzauzc
MC1BAnkRfO5QvsODVJvH7b1hYqnwxMfGF56Fb/4tA0hbxKAzlAUo8NXOrYD73MBwK+7S6vREGBg5
BBBoQGeFB2Lov0QfVrGGnRUU6w2cFX5NjHvR8DqCRrWqiLLZqj7PmuKUnKJ1ft24RxUl6hlL6cTs
f87Ov5VrEOzr5vgvpvVkYorUKrZq9FBHHvrJGtCs5Z4Zmrah/2BYA8hOhAFVvZj4rQbF4GujDjk7
NS67HbMM4oMD5tV/3SYqQ3QRx33HpPEJAHIQQal3iHCc7CMJLT/zf1abPwkCarEO2D+W/HFXi3Pz
hi19tDZaebB1WW6QJNfYnGz0zV8cwxAbEA6Yg2bmuLb2oyLKha2Fq7E2Pqs0v1VtXLyYp1iEA+A9
KBek4n1h/nHtD8zerEdQZtNL53DU8bOuVuwHPPLGnW0gNb4URjV+rO6habCgnFW7Dl7owT/I6a6h
3fwfAzfpA52r02EbClXS2+FtHIbz+hkxiHnjMkndpBUOS6kiJT6wjrmqP0NeaKVxBUmo5NeBtHKG
9SnLzOTrVGfqGnXOwF8ZOXOpSUp3LIJskqWErr28/mfHARscnqEffu5j8mpqF3QQtLrkblu+8JY2
+uRgMXA6J6nMU294GgXoEw9yjHR4kKu2vIXYL+K9GAra65zFzLema6vO2cykI5nOY6WHHCLpToHO
bXarKpUFRQ5GJ2HMGIuu5oq9Y6TyGsntmUYjQEa5SwtF18GuvWmVxAmF0bSZ43pDeE7jOelSCLDM
4mr23t9ylOSXY4Sw/WJ8s1WECj0dV9ydHwtE9HXsT7wqmj7q8v/FBpjJg5wKJk9uMBi0203TCKmT
2BzLcJQ3MK+CYJ7kQacW8/uWrGysjUvZVx8D9/0evxadz8dr6VGIeMZ400aO6MEIMhIv0EoLe60z
NfEpK9RInmArlcDpnuHkBmyRnprXz+hxCovnQzqYF/pyS9cKfkQyN3gsuQ8zpNpOIoKdlsDWzEV1
sMK+uXDLi2gDICzPpria4hcO3MRQzgne8aPpIwiTgjSAi0tyq58wc4MqLGYA0Gn0GvZwr5aiH/gp
vKrwFU9SzdBzDjbBWvfY0yhoIr7gTsLCyhjLJZ9ZjYd6CTzzqYPNSz9ji6PB8JyvFcroQrbv8K+7
Y/+bgkIcu6R2YG74zhXBoBovHw1lcmfzOWEY149OYU77PmrGV8b+o3u6WImrqqtJPl3qV0yxbcW1
IFH3Capbu1IDr1G125BB09tKo4VyohSIr5t1W39O7XvxchrNspWG2toQP4dJuTWhPUBA1vh1H0GB
ZnmYHiAtk9zUZfVAscvWpItspRTYtKGd0O/GGFOeD2Lel7ieI5V1yy84Gft67xGmgqKLstkyY423
gwQvTNe3j5x2TFXYeqDy7dWGd1utryHwXrPylHcbmknos5K6b6cN9yfYLlJvyCCkCraPkpMru7p4
bVC12jz69iliHk8jw62SQpPmNmsO6tYN74rXFw6k2aR0K3KyKt3OqJ2X9FS8sHd5+vZZ8oji5qIj
e5mxN2JPDdYynM7bIy0mPO3zO+yrg8ruLAP6HyjS19NlNjsEwxglZLH1zXcttSfyEo0b1n2xuYDt
sBEaa3W8XJuMPSZ3CANKcIYHbnvS2vQIlM5GUGwkxg3w6BgkEzGctogDM3tuI4l9qk+IS1e6Ml3K
yClFKQTu5E4yBtaVFNmdBbaFb0vfBSahHgg6hTOfSJwXfH6Jk8w2EobRfwxTKDDehOc0ldP35SI1
XcaGzuBxjlLKUpsM2mqzOhu05nIP5Zyajxby6wAjIQ9ZzCmMrRzKHBAwFPN1AxnXdRlHrBhhcaqh
kIEjVBaMcqqnK43JneFx8JzATLpTNwBJKApinysQ0TUP6d+xZCoXGMOUiyaMJi1yIfS+N9/PQGdc
P9KablivBL/TkG4IVPtyqfGQKsotEmA8452DTEyLLe/42yuYnDdmB/fz02Q3mvFOngxc2zy2xpSa
x7V6z5GhBXtu3+dda+2UfFJR7lzCi16kpIkJFrrxmmCv+PzBePb+yeeqx4I593lXu+fhIGe+uBWR
LPUHsZaIfMqi49E5JURDPVMAm2VlbpYN8qhZ3mifY7z/W0XXI03pci25OkTiXFBjXCxozJswdElf
KeIZbSBs+Z+57xLe6KI4sKeD73yIGhdtdMq3urrf7LRC+8dmXsf5wwGn+epixIJsnc14/oDLh/ma
VPNb8sFQrI9DISKTR0nxV8pXLdfxGYbdcL+0r0ZkIb0Krq9v7aHC5Ngo98vco9mkHtkrjTCaKVcF
GWSddPAa3ZeisucbPl3AuBYJM3DW0Wa8fE/r+02lXp1fGy+gMl1UTPQ23iwfdqANeuZf+Y5eCH8e
PuYOT21CRXSQOGG5xrAIR7g4kN8pvO4R9rqVZDDfqOGJN48KSJu/jwOyE7+/TgQtWkc755KhrKVm
g4syOyLyNfY3e3vicsJpmcv6SCKE9iz2dtWvfKaA6DeG4MM4Y3OyIVCWwyWVyfsIOYugxCfUffTv
TNzKWpQBM2c8r9HosJ7UbFoj59iX3iOqUVEndQGg+QwhJJ+SVWrlnHv/7su4obd4GNwKa5bjtdHb
HsD3xtLQ2Uc6f9x2J4B4HhV8XQ1Lzx/eFwnkLKkiAzQSg0jxcGnbREFrCJNXCrTzGNDoj4vbotEJ
nG3gXvM6VDxqbMlUR9UnI+2N49CDQdXagkMmJ41QztgMl7joGn0mh1HkevOfXQvFYW2WzIrGJhZs
FTPx2o4GG3g7U1L8+G6strPmJS0lmO8DSDLDLMy69Wp9Bld0XBwF2AZic7AZFwXKWAhAR2x8ih5/
C9pL4pxLSN9Sp9ruQ/68br48pqfvqS6Gs+m/eXGUUBDtKTwBGUmL8NO4MUFuz7msh3X84ONsKtiu
P8lXa7S+DUeI9NdQIX1sP6vkMlWTUA4MlvTk6l/NrsXwc2GRf9l/u+GfkwkRG8P17ttQFODW/3rh
E2W5IsWitiNpMVJSfvkek1kITntyZpMvdZv3/8E3HnpNfHdyhWAmdcTljyXy+RRr0tgvu4SUfD7r
XunDsRGSbBXUVSvjkUGOkZtIF4ZlwUKksAILc+dDSXUc3N46y5vOEiLW0JTFew+9byj/NzfzUWF+
/RmsdZbJSDon8jp3tfaM0r/4u7wYESEB6V/pKCYAo9nIcJ+sP5LcPc1p4J7Esf+jp3D6zadnQGFo
K1oMbnRXSzP3oXXicAC39zlsUwFRhFWYP4/sFSVTShgzRUctjT3jNxaGnJGLe4uxDMvcXdazH80r
rqOAFyDd5zdxkeML5sky7XVIS3pjHCP8WZmyeQjn6xIV2LS2WkVCT04dwJwK385lhBR9ItfM3Yh5
YVD/L6aLlFXd9UE1czUH8Kq3tLwZimTLt1V/oZfqmlbAnbiPetAT8PiyRR36XK4E/tuY/ownZZ/z
Hl35plvqvBiwAkEZozcsqT13KILDy1CnGsFu1ogiREVxtWIrvL+32lvCjZ+9Qi0UCLOoVKYXkyAi
JGkQ1wUkrfoEA+EEXWsMsvGsHdPNcUkDqcjDVst0yCQdexWr7vLyR3WyBi00JEMo0Xe4AKc/LVqN
yRUQN3pdRjKwdJ4orDPkV1s7J7cobHRRMVujcjwyB2OCFMMCkyW0zqBnjNcIbFott9vkTO+IAHTy
q5riyCEpn7kr/q70yRzJAC2dgrdl9agbdgHJgGoya1L4dbcDiSoNyO+lA6lA6Iq12bSdkFIfM0VG
0NI/QsbgKtLFfkNj6R7jaJI31A6FEevK4X0pcukkIH4tJZENondVsJMhlm/tCaPzmbsnnhrH8aFm
FQOAqdGwCiZmdRjcxwNdL6CBt1rANUNOmwIcUj0Nh/jnnaxWdNMrPJQgL/EwtNze91S+dXjGXa0k
VNj2OByAzPK+0MGA/UphWETgQSuwvYGPJdb0SgCWoOeuSPNs7b6orDgPS+iXqQvgnEsCB1Ep4F5V
dA3T0DdtV1piyzE5YqfimuPXPzuzeCoUB5B/GFP6zowqJ62bQIgJv65W9HAN9J8iFJcojvXlaBEX
wcj3cIHBU2ZBGNEx1eouz6mGaKDkUEgaUmmspQRdbZPI2ooQLweWHuVGs+4X42nnsPyfCrHR480q
histQL5hufhVhlfJT1jiN2tdhJ24XOQGrzgfKT2P95cNqFZkSRSh+Vw5pH8tyLxDltZ27tRGd18B
sexaabl4eJ9FoIDZLFM8uXIWwd9Zm4YQgZNImEDxuVwO4v9xP4cuU76+F5Pc/S7lVuspejUaIVjA
Vge0xHpoM90PihiX1q6Q7J9T8PMB/Np8nIEQYn6YdDdVsSM0pCpJzCLwOAqpL1igjBPe2mqYby3B
Vui01xHAUwyW02ZdixD2xKcM3elEudIJvkyNvmOuMKjbpWeRTMjnWqTYobJa0WEjrp2oys3AiIh+
VLBCtswYWH+mR7GV9nAYovW+VBfvO0h+f4yGmvgfaj6NKT7PwYnoFIgft8MM3GyQ4JrcSwcJ9CPN
fPY8Rdg8hIO2R8HL2mRR6Ij4UBIK5DRdcsuQdEZpYGYLCBjzblM2TB2HoH3Dl2tRVGPXrolO+B5D
Bs2AvtDyUbE2+uQXzhWXSgSieXwJM8yhK9G47XmyJSOP5iINXa9hb+SGxVOi51y/fO0K59Z+HcO5
9wKXOJo4MFA+waH5rZj3aK5VsOYmSAyhSrxxz74iNFlnCPMzH9AjwIPYB2tvBjw/+LToVMggsKM3
47WCHYot4ddk5UUyftp27NgFRdhJWUp/lK8eNZhQ3LZhkPFphwYMnll0/JRhIeZ52VgBK31G18Ve
pV8WjcMFBjWyrXol1a+R+O/J9ZK4weKY83pa48fz+srk97Ppx4JQUX+b3LpmFTFFUsWmYooV276G
hJQL4z5cevcAMY59tGErsIOsk7kBnDAIvx/GBZdlK0iN/XIF6kzU/c+E2g8ZnZpH4q7fyTJSYok0
CbVHeEuFmprYBoJZnA5cGeERJOP1B3akorJIpiZLl6ta4OMvJ8Rr3cYazExCxd2cChJmgY7edKI/
VM0zwpzp9P1V/4NMv230ShYZ0yClckGg63Ccl3tVZoZoaoCV3B5Uim4IpNypxqqwDWxfWjA4SwF8
nzNdXJPsSjQeiNQV72Vj9CRFXHwEPxZB0t79DUQ80DyOmnY540gQKMAxvD/5Eu6rNTtE00IWkwKH
t9Y7YGJPTXLsZSMMBRRXeHGuCeRQP75WR5BPAxZ0kKF1NH2jHWZO+pM40AcR2oH1jHKe+Bw1W+cN
86xbjfdWnx/v3KERENiMetoez+vSS/EqOZQBOTYzHKIyOUMc7qTICcY4oQBClvFXuhegDPPAgJlp
1G+DTBQ011jIDAkGXBwE5y3SljfrTweOFoUp2gYh17ZDiJdcT3u5BXMjNT4E4RTCWeC5z5e3AgXl
AulPgSCorVcsv2opf1L38NrEdqN0eG2mEXpnvImeRtnjGs2QtWrrvxU3+fziqcjo3oFZQpJ7zdZ+
jrm+9/eJMnOfDmkqF0YS0oIbTh6U6ZD6wvbdGnbuL0xddGVb0Jr8KzzjqIxbhRsEu8D8fVmvd2mc
J/SUHTbKcgc6hepmNxcAQ0Os4isVpVEYivGFWJB1cN1BSnALIyOfEGilLuy+8WDhQfZMg+qeRVLN
SZ/xADn8xMyTudcT+BNztEnZ17GQ6KqJsHlbjJTxnMADd7Vt9YtVhg/mdIUXzaxQV27v9UF17CQ9
EPFSuBZoNstF/rAOX8+9EDvYs7RrDeu08TlaxQ7LkywrckwBKcUSSvyHV8teA8lk95zASKGkJnEr
SvK1KpnfvQ6zEEnyRWEvYLjfftwE83B9mR1i0a9MQzHCuX0D318vPDBUCNpCyC7fYn1TWP9JsVwN
URzzgGIk2WCNAXjBQl+5AkPz2KLf1HxEJ1n7cGro0HL/zje2bCfZl2csRPgnlvrDd6oqw9J3KfaY
/h85HAUvQaYRN241pFAFXCGUuPQfS2oL7lI53huDHpLj29vGNzHwEAGeQDMGZzIk50Tq9KhfcQkI
xl+Fv11uvAccu7ufm/mumphoEjuflpTEtiU0kdklZhuzR1m//S+CODdzjtPYGmzeDGFfcHz7/+jE
5cxU0oWp8FCPLovKAWn3SZh/1PXqH0wfDZjJNCbX9HGIMwnqs5YfCPOd7qjLf+uiiTDAsQn2KuH/
OiMdN6AWbRyKOxg58AKO0rjuFKenXwMec4nAiMkr8ZCadz4eyrYj4+q7r5IHMa1rk7ZEZEtPGp0m
9Lncr7N8tv22J/3PzMC5Uqb9fcMaJCg2nfk7kuLK229weCMRTjNZx34BQpwlvL0SKXxuEmxFye/6
vo8znt+glBFkznFCHwbJ7KYq/q2PGPTfXI0Hwz4lC22k3X1WaG5DbIIUh6/IOwkeAQHzqrXt6y6a
f71oB3z8CUKNPmQTmkPV76OKuZDNUsk/8MQoH/W5OQf3GgAsbtsemy/GipUlTTyoaLhk/dpL1vJK
5pm3lYqUrWWkleqWDywfORzmGdeN/2zpFcwpSPAKiatwDF14Dk7bR9odCHmVabND45IgzPa1vLwW
udVkneGjZjRYUezCS62c0xRH75zmlLLPwZnFve3o9VJbd/8xSe6+MRi8J2yJpWW/taQYPoZ9mM/n
GIRm/g4kkCGZmM/ZmGnjyCpInBG9vCRtubzTv2TYbuXH7gqXJRxAme2SjXLm/cHdr4d/8MKMmwMq
gmfDsUgqbkk1WricCx2lYpD6Rp/ALrJm0DxlLv8OId/tguP/da/JdjtnIqRZowqU48QQTOUAd8tW
5CEbLQhqFHHV5owUVtoyKunjkuhvNOS9IxtgKBL0SXaeeeygKbz69bwCnxqUOqiAOBTdvSVspBSY
l3FayKUjuPKbUtAWoCT2VOQz0iuqJNRLjW7aQl7L4Z0Bsivdgeow/cI8FU0KU5jnN0Cvm2RO9X9O
bDEqgbGxACjVM5jeOmheQrwEp4IHYHVgeOzmYaUDkKogTugeib8aR2DhNSJ6l9KCTWs7OMcoc4PW
eDn1ItERFvOoCguCFYbmtT5qClUVV+8nia+EuOZwBw0x2OhMyO3r7bcMgmC8TyKRwRz2noyD1svq
vtrTWoQDsvwrdRby6NfqepowSJLC0MikZgje0e4m3Vp6VAuuHIhgQiFVTnsXZFaCW3q19SK6zSQP
lhGiu6URpETImsIHa5m5BlyvQQFnlx0BLebQ5XkEEt6DRe5XgCxdpYk+WNxFnKC5qVTiV/9aMqwM
3dK2vMfm2sKiK6KDbL/yahPfwIUV8/lXIUT2/23jbRMzf/MBwN3IXBo+4GB0/GEEkNy9W0f1K9lN
1PaHNazSEPcmlAsaoTc2PaJpIuaNPoEraezY7mMbF7SbcdV3E363OI6VpfbnX99367Eaqxj09wY/
R9ZCAyjISQrmEpsWrgbQNjj9V6jkLdAudBVzNWPHRs4yPzmAkUF/+SezWiQ1g7BVcZS6KiLPvFhI
621TUl5J2BIyvkqAYoceTY/vGOL2lkLo+nn2dy1IhDhHzCnCRwZ6x68AHUNo1uxx26z5Lh+DraU1
yeswoWLAv/eQMi6o+t+0hTsdST5uI4uHrkGjpiAW8jVNqy56Zfbc8dzirxTibxmeybLM/apULh/Z
GZC4Fyb/9D9IL9JywbTfdKYginQQwQ/JJ4NGOcSTTsePj5YCXfEbC1C8H00OIaY23c6t20K4UKtG
R1jpVA1LJ7AyuNy9vPPq1kvuxWFFMd1IYvlyFM79EvSRZRkyJx7K2SMwlDV6wFWYqYAaqO4ifXvE
KJzTCrzKRT27l5fgXH941GsujfAwahsIMMpocceTuZzuq5Mf6wiOyq8WaUrI7+9maINwDyOcKvXC
HRIzRYvae4mPWcx/LDr3Q067OsPYVuGr7h0LxuT/L7Uax28R1j9feTI7k3v2Qs27m9o3YElnRM1O
ueP8o2WAKO3k7uo/WrZ8LwkKJ6lODXpUsgie4K4d+/2WuPb6egUKP2UemEJrzqPXZowLSo3mSDZe
gJhEQ2k5+CYxlWFZf5WPzSRrBDbKYsszpWFz5mltvZySSQASY0ivoDQtvhFnB0gaIe+IACe2ZWoM
iOR9w9H3bLciIjCrrdsxb/xjTklOECPcRwwixhnS5D341lQiQ59XAJiNgaFlylXYftCgVPUYlK1f
3z42mEl+7LuBL04mjttqsRU2yXbX5KyXQn3VybFVOihSDYYQ2iQB1eookGwJIgcpGTzvU0QUxnT5
ujMOVZRq0zXOS6eNLXhvPy1t565JIjeyRPoAicLffdYoY9DSW2KOzVpBcoKrfaFmRWs2+lheXlMQ
66rmHJAtUd2b5DtIY4cM1T2HxkHPEJB6accE82m4FPZkY+3Wd46lwF0LrWal0iQJP2/I88cthXTm
MzjZptwHy6jMu0250AkIqBBKsLNMv2IUgdiC3pQt1/4H1Oq7F8lmJ4TX7ssX95DK1I7tcHBh5zDA
lVDReIFcgmiC8v6l3mNfTohR873pinP3i8CUWCOLtgBhdIM0f4/iZsOBaPnZ+FPdMSqLPocqyL6p
rpf7YbZl71QhAN5dCFc92R9Z6Ugmw4y5M4vNlcf4jO1lLyD0EnM6iTORWsY6LxH33itLP1A/vbYN
Zj5TJ7p9yTkhRMRJM5KlGjGmlljVYuE+6M1Aga02lMGW8AAW1F/bWE0IycBTfpDnTsRKOojj0QQK
ThY9XssIqrY2y3SMMgjT6Ef4pZvJNUovVvaVCwk1vawh6od9qI/OaiN0ip3SXzIfcGV4X/YRP1zA
zuxTcfD0WQCa4bf9MGAsW3yun1Q8hFluyisotEHd1g12u5JXR7LClBWmk1d0GSW5ic8fhoF4o8rC
HrHblnWVV3dAmp5991ZOQiIIDgJcnoizJkaUXBqElegPvmV/a2Ua3nJgZNt+RknyxnGhSD80b1j2
DbKgJj6eJXnt0I8f0k2RJ3g0BbiOr1BHai/Ll1yRTQOhqnG5BN0ypHtiCn5dPxOd47ENe+z/SX6U
mDUZ0FBKYb2x20ZsVcZaKmQ6xffHjkeknFlzijrKlECeV0YzPk+3ERduiki11zbOBvjENEa4ntSu
OzVwDzdDEHvTruLmnFDaV4htnKwnOk22olb73ZdiFuYzPKW/FyEd9IMwMVlb3YTXkW3BtMFxG3UM
FaKUMRNOjEUytpP2xCoL95bt4ZM8if4vxsczMZQMpsb7MN2uYo0GDj0qM9hopH5dgFKC/cDU7u/a
MWeMFqhOwSuJM5HGIDstWgMJ/xyGtxEIQfWRlPbA+rn1yEjE3tAeAxTJmy2LSwRpPCsw9pjn66KR
/Ktc+pYMMIFvuQktNJMfE96Hp+cia8NYf8rA86jUNzG8E6rUEeXbDVIueIj8hhSdLn/9gycar3w/
LBMb4mXaexZxVG9HpUexu5AoH/IGk4hMkr4TwfkZLBGAIFhJxZPcXVmM2n6Q8elFu+pGRAUpcexP
17Iy5V6bn06cqDqO29+rG4MHSFgHzGRrwtC4CREpg2Rpt7iwnK5UDZHl6mo1Dq96vW1640RmjNOB
K+aM8HPykdvLh/FFK44mHn4ielokhlpA5XYct2GsuEbhpv0QZwsSICU/YnM9+aZ7fs4WfiPOEMjJ
y7XtBX6lQ1MD73zGxxOU253r9+VgaTh4X7mQaJhz/7IFMk+XuVABJDAOjmYAfAZogrc9d5EZcpsx
+P4zfDOkJPNdp5AjzMjpknJsNntkV7qHX8pG/GJ9G4lD8ufOxM8y6YhjO/dfcGmbR0g7Q43kJJAE
glvQmf4kHsA8s5GJ+kHGIjF0BGf5nM7EcYSePuanmQGM9cevDS2rDfXLmkUaK9JFNvff+vP4/dyi
nP4dtgnjSrhWuQF1jo9d84SsfeopiunZtaIk8oZJ2vlvBZI/Ow29/cfObpZLKupRcJJErwIikeK4
FOVV6xIpt+OlI71hFxWyuw8jpNnYweMGCRVqp+ys0Ig4aIfGfrl/COk4mx6+yAmW5d2yRo4hhYNU
JAoacqEAaYNsKSBLwod4hx99Zg56gZchLfbWxQN+YzelNHj+HDLNykMm5D6U9QW0Yu0rEGgdmHtM
xyJDNGRqc0dp6G1zO2GINt0egiYg+KPBdIxpn3pXYrssVj2Ym6bhe/CHljn2Q9meYaH6gqTuUv6r
rosTd3MQR7v3NouXEyyxjktGsdcIIGXaal0vXNYB/FOAp5vdhWwhHS2/uoYTN2jadYhBki/6g+UE
OHY1xpiANvPPlDwcxPCdfQ6eAhVxItfVkYKaQD85S/JHO+iYJlXh6YpaxgMruGXfgSKQC0cgvafX
Z7WeOhRB8xx3Ga02DmbOg8Z63sWUO4lKdISAb7+mx89fjf5UTRj7BFB9nckQEYebHNyOoJkJ/EPn
1IoWltVFug7ic9dy3uX4XGHKy0Ge9o3iQFWJ+X/v8xPciHPszrIFfR2NMGF75fwAerS32SUM6dYH
dX8Vb3wPeGX+7xP+R1iY7xgSzXwYha1UmwRIhxDaknK7xvCU48G5U+Cx8H/8Zznx5ncJ/l4qKGEU
RUqkvjsMTIwmK8Rzv8e37OmloPU1SYt8MJhlR1rBUaKVKvrOef2QLFjgo4TYZQuH+loGjiNdZw/W
wTN2SFHP2Gjf1xiqH3Uq3y9sopMa1OXI5V1TFdwQ0wYzebvQ23hY0IRqynZoUuT36ivlNd2J9cqP
5wZnOHL6MsquSnLPKoSqJtDrcvlOekv0HTdWSMcBVl5mpuXh01Poc8w0Ug1K8JWMBHO9ony8U988
U0z1zpkRkvSNn1Ypyapl9mHG9XImqHfBbmNC0baKsVPA+8ovH7+coBszy9A3W0P1QvD8ilyttpgi
sYi7S5/odPfUbZXlkrJuxhnxtKiLGTRkJH/enz3OGJ17IVyDPpBB2Fge97JFiRj7VRBKrXwNZFuF
Sy10tvYJliY3ceOrsx7+7b0wmTk+h4CLldN09FsYh3Ca3LCBDKERiv85H4gOF5yaeAIT1qf67pdm
nYLXQmvBUK4H3IMu09Vi2T3KAW0cog5739kX8rjqIr3VMLaXuq7EJ172ONGZbo9fl8qW24pfJbFT
wyBtDxE6AF4a6VO93ydK21yosu0veOMaUTRnc9d5UKF5GEtGxoGAgPwaU2uYaWgWMMfVCOmXmKOW
jpf5sEExQk7swFn4TEFqVqLIa0eOKJNzm6lvienCXPhMK/JtP20JP6xpusnmwGTSi+qNk7/mfiTK
sdakP5mKYKmkTW56qPuFLauoP7hiaHHuGEd6p7aqEkNK8PpXglGwYGVOQQ+0zRIzOgh+zg1ifWKl
m3RyDOf+IjRmdHb1O3q2myDXHL9+hdUVZd2dNntna+9nqpq6FR97t2UxjgTZhakPMPN6wKkyEXXA
s02x7GRsDfNUH+eOAse0F2UCO8/HRA2+EqBlee/XuxGp1PI5Uhe4DwXlEpkMVNu8CYH5TMbJWiDI
hKi0CWc51gdyKiKiIbFYabRUIfSg77yEMnTSvJxXiuFCk30xKh1yzpdJUt0e8z6DWIjNAX2Y6fdY
tU9fkcu3pXZBdak8s++9WWFKGaAF5W7HCgwVUMRPtdg+1GGRosr7d6r0s10dbUGTP5UcpZCymBXh
gWvbPs0Zkcp9nqFAnB+/PGONYoxQry9p2LQLZOlMHOIvm+yrtw3NlnW2TJ1SEJ0+V4P0xrjVaPIc
G6Vyes9SUwTnON9BrA8wdZ+1XS23H8/bZ9uL6GBJ8Kv0fWGpmdtAojkG7XzNbs1+QzMLEpgkdgc9
YhUy6T1rM6O9HY9ItAWf/BFxWv5xWfaf9XhSqFlYgRxaegrlVrmn9rFAg0lUq1VMoOxqJSDtelrr
qZTNS2ACYqNAPybEP7aZGWJcYral5XkiVpwqXMYOeGkWh0ppbxZzJsZjt2qA7wHrBJggIZMISHcS
mRmrZr2jWzDnrkmCgQ8wxPVzFah0FbUzKVHx3IeK2seBsVuqPKbegz/fVx934CrW9O71WdciYTM4
qF24hgaVtxfynPe981QFShJNnZTgJQErA4Rab5UnEEQmJvZrE+rC7AC9C9fkkPZNXMxnBpMuCkJQ
mLw/LB2fVjsW/76+uuFd5AZWYAo2Yiz2JqBov2wn1Xf73egdYn/yFhRogB7lby5HcQbHNrQj4TJ3
7b89wLjZCCvnuQzlzbppREdz+FkC54peYuChYy7UsExyA/VL22wwklC3iqGPJUe3JXTI8w2+Ylr4
jaee2lWso9LFtBd1Oz71Ca0PHx5oDFzBISY7BMFhgxYKmA4eKjEBD1Wb1yLoEYOAtp+4mvHnvcg9
CBbhdNiYWBIt9254nacUNMkYvgltWyGEgUtVh8LnRpUajJvk/7oxypqjKgGzv1mIBt4IwxoQnDVK
9Pfbfys/RnSlI6OdB7rY7myzMbcJuh8ntkUKzy3yrLWBztUENT8oN8tWyvwkERxK2Nw93/aPGq99
CytcZZFAWfCe+5R3DcVOU1Rw+XGqrA2H14A3nF/MNu/7Wbs11fCketh5ijP5WQs/eXOeszRnZvU4
GIXT23HrWRfrTGl5+zNXe0fILJoTApVIKNeLeRIHM2EaafsxNiTWxtNVvimJvSX5n0uuX64xwM/d
Yno+djAJptrJKhAlOqJUat+RxlcNQmHwmQiPOTKt1SHXdFjqHqHiS1liYU4Jy/0Mk705rhTAQRLd
j2yBXckWvtTVIkyQeMHNOeLvYKTtW3liZo5X1NfbyOZeO0XzRjHUGVcWlwKvem/E5P9uzJNdEx/s
WC9+KrdgDBD+q2nyRSvPHeCl6RMT8xn/2JRaUm/M0Oj98CjdjvN2gRYYxVQNAOJYEkXfP9shAy2Z
qFMBBmDW9m8wlK34AXCSM91RI0NKRG3RPc20M4JULmj1RWVPbg8P2kloZdIhsER7874jESILJ6AX
mZuYvGf++ZHw6LSQRNhmBGOZxFrs4crggsc4xAqlwXluLDCfRzSdaqngcG+L18nTaOTAvX/ogXrE
uOx14yxHisEhUvc60HtLvu0iRoS+xGoELSsWjv2Y4x7/7HLk0ZLBqwMcDfkPY4WygkBgomdZUYw2
bGQ0NyxyDpg48+9zs9uTJxGrTcm86mRmXXFGxzmuvduBJjWvL0I+5posbRcSKbzSILST3bMN6yHD
KDuO7Yl7w8rSbMLN4OfeU+65GXDc3IcujLG+/4QCma8gfU1Pr7mfH2VpsPwgVhnCs7JFHqbUHc9o
W7n6FfKKijpvJkWrXu3lMuncvVebr8lZEiKFsLtKVxdS0cK0p7newvPecgVdM76d9uyAaC/RFSLe
JgGqbCO/lc7igPbg4wdm3pwwGnSPwWIW0sxG2E7yvjmSRRUDsfweuavFHh6nbB7BooaIWzuSdEsb
q5HH9clIKVsoR9v1BTkGMGoUDvyeBisxQ+K9J4fyOZcXL2oH19AKU2UVV6VABJfz6PjiR743wDm3
MnHp2LI4yr8vq/VwUEIfmRG1nevrtaD54faUuiGgh/y49Xix+TXrcNllOO7FGARIQy9SzTmbMdug
3Ozl15laTIm5si2T3+49BL5g5CEUN/rYK1nEE9Afp+Z/CrojMhnNiT142eUeglIdvawf1zaaedF9
O5IIN3BvZCxHao/pHEY/LFKQ3315ekZihZ+fv1KP+GVAjzZMJOK/Y8KEMsaNJqD4hXDzS+FEs1ZT
JBa66IKW8XQJp3KYEBJQDIj9NVKR344wjUEk/tE2TS1fyLYl1x0sgqopfvnssL5xl/14RcVN6IMZ
LTfKixJjEp0jWhmOcX1+m3GynEY/JasRjcP4fCDMzmDw8WEe5UC3fG+HgO+usvreJhgl1PbqKiSK
tBVwRlLmQaVRqjQrPg/2QJERaToM0RP/V+YF1d9OpzSEqV8uKgZ3h+Ue1A1I34QIFuP7UztrIrux
uIKwkpCSJfX/hHcHKCuZRFazYpTGL+TN2t0rhIvOQp2zOP5HApvsUZjt0T4bLI0uhjG6TtC6aCYk
BbuzDzWzDKqc2mQosniAcpac+UOonyN1MiJv/aN4fucvSPGwxZmzK/BgrV9gGd0AHdgwr1EjSQ+u
8ONXW1e6si92kb6TyheZ3FgM+MVp40Mh3SGfidSKUrPyU0Tc7vcZz8hVlh9p1mhxjhO2rM27V6Wc
3k6mowvyQSa7jo98Xw7eybF+nzLauaPHmy7ep7TghE6C2RZVNV9Glq7PQ7qlaUCLqCOjyOj0ZPVs
bp7AgsovsOWakEUlV/SZG7Qq+b1cj7+s4+vkse8J71dZ1fcVCVl5TKEQnwCfKwwO0QM5c4K17fQV
CYYUaefPfrDu1oGeiYyvfDO/B9XFNeJsxXKJE8XGktlrD+jbhRNbcjxCVTOmnFMPUiWYklixhTqd
OOd3omYe02YwbGI+rr1XJB6jpJ7k8JMzubQovFUVc+/e3vK7EWgvvHuZqW7Fc/6HaWwtOP7vsfZX
OumhU/HmV+XJa5L+amVTw+InfgPWC4Phn00fx71KS8EINvQpC6ll7b0ujv04TNrLUl39gU6KO9KI
maKOuzRUcZUCroTAv/6gaGAwFkzBAk8wggZ9e8GnKOkl0wrKlggV1DRYFi9feufEyDI5um1wpdfU
3qAnd5W8J6LeZ7gPoAUxzyadDdF2jc4hnMRlpvTNFnQg3144qdmR7EMlIZLSoXh2alYtkxyFYYVh
TYik78SYuUEqFqlrUCU1fHxYjC6MOyfNvUIa6i0dhLWC4RQTv2jKsEmxJ8Q4HqsHL7y0jBp6STnQ
VJ5t2r/SzEriOyd9OEc36B+ODOnnAh6nlz7pAGH2galCT0nyESoddJgWl4CPVDH0DRCbUJzipYfh
3K2nPuNHwbZvl+9i6GVMDQHyf25mqYEW8O7QyMalzbPC+rBfkzlO2ZWD66G4Huq78MdqDn6BiH7h
FGftU2CGMXGE4EMeteC3phWu2wb5OTPF8MV/ffDA6Fzmxtgvg0oktOGaTyX5h6dgrzKkL0su+jdb
TF45amFDuVeq6F3QWzW5lvtNNuGaNIY6vynsTOb58UYroSXCuWyu2ddjonZWRWAYD0hKR4iukMPI
98/FwFMwreIZEEweVLl6z2TUkI1utkqaO96DREhO7nFClLb0iSf8wVlBL6nRFkyaBIyoozYeFlUc
eMa4y0RRg07MZp6j/ZbjEjLG7/lCd6qW+h8mtzluwCg5/9a6Sb3yjgBeOWz+4luti0cQxVcbcHVf
Qw6BtQM9kzn5egFk9D+9O94S6Q6fKJtcoPYzPBXYmaSXmjZSv+LP/HB96chDgkyUUqRV4Fj/Ht4x
CLN2j8n76vmuwnhZucHmUo7hsIk7ezlNN/9zcOd1NBW/50iJUUWHTR2bh7w7O6ZkbjBfuLxdMA7S
IyaOB5YbqvOMuUrlwxpZLrBxQd/hWi3/Kvjga/zk6VilQlrW/dfwiJ/O5XKRSHExu7SXogfVrwKB
lMSTxxlbLGDAq5vDfUXp7wjBY4OKog2+W/CTSiTVev3pmJ305KYrZoyMX6HYA0IQnLn1hsIa6unf
o61uW5XPy8rL5zT1KVndwFQpAsviEJkamwRVPgIRVoZgL5GIeC92nOLzNkrqH4Dw5Azj8DJ5mFsB
SE/nmg6RXBEJaUGfU7hlM8cHtiVncb9gYdjFtNEIGtCHZ4R/ehhcgqSHNMFsJnKvmFjfKotbGEOA
F8MXGQpa6UnsXvVZkwq9BZhvAooaUvAz3rqD6NRnzsFsjey2ifGDEIUy1Nrn4d1DXy8p0YoK3uic
2hvPEsqOIwno2fSiaGB0c9WCIJQugEyS/2hgHA3xyOARk7/pKccIpxYbYYqa03FmsVFSLIow489R
2ae2fCB5rxdUQ87+vfQGK0SiCNnbfMrMRTLEqNJpovMa7aydudW7hOSAhCKw1dVnhSZRwpzSUivr
1sshlCdxnPD+RxvC7ZkZXHgOmNJaP203/YwRzS2QB8Z36geqhP2fAjNKSURIQOKYmqeERFHt+lCr
23r6YG4IwvJX/9TKSr2AXER1GJei7WPoOO1SP/TPgTd7OFhgnJQ9NrAHC4G3XUL1on7Jh3fvFrpL
Z2654zkeYRGwjXSEZY0YqGDP0UGvm/Ulat2LjvijzSQ2HXzvD4ngfvU+Ru3Eqxg5u1NGgV1lVyOS
ETK36sCGrScvrJi3uPDXyg7T8R0OytTc2s4fW+Ipw1Ysegf7MhwOB6bq1bNUQu78aektBMaoDn1o
0eQaETrMaTzmzJ6vgo3F50jq7jVmUV/FeCejLjl3JQf65YTxZZdqJEIv7N+35i/8kAFUqH+JMZ+Q
shcoDsx2ehcf/HhGzVioxdeZdg+VLxPqE9xzrn6higoo/fPjpWARJd+LK4SZE8t1TyoiGLQg9XJY
JjBkNaZGd/iDTZL/JgWcjXvKgXytjVpBiIf7BQYz76/5ExoMAik0VL25BxYgAUJXo81OG4EJ8/6v
sDdqcsb52Vw0UVfLN0Eg/PwSrYKvvPMHq7okly0fLjVufPnPtYfVfLHcd8u73pXIRDpucb19UXc7
WqN7iSOPpRewyIwvr7QKlIwvXc28UijuTOuasX9GaUVNmZpKBu2/nLlVKq34svOmF7wcTtU6jJIv
FqB4CHdI6aq7lsOkMYeqIS9/5MJwNPRGwwDChj8wF+dRpgNrG/aY8xjYPrrbnb/KiZxJeRa7YuJ6
Wvdg/EklOg5zAN/vcmeHFHtMk1ektY76lOYbGYDBzEuJGldZijek7gJH5JspgOSFIehcMmABdv6n
LqGz/W5G6UWAMGENhhXkAn89NcaeApAuFLb1sYWl8H7YeUYrgZ2MjEE3WueQuCCX4j5UGq896P5+
Hz5+5d6T4fApYCUC4m6xnjGmTvG71VWG6nUXdVdCl8kSi6wxyeOYeL2vVh4rCCla9VYMPgFpM/3D
0inEgU6piq8VWWiDsjWuds4pL59RRblQiPWKl4K8RRAvXDeWCS2dndpfxh8z13ARX7r+w/uvhBKL
lLmH+V7HkQtwXfF7jyjT1WWepenqFWJ7pWCsBCTo9kio80MM9bBfopE6Z+FTs8hXXh5VLA6Nf+iE
HO16VIH6d3uZUuRJ7Y1K2apYslVgn0p2QmzaEVZ9cDWAolBLlVGMSgmIRUUmvP4Sz9FDvPIFEv/V
V7F0JiEJxxHKL2JWhYaMt7L8AhvIjyJqCsxdr8EF+ycXPC5wMPLCDnIaP/rgixFp3QYGVhiAMFRI
hbkmyHxaENcNzsgE+HyXQgyjSfUaxgkfOw/63Sc4tf0GapcdOkKphOZmA7i2LQ3M1b/P0EkvpF2F
L8E8PhfkaWoAziwvKwOQu9rdgStDFYmcUUXn2bYNVSia5kbSEcyVOBWQ0xID/btF4woWYEJp7WFQ
T1htlqkjg59999qPpT+KWQF1KTrc4zW1sYQsfUDLDCojtpWxNcCEt/+j37EHrr9fqORw6Dngg776
xpMByk2KmPhzNVY6M0KcxYs7TCO9Ozgp0kdF1yerx5YXjE//oHEf+vyPKm9WR4FrRIBsJXHLDpfa
XJLL69JSN1ffxcZS+Tf6JtkE8nDwHR4lo1jVdnszPjEd5Ge7bC+zNZrFUqG+zRUSsjZzzTJnhVyo
4dj+3HUdt72UUOpgjepXyefk+NQ8VTwXEjaTsrHciC3cwfg+09mgTl5catmzbZLzRgK8tgemXRji
FvbLGZ6yJguAeg5v2yqwlDRFsB8ZmBs267Hlsmsz7Qjb7gZ7b8rRlq/+RBYv1fxA3I59h8CRTaDj
PdSJdEjqLzY3uE/hj7nu2rPk93p3pzZ+CVziMKco+9s/Zvs69cjRcE/kjLBpQK5vxHwlMzDu+NUY
vg5GV7aFCvsXVDKaA+vHYYVb9kcIphXe8N6Ai7dcptHbM0hbxRXUEGwVDCWPcDyzPvo5ex+cS4aK
/1+BZhCcUPa4Ck1gL0Rk9wpLgRigwZ9GlIMm7U1qg+kne8O8RXNzWnIlk5e5e4H7+/SKpWy5T8+0
M+Z8yrIGq0BlbZ15S3/VAY1+fAgvWLzsIl0TFZvYtT940wyMAsQDtEpV4G3PudAeIaoAUdNBsEP4
Vq37K6Vz9Jh/CZFOAxVhClgeZkX5zcBqfcInSXkfMfbjJTKurSkA5g97pp3ZnrZ4YvO5wPf28vWT
9w7VfFd1R5tPvd+8LWVWpzh2p77CSQe9wD0BLc9kb5yCFSTBa+rnyooMgpNi0V5q5tCiiAj/CpG3
4b8CZNaj6CzUeNrFH+drXfm23FWhyfcEhzSJUd49CNo02wbCRXHE/DYHZBZn1u/MSKdpKP6UWH/7
im1w0t/81UP+bZ4XH2o4BbEFlwoPoV6Tlt2Zve5Eg9rvHKIfFbZwzZT2gjytM6CjPPX4R0TqKoZ8
1dCvcKI2cilMdJ7ZM5styRRWZV+VX/LgLxO9OAc3FE8RMIX3Y0rSelJ7TMnJ8OU/AoKDsg2wjClv
V/FtyyXsjQrCH3x14CClldZv5QSLDN11deT/yBeQeG7ak9fUdwJfKBI/SMlziCAw44E+u1yMPMT/
GGLfvx+X0enVw0anRVaZTuMliMTcIv5m0sWGsGsumvRUvjJJQ4e8Y6ursyxixYXsgjNYDgRzGl63
0komfFdEySsd6VMXtLOm0qIsWP7vdpp/AvFdfY9zOKo+hxVJpLC4leqwoGggfoKPSUsWUrM71ya7
yO582t51N6/iSzZcCeO1kjDZLqfVfbt8zgSkY46gIW04Rs9lvVv4q+fdI+5/zxLhfvNgEdLp/4+g
5ObagXWCr9NfurBXxllFrCX51hR+yLf0sjcgj1+YYxz2lxyN5ZaPUlgPwicESkozjOsOobbo4zXv
j5WZVEFSeis8HP4DWDlWSIiTTXi5YUsZMLRl2EXWrMYSbFySD6CUfzUFFBR36lEjnbNERMWTNtCG
2ibqj2BQyq2iGUKLg7eMd6UHtIzEYvoBvXAoH29HIwb7/ZXR/da65KFKG0ssUirKpvS5IBrUbmx9
H87yFai5inFOLu3vncNVq3W1qz0hPpqI4qwxOfXo6Tjl9F80tq3pv/ByDKaBIznQG+2TnLMsjD0r
8pKCFU06ohi9kh+cjBG6E/qOtZs26HLeYF3cbcFB4tOqEw48+DRNctaNLz3ddoV2bXD3L/i26Feb
ouiTcm5f7/J18i7LNvlDKf2vkP0sXFJugnaIrbiDqwa7e+UxZadXL4p4aHrvOG6iSiqOJuEb/zfC
bdwRIIF+wYWyCwhptLwHG0ayhHHsX6Oo+BBIo3XhAK5deK1GpLI/3xciXFY4RhsQpk7jhfkr6FdH
0Wr9KBmQGiIguNLQWKdX5OFhv83ZG6ghjQw4KU5BbO4qvGn0rjOvDvwjEcc8DDQB3b08LDJ++wnz
xlg2f+Ld9erH8JT36GyTHmX8gw0cdyv50FJvEUFOvAnfYelyrJuKmYxr/x3ZaPhoQxONc/7GOi8/
Tku3w8MsQ85TDRwDjbnZcigmUSTgHQsvXUPYR+oyZRp9qCQ+rI7nL/B/AztIqyLjXSiJAAQZ3fgD
Ck20Lxu4apabWiBGqmZqYdohUWVLcFpNwkaBjcctxXS3s4hG1oQ140vKh0Dy45kK5Jeyy7A0JA41
tRVNC+cMqaa6jX6wk3mWUz2QoF5Xk7XqmSs1FTm7Ws++9V3sMRWH7yxgKhc/F1jO8zJbNNwQaJcV
z5j/Kd5bjvCcN+tNEr6NHw5ZKkIdiQsPDRZXxeAQjY+t985nhBpAjqQfeeWpPCZEVaFx/i6fych1
lQ8WD3sQmPkp/SGj3QlcokzcyJ7RpFSaHDaRTQEB3kCg5C1UFjv9rZc8KiFdVQjh3TlANgrFczqw
LVXVY+rdWi2/rzvnoVE1l0z6JxbeDOML1h0+HFTjbJm6en451fmYkhPvsIKVn+vNBKwC6nLe0bfU
We1qpZJBQmNz2r7IzjB06d7P4R0wX7MS27TZqnrjPE6aufR42pgOrw7su4YVOwwQfR+qChQbJKbi
ISTxg1HUISyD6rWzkcOSckvQ1SAPkecw4ZNQDj2nv+QHt2byA5/+0t5R/b2ot6xtOnW95082PfaU
B//K4F7QrgwgJ5xZ8X6J8/HLtQV1JoXqk1yUwe7CxYYdxe4M1KGgfOdQBcqEJs3SERdZRD7B5Xbc
p8VOyzKkxkFU32npdrlqKquLmwIbDeMPZ5Wjdx0o0iyZtXkVFo3dWvpJHsZBczc/BdDSu+PqkgBa
ZvwzFvk5CnjFQd3jDWhI/TfiFdZc263xFdjpWIsYPs9FMBrLEp3dLdQ5/r59Kr36tImbK59Upk9d
9Rbw6YZE17nuszi1pM2dF8ix+dzT7HfyboXTvDFmAf9AAmvFBB9Zxgie/63Z1rkdibiQxa18mJ6A
cgGbqlajO5+5vhg4tl0vIQAQYTeM6BS9ErPTijz/5Z2fp9cgNrI9zUsIEIMzI6cgF9CqiukCy/kF
fl8/w6pYSYBJ1nog55NIU21AxigavaZ8/MvWolsOkv+UKb+kqMxBBFeiS6/LHlYLRnsNKyo/Tjds
4wstcQtNdzypOBJ79Ro2joyOEtHvE19DRgFR4ng1iTV9bcY8dcBO3GI0vRbFwmEV1mbBKK11o7DO
edTB2i2VtACqHsAD+N4AHPqNIe4aOIuDAzR5wqzP4c3k0NzS11ZEkSgQb4ZnH9F+sJGi70UBh9eF
coc8KQPJRSslvk2+GVv8qja+lrYqg6Ja2+qPEEW9LWPS3Vd8DXfU+sSkPGhtbzFiN/yrdzLbbAoa
YgwYwiJaOwNfJciYmrsuZ5R3oVk+0Dydsg+8BG80GHb7G3I28yaE2Te0onssYdIJS39nP+EZYnPh
RT7N/S0xhdHugt4N9CRvdVqUwHM2bujSLc8jwaN3bbbnwHBwokiX2xmKdVtWSsOO/rpou5sCBAO4
0efPBrDejN3rh5jzH0AJYX4pvOiY7bo1tbc7PR0BY/6wPUDsxSdv80ILABre33ghk3rca+RCLhgg
PYsMhVExZUjhHxVaGsJvOBgHbZmJz9UZXrJNCNx3AGs4WE6AWtGtZn5fo39dxSZfK9ybwvasyyxj
vinrLee4PZYto25v5pTFmiLNZbRngZ2desJPeN7aPTJ/i3dELOcBuYMhkwg8FsdmmoLD50sCoQ4q
3zRzxWH1KB03gWjN7ivhRA0Zz8Dp3C8LaCUntNFnY36t9UR+a89OjsjOo0MqLTKeMUKDFp68eBTY
eds0KOMcqPlOPv2pLNpobfRMMuDLV7kB/U6o/YFCq8HIBAVN+Ud9T1l0HUsOC0H2OYp+OU6FT4J2
KsVZUhpqROPs2qIfyIcLD1j6IRIYbmHvDrdMHHzTDQEFEuKUi9yOUgS7w3S87BlrjC1asj+67v8Y
3Mwu5MElwKEJFZWYCLmNvmqUpMZur6YUdeAWrgsuYoQAA0u6yyuprr+4AwdgQDZufqQ9U8vm+pNy
AjPPu6/1xfMzv3lrRqeHfPgLyM2U0jv0fb+P0zuYYM/CxMdwnuu5km14l/3BR5h+YNgztOszvMwI
B6Uexpb3NsQ2O3xNJhh5lUeF1e1+JRuCAae88ki1h7cH1jVnGkjjgKlP8WEGMl6HAKnZVMuarO4T
h0kaxWcnRyTeZNyFFgcUUszyC5Gw4L3i0YxJ7nKX/IfiLJYiGsNkBskKDQy6oGSYnCfWnbapp+/x
Q3uiT+0+zgQRluyIl0OqopHR/VduSuADljwsYeAKhqk4hzGyv2IfvSnmeq3LlGaK56JvgmuqcWXe
X+tTbZcveWdiNMlhIaDTDNdc2/bmJB3Xzsol4JV1XIiXtuiW097NJLJYxi4vCNy22R4N+zeHRU8m
8Dn5XfCV97cnlz0xjG3OHX53eyuMpeN886tUrxI5KhyVzIngYP+0L7qN/W2+d5bgmx8UAdo+Kis9
Cf0ocK0csGQL2gaea2YtAQYA2pfQcDt5FBi/pCbTTgBb10GUf6+irlMcZKBYgP9tJQn32s/aR2of
Vd/7LW6+mxo1n41m0rakLudawyu45x5/S1K6+fZ13hnSMuXmomWmT9TFCx2sEAmMDXhpqz/goRry
bx3/EWZ5qkQwVKGEYKeUnE5Bo9UK4g/HQQyYc+CcBFmVMvvgSi3zKQh4Pnnsh9qvppzn5tAGcG5O
08b7bbT1fDz76c6jNSqlXhaUws4k2VYFiTJP+3Yl9ihQ5tPMOkvxXLJFO76sZrteG87BR+HDce2b
RtSrT4KhBlRKot0/sM0qV+sA4pQk4Bnxk225gdxweyZ7/QosMvox/ITwdsb+wVL4eKtyZKrOTkzU
BpLLqZnRj9NtROeTLW5nDud+2MDl6cqIVM7kdwCDUrpe+f9o/oqQ/FsVIBafim3WgXggoYm+2gka
PCNOFlBw3si8Ogn+TKpCpttDudobRweam3HsZ7MngdvbbpM64ARG32YwalkIpL0int1Kg5sAIy5A
Om+HPSEclqlakqk9RhKeQir2VjM14X4KVTuczY4b2cTANLEbxHj/MV104YYb+BT9V7PEn4XLi4qM
MUAscGNBJtBFRtFc7JedbuSvdadpy44tr/t+IFbVQ0sFnVrglSzGp01bRjwIbJm6ygvh2bteyM/6
NQ+0TRJDEK8WSGcfGh3GmF2wTpZFfKR+7Lm310aNITE3g2P/sjshQ3d7c5CJAJXKEoRCgahUaFX1
RMr2gJyy4zof8u4XpflS7xHEkEuxYfNlw2gIlxFoHrNAOxH4n6/s7SnFVksbmrAs840hgBVZfUAE
uUeQECqjlRXWxSRGgX1m/Y7y87/TrG3RHsk+AN/xigSvBcV1o6/CAGJ/rPN+9pQsfVYliJ+/Pan0
mgCP4+9qFYdh0CzplgKGK2cR2lnnjAryPQYqP9p7CqcuEndYewAalUzL5NywN8mATDc3ZtzG/J4J
v+YlylnMF3HqEzaOfueNxTPeSY5Nv6zlnLP2S1Cfm7A/pNySTZPTlPhJmmIhug+jTTxbcjByN9SC
vMslXOP9PlVHUJ40CqI6pUg4tKiTtlWC6A7zr0BmXQ2g6eA1CyZ73i5nML5bU2Lq43by/+pfVBgK
zoTr9yTBuiDL5/MDir6N3MQcYpNvxTiEaG0/flEQqcqj61LfM3M9bxtbtWsGL7Xbo+YUbcfF09DR
ekDaWIhnmjn88ljcbsmNMGt+jHEDsE4za5iNMhYsz3qGxwc2I+hAwHoUW3vTEWghdWPguQGtfMPG
Nw4jRawhHD1dRot2Hwz4E0COWZI3FQVD40xlL+U7HtALrHYFOE4ARCBKyh2TeRzOppFNWzpep5fs
Zm0vyDMKPYEqWIId8pYoazVA457oBVl0LO6gM6ZdhL2k6lF/2oS6RVr6Ojswyr2Bi9+Un/LcUXvO
0clKwBV61l4XmARRKu5K3BYxR95iWNZ9MHcYa/eWDsdN69SMWme8sklIrPKI0xiK5Ki/hM8mLJ7w
QSIoBRW5RUD4IxTrYuAPm7w8TWKqfvfsXI5DPDw52Z+G9tBPRhdJ92Nsd/oiHxBswNNwhYYczGJm
wy7qzUuq7Pbv0ApxBLmMJ7ZlOP1HIBy0nNsIn+vEzqRlHBRHBqGYgYjOSyt01jWECZBlnuqdh1CT
xc271uuQSjm/y2ir2o9TDEWNPAqQhIP7mpIk28Qkgt4rzCCG37gmxvNnAFemKRqwrkiA7Vgy2Cd+
tliKbKeU9h4HxqdUCZMUlFQB8NZRv2B5ajM/tpx1xg3FJpNTkLZ7C4KyRui2wnevh4azrm7G//6q
JTChg3/Mx4XirKYDkzuyLJfF18Ze8otstsGr5XLqm8B8JkT/65gLyuwvRHzqeRVmGLGTpwS932Xy
6X9Cn9kZFQEoaee+kFf2rl57XUM4LhLF8FaIrOKMlpFHFqZqP8fgEWX3+TU5LWJMcwpGh+txNa6c
OT1jdFp/UTsmshrWI4f8EAQmq+wlNAbMdwLoLklKoas8PzQVw70GMAiQ38LVCHtZ6gTruX3a1Wi3
jNzIPYSu67VNp6qkOFVQWPSZDJ6LQBYFaN2Xv1+3WVLbd8xSGsYkh3bLVOOlkGHp82785UxIY3uU
50UoE+kwmEx9ZAXe2odRs7f1AVdqwuIVioj34UG9N7oAevP9E4W6p1U5n55vsenTAD8iZTxzmgNS
dlNbvLkTMqVWKPBmcJhWK5LQDdidl0z2gd7o1Rgk7IDvjvXHGumcTwENvu6M2Ip36bdUKslRaSk3
AFcjX8XN8RfCtS9C4V6xyatdMKqUV7yP3tAkO6MroTeYzGDecoD/0ibp8L+8QEIeiRMQqLw/96Qt
ACBkhvgEOxiCNDEBbSplfXnLVpc9JdT/gvwIeFUp+KnBxsAetIrsyeF/go/YPGYMxZjcQqByjKGC
bEbqKDGhMDwxRbqDP6uxDMalSUC7KkUffPkNp9sURQ/AcEwQUPCymWLMM0szpj0gcLpjymXCNgsA
7hug//4BIyau8TcCweRbktGf0UEngYE7D1uTBABbVR7Amca49QRdlUydR/F22IYDXDRdqVjORmS8
4ifmfo0OeEO+nNM7sFOZrRHRbSerFDXbZWoVdCzIrn3utLuAF0jx/ZNly1rOcCgRJP/BaQRd+UK+
5xMQkgzf3XbfuZrN2KsBUg6JHonsdc4hBmuDKSfvQNn9VUqNz0jwVVieFXlKBrvi8y+IZMOq/efU
MxDs4UaDT1SACxH8h6wCN5MFwUo2DHWz+9jaa58us4vrczYS4sYBrFcwRXz8gqmdvcpu6M68N9D5
h04bwlsQohEn050OMzZWWLxitwWxBqlIQRuscxQO6mx28ofhEGqioHJX4TwVLG7R4xB6YoDx5O6y
DHTT6QYQfEuqrenMPv2jjxzItUsnXyLQSMjpsBCjqBmpQcpSMh9zqpQPJ0QN6dTcGg7uGK0QdTAZ
H8idwhkWmOodRQpeYR1DFPYmI+bDUVEVzq73fNA1uwB8WiWxQX+WQTsbphjkv7WxyGNGDeMzoh+1
4yEaHivLdm6ghnRvLCAznSiqpkrtnITo7rj8zsXHQB7grtLLGSUiOBLr2G9VP5G058XqdlwKQSfe
oW3LwO4hwkUeC4DlFZDU6ikZDp4aEoJ1O30VYg9Y3wjcMt8KhDib7593HmiHZfSLFdx7XRnS1SBp
Mfur7kUV2Ho0WDe0SEr8rxVGHcDFRn34xTnY0aHaBsBEAv2LMqmWwDJEOC5aSLrpHiAxCA+0czXj
V2zG+1TrKRc/K4DwVmB6YCDyb3XVdG/PLpWOJdEMqjBjxVCwYXyx57Lu9KYkxrLpsCviQoNvbT/a
YAI8arVxShR+Z5HikTxMlhWpai/U/tNloExrOgGdI0f/ZIK0XPqCM9biHPWqrBS46aBdw5I2yl5J
AX98hdKNwdPP5U0Cuy3xVjQ38X7HOmbslpaTFQMY8e4wqIjAAjbl3YvGWRisp+uhOTpXM1CMQd/Z
M3s/QTfo6wX6ov60T1w0pCxbxVYABKNyNvJZtLdEj5D6UGrTih8yRnVR2Md6l68xyi68HR83dqz2
mibRl0c2zSUT+AHXet381wvX4A/fYFlkWzMMCyJr7dW82cYumCLA4wvpthY1ERTsrFW2dLXui9Xn
kslwgSdI+aEnjutxCUG9zsDmXAQ7/X96Z/2g0uBuyYYcDTvInPEtFFsJfT3KBJNN9jT2HwPLZim1
uBCihREJGBaNavUEYYenbijJXfUgRJX2+Y+LuElDCkykoUfVlHkRTxLxzC/h5ToQ0nUx+pGHNrpi
9+SOyFkKa67Oc/bqgX4MPiOGgOqfqDQxLgPGkbV93ETb1hVITM/IjKccsiMvNV/ENv8o5pwMmjeA
Tvr/vgyG2xbaWqttl8i92e5tJqe/P/GLMFzbnrPvJnz41utGBH/uFGuuxdQFYzIJte4cx118MHOy
zVF8tSQOkaR2XkFMuK3p70AvhMhdEJ+zd89mj8Lp9lKi1ZtHf6ucW8wO9OfKx4Jot6zL5ucKR/6H
lD9WaxywkvYfYzyGlhYKO0BSIrM52WOrCSTwoeNGUpXI9ciO5Q3USicWZbsga44rrHdhvBbmwQ4R
SW7YKaaPTukUfODebKiBmUF/LbMeBiqfECtc+fiNgr+SJeEfyV4nrQDolir1J7XR93YZVadOYe8y
ONbRctib3X1jnJzkwLpyDVT9WZ8mntPYzCTRkKXi7me3tZvy6unIW+RqugCbBWmQ0xdyBvxzsVko
LSOUMfrOy9exszFvnkueMpqTu0px3tYiHckZf2bK/mC7J92i7oQlWcP+ttxGjscPQ1qg29YcStB2
uhz+hRQK+eyf48BqvHlbLYvHwIV+1wIAUh4i9922zwQVF0PVziTMKNoryZdDuKQiQkZOxaflG97g
Qn2inx6g2LD4SSJGLfUUaYcztcQ7retu4q8JXvEzNg9pNTWYsD7kWR54t7x6v9DKEm9Xq3bNLbme
Kt1HS+ErWQx41HjwaGhwFMjBZFCGWdQ0hL3PCiEkKOzIRMCUeMckb3TJqVuYPdKvOHy8VfqfXiEA
JM1x70cYY+/AjbJ8851wziFefWkpbpSmTIAd6JIx4k0/eOVgCLIPxrkDk6lI+wPnf8MBx4bPxRyo
x8BTWhUuqZ+FulJX+Zx4QUjkfS/GR4+NXu14CKGZTKq3CaN/5CW5XlgyFBIbeXMCWzyt69o5nXpm
UaEtPzQ7ujM3/MvXn2U3TRR1FGvtU80ncRggisdtbNEXcTytZhhGH9oMzkk1Vl/jZ+ACRlN2bDkM
+hlCI8IxDrHEaeSbS1yjJBaZx69nAfkQVWSpyrWxd/AMrt31SYgSxOPbwmTK74Rm2spjZT2SBBQJ
rJ/V4YokXxfMtNz9cmrhTpknrVxdRnffDrnuSTiT5OcPRbTNaRiK8dWPU6NH307q8k2RwUCo9JRK
ipoiuKh1VFQjc5RKfx/45gQpwkV+pi0o4bHfa3BzI6FAHfvg1RVm3WbbMdaqbcl0hrwgQ0tfjIRe
IhrFMpJuKp4hq/OKjFWqcrxcvBPVnLbO9a/+0It4TxHOgDrFNiv7Dgg5/GLAPzzhu1mynTavdOYi
vrghnTN7bMuJUzdJHxt7JNh7w0GpS6I2nIkR+XdY2ra/PfDQMJLQzBYj4lmHtPjRKOsXKgNB7ctF
1XS03qVu6xbgOd/gT/eVGUrtne36ZMPFV+wZUp+HJ09FGR5HiOwiso9rAtjDMKs+Bml+R2ivx8Vl
gdBGNIuKbcjn6OUJZXu+SkzB7HSnYiLiTTxiEa8yYpFfDvscyXJBkGeqlsV5L1sTANHeLvN4STfc
6/hNHUHmOf9FhTOiIdZ6BfobdMwE4YOhQura4zNWiXAFeqBevWw4x5KMRSY2APDwnHA6LJndbuH3
+T/p2q7dVECBlyrECn29otQ16H64Jox692c4tkaayR/HGZmGB1oenDxZnCzqdh8Dz+CLR2CDz8GT
v94EMNd4k/ArEAztSUtFYSEFFK63usJbFBLCMmR9KgjkOIDMWqoS8hVL4IAAWA47PD3fhgXNpTwt
F2l61ggeW4kpPc/SH//4FlTsZClcYol+Cw6kZNq9bDMpQlqJ2/4fViVgDxIukshHYY7smgnj+oU/
mwPxRUdo+b3Vqiyr+0wUOaFtxY23mirIE9eZzbB64T+OCXFaqHuSKAfm5gU3iGGEr6R32nvyV1Rn
7iULtJY6ywpbPHEFeOmRoNjZHhGSf4pbIH//a/92+dpZvj9jW68+UWYR11hlI21X9v6o0dAJ966p
/zD1WB++iuF6sUyWWCw3Bn0saT/3Xt0dusjDMwMMr+WpicZOndtV5R0gy6ZkKjrWxVcE8Bf1wAEZ
PlW3AD51GRaN94h71m4aNRWkVZ8PI8xKsaO6KSsx+T80A7l9ZXQHfAzH0GhZydASEvu/sJjsIrBi
l49leqdsG7APHwel0fJcxdlS+Thz271h72iIYZWPSfa48ia6vQtVTTMLvq5o2f+c2ZfT/eFnSmHn
ongolabOCCKRKppka6vHv7o5HRCi2p1Qooi+kQSlHUmpe9ampGm9XZ6tdqFUCrSyn72AstqD+n7H
yLuVZKQAnBUIN6X1bKLaP6XodjI/i+0CNm4UzZa1PC1j4/+hHSEP+VcHCVYTYBs+9msWBGYm9Enp
2qWHRi7DcqaLsZDg8k851moPQnutBUpdbcTaRyVM0aYjwOmtOB1VetQ9+C17an2ioF/TjliGc1CK
Y7I1arLGZKVl7/lLnyuFDGVkb9JOJkMpGRrWGlvh7rfGIHjq+HcFnl7Gm0WAGsCoAphT6+LoTY18
dP0uOpn+DdB0miLCwTAZmVWc/q4F7Edpi82eRvnkXi20dH9/FQaljIZhN3WZJG3ZAgamnMQ/Y/+F
+k674bgjG1/mShp/IR3N0lcr+BMiawcJyRExLIoZ56J5l6MHKxOYLzxKbNI8PDB7ZRdfk5g7TOfW
bbqBcGPIMiR/Apq+zTUyfpFujw18dY79TR0yRl/YgoUVaBgeyHJYEOFslz4yu8+4SYagTzrql3hu
/vbFUgh+WICO3oOOBTt799YjJJKsWI3bPXhtxDWPW0Bk7ep7EXk0d/mUKqkgGMQ1S8szHtkjV7b/
gAR/+cLvcwpbF+NsLd4rVYmmz1x0RTuHPIWNa4zV/1pGEg2fIY0u4BGtD8SA4kV61OOr5AE6YM+2
QVn+KT+RwISe8WWWIVYApdpTZcZwEaAHnO+ygD/U69kVkYKingCMhVRogfDCT8drEkY+xYpsnVjt
LSxKCz2LjLaoQCqpiPbShmQXUprzf6eGO6GBXpejzMP/GgiD3S+lL88JnHfw26lcBIqtpZJPeWu7
sBoMbYyq8FIvpUdeV5I6h0Gfew9DVO802iEnOq2Kzk0AaSllEhAf9v4AKk7JlYs6XAJJZo1BnO9D
JzjVXDcaVJVOA1LuRHO3Jj4Xv3k1CLk4GtDqM1pPsZdKqTMn78BnHTaF3jTmiLc/2j8YLLPNok7b
vNuOzy7ab+WUaQdtmWIRgE/eP2UhCCWrSiIGdTrIMjRoJLOLdHffdKAJLTyHvk201cnQNIwzckfx
1DpjP3B7NVjD8kwTYdY4NRHTMSJzfEeHrtg+aClBc4OZuRJwZKpBBYeEFYa3Ag0C9j8sdDffbt+u
8F04pyeOeBrGAHEP5JxWYNR7vsSMwiI85esxt8jLOX5bZDELZH17r324/hp0Abd3cl40R1tbtYI+
A/SfXk+2l8sLmXF7EZWdYQ8rg2X9NyA5G95qxMHgJiRYuBVL27xA1OkLZ1t4IpyrpDOsc2qe3Ebi
ABSr8+bvd9tlryTDqog+3b8Jzjj7OE5lK9YTXeeOZiOx68wr44W1aINRRz9d0tPkIoi7DCP50M0m
1m4idkFGlh4//2U2E6YNYIGjS0NZXGo+itjMsqLQULyLwGBzoZ8Rz36F2rnA7S0bH2Eap+o0cigX
I9EhlFufnPJo0eCGG6xRK+8mAinAqT4/9isKAEDE3NWBJv/w3GGNeXI6BYVr4zP/h9W8hLc8sN5R
K8tF9Q3T51Kg5dcocf/xtUOiCClV0/FKERa0yRONR+xyTotDdigJpZ/1A28Hg4ytqZAt3Yk/zB97
tJPj8o80UbxXrnVSH3jSBTkHWpg+WVcj93Qr79BCEndI9oB5n65MtU9DqtgPD5VBZmqodtFs/hUy
of0jLPXmEi94VqDstZxdOQ0oIshLH+c0Pu2ChIwztf2YFfRNJByrZOHjP4ftMP9heBG6Y14DDurJ
0Rk0ZfMuhTY/bSTPoSmpaCeatFJyR+n22FXPoMlj6iUStHNOKMI6pcv4o2sNPhQHnwtRBYDUKB5f
wgpPwg7qfyve6m78KIfe5fzprM73GqqK5tY0IG0/k4BTle7NeJdhA1zPvqsP06OyhmxgOrFEBggC
Gyij1BCAyQD1cHO1fxOpsVYTzimTIvKhedwdTWaBLgxDhM5ex6Ytd7VAdigzQBZwYz0+TD9x2vRg
sJRcGz11Gxe59OTWwxQz/xDPBYldFwjJqkDRLLQAXcSlu1J4pLAxst3a4P9GLhTtjeRCUziHF6+Z
322ER0RE4SGXaiVlYgWxZdM6hjSQyYFP4UrLb/TbX8E117A+q+gmvepvHTFh/qFRW5Cy3W8+kpYd
Bg1CX4529KBHEoOHJ7/9AGD80tL+Ek3Z/Tu0sCjol9zAfRh5fkF64Js9R1aP5t99d6vUAQ1udnmG
wCVzHWz5PPKyOWFl8/haeTfRtmEBZ4F+oHdlVkTj5j7H0ywTGW94iiMGUtEC93Np3txiTmAj/3ii
4twVpd4eArr14lXpdLagtxHM3Ywpi6gpPXKxVUMuiL1uIC5hjV+6U9dqOKwR7oBpb6A4vylAFGp8
nDQ1NrenpatOicG5kTl/hXJQGu+sbC7P++KD23OVWKtS67sK6ixqsHBmppEun6V3Q7qI3CY57AMl
ZlqzXGWTEsCj68BnO3peSk+ZK5RW7+Y3eDcp/kJFP51bfu3tpHmNz5Ti6GQfQkfBu/PAjEv72xpK
/OAD8NMZdb8pvMdIpReMSkd68waU+q3CYUPzyXo+hC8IRjdXwsx05joCy0sCk47xeIXP5gafy31P
rnC0AqIguG61pwCjyBN47+XTHRb66J1wa+bRq2jNJPvPlGt1oxqucnidbYr6gdiFMcEsdHNPBdPc
ZfIUaQbSDnrHqWhstHWhAmEUHR2nlMoXZYJjyM22buMRpjwTVZKtkaaUSjCoG9kN6+MkefRtIsO/
ADTPed6/3FbEtWGHT//TQ+TAixyNqm27dL5RvcpbLjcuLsJzJRxUU4qNkhCLBbtFNC9bHmTyf1Fs
pyCIoaBJucLWwy45u1PN2wJCwB2CzM2rXxLGnSWty8e0QbtLCyK1uNgBdYoVyI5hQXDE8bp9JFry
SlReOIksVExb2rMhkh8dL8oLuEZtIIZ/63gpNgzVx945AGOOBt798wGI8Jba5CSTL20vB78A5mjR
eS3st38As6TbYqzs2KeZgD0L/Z8MnGqjFY5pQPNukg7Kr11htmBHx/6jYI0iQEvCozHCEcn0CzOY
mNEPnZEe99EKCYlm8wy9+XbihkzG07BWfvCMbhKSEaYG2DKQPD0HxkZcmTmwiOVNJAlJj8FFr1oa
g8GuCgmViGwNWq8fj0RZYsuMXyyqdL6ovB2DOkgFZgK7/AXlAo/zC9V2bldm0dJcI5DzzziM6Cc8
6ZjOlwY+B+fOqZLenWc96oJ2/K6IIkyIUaiWVgzzHOvuKV3qynsnIYEgs+1KIOhvoLJlrd8aDeof
Hz7cxiTcRU9QdJN9ZiJD3g5fXi5jfIw6JaVtsFewZ9/8zyrmzRaMj7lxR1cNkZIzOJUjpmnQ6yyL
zN1gKN2mz2TDmJdesSOIRwDIf2q9YKYQpStSYBE77ycXVzmrDK18ST63CZLdzLzgSAzgfyiipMMO
dqrueORjknCW5epED3bIESS5YEu6UXO7zvw+1PBBA9kx6vZH31lfgJtapGjaYoXtxiZe+omPL//i
Hd6K9iyqUI//2g2ERg2Q/+YxUjJgYFgbX8sJuxROpM/4cqFmIkM//G/VoaQZqqcRTJ5Pnzp2DpaE
qogoDNolj2L7yxbA/IWk2rg7avhYa6mYsbM2nOMbqYl2n8MtUANhnOxgkV2P3/GpFpHtLCpdcKRb
piVAkPeJTHOyQzo1yo0PG15IuhsPIwBacpeJ3FF3D/ToDZfvPhbwqarphNhxyCXCcVmZ9GThkj1g
0DaBpW0lK0N9fDNd/IAsQw2lNQZWvTmYiZ5oYb7fKZJPaz51cd3wvKjAiTOwvDQzPyJM4fq5wIwz
fF4Xw8GJaqatZ6J8kC483TtsOrDBIW7bsJS64+Vj62FjiXixC2C40ZfYSWTBcd6rJbziPqtVuTrS
ecpLiOq5bwQ2VrgA46HKNcq3qoB1NkDpizZCsZxh01NpIZySkTaD1Ssn4tHWCE3HPJzhIoIifT6z
/LwXih5zdNwLhpRu1G7a5ZjWegkWIWoQPJxXqVe7a6MdL1nrBbJ9HLzz24+t/C/6Uw2XaLcGqNxl
DZS8VqstZr6aZi+OYQuUblB23iYhDcOS/3NDn04D1AMInSAQ4qJekAZlVEtwKfgPAQS5ADcq0ovA
yTk+NcVYmZIhuzYBR448cpR5I5LOa1XxF49FRALyBVuJhsAgo/8pmK8nGo+B0lPS2dfUdJJ6VcGH
q3Y/f62kAkUYHUzLJATT/NF+JhnrV1tsUyIs/poRfSZcQPAE42FZPC10M29F5VDn9NHzYGoa9Wl7
8+Z+J3Xn/0A49oR2/U/Ndk+9XJisjCAWP98ekIcv/dAPkFPj2sm/r6T3oEnr5BQwXLX+tD8LQbcx
pBVYLHE6cyU6gJA5G0jUIYIIS9mCgIEc8XSFywAS2JYX73fwpHtRCyw2NRPDppG04gOYqWF3Ds4z
jJAbFcSaj3xUPSGps6I/kLJBIRqP1gU0fyESYc1tDXxbq/oFQtqvVeeUU3RpvliKBpci9DfbkrfM
5RKu19AKPLXc3Kyr8OwLzafIc5itd5VF8XUrhhBfJILzAquZprFXYmmew8alybJw5vdDY8dXLwBV
ikiDA1lyF6B3zGUcO+1qh/9pe0zolkJpgG9bbJXV7amuhZY270OJ7DPgkymnkf4DP4T8pA0AuYgh
Qj2LRVU+t9aRsonJgEYH9WhkOqB4a2PbKO6kjK7ZmElCq+s8BIx/22LBkWEwq4KY1P8rF9i9gXm7
9+ZjnlqWlvaR1TzqL6nRFYjt24+KuAcgI1so1wRe8wkc6DtB4+3tbYbNDuXxV3qgbawZxDqSyq+C
xdL1gZIVhyrpaxh2UNF4ugTzFgYBILskmUy8SwdnKhnmAGPNHJiyWo/SmDq2syz9aWWFLiOws91W
TCPF9ectMpMQeLXQV8S6IG1QvKWLHXxkRGUi+xzY3VNBk/Cd4CzmY4ByoCFSxw41zBXqLjQxVq1f
qvSHxrF5mPNEHDYDRFmUrw92AMivdr5xjGuRZVjOu2xvoJD9u3DiVmaDuUZBsoL15XiCGC7zh7fk
AFcLqApIarsuqJh/rfw8L+YTG6T/aGyvsix4gBaAtAYEJosdktZ5C1nEwUHshoh72cdY2AyvLGLT
sS0Hp+lFHJBEMxSpW8fjeRO7vVuxqHX8xd/6qfXLNtmvVdOLvq7ZB5oM5M/ml/chMJ5kP/+UWdGV
llyJPKKIFccxhRgkSJPtpRAL1HRihbhLsOIqYEJOWOv2ty02aqFMhLW5AL9UVhsfuyKR59lDz+wJ
JsBQD5KZ/87yMcBZFP8gZ1DXAjUTJn6tEf0mYUKhHTOJMoT9BiMo3nh2khWiE7aLGyTKCfo0jbiS
vf8o6tTDSLVWXavjaYn39wfvYXP9QW9M/e1vvCzilDgcPbZeU3kY7eXkockrRrlMN1mzFJPDeCMx
/yp2eJUU+BxFeCDiJosJJD4iAlCouYzt2v2IJDgc+5JW//GRNqXYzP+wjqMqnO/H3ZH1s4bdNXF/
Qwaz9lilWBEgjG7GZj8iNYIgkAq6Y9gUhsgSEJM10RqGObkGzEZQU08+CgD7dLWS6HSDrkdqPHnY
E8PIVFfOmMFeE/YrGYKX5TlilhgT3x9ZMXgZNa+eVvW/JAzdSDaOw9kCb4+PU247sVgLGQteDaAo
C6pJHDebg0y9XUY3Wu/4/eoBzakF/8aZ4LpmelCbmImiNnl1Afzdl86zUEFQAoIg9+YxAo/m8Mjt
RaXG6d/9AvYCoO0ljUgXmqiO4Q8r1GQK7dS/ZayM4v6eBdDA/JsMiEBQFqnxei/0SQzhFoKwJxNU
FjtC6fCzEA6DTC/82Fs+P8H8Xc//1zKDcDYgczyJUHW82QEOtF/+dWQ2Ar3BaERpyCqezBVH0xwg
F4kk/xmZDfuOk+jkGCmGt5ZkkWGmqb99R0eBQiVJJ1ojy6pxteG4E92jSTsSJswEtMQuU0vCSL+Y
g2KZ/T+GGY3op/bU+UbIQhYFuped/6GwRuKfo4ElJNPDNvXix5U7iwqabR3cv6VOF1CBKhKArB5y
q1hkA2aKWm+iMKB9t9SDkJWUimJcFH8MblQq9MJ832NLIq/6/ALSkjcKIFkzWNEb9wJw0SAfHTEe
4Y+yx+fwUOTcl2JAn2gRhkzlBluwAulhiQXvzvQTlrmiMgxkECNHDUq8yMrs4twtv/ZNJa6LMgJg
0mQ/k1qoJsY52WwAn5yvW3+XsuK6G0/tgkfBGp6/ChV1wgx9HtOI8SNhrcGWqS/rrXFsUfK/Bfjs
EggCSwOYHPLjg4mtRX5k6QY0hYFhX+vfA2ZrFlKLdzCM5zQ3m70YN/IcT0vP//uuRyN78JUGzoXo
aoDmJ/p3K2MW3PUt0vbssK9ukwk3qV6CEbZX6maw45lBi1Py1JnUzwFJgdL+ZdkQ9dnkhSP+AtM9
h5Ikd5eIhjPCxFfC8LwnMkrQ+J+WRlhwiNyJhRnSFX1icqxeswDKrK/BHAg4tfFDWwz8VNJ71I3F
SgNaiGCpOgNizBCzYBIeoXtMGmaR0dJH0oz+WHbD7JbDfdG2epzCQFKlu4iP4CRzVqbkDnkKFGWE
u6pBB1gV4ch7Zuoz91Vuu7JwZZN9SzWeKsh7+A+7imDM6z7ktUmEeEkvpS/wVs6jkbiJZ021pE0p
G+9r7yQ7CeObeHF4o7sg+t2xbwVm62C9XZ9r88SjhT68Ao+ZS5GQsvyAi8WzmcrEUADw8r2Pdaqr
GadQ6n2dBHZtCvMU3vjlfACvy8a+AQQ+snP9bZ2ZyBi9JSaknIxMT35XgmAyMIZ1vay4sZ9pX6Qi
yaHxtJBT4T2l1fSNcl6m9mAhFvHTfOqKCFbs3S3TqKbNxURc039GlVP8DE3F51Zl1QqCT5jL4c/k
c2ExLnoFzzBXWr20hdBGWZhedWGpDZZtECgagPsGd/Ri8iq7u5/kZ3sWfzognqBC9UZi1JLkPc8g
t6LTeeGqOpJehIcJJfYQa52sYAqI+Lu0+7i4Afv1ObiNm5Jh8kSjq1OFn46KWyk0jHKF1bj6+3RF
Ian9qQPWH9ROke+MEGqeWn7zAVJIQ64uutjTG6kCsq9J1HReGG7kx8yBlClyeda4ddAwfHa74dkV
smq3tHiuBp3yBWJb5lHG3+BjFPa9hh9E8fZngvhnKdpq4/i5OIY+sr9dbDMioSFmcY3jcRpqD9Zd
rN7y+cKk2pR6kwud/5mlaMdrvUWEiZxZ3pmSowKTgyjOZ/mhUwFZ+zGNQYXQLVNrbWz23i6Npr9B
iWUtUI7DMxiLZrpp40JiUqvPP5YokqM7PzG70rJjEaZiw17cdI/bR0FMS1IK661nzdh4C8xQOkAV
zWBkdLXapkKC1GatL81HhxXn3BRqVhhsJHGXC3dXqTBjr/8Bjse1fnbFyMSLuH+9+mt7nFXgjk92
XqMC648uJeNsKUMJtEUvX+LxlT5IvjxG9613dKy7ZK+T0ips13Stf6gnJLGjHnD/12d4bYLTH1T+
cAnehRBerCm+/f0OmCGsL7kNpleYJY5+KaW1S+xEurkUqcv9oN0P4qBEjxu8F+EKSNRg2k2dL5bs
kBAyiTxXH5K7k5FwdBF0CUp+SrUBJRPvGlI6RWKdUO/GWGDMS5VjSOvOQt+mEhhy2Pd3ludJPdOq
JxvbACcfGGq3N6HrQKNJNy9pD44OmIPH0InTOcv2GL9mvjbjBc8SjH/H2lTLNmTpXx9fU5A4VGxM
WJelM6wcM2SQwzXl/xvEPm5hXqpXDtk1br/wSmAFvtpQXTdvK/oFYMv3AM2MfsizpHpsFVuI0+pi
xqQgadTteMpL2jYEBf/hzv67Df9UGcmTpSiYkcJlX50weHevlaDNmMGNEncvfeE80JYMQEUhRkx6
HAozuc3tlQdTDsEk8sUJIqB59xD5pxz5B3pkhpVe0QMh5i842oAf28zGZC0AuNLDhD8/t4zwJr26
6SPAlwOWOw9rcmXwqHd8Ha2tiUTdJW0A8897ovU2e3q2GSnrhG+7NMF+QGzT4mruCiokXtCv7/Zi
eYZW83/obrpWpG6/Hwb3fyNyDLy7P/4sT83y7N1+JfvuB5r4HkUyIIu8CP06eKjUzjD94N8DjKsT
8PQ8f3vVLRXzrfXk5QKNyX3dvioCeKBzPFwobPirjLujsAhlIHTVdhlVIRAeelDm8Tp1NqsOu75Q
HcvxDdUSfLD6+z90phcgEPOgROfJWdY+t862GcpaOtbjQpWxCJjooSr8hVFhbApBRBGhJuPcBBzr
FFHHcnWlLWRMBDxMBQJDK76ckoJNhLQpq63LPKCCEyiOaH+mCGaTAVxCGoP4fzKCV62ZzR9JwdOz
ZBwLk9Twm8KbBZOOShOrDOVFl+aN3LJZBw1eyrdgjoncxcqKbhndJAfi9Mwp136ANsx9yc+1Zv5A
wmWHmg0lOwgQ9tSoTxlyffTF3Q+dPms2tIOurFxmd2ApFAytZBhs2eSEqXWPnTh/fhfY2Pu/8nxY
CQLncdLRqwDa2hH2/nE0L1XKMlWW03319qKMwcDaGLPt1/03RC6ULu1eyjsl+A+F9KpVbEQtKi8K
phYLQPCXJGDGjWM0jXUGW7PK5eQV6ty+EpxJhZhJtVV+jfMRW9R9ze2VhZavZ3p3bLcnVjOtOfsx
5ocKq/S67rQUpjMCvkalGV5s6nsAwNx5NJSOWY56Iz+OdG4naIeCYLLiVtFZYlvQbQPmH5kGYmLu
FZjr1AfwVgpfwDalohloiX2IHokhzgQal1tDxBEtMvtcxllziBoqOMJFT7yXsWfpb6EdO3p6bNK/
RDowAbtWhyDB95AqHDZCp/Gf3toiKRvIsmdsLDxmMqzE25uk9nCD9NrCyaTC4ZIdvclpwXNwtkkd
eTYFojo5b+PPzEntYqGgMCpmzIWq9WNJjbgMlkhFK/U6CCYZlo5Gpg97IJTry13qIK9+2OE3Ol/U
GvRxakEXHg9s1bRcVo1SnNUnA2+0NQt9CeLysgwSrb6bSmXP5iIT3c4hJPXFoyenoGtxnCVJzml7
6gejDjKz1/16JMIMKM4rRXLSDNr4CyEQ/doavnyNCGOz//lhQ9dbtPyiJ/d6To0aq2X+7CWmqYuW
d7vIlZOF2KTvUgsxvyf+WB6RHdUbogu05mW1a0/OfTnews8ShKLhziOqV9ll9qx1o9MIQjlXdzjG
PtxxuseVnRdywLhJ5vKdk6SNQ1AEWWP4X/Bm3OKIYEudZrO8qIE2WCa6eOwzRg3ZPr/puFzsV8K7
TEOq0RHaWB9V+jSvBFKEZmnvu/PRu5YFMuTGpubWqvALsiM0UIwbPWmEmbXm/zHMMQbjLNWD6Ch1
UQwMtt/v5YJfotTbxn2kStiuCy5dPTHhmP1ALXVuKIkHfY/hv3dB/4IwA1b/kmqdAtZIHnRAch51
aB+mBQOA6DW94o2nix9FDcsf/EluU+iO79QLqSGZFwGeqyDhsieSVImW15Iuo36WRFEFNQawSS+A
qypNfdABB6DOgijVZAV+mgWFEMtcCG6tXKYF/uCXVjob3MuKCRpeqk2B4+u8q1jWExCcrT9JNZyC
a2wRf4vHjLRmrx7VwPzGo9M7xL/DWx8cnw1ga6L6Ys9briqxmQmD9fZBpddJ8gQ+6Fe3+K4Sf1a2
A0hAWtqC6wFzD8CPV9H45tcu6+AX23K+TyFLJzyuf2nwA4rcj0M8suv4lszW/00Rx6UjayqTbEF3
1EEtjyC7dP9FgQ966YVwNVG0PDW9D5Ge9C+W/mpB5g5wZZZ2W7SdQG4VAPYg3wzzPnTW1dUuEw/p
/C3C4sF3LsJ++zJW/8q1Hqcfd8UyGvDRSXQA3ZsQ/9dMwhJSPg9Vll3YeTOhUYKO8IjoT+h8tl1H
3j8qcXf2MnPIDauGnsy6I3yK+IIw057lKwtiYQYOqPPz7PK5X/eMgecryMNFTxWZJ27Ort3HZALC
O8aGBc5dtqUTcjMIHvbdjWl94EZqBzAfgGBGsObT2spZqpS2FdGObhgjcJ62ZRTyjnRL1k55S7Kt
SJ/lVUKKsmcTIQou7pGc0RW+bO3LPE7fj8CisqhiKJ4eb5oOEtTn0PAGd1NOK5oluHOKjGGuiqQW
+6JyleAF8rqKV70CeYXpsPYSInFk741dlpKsIXyc/Fo5ky5TCDP7tPTa3qZvAhU3M//++SzQ2IV4
9aLgJiV7JK5yKBDOEBegPq1Gy+bvOj20/tFokjGzvp1LPLfuzzFP9jZeG4ALbOhnS7iT1UNEDQel
D2zZA8IFeIfW6YL7cG1gdPsqVoJayrvxqskl4UzO0t1iVAohxjlg9nIBGJQLhlbwHVHzaEvv4Djr
jrPo1IbT0GakxYiOh4A6dKmoL3QONUuwxKOZdrqmlTAvxocqgsguP8MAsBJESuPLjKRebHLr4Sbb
bAPdiLyaCKygIBzcZaM8u2aR4kQnR8nBRovurT+h1eY7OeqHQ1AxWWkG/C4UoeD5KwpqQf3RVtuG
Dq9Hw3+F5O8o/MCc0GrXIyTJQ//n57LgyGi4th2N96UGQL1MhcJ0io8OaBWOpwk6qxI7fmlG0Olm
oWikm5mXGX/ThUkmy3D9MDF+EQxZyCcU53MP/0pK3SWNJji1j7YdQEh9GNF8X9hvBpmnNLyr7dAw
aoMVRUmK9FNQAO4PtB0c6CfY3runlTnvErBzxNboQZFA3ijVv94eySgTNhDIPIOpWi781acsz+YO
GjAmEOM/UZLmb8nCduI7uVZ68GHeThhfyLES0AlMAMRgI6X7pnLVZ0E37Ei8fCTrMkxuvWEWvwQI
caEE+iqdJQKUxJH/j98vsQibGBiXImuLXfn/3qlrkUF+ECaEE36JA2l/aKr/wRslIAzP74tx1DxS
FYY6k0FGGYOGtk+dhG75MM0qNLNN3GceVfHsMqrA4qKwAWV98J9S0NLXRy6xD81UkB0LQGN1ftX7
BeyYeazXg7reO/kWrDK1bRDETlQ6uRWwD+JmqXo43cvdLZpKJPLAOPEVJZ3Jg1LlKnPU1vP7dt/k
EeTAwGth5i1bXYiTfH5wuog8ejyXp/hM2Md4ZSpuOj60rhWKw2oOeQIlsQNUF+N0HWmQUfTDXFVz
3MERQV5gphSygxmyZiZBmAOzLn88+va+JBGkzTYfV+T2QXFTmtfIUnlkXrqw7c5CExAw6NE7oKni
yDREjTplyNkdWLoNxKR+FNA/4Ch1iVknLuyKsDGKo7oCHGX8Y0w8bmqYmOXzGerPJW7KsslqwPmG
TvyN+RWJeSV/8vZr1z6bAdjWBktTAH0AwbkAVN2KECr/pehQl5xFWgo7zEroDn7c0oiTlikvQPRW
g8PteWoUEOwafsRDN5WXRLbgXHcS2LCrazTg87u5k7VycVD3TE8z6XgnIH6UXgU96h5gMzCBJpAm
QQYadMko2b/9dk04rwWdR0+Ha9bSpigmmiPl6eM8JqaeW7SGlxr9uwK48Lv44bUn2NVt20jJPJlR
WuSkFxL9mDd9lGkWKAuElp9EsV0priSjiX7C5z04oNB3neWJHMQxD3/bb7bt4l2CJXm4+8lyt2HN
6ZRACIprPCwZHxIlrpOB98kbKxKzGHwF96wNWw+hP3K24bh7HGrbqlM5tm45IHyC66vHUWrnE0WQ
vJrrEhZVvyUv00EE4s1syGi0RHQqcy3JYvFpwZUcoxYZA86SfCI3HgxVEO/MxpxRHXS5WVQ6j40K
+h/yYSD5LLSBxqlv+Riz8O3fDnYODrD4HrjF9xw8Y0utV3lkS1aLRcXnVBDLHrGgP2cdstgL4CDQ
l24Vr/RK+KizwlyHvi0dWy/EXHGHZLyhlYJpZd7x/AqFB5IsenT+GN1w9gwX4by5RjApMbxMREsu
MtLIyXQAXSi29P1ty+xPdpkqCDMZcrzuoWjCm8+lL1CHSbsnMmr+uI1Ma1dvO5SW6aRFgum7eEVM
4tNMoKorgePYabRMLMOWbWWRf1Rhkb9aPHyo/uQui1SKX3yDPOulLdqRp2Naf1/WgGbhfrcbQXFE
6MnjTxUD51pK5dD/0hX1NZuNTBrEp6pDhXUkeP3FT9+Ac/xjs/htjvZPakRiEDawLnDlaRurgZbD
HrjKlEnlQ0mN87uBiwV9LIAaUsNnMNWyVZEn8LIMWYTQzDBxkDz57qsG3RSkyNq+ytXEQ47vxtEb
EvWiwlVtj/XYArrx2AGWLJTfN9BtMAtOEz+Sv2Jl4jEdECAxjjVPrx6o0X4uWBYXNonwzy32y5Kh
tCUQFFYeWwl428zDBgsDyoVSO3iswzgr8q3mpd/1y5NsRGF7cUtaC14v3L2tGR08GGiUUlaTofzg
lT+1kMURJb6W5ii2aCxnZWRR7Dqf++QuDHQs55LVkyqaLDXbolJZCBEgtsveclXx0hH2lJLRByAa
778nDi3/nHcs+gUwdp0fmtMZ/k9Kj+QzV8UEt6/Ebyual9Gbf3hXtjXc53t9EcTAxh3i0JXBR4+4
+MrvY7CttB9NurNZ9YbRyYDTz+2oK25WriGYP3QZhkvnEqgCBkkzGhTTFJwR+FjDM0goigOdTVx3
lhwylxYeSb1QvdreRN664yx7WG7WMNYZoJ2utKbTkNK6BFUdtivz5L0pAEeLXBdMjup+coW/zL6X
IJSk9c9UhI/UrXKlexk0Yu55thQviH08HaSX1uVMz6ycNSOh3XnQbNd5+Ofdnz1/ZLqcd5NgiMgo
CrLkh04kZKPHQFhwzfRpVTp4uJzy5jTbSUo//UekSzQZZEv9y6E9LnQgKSgxE+W0MhvzXMxwEiAv
JQTynme/6jQ0CbWGk6BVftyOX9moKtxhfolNXxKEfm7VU8KdrRsaHOBKeRytmNZyGacrhE60bG8h
ujLTxbsZp8M0aIJtrhYxLnT4jV+3OVEun0/8oRU/0eR+yI69gXsWvmvSepwlPWUw6FtKlKUvVW3l
lkXT7683plx3dV8aOOQ7HRnKjfMaEtFB31REGbo0a1+1KhWyrOE0ymqg/l/Wmq+pHgt7Hanhjv8F
KYO9qXiopG2TE/AsTJhl9zwnbC/LWLu33xo2QhX+7gm7D5L8qdH/mgJKoFqwErls9RJ2kpUtr/Rc
+RY/ME71lF5fDBd631yACfe5d1jdhfssRMbyGPOwyUf0qM7z+hKT2MoNpQKmBxF0GiISe5RLrJH/
COOhMA7KbeLjkpAwL9v9J+g/0idI9YmTougYBzKQVHbVFCAEXMlXXUIaGSuvTNArCqQXm61g6Uf4
ee/LO375MsjzbAS5xbKn3rn24uscNfCMm3850kFloRpWIcyBjJFpVJCyYnegENm+esBs9olnk0m0
QPbMRTEOF6JQGbjpqGoIh6TeJJg/7Ymt0wgUgaSms9qw/v+4bRBBQ1fSUiycbLsNbv68zFrnMQxJ
hh3GGQxxAB5s0ebESbBZMXPBT6ni2gM0h90W/cJ7005fDuq5zxPeZ2+Hsbdcvrj3+eB9GMlSkGn+
n2lxjn94xGIveL0V3PzE2OKc7d/ynOJsLC/x8zKkcJ6VYZptBitJZ8wswuSERflLa8uKhxeU9w1i
2809ZsjMMKQuefx3sq4JLtBLHpEg7DdZVGyy24JAbL6sWiXBTU9VO8zm0JW6EeZc4bLqjcp/TXZs
8VyxR1r77m2c1xUxtcIgsKEeiX87r2m3sSnfnwpe+qtxWJ4MGUjYAZIM4l5fdPas9kFMtu8nuK6n
C2fACvZKknMcztPy9+5nWrhmcJQ5VMvPQME9qBz2mz+LZXLVCC9z5HOi2uY64xlVvYZWv/12qzIH
pGwPHd0xTXBpdQkc9HnIjjgXe9UaEafqSucgB9GCQ1hfl1nBFmBET6almZaACOymjcURG6eJ58Qq
xyZiPvp7FINurjIEOMHBzx0omz4ewH0pvNOzLtgtxVn4abfjiVLUQ8+MxutQ1r3YyatVqiyZ7f41
wVOMhFeKaFztkkejnogKFZcD6DWg6qA2D2O41CYrIMhocuETYqjQgARkzF8Ec0fyWLWmm34AO3zD
hT91eveIZXMNmOF3khpBxkmiGzbsXU7pRmNUH6Y7+0IgP9x56xDNntP9KnkijdgIlFPZ2jZxgh/w
xr9nIDcKYm/Rs4THVdInQnNK8cxGSbjLHHSnRNilCg/zgCgt1lLiURZjRAK0SmKRd9Xyrxtz9nAV
hywu6Nzny+zbDpyyYmjJDuiqgIeEtOVqSxQ3bf7e3W6Vq+b8r4O7cjkFThxGieOe4jFGX4nIdUoC
INwCPbaTCj2Ms4OgoSx0moX2T9wzWxmAhDthTvF5ZIHH3edSJX8lv65axy5mXm8Ft0OiDm2A6wo/
ABkM0HYJrxcMOdsSQv4MB14cK/uP3BemdktFesloP3Xi624ADsuuheufkXdTLlDxPoHJBsFlnr2H
CyCTlwVu17FkNTNZqaPMoXqYJvopWvN51TtNoWeJgqHtnbAWrCPXdXYH9+ManpEHD3ptR+3T4zxr
XF8kuRwKim3rJ56HWk5kjAc7ITYzx1FGXGG5pLJofnFUxRDJ+azPK3ZRyCsog9bbDfvIhf8iiiGU
Rz+XgNrQzjf/aQk+jah1tk8nXvBLZUhboDO/4CDd1QlU6ZCRwpNHGyNkSZBhzxb+RJwtKuHPRGhR
wOdKWa+V5m60gatOPQ6Kc39hFPIPx0MfCKMWGtFAL7ppy32S5hGS2pAMETUy/ruCnA5qsUXZX+UN
f2mKAT4yQZPsLijyuaXgXNw+f2HhvpkgLiPl1e6G5WSeEh9npFtG2c1j5RZ/f9FfUd2Dje6gzK+1
pMeltzVscMe1nBe2xpfwWMt871Y96q5mV6kA+MlD4Lfga+N/DtKV3+W3OntZlM9Lm3Q6mpJZ4+H8
wGWoZhfHUdrD80QXgPEu0i+MZKa/G/bfqATi70D8pavv8hbHKktsylHr7tXhADsAecmVVpk+7Ufh
0qqLYcDjY+CqbwZQg4FDefEPdQjE5YfV1FMQHxxVsg/sXoQQ0uWGw3ilPnOftkfx3cOUdQR6RzHs
pWT70WMtfI2f05RmYtdenhay7ziK1aOiMQiKtThAfPs+XStavLDg37R6R7ztSPAubHxhhTGCDBxl
JHtykkl8AwXcQCOi2GYinEj61jy8jxexacFBHTSSM1Q1q2SGDXL9rmSmw5LIgJW+BcDEuNTY/vJ6
6awl9Ae8zqQ3YDXGCjY8BBag1391urEzyxr5qA6kjZH2sNlvXPVPDR02ZNKmhN7Gzp8zkTjjnSbl
6sYTKIk9RXPqQ/3oqmJmnKd331FPa/EuX3+h3l5i+XCKVY7AtiMZ9+h04BiVXVgGMVR9rOVySjrG
GNWQg1oR2q5lwpiEmt+6jlnbUCNp6sqIksEPvHXEAEIGNZa6XSBxhEGjg80bz7/aN3oyOrshVnGk
HhRlhAdHz2z6Hz/t9beioJ4kCE15ghqe5GRrL1FSsrhKolOvoOfgyi5PzyMLVvo99T6JtEXr+EgK
3O3rRZoTTdxI+NvcplH2w4mWSnXsE5ws+W6Ob00Ysn8SAvC4tVTlyegPIVWvIghAv7iHnNdRpcGZ
syGm2WcB4AsCfV3+qRCQHZNyRzhHr9Y0Nzmwpe2j+Ro4jrrF0NaMiWT10Uuh1LNQSp532ZuPs+wk
SDp66GR/jL0U0TlVG221bEDZ7QFWUoYV8ZdvVbXcciH5kRBeh9ZPd5YU9dyaYnP0Mku55Ax5Ndf3
GYmcdgTI4hJuuvD8gddNtwLp7miztm9nmjWqSKj1cjsJrS/jYsfLvePISGze8ZaIQKFVYEmKbr/y
Puq//g2mIekdgJT59B1gdXvrNuTCmnkxMo03knAOTCNnhPAmPSNs7eaMsWpaGmW2FBtgtBQkQVZu
7X4ZYFCaqQGqybo9DsPEdIdbDTqXYjlXvnaqh5vNHKxWZy3Caql/ZVWX25W8lnnh+x4PWXCMqGEM
+UzE7Wi0lEkL/+z/1ffpXgVdovHs5OKsHtcHIRs3GAo63pNAj2pL8rgnBBiutJPJpP4SGKpyJyAB
i6ypAFtzJZnQ2/grDS2XiV1/ZKWGUyz7IWvV1D27Jb0lM3EfPBFj3yGeSQUBibnycxeXhjDJ+q2u
lA/4obIHejNs16BeI4DRzURVCFR5WtxXTVmy+uLVh0fFjbVkOUQUSViKuclWngMfiShM71eOpPJE
Bo99j4IqN9PHM+2FRsr1miHMme6M/MfaYm6DvDazFC2UbaTa7OD1/2XyrvB2poO68ZMBmPLAXbp3
NcMhCIuOo9HpALaJWMorNGMPIshlIUQuyTX8cL2he/moghvADW8su4PCQW6DNQJsynNN2xlCIG16
RPYhnfXfmL1XN7kR9ElD3neG2QYpzeZse2mzOI9EnjTbkY5I4Vons9zwq6666JiDtxn3ckJThRIH
vali8W334GCDRhlybrmngZrU6t700Q9lc7GpAnNKG3d3jWcfXoEHMFY/zcwr4Ihk5ByxcsWsMFws
leeY6BkZCjj76MnXV8aX9mw56nDFf1oizEhKXgjGRAUeY3boYZYgwR4Z9LghSasdvQRZqNLZbMSm
H87PhNq8vGVazK6zFWCeaDxIYvwWntKSdi18uZy1zDoCRhFHiGsXMSPRZtD6iOf+4p5Y2eozPXoG
Uuq468mxcra/lMyhVjc9nq8oKj3gpfpPjReDHto40U6xcpjBqhTvscULlE2YfHGtup3xXTMaflKl
NsB0Vl1cpTa4y70FAKA+LP0atzzIXxtRIC8sWEOu9pbO9+JyabcobEUlFxWt9kUqCXXQxvDFzdoN
zzlahpOlrLCi9dpGfRU+JS1pyJCVGZdnAfljzfBDzy6iRbWwGY3MrU+DftAOWtCzb8G2oreUye+I
+CCaGbifxZ3RPNws7skM87Svfcu1prtWEyoAXSeoPGmjHnRhk8Dyyn6vtUE/xCMmgMduLhsDAnAx
WB75RyzwpUUZ+V58qenKWwCUCIKfg0TJYxGbz8SdM2OeppWxNjMxyIHDXSbuHXlK+qsWXgnlS5Kn
AbXL3OUYgszTjaPV9J6Ff3LY6Kvb168YffXMuo0Dr887DdqeI/hVLoHTSZbEHlrKcFZfgermgEC8
Q1OBahmvdwvE6+n1BLAWx2LrHZmpjh4c6Iuv/jzVw0m/QIcYNGKBo4PLFf7mVdAChOYqFoymqlSQ
k6pj1arDEWcdeCJ6LU2fkRS98W6jupfx9fRCEih07NH/JsKphsMG7gXvUI8szcok5OJBqT7bgcfC
4mjlclIkCQeEvQH09qjazY/nfJdw/uAcFYlVW1wktjkRG98Rc35cLvZyDd/zhfWMCQsEwB1drO2h
ZAHjprD3X8fuXiWyayzmQRq6a1A0/zTslXNdp02VWMCkjUiVFm1qMd2vA8C/z0zxYCCcKMnfQrvl
htZutAH3AGCfaPFwKCnPKa+sYDX9QZvdLBVMHxCVi3pljMJcaUQ6azMS8XEjxPm/bzw7qWTbG3zd
kSfeTA9SZACx6Jj72juCpMahgM1N32oVeOHxPcp7Jx7IQodcNHHDI8/ZN5b8S9EVhqi1+Te0yYuU
JpCF781qpJanW/clD7R+bZxUjqo/pmHqZD/MZa6DmBaC3AjSgvO3PoA789D4wGVwsD8gBG9KyA77
NDTKhBw8CEe6jeCbxBK1xAoQAWEml1F6LUjqmlsor5iTrvLB6aIm1RxWWDb2FjYIaNCAkCaWXlom
pqT/pS6dbRY3FrQDk3B+S6qC9Ls0eSpVRoyu8jMXJTiBBmb2SInTd5KB6Enmv4GcCOmQG9dIABQI
xfnZug8lgfoqKYh2s7OAXNjcsrz6dc3t7NwuonmfeDKRvH03bQCXzBDEDyRcXzXl1QuBq3OjchjB
j+e6Gnyeebm5EPiY14o+fbYJ4w2iTqHOx/Tb3r9mQwoCbloP0dUeMJ//BB/oWU/J/RhSM3wqVAYe
ZngPnmaqSuFFvyVqctYcqSqoI6S4iuV5xquxy11SCHrs2Fn4QZmBzV/VoZA5ejCy8IzyPwzGlwrr
RYP13fseEAWqRE1LKtTpz8HUFd8KdAbpffHUi0oOkelmHzto4Ds5X6cvkKTPW6lFwI9E7H6o5fX/
DXb8NSUz+i/MgdCnESHaXJ0GynDXZvr1BmxsqR/Wj53esbmj9b1EgjP6gRYQDu5q106oSh03xho6
knGfVcz2MXMmvFTAJEawfV8Bm2/68mto/+jHECB0Ka/KEM+b1XXGidphvpnbCbAab94/5/7+v2Ix
XZQx9OJQC6JR+xHB2jFjevBf0L9ZGv+dp32rM46mmB9wB8gVtc8Lx7Ft5C04UjHIfd4atTfzxJhb
Gl9/R4pX+/mod6WLxnor7MDRtUgRDCi9JXB9hB9+fyBkS+j6UFQ49hqbMQGM6LIN0fMb7nnX50t9
LUC0paQZ9h1rcizn5f3fCPneXUo8iPkxZ6JBpLbe2/ATSluQijMSwm5fRX6sDswiOO06hbfAgA4i
K0I1sLgbiKO/1WYgQhV1s0mYyKpG2tc5Er7UGhlBduzu+VKjLQFE3mJHW1Sa3HQQupJiRa72pSKy
LlWwWHeXYMc4/hrX7hLqoxKXUs2SlWjJm3W6oxRdE8GY3j38v1w3p+8O1rE7GOzY4I/DYhzhf8N9
6whEELYRfV5GwOueMrpLUeFmXy2TpEvOOdEAUy4j01L/8iSOnwkdnv5SdvVPg0bzbgDKeXefwKMY
1VjSeE3Z1J3kFuX2/HCNt2fwmW1Jzi/jbOin1Yq0Pz1fekJE3EqwAONFzYUaXl+xIAt0t6sqRdCu
o8jMPsLn1hit6sEe482zAYjcTxQx7yttDlryP66tde+FV2RLuDHNJON+m6ysMHz/3RlTGIlnfj2J
/nftMC2D0ddZNLtcyLHml6V5Nuf1dxePDjZpsD/wLCeATrhTAF4c1Tsmp9LpS7D9ntdpeKibvw0m
dDI2HCPfzYHIQ01hgyjfe4M6lFxnXceGbx3OV6K8Xd5mMvNlbXibvg5xoaI1iun9ARGkYdjlTdKl
bUaAe7ImOKKSZRw7Ufv8enO0WTt9i6af8WdAFcxuH9wIGB1VP5wMXhSQjP2grHbWXUEDTc+MdUH2
RYc0AQN7gzK/Yvnvir8IcURvSmBPHIzGbBN1Mscj3fsIBFu7BFSP0luempXcpyQpbS3rj0cnarvi
pwcRY6TUMht39pxlNvdBqWwBM5eo4uTl9Amh2pvKCIAeO87y8bMTce3zEFjZ6XngSgtID2fZ+5WT
o+HKesQ//WmRqMXdP8duN6RJXQv0pygucBJNWeTesXelJvaojivazuBg/dm2Sv8tu3ArDQj+EixL
VKlCYholBiZbbGmsu5WhgTxg343txwVWHGq5udBS8C20fJHc83NfnB7fJnmS33erHxrwpgi5yZik
mYFvWDoyJS8W61l6CbnTw5QcOK06TEkLquvCnSV8VG8MvpkrUd3nANDAwPeH1S0r9tKsYULCMT6z
JDbYCrn5U61QxlyGeJwyYnD07uDqX4+AjKYkTxeUS2idBH/3K2aM6jkSwBOcdAEdndp11lw9ZAwi
sIiUaUhRqI+9sSUC2eT2MsE/KXVgKbli3UYl5qUuXDcmr8rrkJwoLChZkdsboPcCPoMFHxL5tGYL
6W8LF09M4rBsX1WSU96LsRkY2DexhDwOQyZYVhoAsvjLZarHJIuyeTtrb9MAOVKx3x84ugOL4yhU
IRT5WgckiX8EbNnB0ypC5prQz5UK2o/fmmSQQDwclQ0Gof52C7qCZkZKJQFe1YrlfpbnWaAVAFNJ
JqLh2c+haH3L1QkZw9VDj1XsiKtVWh6DKojdmcjcnkFQXId3y9+fzylxOrj5UKrwqnNVLBw64dd/
/EDPs/Zn1enmKS9m0CtOBGsnwOWs4PqXFQbS3uH3VcUtlKjwU2PoomifYbZTaSo18u7T3gjBrFiv
vHvuFsYyMkqE6xShS5yvJG9SptR5sewubarG+++R5KMXs2/1SsAjt4POaFpbVyQwgtv3vSYVt0d6
Ht0iCGzYQXySBj7aTMeje3U+DPH/bD6PJK9HkqNi8lIWwXB0DEIz9slVDZVgo7Pa3mpfm3nIehJi
8x0aEncO4bzTQ1/7Vw3GXyN1fbMJ/WtvLijOvvOW1qNLQRyL4s0eTXf/M+nBxG0w53FnPbMI4eHf
98Ps2wmteAkf+BjD5EVrESbrelaNmLIEkd7CjcuFdBbhHRUdZgOsMb6Z6/Ali7DJYtGyacKY1mHh
GsPUn9ndVOXf2PocuFql0lio8dWdBs/QYfkqIf7wTSugo9dkl3iW3pfkFVUe+o+jeI9y2C0Lcf0L
6uH6mpfxfQGocZczlYAUtQrQS05kcj72faB3kJTJCVNaJMwxuzG55fkch7QYsOpczcWYqved9Igc
FLJxfX6iTFbJRz6J1pL5EY/QCXo7zliZrxG1jYS+5oThUQ8gXtzpN9dyOpuhRaO6vMz0vucjl4mX
WAdr5HgUJBzGjXKVbuBrenAWQvD53hTGe81gpgNU3HxNRYY4lPiwXNDxX3IgSwGThRf1w0u84PJN
CrJiP5RGSgJYbD45YiLnAepOwrCPbVD4NA08XXjp6Lr30im++QnsD/W5eEY9DxgKWVpIRcqfByjN
bms2Q2enRmInmYUWUsmrNpSfxOXX3WkRJmPV/76JdRX6OujTo8+ZVmjNT6cNqhZsGHp8+B1m4vjB
Rj+Rp3z4pqDB9SmlnTnsm35FI7ubRfTHfn+uBfh1eRyL+8FR8xXq4sy1VvwLEvERgw+w+0CAuIBC
3Yqm/4/ThSlViSDY2RwQwf9uEL66j6OvLkPiunhEsLXlixgTvlL3KTP9JYrsrqJV04Pvqzth15SA
CUnZbQcVCfIhT1zAhai//yR+sLlZ58dkCW0pRRBNxlm4vIE52VrpY24j8TAaSnJNIKx2fnM/dl+X
C16goZ48UfPGLDPPdUvC+kUskuurdAMJSLHBU/DxbcXhWgoFLqZVLXpm44ovG6Ix6HWar0bY5CZi
eozraT6y4sxRUq0Fy8Q5TcSluRz4M5er2YJVUJ2W5l2vHEJ25G0XfNnsZZAN8VBk+6ecuOYmaMpV
0fYUPSIbAuizBMK4uhKNFY+rwz4CK6Om7i+pI4wnz47QQ8lCxh1cQKBdsvz6YFN6KsFhQudziS5l
rl/CPlWc4u01XLC56E+KS1Lu/LbmAHXbUk3M4YDSFVIL90/d8hKUmA1RP61WU+Z1uqHVeuuGh196
F5wIcN/Kk3Ua1J5SGMcNS7lvgHVHy35+TnbZQj8dAz0z7GliN5s0I/D1CeRSobQmGvZkWC+6J4c5
aY2SzVJeWMPf5bHKpYxutoQFQDvcm2Sq+B+MPK8EFF5jmUEIWzNTqFtinPStDPl45DE17ZaGKs1S
t4fGoP2F+UeQcCu9xdLq91gxTWXpHGWf8keH6CjdtVGAbyq0yXQK+v8cSuIFh/fj1ypOL3ClWqxc
7SLb38mpqDDgKuO3UkVmriGD4cVP8bcfBijX5e0k5zCKw+1DLLx/s3QAhWUmpVXmAXb1TbddoSEz
3W5xik11pbyPoZEW9XIoq/J6w1MMPU5Ij/BMyEZZY80FTf1pyzcS/RW2TYihoqwqWhTP/U6OlqiV
JjXrreoWZfX4hDCohj52MCDdRr8Xm9CCy8diZz8JA/8q+yGj7dUg3pmc0QR9C3YsbkANXCUMEQw1
0A+3bUmvUptqYU1MnX/vZa/cRsiTbYk6lHa9an0cBzx9EmIQd6Rbq6mrd57bGiM1JnAF1MB+FMAo
quMNWZOQJirjo7nE/UhZ9nt4qUGkqCtFMZ3y8S847ivrQbDo1EXcJUjqAnK4r2V0xjrlUd/jkytB
lDjKrLrCE8sABfvJ87eG+64kts6a7/clLiMs/96iHjZH0Y4HSv/dz+TYlb+jDoRbODoieGUP6uSK
bvjNf4KKmiWnt50b5AK7AyUzCRhCVF2pbOyA12pzw1vOrWn4YxSMcJVX4ldjQITHyxucm2LgwjHC
oOa3QjfcBi1WPPJvcqjY0Z2fLrjYwbQDiUfAxg8cr9k5WwC9J5s3/m4+lnHdePHMP2wh//JTQbc5
UXCcZJ6RgxT9IYnPx7Uapa4/IksE5IW0wSjkFKdaC/LHi9H2r4YzvdcVCzRyGH4TRHO5alGsMErl
npdcN8EP9hH+uUpBndJ1hZ6iVWL6CrKdfr3NXYiqb3lF0cmuTiqx9Loc5o0JkTiyQYTbZiqPVuD3
wufowWzCfrjHY3/OVxPP2s9XmHfewwe2WlP+6FN8tQUyfMDRxdJaPo+6/DHLAM4YztCeEBuE4rwT
016Re6C/uqY3rBvgxBZWG1kRpFgF9DsBhQquOd1v6+7/nzgFsVEWnuTzieb4dvHcgaIm2/4DbAog
yImnw3/NtwMo1tinIVBYTQFKiY2fwDOY92fDMBOQpnKpX+5u7tz+jK+Tw9zfaQe97wDki9JU128L
ToPOu/d67TspQBICIvuDVLiNJj3Fe+6fl+1E5WImBqnwDGUwtFXsDhUQN4fBQRk0zG2o5jR2d3lc
iR32Qj02b6f811Q7YqITCJBDj5Pr1cToUQ/SKh5ow6Hc7vOWcmlYhveIg/q0Z0etSXRYYvfHPVei
a489QUnqPM07L0VdVbqFYf523UtBqNE4TaNIIvyanfJKHgWPQgyQxAjTWdmOnyvjo0xu62nk8ylU
odbAMfjjQoWO9br+xPr0SlcgmNF2U/rugv/qs3ix4aAY2wS/kEWHd6hdIG2yOO04YOTNhNBiMmdy
RNiGZwPJfiqkBFN1koucHloq2xFmlqw+/iN4QaQp0BwFIj47WlNz/bF93Ejlq4zMzjQjardoW71T
AZ2WjalRjrGALucJ8/0IMcUq4/vFTiPuzHapZ23w/48Q/WHiuH+3xS0wmSWx8MOhf8lZet8JRFGi
4wIt5qM/hA/mAMakVU6CEjtX0/grFAKr53zEo1ux3VCh2rcXpCEJmjtY3QRYC2ULzu1hFwWkmKEa
izPNjQWa/BhvG3T+x7slbm65+0Ufix6A4rTOlk//u57pfrHkR0H0iRsr6+mG5hciINf5MTn5exsx
HgM+MwrKprnGl3gICWf6zUp5bgO5stzu9Yjjn2PbuCbvmUTqdfJy/a6aw7572OeHXfR23STSF4iD
8ZwP57XI7IVavxaEs9RT6lwXXuAjVG28h9xkQvxewennKU6ykaHNlAYIIi9c5zel04BUHVoXCVBR
IVFzeu1x9teQw8HSO6Tt4m3rFd8aSKGlOso0qNAmNvHG0xbDjhlKf3UneOrqvBzoWEhgJt51jDtD
NpbAoOm6EHZxeakXwMne6asUuzuam9CoNyTJaYUWEk7RpWRQstlEgqpAXL6YxmLCojj0+DlucPg1
HiGZRR9TkyVkiZnsBlV4k6EEPcYGwnw//MbFwjmRxaZ8Dh1rjfOuvHzAy50R2EacleDmVQe/Uy7E
zPqKP8d2jqAMhdFGqNWnqi1653O9L3jCcWPkNo6TxTe81RNUAaHEe3qL5Iv96YqOAIHADIbh9LFv
VxSCNLoB7hgL6DJqpq0TSE4tZp8IwEFkT2Vm2CEhjueYY2a0fNSkGlrpxCscj6ChpOwJd+a9azYz
qsgdKam7whlwUXuwjtOtSBku4UzoTZWrmE1KI/3RE8WO9RgFmHfYVRRb/3aR0gvELzGCLLnxAcRV
3UCqwsHq0ypRu+Ij2q8PiIk1rw2O7wLkajrq22TMPTFwRVmi9h3UzAMDFI5OjqtT8TL5mA8i9Nn9
Np52oFKUioHzMcG4ZdXAqUH89j4NN+NuGLXuxLDrGwAmDR4Y6aZPAxyGbOfXAf3OCgHsDP68a5Dt
HK0UOL5WK7C0ZQkLd4zncVVaTKhy/Cx9pNL4GCGBVl/gbkwqGtR+xrPDRgNs7fhQ7Vngt7U5lIKX
oK1Bf6hfd0PtQQIHHHLvawl+a38VPDuA5uXgCvhAhjSCCjX3cwsW4iR0pnnn1cVz6B/aJYy0L6hM
jZ8HYlxXOEG9gRkdT+RAHMO3efK7FPjc9OerJOEOcR4LcsdyxdnIC/V7ul5us/KH6qhgX5di7n+i
dWlwnWgFT4cU8YQWoepK7LmyBIeYVULdUkEH1JG2ku8HxMET4MFna5nEu1xKCC3HemA99Sl/vfj1
xFxk6cCYWQ3Rq4lTqPo7PvEHQlK77GPrYGtUWfY0pWncACEi7Dm/4RTVJKT5Ww1khJ/xXDDuQrQU
ZUX0gs2gVb8POV31lvnualjULUYhGDOvMgrG6iwb4wh4r9pWjEcPtCSdZ3s1ZxNFhP38KvIYHea/
qJHTCy3ZV1yoSoFIzF4Wk37X3ja0+/C5Mj+jNpR1PSzGZV5S7G7NtaMVeEFWYFG3sXXzNL/20CXl
NsOWr1OnCNOItOBnQwlKnBOp9KYxvCzdvTgemYKRxq+SVhBfTnAg6eImeIHBgBT7h5qYjmXVSfrR
h8PIwdPw3UzKsvjX5UF8IliTCawmliPztgoqPJBvFoaCqbGyhs5C9p9fPbMxa9yDJ5JxFEleXlUy
Vv1Wvpub8B5xKSoye5uotSqY2lZn3BaLRPsKkBwcvDrROifA+rRr8STMYrC2fWqQaQGnI/+ws65Q
MrjuQh1g4kyesvbsxScF1FGbqCozxDepJ6+AP7ukC241xFX2n+OkLJPYBKPT6Awhc1frJII7NUxI
lYzkpCAYZuW/iTsGOiJZ+SNk4KFreUn5e5wRLJ+MG+vwzyCK0o9Q3aYEw62o3+uPpotXzpYOMFLj
YFmcmg95xyTxRc7AIUwrSzizBbzufLtR60F19hyTk18YCjnUOBcSguQIzLJ+H4j1NX/8gLGBrMaW
EmB/8DR2TFXV/YwFO8NDv+kUsDGkwzqNkIWhv+GCOkEGKxgkWtAKHm7V3lnT75zNcn8YdY4qykjn
BoBJWErEit2ihTWQHSonvbDGNkpgi6K1GGfBDqKzpuSMPA6UP4p9Nj9L+akXttdE+F20nvUBg/Pn
cyi4uYs1Ovy0SazMgVI8Z0pEbInAe7LRv0GKptLcgj0/JtrI7Wq2hYv1s7eo/cqWbbz6GCyn4+5X
HwoT4V2xl+A8t4+2ddlzrGMLa3MUDLLDHYSfHZ3/4IfxcF8u2n665kvLfwaDjc+hcFLX1C2LDCpS
44rg8/RxFAhtNzXO/FJdtxAnRGbPcjDqmC3BfYmp3TyiGglrMQSUKei7JqAq/ZvmGFIhQz2n2f/E
K8aA+RXdkVshz2XDkYvkU91HqFxk3xBS+r9eQFuXIu1lJq7PZoz21djEDoOB16xCb/kiqwn8Dxqd
C9rryNN1mQygQtS62T16ATP3T1a3egrnXc37N5gxZK4nU1cWTtmXvlpeBfLq4wDLnnDqSgYVWH/u
mWVdhEtG2a6FhyLJ07f6oBKTv4Aomx5lHr/gAY8VkvgQhUyZt/GiMpNIoZvGU1eU4ZulpSSRYSFV
8rucYBVul9/BQ1ALzI4Q2NciSr4wiSpKuQ1YfVc+YgfGNNnD/OW1riCLewbcnlGbSzwnGUBUpTRb
472DKmbYA1w+7rVDdi9Br3OhFiOhoX3uyDj2IaKd+av8EhaaL8NhUiWaLvnRhYCwzRjqLAUB6/7D
+J4eSF3NKCnxwILtQPO74geuQGUuqDEbIlMab43mZOe2+gGG7sSCLtnyA6xS0Ju42gtscQNrpc4+
SBiWIXCjQ99Ul6HRTP7tR3Ez08NBjjajmDCTBC6RfO0Fq7/7auaUUdDIdFcJJtDstCmeTtIr1YFe
k7CeoUmmmPy+NblSpk2eAAFfeIkZvYHWHjif6UnxDzJTbtwtwd2cAdyn3UMHgCrZyvYBOTqly4m/
GuzMZYRnQKNth+HjOEy1PNBYln+RAJrwR8BumpbgMlTxs0+7QymHGoYudf/PHhhWnGdhcvb69ITg
dh17fVyC2v3YGZW7U6ydgpya1ACI1U70JeMVytIPiYYV97Ig/WNTVRAEZEcbVFUzQsGaJBkwRTgF
Xu+zZjNun7UBapwUcT9muVGqh+2c2fkv8cwYU65UMAcGrGsvoM4wpXpVXxlu0yW+7iobEgqqPh0K
leMoWkKHKfr6VuxgOMaKY5SM8B0o9QTZB2UszXpq1FjbVJlnLGefQJrbRTGvDjfpCpCMTJS/yLe5
RkeYcn8pOTz5Sok1Xutj25lDqFYvzFfaN02nAXyaFYbEBfyNkz4RmXkFhfyaMkIuyhYf8EtJlssg
G2ZT506TOSf8piIqdO9CGVy/Yu7dnU4YmB0QEOvMlkyliWKCDaiGWZl0PZtGv/aPXv99seEes5aW
Y4qoRcSltdWPXePbK0jyvYnks0P5ACtvBXVzWeGfRtrZizus/gDvF0PXqSAQRVblXQ3fPyMe3v6H
61l2YNhGnIQFTl5OIYGCvbXx23NX8Gxtn6vlfdaSqcAqZHc3NgKPFZ+3yZ28o0A3m7+i/3K5JXtK
O59KxX/ZeYVC9KAGPM4OiPRK6azDgkbvDQjv9NJNElHw8GkYKBhy6N5jpK3qpeBYaBsYevvGsJJj
nU2fP/X+6AcUsZR/XJwcLcc208bt4+gu+zEhj4hzx7BdA3FmVPiPBw2W3oku+OkuRRO9YH4J0tGZ
5wPA60yUBn8U52Fld4uAyHL74ncGRAnqhNLnVT7noMfpKKXsNi2Sp2oMAtLZsta0hPLs9GovrE6I
J3vTDTaP77c1fWNZm610bg1kQ3bpMkUo3T0nTFY3fO26hu2PMtA4QE17d6ADULhRydBrqs0dhouk
WKdmL5hxbluW+Ve1jjUEWk84fgQM0LNaoDYpdJKLyUEw3vaQCVTU7O0dBLYMO64igq/rB4co4YAc
BxzMgE3y2TVv2l8O8gsq9cWNEKPzsJXNX6Moc7NuWb8IEdPFIOh3tigY0uB4Ooq6M/Qr/Eb/U8Lx
nEncxpgPMSOiIVYjEkYlWejWsjR2Vy/EzoU7iKBDyg/VDCb/X2dj/cBrYywHPiFOor+869SAp4Vt
RbGG9R2v4ChKDqbz6zpIx84AXxVVrujUxp95uG/J46LDhPhQPVmWmiPZFPBFxqJn5UBtKnzCpUql
vVpmP9bG/JAGQ2dP/l78fN1h1WyXfeOxHOCzGhk8HEiVPJZwpranUrtTKZbiMxqjcjl5JsFONR6Q
i8654PMTQ5x6oDANAqRqqG6HPgn3rwsFa6QpzGyWEp5PMhVfT+xIybbfy/anV2wwIWrVJRbxoQ6e
8GJ251HBH7E3scD82KcsFeBrISvD2CO+lhpPwiFX+FDIYECkXTiQ/3xoTOuXfp6V9uIXhsIipMGj
88diSNEpeNjAqbhDX32Y4mjMW0GPuQHzSpe/jiSDjOLtA34rym6x3SCWVsbHP5GmDJsExRj1DTyF
3fdinC7IrIPDrZ8+XOq1BzAP4FEOz5AzquAYDT3fU3wwGIUlN3ZnE/pAPjtY4zaniD29f96R1n5g
cVJ4WqsMQB5WGYn1dAwoprs4og8qYVU+6zVmtqEjVJcQSkYPSpWFRD82JwM+q+C4+jFQOro48j/d
P/ZkH/x0lyrVrYSqsJag4eUZdDUDlFsfKyMLJ0LN53nnIo7+epFpuqBXzzUHkHvFqwcVOpbgWUDR
E++N4Jeh9wB45FrPS96VafQLKSpOIagjlMIKlSEN4D5wkuaprfFssLCO0VWFMvYfrowwGpf8AU7N
cx6XLTE9X6X36Pf0yCN9F9S1m1GTItnkZj4H9e7UBrpA91Az2oEsOMpgjapkGwew4QvkwuOlJhX3
GgF8ntZ04eXK2n9w8sQOYWK1O0jNHqlB6DklfvX8j4sV8ShIOI+T3xFdMvMxih5mta4JzGCSlZ9L
yQ1eR+3tYkQffwgKhtgg/MW6A1AAR57+bGl7FbVYxkOyu1TnsvmdrEpiEAJGSCfJgJHg8NGkAl9y
/vPW1DOp+vMRuJgSD9mM4RmugztPRKFO+USpd4Mo/HtajkxqyP3ihDVQPQ6fkhIyGMARC4yJgorY
c/ISVAs3I5vBx1VaOUVYZWPWzdduSChUKwFm1KcIle1G3xAdqfPmHtO0etG8JC8Z0NkU2mS8AyJl
AFaGGHR8ubj1q3qF12HDzcv0a9hWhwhDstfZvNY7NJriqzQwypoz5BSaxUz2xV7D8r+tyGpeWNYl
RWc7QOx4nkE15OjFT6x/JlsoVz+avrkZJ6H5Kfx4bN0A9ltvv3aAOlah5Q/rzeNCJLOZ0cExAiQ7
qMnYpyv6YK5L/NFjymvbZ122dr+z1afobRaIzLWxe/6XY2eOC6M13Kfr3oQ4S42Pw5Cp/B5W1uEq
UmCokQ5Tjl+tBu2yikuq4R/QJFuntMyvi7ImFD8A4k1s75/dIYD9/C08KHxltPx1r/qqbOWLpqrM
ajn7GyEFs/EYbkNK8xT4yDg7cMtCtXYPH3akMa1pmda69yzkQ+AMNQAAiYWsCISP2Sq04j7v8BIA
a+xiiFc7Mdj4kQYkmeJV9sPU9YofYgyXgulyr8o/PbxStSzhk3a7nWbkgHamVCS+lSTKTZWlIRyC
dl6vWKCn2DrsqDVj7RYgK0mBCMO16OfW7mhSX7jU5DlIuUsnAl2GShmfPl9cLz2j5PqXsmAPC4qD
QuR4PVglnSUSjtuI+cskbQ8qbQzngu0Z8IK8Z3ktjPEy5v/IXP6XTJ7IPG++voPwVwBwUDmdr616
RQfe71ZsPovlIUUZ7EAAHMvqcxL3o0OQaUHZ84qNNAeTp21ZhFD8zib7iOTG4Pl1oFgeZfNBvTtP
vfk0e2JcwOc1IiUOtIgkjcMkeWz7FU2MJRuw+qjjg2MjmMzCbVYaviRiZmQVr2SQzgtJOZ/DxJ3J
+cWFxtaBc3zgLgFaOYNdIB6OrcBouNC65sujZ+SlRi9xURO8/5e9gvVAo0drjNx858drTj60vFSA
pmaLOvkhoeZH1pRsC76lLqsNlk8sJRcN0PVfoSJ0jh7AAyuW1DN7ayt8+QzrPaUICzfsDjnLxtBM
Bnhorejkg1RcLrc9nl2IfNyzIPcrOIfSb4Hwu2X8nJA1/nXRyvWEut9DS72LArbih4xdL8vvvG3y
t73eZeZM5wBxwvdPkCTOGSYumh3o0xVBtoVxy4g/FbTY+I2wTba/hodoMrAsrpP0v9Lr4FKijYKR
/WJ9gwxyUhOG6GacZNTUcV7b9YH0uz1Ofvfg1q3rnvgl9oKrZ9LNYuRrJkB1UVDpKqOkk/M8o0g3
wh+X6xyg3WxT1Q5YTSdZiys62Z8iJ1OtIheexPIqzXr7ILQG1oTsXEqJd/7Pce3R8xzrs44mzAWE
Hzcq0oc68F5civb2zU950lp1g5o45O4bqDED9t7dCmiwRCEj6M4IDEJ31q1J1IhwEc1xm1wfXABa
TljSwlmBVUrpuOWUzeyjoGDG/gCofWuoQj0nznXKLDrycSWIyau5VQKxylp3R7MkuS5GInSDz7nf
sY4vuM2B/cjiFv8JtmdtfqM8FFrfXraJW+pSXjK/d7kCG7w0qG6qzc7yGirpI2RBTFmu6v/xYclu
bksawY36WDHACMobLEXRIoFPxjJ0nzhgWPjzizSb3rl3gD714Ht+p0po5UXmWiCskIRdHlk5Xe7T
NJaUqMgtr9RanzMEOEmciL2TzCWGBa+ACa4n1X3h4HfhYLM1Taqgzj2u0fr+vEViiLxe+bfB71E2
SfCrvhtAAUF4p0P3QiG03U5qqZCjViElKBHKZ0jLzcqE6R2PP8S9G/ZJWSO20nEfyHlBrMr12iZL
XpXQWT05zSlVYWqRd/cO4Trv7H4gNuGR86i1+p2Ag1rCTXbK65+xQKfpWeQU/JhNde2QEVGreaIt
qoE8O3tTKAw2TYdllH4pFTkEuMukf/zMB4kYwAHHMlS4dPfjHvj6WPs3h1eQ/1PuVeEVK+Ehrx1+
0691FQuii0fvbixkbIzLknB3/mRGczb+zv4qdCGSR03+HTpBT8jrlTuRJaYeR4TWaOealNzqZTLJ
rJRmjIZslTydQoZ1BoxzjGbraoC7jF3DbpKZcIucIl7h9P51qeHOA1i4Z2il2gVVoLrRaakP7Ypr
F0vlvm4Eg60sl+oNgJ0H/U1Lje4JMaTzYDSigYx30Iu+w5m3MNx1EE2DKGz2k3J3vHpuggmprEhu
E19Xsn4YxWprd5CrOUMdDwHlKIFTT/kbx0XqadhjDoUq4bj0NY8JF00ZC5psGkt23IHxGzEd/LMW
p0TCvKkUqhdzxswgFDM9nTvs6DkvxGEFpEhl+VFM1F7Y1EJRu3GRTSTSH+EgF9EBXd+cAOZSZd6C
qG005HohbBtdtuBtpaIUQR+R+m8yDMUAFUOAXp/pnCL3dSze457aKy5ReQQMZWR751xvdFNacc4e
SRK5p/B2l/2/asB/S2Ktu5mlXri+9TClCQnE2A1GD2Cj+nQ3/9CxsXDXwOQ1yaeGLOlL1V+WkdJc
G+omYp5qApizO2AldHvQhBn7Eye0qkhNnko7M/xAEg0KE8m66pi5HDFyf6OMZITnnkNYCgJDsaKE
P07uDjLf9WMmj3/xj10DWmoEH9JBV+eZBeor+hDNisI7yAjRL6FEp1GjPekMwA8JRb2nKMgr5idR
wlBMFNtHzm0BhxlN+Vi3Zpb57meawJh8nLU0a7FpFqih9iU1T6QfVbqZ3N9o30RYMFo2tP3so1tv
G/MdhUpizDnQRHmEZ1+OzzzMpSVLGOgiXQpg3bZv6GHQItldFY46L8K6M/AD4Mzkjnuu+8DfWJVO
a7N17jb7fwvHhS2XnE3IV73B5Eugk0n2w1brR3Q6PyBxpuNYAL2TTB247OR5hahh0LIclL6F0ni8
ArKzWSYmx6LsfOymnUhANGk80h2nJaRGlSd98Wa3Q8c9sUzSkXUqUpArUF0jX4JvVOV952A/qemt
2pWFPTByLCdhInEtUHv9YhbDTPRnYfA3ujqb3nHHzNPXnVylf8D0wXJNbpNgm2uUqez6GCAU0O96
D6arInVwpTE8Ps8X0mTpD0MmwvBWP0zjUYkEZ/+MByqtXeU4htFX/88ALohgwHwHCwOuxdHx8cyF
fzwEct1e3drAdnIZ7wToUpbVwt257OT2bjSPb22LmtTBz3NMVOCrJdWP8H/pSUNs4wYEMfHIR+mD
303L6T5M+BGgjJo8GI/fju3coEr+KPJ5ndui83sKfnFVnDz/E83ueHDXfqQN+WbUhavVPp8dViDA
kxyIpEUXJ6QghdpxRA+0SMHE09+fmyFrPLpRNiKDu1PjJmdQUgaa/S4UKybsfGWKN5wettX45VxQ
SLGWxaBkZ+7WK6AMyE6ovyN6ziaRQtPLQdZT/ZhTuDruvOXoEvHM5XYlz2zRcS++TVYOgbMlwt3F
VzpOrWFlNA2cjnZQ21OzLusDuVt/uoIGmHKwd5vH4ISAK6vABAEdk6NxH8ecuBuILiIDsJ+mp95y
f/K4y2ODx5twoZiC3aBv31dLCKJq9nPHRr1qzzyMchw0hVfl2PTXFhbHugPqw+ddc7AAeIhsNiWa
HzeYMb2YQaxG/TirUkF9Kc+g+LKatt3m840N8qvZ9u5RUR/yfYT1Xv4u4wVuWQIVND1BR2I4AZQz
6cBbLVaLyNcl4QcOWmxlAeAwvalhKfSoPKrar7dyG1MtVhfhTfbGFqunm75hefzM8O1dS+7pwNih
xZQCYHRAlN76nYaUz6x4Cm7dmyQx0r7GlNcDT4mWirq/VwY1EEZ9v2iKEVHbN1cSsquvArg/bCVt
PqRkuLqnlh18ti1QkuxbfuPAaaPFocijC7tUHj4b5Sv/oqcovJANeMlYjmoZjr/6UHQKucGcY/1B
5LLZjaUfTm+Z3dila5ZXYtASR20uL8bVCYlnDhZKfXhh/rKxh40bs96ZdQYhR7fs4UzS8yiJxL2W
CduXLaJt8Yh6GscZjDaXB4TMmVcXDhY5rPGCsE38DVDrcEnJCHqILPrkpWBbiyXctOoMKrlwUP0Q
ZO6FoDj4+XaiqLEjMozmVPW3dsfKkuFjpTjd3hZlhUJq9KdA7uI3WEkaTpEO4jiCa05djHpxazqP
kfRwC8AN7uvx7yJeeXpBiLVfDyRuokV2N3/umOMX/Kb3Lltz9zNdJxVtZsAsE0v/d+GD6ElsqTzY
h3wXtT98sklLHyrR1uPDwBQzwoU9ke+Ku2lY0kAGDh3PK9TO7JTrR5+gojqCzkKR304mMehMiAel
ev8yBHobjLhw1P6AGQCRyUIq+0lzhYaIP9fV0Ufk26nMniGkyZeO/1sdGgDuS1lREhvOnvWW3oK2
th4j6LFF/4p3WSgXROcHWCv/RfRw5bqKQZzdO5Urhn9oZVv+nftIQk5lf5Cj2XUOX+h5zZ+e6pEa
oQ2HOtZgfsoLdIoQhm1uZP6u5jXDgBRf+pvPgKbJq+NWMgGsedUTVhKAZ71/+saHvPf4QPk8BhRO
ub7PL/hGlyv4Ws1/ICxGdjBJdxHxbd1jHshPjzjzXr9VMeA+gQzd5OVksBOZuCuG9ALrgqsO2hYa
QfXaBkTVyv9SiJ8hrL3Y6RS/KsX1YLYUAvZfwgBoXDZIjPMheVA8r3Nu1hH6CJ/0Uyka1w0awMxm
wxj+kqWt75xqVtr+1ITELfjxsrtdnu6tYOVdEKheaJcRa/q5VDHF1rxfa5v/BfYVTt6c5g6tQ87s
cfiC/aIaDd8pLSKU807MxBZkv/nS39Iqc37Q+U8gaoNiQMuThB80+wDVdHlsTmFTj2joJD2sfnsG
DQqgzPi7ugsP/xg1xM1WeW1eKudHgC4BxHkUPgL0vZuyFDvjTZq/ADrTfNoamKo/KZHqsfbR/ioE
TdNtHY076ZK6xV185FVdctsdqVy9Gfk0/tm2f2gQ57YH9/2VWG/2arso9LNViFA4SDsr+ykq4AFt
dBoZxW3xaArFtJIyzJ0DWSLNFtEhjpA8VQ/PviYv4OKefynUc45RReRARK+Uz/CUePr98XPt1z5n
50qESXSnOvTHcVyZ7h2DYD8QZ5SSLdIczDrdr7HaPVe/0wSVr4O2b+R90awHQaWwZNdmkYTeKmX8
zPV8E9Tl0k882HwbNzWQUAIFbuO3uD6NIHrUBBjPMSNNmkEuaNW+ORlu9P76Dbp7haIoG32LX43w
XW9m3F8ZU9/1Zx3L6nbWrx4sD3xxJEj+LokR3m8cODmBtJHMeBrgEoygRUOJ+Spp3poJb95uZDyZ
gE5pbSmXGIGBONJZ0I3ACJJVIFi9zhPs1tLzCEt1zQg663sjgBu9j8wxhQ4EPcKV9yAiy2cHTupL
e4KwVaWhOlsEfh3EVnxWtkhrhwTcyJfBUnDhx8XRD6T4+vr4xnrIPTliILY/kTSysCuF14vcYZj8
/8aixdLCB/In2c2TcufBHw7PNwQb2qVsMNt3xBc7Cmil09BFcjB/NweWNSgT6lzhay0QFOmA2D+B
YjBiXpJ+0t8Ce0YkYt3rYrCbA0thzAmtgfiycnvJNWc1uBeCn77/B4x8XViyYKfSmGipqeNgmANp
wtFAC47mc4NYpb0hiBjmWNSRMBokIQvzK+N1lCFkBTbO+VgpGoph+ZmoW3pQSLuu9ywuQLMugipZ
/gSJTQvmzj9v9Zln4CZupZj/Dyqt1Vr/XF48XOd95afoN3q3qKu0UqU3sSjvQSeaU7NIuCyWeOa5
B4P7gyOMOZlzb7fpI70UZ55ibf6/n9zT0Bzi7IB32H6yUS23tTYoOp1WXBNKETwJcBJ7lfFlV5hW
n0oFlK0dAHe8o0wPTuHaVKB71Z3Exwl3LujuuP+kbuBBFIiV7OW6mGQn41pI2ElLSOrcT8WkoF0r
40cJWk0QT/7Wh3QMsgfdKYef9+M361WiJMJBhzl2ZSccuKpqh8h+Acx6hAf2MyXop4q0MMdz3LOv
6I1P20YFV1H30MXNlvwATDmRIt9S5eGpSuBc+EnPoXhyhO7mqXEmekJSEJOikt1RZrJoiLPQVUqy
NwgfI5yKjagkbuETmIvlqjPLPOvTEONuXAoSYQmSGyQebpyYub+Nf6f1qJwdu5Jh+1NXuXgfO2vN
6eqViA6h1al31i2HdfbHMsMdBLFi7kAH9lQmcsn863mp1VHvQwVcmliJBl7RcQUR7NMA1eKwKRN3
Li5gY8DKwNrjqpME5JrSpf8NKX9SBYEA6rV3WZFBv6pljTqz17UXT72xFt8wBMQs4C2b0sTcbyUV
EN1dg3S9D36AHKxZvc4Be8YAp69HRsqGKfqcn/oyeRucpeSs/4/voqJYJBhQ11Xdw4fpME5PIIZ6
nzGJb+ZUmkKB3Sp9LnUXFWrpRjgYopcOdnenHnSj32E2xC0mLNpgBvq5CKHpTSp3lJTwpdy26zm6
JSDcNBisqKe/nlnxWlEgz24e8hNpKaGr633U5d50LtqmoNLVXd7R4wmZC9d8M3Dwlf5FYdXl9M6J
JgYTjPItbqQ1X7IN8RlwKvE4I+FtYcjSJM3q4MvpWBUhRUt8H3cjHZiQnCZ1Z/LV1gnlvSRAxj+3
NJKpHWV/x4Caa/ngdEppa3bBFL2eheS2nY/+yKZJqcXiGWTLH6/3WSpn3CfFrjNFVZDHVEVK23TR
t/0tcvRetIf0ZRQ6qoL/q6PXkrHMFF1bvd74QSlqLKllYQhQq5e5iUMuimWy4gmAvAZgljt6B1lo
BmEaR3v4kiGpCoSXxCNZeXGPQ7j5kNFl4OB3ggqihQdkNBiH305Ua2UPtpEw5whcOeZip/wH0Pp6
POv6eNaV4OMSkJ+iT0JNSm8qjLYrm6GWXeBwbBwUaqbFJjrG4x4uRmGJtdTWC8KkxKCKmq383uIB
2PEWJi19EAT2UyMkCCcUpYezZNAD7Io6VUU16avCDYYj2Dob+xbdrx4Bkz48AY/eDSr7xJZuhK6F
I97nUJc6V5LOhn6ie2Sbz/CdYHX9knErL4q5unpm5HaKuhx79VI5v7V/dRa+58zj9oibdEUI535r
Xcdiys8fCFt7/OPOWbKxc+5rqtbtwt6WUuwur/kN3DK28LZlSYIdO9SGth20e7lDf8ckxYus5cch
YZtRLqpn90hndLpI1Bjbp0UH2nzY1IhYNl2uu8jrkzkn18SvovtrC0P19j/ysQsVsQGEcMzT0FLM
Oz0moFOkC/InHvKUtlf3GDCVOYpRDJncBpHDhyxr3ATc5+cDYHokaldedSucdt2mgkQCbCimcgcu
gYQLSECQfEaUy82bJknHqteavwSJc5IucmPowGruHKxCO0QzK8Gky3f2ywnlGYUL3qOPbJpSUpAC
WEN+JP8nWlu4KiOC9mK/jf/KD7GvaVCnixHdqRA5jWji3pLQK0mikoN7DQGAKu0yaOQqZaLi+249
fw/KxqaG3T8srdOdEr/RpZrviJlIH8KSW8ui78g5um7eMs8kWV/scUNw1bJUUdai1GDkXjA7mTcM
RfqcqtaXGl36u4LhqQSkfBCexDsfAvp9/eSjGULLRst2iUjpSpxx+dVCqKzVRQxU+K5Ha1RDqRYW
OQE1M0ebjDIyDgU1xCrCa+MCgT5Z2KzUKAF506jOO6kN9jm1Vvnwo2O7VEJymSgZ8AHmM4YmTJM2
9FhXQj6NBjo86NarA9Wfu5aP54pjIZFRRUiWCtRnUDoncknaU/3u5u+hqgN/4liwUy9FhGqUXdaN
QGi82bcjzb4TkitEoVLRixKeEnKIGVV0ZxTHrXMccVw/iTJW56SfxehjaY2t/v05PNfaoSCBwEDu
5NZGFWWfwILYDzJSD0ikKf94uEUIVe88/5OZqJ40cuGVFAFEBMMr0fZcEQ4g9UimlSq/0jGvnH3w
r3HztIq+b+NQt7SlLGREfe3VFRWi66f9IJEz8m/cbmZ+a7KX3DdarMcZiEhObObrQJ19ZGXE+PSN
goEqTBwJE3pI8vyepP4qLsZLMrAMjsa/QFbA+nnkwHz266+AYfKNT1+QCAoboKP0X3KHlP5VhWK7
IzuNIMeo3KlhPK2SajrecEsg9izdrZ5ntiWibmGb4t6z9O8rMZtiMBZu59uPQnFBVbbS6Etj/yWn
MZfF/4lSmaY96Lhj6op7j1Fu0nxuCWDDHU+WA6ISQ3WAc8smPYN4uDKxx+KgriqoZPk4fHF94gwt
vGkcgkGN3QXyIG05wn2I0D1v4vJVvu3/3UYgPpWrjzTy2zxMcUOmSQm+ncEAvblUIOYwkbdKQxy4
nFd6pIh24fvB14ibAEAg6qSgrW4y8PQwygPbdDGoSnd2A31z85tW5I07KU9xgkunzZsall8OyVlA
6KChf4o/3hSViOkvu6UOTecvsLXwKTxZ3r3pbQZzWHjiGEsUqdNcKMdmv6si5BdMxUy3M3aTagva
qEU+O6ptypNcIoEITmO99/mNNBZZMQWrulchwZ7505lfRMaaJ2u28pn/X/ygxPtbV+tZv3wIIVNy
6HJrXK2yatdot76FaMGOhMkxnj9URRMs0WOT+I4iZDEFwHLr+rOj2BW/Eq2Q5LCu20v6WdY0NBje
KPDmQ0LvNtDkMj5otEjm8B17BNuqgsHpGLJuOTF4GYLGDkzjBOYzyCoXmrCbh7VXmCRNWCct1PLo
S9c2rnYm4hlLCjA1Sf/czBlMDyUh7eg6OaVmS2wnZ5zpyMMz62mlW4VtoDqU8lRsED9tXFMNBUt+
AUrVbUgKL19qhfqyuGYzz0gt5kwkeEPUrWKiOFD4cTzaU0c41YiaPjSjr8aaVpmveDz0mvylWOcq
20hwbhcesV6lnc2vQWiAXbFa+BKmBkb9UdigLWzpBE6aK6fSOrAzxB7TGLzwZxYRw/9w0nOGoDLo
9K8Lizjiwckr52Q8j2in+iRd+ldysGjr3RJCEHnUasIxBb51PaZxuEb7qvnJ374JejXrps1oF0ly
pZiQ8v5RjVIZVtTZYERs2FbeN90hTgzZ2VY6WVgMQAmEdvQt3n4rH8YvU8s3/gV4mYhpEOrr4c5M
nO7vr/VKVF674s0lCQlRfrSiFgvyGMWzNQBr9BO+UWpaGPZFvIKKpnIEKUu4jilbBgyFcDLZ372d
bJ+95Lk26W/eyt29MrNY3xQrlw0tupCkPsD44o+HToRCXaal+SXdd6LYOCEIHJwBUEEYKmlxM7rd
PJ8dtmx7uz+Zcwrtewff8azDfqwo72FnDHgscIceaz3yj8mHM+ZQwIJ0ZRO6DbAKopZAohObLSoY
WetFWjKD8lK2IafNV08be6hcbQsaUdmpkR7ul5OZjcYcdE6/DiKzFQlmnakBvBw2kzDXpxwbEyiS
jDVWBpQVsfSmtPiCwdAiT1ds3qN1zzUbc2QNpWtcTLcA0bNMOAr5RFf53RXklf0EsSp8b0qm4sCL
PFSVNCqv0zyCY+39bXchZxgGBzGoosM8f+J11q01AvakwMlGH8BWJE19b6Hd3Xm0BJuBKMJCKSef
VhhQPTV/ZpWQaJBAnZO7JUQXr2GTgFIQ6usTEIfEHdsO4zGvvA2wDNuKIfzvv8BWbQMAvARa6rL1
3RsqpO4mH6yTXf5rXkoghu4Fj3PYEOCzREMZ/Ya0pPWFnb6340Z4/8j6orC360puX1ADRyB9A3GT
L5+TDEithcJkfD57i7M0Tm7jQnJWhwYhN/q+eg0M/mVTruWCU/+S7ckBOFZhMb9EZcM+lgb/pDSz
p2Lj2xIeXT1jjvcLNZ3hPQWEbGKPR6jd5iky3xfB57Osy6pkcFPDihUc9myWnRncQ1wr8eGeyfP1
1B8sSMCvDH76sfkAiF6NdVFC5z/LfdtvKVlwcWoHbrt/03tWjA/RKMMLBo7I+hJEu2TAR/ShG1xu
lhHGnoemmb+Y9ZmWQ+VUdrkwOtd2BkTpw5kFi/I4khBqfE4uS57l3IsOl4ULOz7oNn1xFgoOUDCd
fjE3GxjgmMZ8eWgj53AUYwguP/EhkI1NBXEVLtU6FBMbdL6wK88Wi6DMYeXIfPe+s9Q68c51vG9N
gJ6cNtqLNm21tOrZ1M57LJ1iOVUI1dQ7OfoBW2BJ17Milo8FK4egFSq2CfIlp4vmvUmnZ/C4XM/a
lXvavTRz56DUNPFgx0XmgvTfFa/DpZrRRXRu75XR2jjjQsouN7bbiOTWIFK9VqJgpIbK2Nvxpq/s
dQS86N46i9/X3hrRIaCQTNi0MxNnsQPrTITBRzh1Rg1siK0cdA/qS0wRSBmeze6QpeyU40RuOvvO
MnJ7r5dEfUfke8qDm476tnef/48DvWl+blgi3rN963dDDKZBJb9457VdcRTSZz6HHOYfWrs2dJUs
ZcELdZuxdTo3debUO55K+VuWMkEfuSCBtqc9HHiuFMRRCBFjgRRcvCraItf3nhbQ1qwPZ4Opyd2Z
YEl+dmEV+WQxRIzfrhcFodmiol848bxzi9qCRKiqu1VVYWbyB9UoMDzXA66ApZt6A16vePvinX25
5oQzi1QM2e+y7jRcVe18QlNtVCY7FR1vVoBMJ+LEekw749lwN09TD5r/BmLtktoOG6LJzzw9jYr6
2bNd/moKF3jn4FNCV8VEkW0REUJqREpVxm4lPTi6pVKKxhLCIoHM88Grj30bSRnyrDOSadKWNvQ1
NEtbDbkh3KBpSik1EJjNVR9W5GOKvyOauz2OZyaWqqURZ4UTlcT75aF84FmgejiifD4cQfIu8EQd
sNksTVkALoYw3oSn5uuoE2UhEbnoOif18LjWdGSAis6zdBw/w+0/qZuXGYRfbuqzLifrnXjpN36s
5SXv+sCLJnrjZyvFyA/JxJCFiLvB8KvKEoy6nQGnX/S93aLoG4OIw3ABW32+qS7ntY8wPRxR7LZ2
j8xuIKRlfDouLb7jLw3X0UUH/uZoOypyIe0Kqni50AkczNykZVWovAEe1gIFrfwAr7PdATQ3xIXB
t1OR05uDNr54dw1em/CJgKHs6JCPLShBMJquUwBfp8oqcR2oc8JhVQ2vIH1tKBp/6pO5NPlj3DNF
lYhytIoDGCMyQ3d14aG1sfrbKa3CyPOMnLm4MDk8OGYhcqJmicsk5UgmKYQRRpDa2/KZlT3c9a3h
2Jj4ptjq+9FsWukl25kNWm2+uSZLbT4rdaqHxw6elJxqGwd1cvog/pdxtuH5XKJ8E47N4i74RSLU
1eZoFqHbx6PV5gCFVFU/fxQmR8Jnj/VscCv7Hs1cD2I4/9HZ/sA6hKFSoMOyYaXwDPElKr28RwmV
BSrircA/fA5Em+6dZq6kA4cU4SIHs5sfsQYn0pUzeLDsp5sBMRrfhAmw613zh8wnekcMnuNe0qZp
IxEM/60OP3w/P16SutFvyfE4ZI8lilBk7AuLtAungGjql+mm28jgp+Z9Ddk097sg/XrXVahRPRWZ
FIW/edOVCDTrOHqnad2B07cDF6AwyDArwj5PYmPG2J4JrrLES0b2bkUWh891/cuWxV3n103qLKJt
zG5D7pKrf7K61iG1Twdfq3eFOGjMFbuSq73XwROAiE/YzOs3ktnhJri6KgjBgc3NHVuSaAzbFMdC
dh88tzvpkDKUTOiiJ/P7wfrtUc4IkVDcB7YfnlSNq4NpsPj7Lv6221FB2yoNDj1ePvZrKuH7fP8g
jqJ8FWpsJU48IpsNrYUSlc6YloH7J7vXF5lRHnIkb3m/PI9j3ejP5LbJnFtOn+PavY5nCcHdcQMz
TxFYsqWsLZv1RG+cVHjZ//odLUfCF120e+KDuoX8ANKscHw7lAdObN04ju7MJaCsQBU0yCw1giqZ
4CBHNP5lmDIYmUQp5j6q8abaRuvl7kZ0GX+HBV69Pi6w6QOcosOAlg31rVgS4QIbblSv2Tf052Y5
EVWdb4eLQnT19KU0tCyBTs2y+h/SOtBt4skeVxw3/Oy/prwBsu29Gz7FsYwzpHIB5kk6ZLwRKdp8
hXLun2C3xpDiK7Gt4zNeG94yg4pTwvnUDfII7uCXnD4mHo0mAlcRo9UOpPuFXOTp5gYo65WPtdu8
cm7749fmScxgaOM7VuHlPCqKrfvK2VcWz06ckJt5eJpUHGn+nRhXzO7tcRGK3RJcRyJ3cGXo1Tip
v/pA+mHhqkuhTzw23H3V7pJiHG37AivmujQYd7pgyihzch6wea1yIMEmSr9fzZmRMRoiKHop76uY
J/0YZ3nQNciHKSk9JFeQ7SRNOaWPeOG7Nr6qsejuWZyoinTJz/aUouVt9YMT/BNFIu3Sbq4u/Z/3
WrJqCUFIN8rgRjYoPMCDQ29vKrgJ8dK7Pmbw5CiI47G6oiPVaXl4SlxWJbjtolLj81PlgSV75wHp
dkdk26tr6AxGaRSyPP8aGLL+UDVTervQblwryv5xIZmrniPe6c9leGOioqPq/A2Hkin/hXSoMyrx
v3WjpQGYN23uopdhhbwR8Ko/6h4Fciy6Rd1N8UBFhfDaJl3bmKnuG3ujYl2vfq3uSoIbdUTmqZB2
meYxIRCrpuRISEtf0IksUlowQVGZpWuKmglnZKtD92hO67q46/0xdPSx6wM+3a5gQE8LVEQ5BZ4w
ijhKhisupWD8thc1FnbB0xoYFZffjoA3d0imheizYcYkQxBsQ+pNUb75AChNxRmY1Azd9YVutPE4
5nd+/5NruGzZCVL1uZs60ETTBsQdQBe7xoSN6kfxBJtL2XCb+UPhe7nzd8/Nd0rtQHPKUe6CGOKU
6pW+n4qQeNrZija6KIwcEPgQOGQXAp2L49oY+am++a8aVckINMXtE7kfSg+WntJKbwu+yoRea2hn
IfHPMU4+RiMYmLoFfnfNor9n6WB++H9dd5ayHdaWoJuoZ3pKkHYuvJmMJGjjAFPoHK0vlib8PvF6
LXJzv03En/qUR8yPfZb2PVKPqLmthDE5M1efuNhzDoOimFF4w9BopcAIuMc6P4r2PP661ittXGnV
x/v7U0lCo+viG0D3hvtTn7ki7uEJJE2osNY8WK3Fa4/dTIKm++nFOrSOEzy4dRc6kzNREGpLGVCD
O244D2QXvlL5liDg9rqNKkxxKqeOE1O+kl7c7beJyZnH0NN372neaqeWq5411z5ewteBFNig3qTq
ntk1EAi0PoxEYKZW8Ds1aPN/Q0/HoN0kn/beY9Zl7AlBMhGJ6ONlufgcCTNrnSbhVF7DwUuOW4PT
IhFg7LubVFzt7po41CLTQzAaG2z2WCVMfH0qPuEqgAWOzpCPxERfbEDAZiouCmVWqj7eyEje22Iv
p21jqgt4FV6++NbbRhEq5gbw253jwmG/0lKfjFxU2GFek7G6tIm9zLd29v/f/6DThobNYulU7Ck1
1oz0ZDRspmA5RnYD8yDKhGHqwhyNXifauUJktsvicrGxCtTwVEQDmp7kCJUZ/b5ri11rIu0Xcgnb
rmDvPOdA3hZNUqs2zx4C53MOrvtTvH85KHycC3BG7eKu6N7Jco1f+vGgVbGF21vDn/LZnCtCzJDo
TzFPCgnppAtrAGy9sVAr8uM5nNwXGL1n/ZaZ72xfiPG4w98ORo37eN1kPSZJSIDLvjv/S/wFyFNH
zzZZGu8LdgoNagvPc3mTEnd+Yk8Z/TR+CxB4mpYAGMM8uureIJWwgqXsk7P2u8OJUZJgbLzKWQHu
2//YLmb0DqtoMnBzRI4XO50Kwn2E5uSY+SaxoFAqqvjuiJXTTtgEHyQZDorvf/dWHVltt9rsQMfQ
S0csKtGUPxeSzoPEWrilcMnk36ikrD0ThTRBs98xkfFrNZUO4hc6jfk5WMemkCm1u7r+MsqEfItA
xL0/YWAP4Idu8yeMw69q/uclcdvf/1mL12fN+7Jja+M2XBrGC+4gaSzRikfjWjWnEfDe1tDELOt0
EMZKPa5utczEYDOuutO2wp60PzLOGr/F7tgVg4YVzaFmmkNayRzwmECTwXPa7b5DXQp8t9CmauaT
mRS0ChfJJYieJXN0tCcanMHk+5llMdGNSv1tpBspom4ShHmiHKZfIVjsPV4j59sK0Y9WBdPPIORP
Tqr807OcAADZ0v7v7ciGCPFzliNdJ3fcgJ9rz1FuUsV2v4LwGeI2zruGoyib8uWYOjWyk26eL/fk
Pk5Pyggz09maHHGzcaADPRCHY2U/lFa6UA3X1GVUVj6nx6F3vW5eRx8WjRX0n9vqH+f2siqlP0Mc
QYKTVDCQsDICk7N+Qsa09jeuBRbHqnrcpoF/K9grUy+N+pqg1U44gwTXkjMxunxBTgJswAvcNDgT
NR0cL0Y+5QBCs+uQhHVfeKk9s/TDgUeyGNQ00WYUp5zVjeQb80VfPLWIz9QJ8cKbIWB1v+5gBYwc
HtGdtGj43eueSXr86Sn+MKdjU4xi8P1XeRbD8+f0r1ck54bc+zcN2wD7JqHX4l4X7tOEBk3aNiRU
+6pc0sjA4sR/ulFm49FZEaacT3wSRyNaGrR0LxpfCZ0B8BRYI5xA3yHxZkS96MZ7iQ6wOCALIFCJ
gPv5BIHqzr/ZaCNRye4BzyuOdcBXgywu/TS+B8g3ytkGa4ezFjrCkPbchamtIbrgXGhOvFTGTyoO
o6kt9EEzyUwFDl07FLneSDdcYwXFy/VRm+y04n0OnU70Q2+hWIGuNXUm8fO1jKBoJgiGU42o4e0g
HHg4lbX0n0Lur3saIndOFAZo5scc7hBsUWdE//ShTz4LCUTXsp/qW8Q3fWK5rWv458Z2ukLKmJf1
eNXXAYy14mo0Vb98J7vkmkpDFtZuXdypvymVTc2QNg/fI5SEv0F9BjxVm4UPg1F2X0XOrdJFj2HI
+hGdqxXrQI97zRGxkUZCLme0P8W/xxt9NHgBtWbmc+EhpuzMoZ+VCPhoFVMcZ2q9Pz58b6sSLvYk
lUhRnarq0ugQ4qQdQbydvM2+QySJzLkrcL9DsQQVbounWMyx3pDQtdtrcjTkGKL4Eqr9yLyhW9Pz
KZ5te51Tw9pvcXmTeACdVvnugGOKGh7pN85HVVGVUMIzn6K92DSgf5gQVros72rC0S63feKVnl48
00hrC3DsfWqeiYB7IvsIfzOF3qgO3iC9Gxd/5PHw4uaHxJPpXENDrIGF/3E5ZcxkaMrh+NcW+hgk
me6PEHTxZyhXnlbqD3mrpD/WtQUGSZkwAj6895kRd01PeIpnrYwlWs/qPq9A2QESvuFFn0agUwxB
EKoWr/jc33cxfizRMXUrD8FyYoS6HWj0qCw8MH55/AhMizEu/OjCc7GBNxQ1bBjcwj5XD3+NY/wQ
S/ZDo4hMyVop1lWGuO4c3/RlpgaLV0vp2J6RJZ5XlyxfPRzp3qgZDTtNIgMxus3sE3U8bZgRcer4
W8Gcw8yVcMYkv+GbYhJCQUh53mdti6ZJwkyGZM4gAJhiRzuQi/Sfax5TO0EXkZqaow/h8WQSoQwt
OjcxzmMelcGJ+wprRYoFg4qVLT8BSjWWTUX8GpCdmStte4rDUp5qREwZogSkmjDdsg5hBiF95WCf
s6FRTHtV+bO9l/y2XVLO9iafxbcwliI+F3ebsnoHhLGVrAMrh2LJ03eme4u+wPStnQ0xl4ksT3so
hUzfw0VIXfsypz5EFFkW9EUmJmVuGw04Wa3n+jCZf/0Kk3bQbM29uZWPQoJWP+cGXI22h9xpgZze
B2Si8sPH7Ehb6mv4vTILzASHfxwNiXQ39geYRw9bI0wBlK6kLKH0WKAsh1cM3ZLqGnQPQwMXX9xR
e+WRK9KiOXR5/5T/e/6tQzAvYiEqFGTHhuKWpOrAxRh1fObIA2+7HGddPVhwThsCF/Gzi4AR+92r
piWvZJrsMfzRqO0ZLk0jq8nOpld9psvhaerYtBAZgCimrPoowuYS3GrElc40ClsGtdkSTvq3Og5r
2jZNS6jRoo6hU2P6qkr5Bx3uveAL8IyoxNTKfoYNbQ5zgFVpZHW7AQtzHPJf6JJ0vCJv71FygwfF
cGzZONQ8rZppw9xe+mvhdiKGd4lTaTQY9spA9moESoYZWnCSsv6y/umsIzh4a/uMwRloJ8HyVgCF
f3RUwRdnAfb5wgfuGaV8OQ9fognkYOBCxreVPwbdHE45YXcjJGi70AupXlxx8uSaALyQh1j/aW5E
BJlyWC7nxbqAHIY60T/0744tmEoqRWqy+9FK++WQFR/iZpbf32ZIj3bxfzSUBt6WH6SqdArwwu13
Yn4rH3Ce7VvaTjVZYg6wC/rska5HtDJ+0UkS1Qdlm7iKZcMu27RyqtTjkCtF/4TQQYXU2arRXTyZ
/R33Qi4Pq9JBWA/xXa63eYu2lutrQI0WZx5NZcHqaR8hFP3jqF98lv6R4uMtPGcuc8biroHy01we
+FBKeankiKfbgF1QMi+LYbXjXMMRFbWuhEwmRSJj5kWeLQvWQNTg/WUoC5fOKE37oLuLZnvAv10T
BafcPm79ZgYzaGjT1hlFCw8C09MYz2kjgBjAbQp9BONuA27oQ5M0+LHIzFWZNlZScjjyihSbyEza
b/nWcJca45rA9Yy7rk5+gE2v9Np7l7mFwkpuYBTC1BbM4+o+KRK/A8AdVYj2TKfWElN+WTlBGMr1
OPHbW1KVqsV1VaEazk7hWoZKaXM7wgH+5wQ+kk2ok5ado5M3LGrx4aI5QEoHiIUUs4tNnVHgTqDg
6U6/uZJV5q13rq9U8ZfurblBtm9jvLZ4XFEq/4v7hehT0RvitaR1aujO0hk2XNEErHIeXv2WCaHy
IviLxl/UYjgJUzooAqfroAgux5BfVJs80EYXBaIHrFnkIisK8PIN97dDKwukfvSQB/13f48JNp7Z
SD6KXw3de+Q3Gmucm4MMDdFQuH2091I1kxTVtk7E6ONNUq5lwvX6rxbWLRlDKV7yCT1+ZPRjxv/W
PqB/Mnk0rh75CKlgV4NgKBLs63zAlyPN1QetWtZsIbdffzPyCHStYVYH9otlXYgUNz0jpv7rIFCS
HJNYWq2oMKPrN7k6RJhuVc9cRBfYOIkd9NjbrXDpTFJh2nE5n4qLzBCRz/cgVq3cNxpT/Gsl5n/0
7JNqGYjuFMhVGxzp6t06XrSw+rRvVY14y4eIZC8D7pBEWzH5SnTYpk0oDPDiw80XTo5ZWLmguo0u
2RCTux9lZjfj8u5gUE32rQTo9Dk5qvnE5Ay6u5jYbkonZrsNBaqhR8FAIcdyXhi9gtBaOiX/Dvme
ppMQLfe94W1jYvt5SBADnJna5xy/badW6obFkXRZA9IuoLjV6ixBOiRGa1QtT0+/Gx/KKKm39RyB
iT3MrJl7Y+LVnRZQRassYrn4eH66ZRVbjeBbwXOwjL26xuBXZGRht+ATl5dkGHf1uHee+Zmak7K4
nIIZSlZfddE/jbb9nPQa1YOO41GFIJV/PpoFd6ygLQA1hQuyvPEBvnavBmCcx/ZykEd+XUk/hlRA
hmYC/UwK+lmIt3BLQEd6DX+MFZPJFgz33YA8cMAsMgWFT14UUE1BCsrQrbPiLzrtTj+ELEhEYnrT
XtU6NR4+44yyPhAzJkA0Y8ecPr9EZBOMUa7hJzvzWTs7U+8hs0JiE0n8aHaJyIlnk13por758J5H
p4C5qwelsmRZFCaeDagNQYUB+8iQ54C8Rdqk0J++fZ+WPKdVHy9GwEXbYIQiAt3zmoI7MrhEpiHs
Z5rEJLCGT/V8vjzPHB2KFXRFlJfunAAqbzjeWYQHJmPEH19YWnSbLBrytGvx4W8bJDCSnS8wQbBu
MN5Pu7c4Z3sUFej9V70t3gwaz1QCK8LUvJOSii/Qj/TTq8RWKCCChtVRS/E9hHC93B3H/AFzDQYe
3eDUsK6npvBDiUMMkU3/rcVI/T0i6wkuj0iJedAHuH9CDEtSNOTY300khuryC+Miutmtm34/0pdp
oWHibgq+M6SspHPwxGsmDAy9sIKOV5eFl+9THmIvhHLf81bq39UYr9mUs676N+F2VCWCFH28Eo+K
J0Voi0oqNProy228TcjKWMlqTw4Zww93X7GakI3Q+51Gm8UzUS7PX5QDrBoOK8f3Ko9JKh6pq4sI
kcDgoP+UeLq9+EqC114LPwX3D+k/b1t2Itqts7WOTppZ3uomoaEJbZbpzMaSQ+N/Szycsv9tVZ1j
vD1E/GeUNYn7FsOA/SGVx91h8yrPTV9e/iYevYTKoR1EhXygJwipeSpqoLqxlvW4oWZ7HmZl1dqW
mC74kGv57o6zueVkbb+gsnDlll4i1AYHhSelgNbbCzXFw3VaiHD2D9xO+5iW8sH7H2jfBZiaIWf4
95SL/aX633X/pxa/IHfIhpV507C3s3+dEbBfLZtUDg49X0KI8uURYgMJB4Mv2Rn+CuRxMHzhAnWM
n0KZ50FeSG7UgXL0i/baahf3POjDOeulYuToSUc3hpwAisHkxE63vQ9EFUb1ciCvuvDJlRgFpv3a
S0bVpJW39TzuKbuGsQI3sHi9UwG0vJZLD748/nsUiaar80Z9KW156lwlSq4GuDuT88yRo9j3nqi8
6i9mT9Fa8HV69+AXBEFMLKMz76ojqHCNfNlvs4sTUEupd+Hte5rV6g6mBl/+5+74cwin2ni44TC2
IlsQaLXlsjIMUCk7G1GFEgCabkuKS1AU0klIx94rqSJDwQuJhRA0jrFz80Ov/EZQoYBj9dFN1wY/
ZAyTvr7MO9/LQ3ZxFmayQk8SY1Eq1fMQhofsujGT1aVyRR0oQ4LYSRxD1RLMblkyS5Qvj8hoo7Ya
Wt20+AWaXNpEEj0xXyTb8BBXkvRk4OlXrHWOzHDbPU/LhftiIeVnkEUUEOgZqw6B5RxH5GfqXcfw
wMuXNPasTOME3YdHc/q8aw9yIR7Bf3RoFYoT8ButGC66MFoWEaULmKbSHtYI+1w0WDKFYcp382GF
8r5RIXUSBpKStDSvhOWZq9Biaskic91mJW9euydeq39RRty8qmhTuBLM4HtSfwqUfA/XwoN/dnxG
h8ib579rNbViWPTxmBJHMOa3Jsfp8kpnW0qvoTgvR95lZeuBrmvIkSb6j/uCyhSc/+HLIs4LI0Mv
J9NDUP+ZX39fQTzk7pnFBWK3Gs57aFPKFOjyQlC+CLVOsyosn2IdE7T7fQBxs83R7a10d/QHvtJ2
jRd06iBN+J9CbvCEuYxjoUVAbMqf2SYsvV3mI94gA+Tj7FtzHzSzyVDcmqREL5aiLQe1t9dOsBGF
TnbawBpiK3Tmi4vODca6Sge4a6G4r1xJvhQtW0bAeaSimcRkiPaBRED+PlJTpbhVfPqbiZOaXlqM
O6WIqsjFF4tJoJpV+9A/jzegpT4KTB5IDWQm3zBO7Ti3hqNwKHu3KCRLf8pSAY54BYCK6h9Q3ZDx
ANGBIHGi6eblviTkRhsVE92HaT1UO8aAZBgaw2H4ErsNk3MQ1wPcx0dvjfLbIh58GF7hJyw6n5iz
IKsW44bBYfZo/UAbVRC7i013yKoAzsueV1KKivKxdKfJ2zUlOrM/9+T9pV+moc90ZnSiyISuMRvh
vnxwK7SeQJBsSfgqeWFx/HxbhUDSY8tqlcRSftu8ipTa5VTT3CL5j5TYZwj6gn9o6laXH0trS7Jr
d3yAYS/c7D+FEQ6aNaHSgvpZW0XXDBbujXSlWK95xYJF3IFui5aM2nDaJRbtdBLYZznCpYSEHMz4
Zc7kow+UVwILPcw/tWT/ZWTcozpCOXKkCUIry78sZqPc2xtDdLeDJQXfx5puu+L4PAiqU7A6GGYV
GNL64sulvjkHWn7d9gPxIgBFZr0hv4Jbn6f0ZqXtPsPLXPgnPEULJQaYfNyCKWP3yhJiTwjexkKb
UILwiCg8YXF9oyb3SP4Y8m96EIlK1MQYmJA8LJxGq85gBoeBRa37ZvyEGvLoInU+hvslPb6A9v1a
9TDOykkpL0xqW/WsYpmY5KNde73PZT5J2WGbDqg78TlUKW/gUzYuy+Zw6qnVtD/ldm8r6YeLQtL+
rej75TSrL+aXAuyfV0f4F9D8vRO2ik2uZTQzTy0vVoAjFPB8XZYQA0kRh/cJt5G6F5WSXfViwFP3
CRjJLSL7WWb/+QqqIV/vWhzJFAB+UOOHtCF/z1pieGe/Dyo2JzwOf6gwdSai0a+GBg1a8f3khh0R
T0+/tyuvDs8QsRV7JPdIHydIQ0bzkqa2vXa3GhG5PoMrtfLrSWJmE94R3SHK1jBb5kIpxTbBbea5
3BnASX9Or8GgcCusE/rTglw3CK/FSM8D1nMJgIfxvIII/5XbhaJiQngaPopgJOB2de/DbiTsikrc
5t/475Y1GCEhcwmAbGkJpO/XK4e/y7y9KkarMieaNsWenhe2jdS1yk/FbwyV2STQv9dY69pVtj7P
a6/YQflhhsITnWNJJyUHSVHNHrLmoI+fHigBk5SoeN2qfmT0EONwyKKhq2d5/bjl8boZ7BFJgzG9
fFbAbaCyxcfIhVm5tSW+AiFIXKgbdyeemw9oDpYPsEEeyqhfDutNUIkVqoK12XF6lMWTtLXQXX5M
3MlszW4JZggiqonWeLxktB9BRyRiPm0112KTYHBbRDop8lwvndG+tKir7P7rqZxP+KMXZndDNMDG
0J59a48tPkTleh6EtkyLIZpkqarMEVjkhZXbgKLfWBWAWziGzSsw2QL8nYH6NBAIQNOh+Hr0hGyR
DOGlf3rVCAI54RgBhswSQWXyotMrbigHhsWzIX4h8Uc88Jgx8afQubvKKQAw448ik1MhIVt2Icvm
UMf3SEeQY4b8DIGmXJAnb9G68AqPTESvDtQda8GgBop/eKaAKUkbehLd52lRDLMkgLRX9e1+F2b4
Tip7QEOV8ZzIJylKa4uNUfM1qRLd24CGxNIcDyU0bvnpYWgOBI6lYJKYx94nojIBau1hvawyx4Hq
gF76HevOL47uNfo4KibO18rRCThbt/uPyHMh8IMfGoF3/1Xt9EtdK6QKSz8JouBZZk3qgCzhodu2
JJKIJoiXfU4UR8sN8L7WXaLua1d5PzUF3h1SPOBaSeXrJF33aSXQPq/93W9sotGXZPPZsl9wpqPc
U/5JItGHhR0C0Ln2njYeAEKyfsScyS0Cv5LrxewuPIOA4XX8K0JXnqrP7hSQXpP8nx278FbOl22U
ZWA/O0bd7udyBu3jmlTyBse059Iuq142fsNs/jQ9DnTdq9QsYMeU74Baxk+Sh9u0qBWiHItHqZ6d
2b9OeWe+eGSQ26ZOWkME2k6mYSRQ3HFpnU6FxSML9+FyyP38eAzNQTy/DUiN8voBCz5G6MvG7q9M
Toue9yJ9h7qLoq4a8SZtR2Ox/iI3GimCHFZH+y8Xgir/pWXceTSXcIcNnWLvFX9a58LODtIXHgmc
BplAIF6RiQiip1wiBzYmJ5aJ+5CfmHcfwhyI0OxuTmNUXUFxvG/bIg9vl6/fbpiPH3dzeQYTJGmO
T2IAqtq81sbB8zWvXF05jYCR0KcrYBDGryX5DfQfIWJuXp0eKkrJvk+1eVzt73pmMIAQWcxSmxVq
HIvmygi6C7HTi7M69ttzYvirD3AHWIDdJaBnn+z02EA2JbCeP8v6z7io8Bf2U/woMJUnVGwZ0SnH
nd+c/Y1FXzUf9Ms95mXDenB/wYbBU3RRg4YR1CKhi5NHBqUpGsfZYdhm51bQVtSkGQqiyKkq0QsX
6GFPdXVkLXTGAWN8CBMz0ctyM9RiS6jMPzmJMCinNycYVtkzyuhuzrFrI4L/L97LzDfMaJxbyk74
NtDCKgX2F8Zkep1/3O76B8JV67tcivb93ToGsFXupQ7Jab+ZgNtBOKHh2uYN9S42O5ZpJtDZGerJ
HcJ1svJl28xQ/CIqOaygdFhCbzi/ifxPK+aIrJkAQCksXlKNrX8v1YTCvqetf4CWFQhl5A8Eo/yp
6F9aPN0LjXFLPH0bhOZDaEwjh1foB7h9sk9On5IliQ6QEaauDtrFeRMdnxf0fib1SPoF6cZwibW4
dNuEL0ZsxAls+w8fgjsFkYkTKLmqzdTN9OyoVT/HfqyIidvOw604aM9nq7AISw65spzQ88qcmzLT
ZthQ0V1c+PB5Xf9A2JUdWUNHuRAF6/Kq8PPPFGifMO7Pc2PEqaamWLlKAUGIdmhdPVK54ejiJRL1
YvP2qkrnuZVBl+M8BJLgtC07+SdJpPY/IjLIBawISMp1NGHcq7niqOW1GzTyc3ARJSgpa7V3nKJd
MuuQChrnZyLD5B1MZnchVBszEO9z/GpO2tgbnJMs2H0lmAD88LXXCAROGyv2ih7mO5wjP0dRaBHi
C7Ly2Tbe4zEyIF39K/n2hwOYEqNOsHJqj3HBdpjJcii8PJfmcKph/EyYNKWJ3gEwfDOWffhibW+K
fnooEKQQeYVXeTjscSSsBDJ/LLxCkfRqh0CUss9eWz5VKDb4e6ahO8lHVjlPAMQt1vAD322bv3XC
TAQLSn8Za4E72X86F9O0EXM+qXhoJBZKOvcrk6mMiZt6vfCEX0ZSY6O4jIjRxvSYRltEIm88Y2SO
A8JfvXCbZos+8R2nWWqkn8Y9F3zjuDk9cwYH2IVigkak+Ft5RmfKEIxhPIO3/myMTwBNgFzPBKzZ
keztsqI/H5ScjJ8GLIwitkfiZBXnhJ5TBfmgSvjb/GZGDM7uR/6N7WsNIvUWCXBP1QEpeqKMPtD6
Yn0AkBMtq7zpMchHmZH4UNRrGfXqqbtvGVQlWQEOieovdH3uTzI9YAIxAAlXOrk92Q7YYI27t3o1
Xeobx/pMkzVBqERx44rP2VQAkuerPO/q8+gmIWcPB4YVLkrP3yjagEVRe/JSVI2Zs9HUg90fh806
gcKqM2Ymp2gijCjB9p9LjGOKsWLNeHRhst4JC23vXiZbgElqOIYBDXuTaNgc7nZIIGSwSEl6REi/
+WwC8U2E4LI4Eq3aC718957ZXUXTMXVaElLmPJX3swuIVHMvUVg8GNTwXB+x3/Gn6QzPbzjsqMun
9FYXcyhhiT4CWj5OD2jd69cY2/J0cGcoSyHhAT4s8tAAL/R01ef2ot6E+b8f6mEaRB1UOSeH7B+8
eSNhKV3S3LG05WZ0Xj3Wz1geHjVYCxZS55oHDDK2U8M7Johchii5NdK5aTsWLbJ8QMi3lbvEZ0UP
DUQShU7HwTDD7l2ZofS1GMQdNEt4v9sem3vAMMJ5fz5EVOz+B3d+G+4uamYHQGRziEAgtKxxBiEf
AJo8UvR6al34Ls1ipwXglb301NU5k6Pq2nH0IyjZ7mJeJsPVODzmB4oI2YaJqdHPwdWE/D3ADQ2M
Q+D3Pz+iZlmgZBiIVDbMzQZ0WKE598MGsx1kH7U7ViQXjAZgQsoKnDLrNcnyd0vwI200cylnf1UG
ZWfUOyVqx5aNomyrTNghvBTc2jUOd6ofPNh8bWImT5rHY7dgjqJN/UTZcwALrIlkAaWHsCV56Zh/
rR0Va4kb2sLDUsVrotPakxt2Dk48f4g9VVMijMFj28DdIrHL9Oh0zl3SO3yNit+1aG90LOhzlKEE
X7k3NXCkMKVdBOj6wadA2Tn2bK3xkyBmeE+Snaoq56S65ApOVC0W9BdmG4pT+9cBZPRilkHAxsMa
DIi3Cis5CMDkQj5A8BHVGCq2jR/wN6/k+y+ZqoWPIsfDCxG9HQ1kUFWW2bN71iIymyDfFpdrJpuT
qtTLBlaVgI30CirJm1V/nR65KuhY23hQD2FFnV/rStmMQEs1QLL/2NsXUexTbxMgI12Yh+Cc1Gnw
hkTbWFBp5Sorq8P1qY3U7qvVrJpykj85G8BSX/FjbQdJMDtOY+GefYNUbxL2HQV6iiV9iOkJgPqE
Js2G2pN7ErnuLEqvSsQfwVXxzWqhZlglhBqWc25ZI8TjNm5k3YyD8z6iuHLR+gWqLwn4n8K+mCF9
Z+ESxqR6QyC7CsQMXL2lvlM28rBDqVbzr+pBIYjVdthSRddXn+WL3NqIfwHuAA3qBPwFUfTQQWha
xW0p/UWJChhGj2111CQ9IRUWXapJ1Mq/oeSmihugDfTAA0nQauJRW454bDkTHUYcBfop5QJK6sZn
NA7Ps16toYK9U4ZREC+odV/DH6j++ZVrzHz1MqxxSCmsvvri2tzeug3JmBLWhgZCvyrQhm3Heyoz
cU3cuvd4NDb9ZuC4uYtH5q34LLVNVn698CaNQkKexDLvsrRs/Kzpz0Q1fsu7cJFcn+4/0vwojpCu
5XwNj3tmcH4MzzPYHMc8WUHVvneVbCsHWqSJJSXUhU4u5THYqidUXaoIVBR2+ye9CWV5hyjD4ztv
3kB71nVvlijst91xhFCxm5YNyq15cznGnSr68H3Er3RT3SkDarSEW6+TK98zF7kbZ3EejW8txUV+
gIqByK9Ss4TA2eBiAU3qcPhjkDgcEvRMcmiN/xNrbcLd84Qkt/lu84IbDV1EKJac+zVhBPaCxJXO
ZrtQLumnw+wzMThc2NnGUhpHwrpV7gayYQZlAVbXGgfpILtPZ46s6rzOlWFRbPXxHEvp53XU2dsl
aqnv6dtULXe59Kzn6VigY7s2CJbLMnvLk27mouGTrooFq56pKrmFJEhy2ieF9VdynDc/R2kvuccR
MRBKNmqu/8qDmm9Zil1yGlPY2Dl1p3et4vqydiSajYHywSqBMhSYOcvExm87vnHeEFe1gWknrC7K
fk9OLMCyx0BaM45Ge/WP20D65HPlWCSpMGdoKMjtVphtTqaVQ6R2Bfzz2tzBlLkEhX6polSJD2ks
GUvSmtPqJrfE1O/9EvsThYh9UGmlMZxLIzr9JSacfDj4vlqiA+ergSSS1gXxq5XHusBKH34kqPux
vo1tfgziAj5tCN0eMMNbrtj/WrKEzbN+7fdNKdChuBfPdqyIieA01nC5ChTy8+lS+gkVw9KoDS6u
rZG1Lyh+gGTakPHuw7qe4Ijz8M3WL/EgGvZRfkCo6OmK7Kl3nZwQUaKllMUEnG8sFEEbeCelHaUh
JTPx1cZB8S4i6xL8z+38WUIGKTxmrTGmSoVFgYn3l7+12CxLOzdeWsGq2tsJO2ZS7dOyQmuyYIJ3
YqML0nqm8I/zuSpMKknU3M4zvx32PhRGRFQoYw4YB7KZ3wIvAHSV9YZNf7kzZT2yyLtjczM3hNLI
lXLhol+70GzDEaBDmtGlP8/jGRgZY+I8+8o5kvACeGF59H71WkCW9Rzr/wqfCqjItJqoPlppyMyz
lLpDcsmtl2WVIO2t5f842/+wK55uJ7ds0coDIS/CT905d4Iqar2+YRDTRHegnl2Jw8S9ihhNcQ+d
NDpxRkjrcM+3s7Eva6p+3a//UkMKXR3o9mxMaseZtrsoJbTLW8f/zZ/qppfUqQ1Zx+d51x+d39MJ
ACJuzhmw11dAaCmE+QN6aDIGCE7qIfe3+x1S9ciX5iJOZUZqHmB8KvfLutv9JQGgm0rjKjgzOzKv
ARlzM8f9b3Rbkncw15A3l07CTwRvsGnyFj93Mevh1gAse/1+Zm8qx53PXI1NpHfLZalip9DNrD3y
B1EAXQmZ/uQsRcFh7NvrwT8E3AiPFQ0ChIHpeybYyKiJrBZekz76MwqzwgmX+EyI26oOo48TT7jC
1MNt+tXaLM6UQ+8SzZV+6EQHnBOrijrkDKqbYCZ/9yY7INHK/5BviXfGshnhRJG7q+u5hnT22YEH
HtihLaig4lZyyp5y4WmwWD6xjBfNTX7/UfCPQ+w8PK1WEac1GuojJA1vcwN7WFfoFF585pfFd7yC
dlcgpX9X7yH6AY0VyXKXYrjarRWRXzjfg9eq+KkVvUCiaWqT705xY9FIrJluqzxpGfsaj2v5D1wM
4U5twpsHPstpHGMcedR0ksJzyO+pJCe5lwdE91eKKl2AlyWg83r1lSw8NsYsZCkCOz3+sCqvqVQh
26GWuAItOx+wq/zrwWPzP1WSAPNRQMvw9MAUbYi92kMwm8uOXLMa1dlSCIhiQjvr9nja7LEiT9F2
yc/Mv18BYX3Ga766XXkZ3zSG4GnGpNbpF01prBU7ib+D9BTr4a3ajIRGB4u/qRsuuWJaCio51NME
UjWGJu9Ai5nvHVEQ7fwkYAOgnzMxubNyGmJyatMMLNGmKTbhGTuSsqcLBcbokE586P+l8GghwrRt
ulER37kd41Tn9oxcXqnkwvY8xv1cYuhQ3Jurt7JDs0y5+LfqKTE0XuwdQFzJKXFNRK64U5pOB6p6
nfWVXIw3eBCe8/ZUUBWxlRpLHDuYMZE9XydKzeJnME5dc9xnudB5KbCsTpK74ubwLs08UHHN7PJi
nsdzJPSDuJ2t+lbSl6FRpiqxBU9lPuN6Sa1RkSPIORx4xC8ZYnJUPj5VCIMPRdwjec8JmznEMCRD
IW3iIbzI5qB2IsJX3qLiKx2lBArhSIrE+pJNlwEr2t82u5Pu5uSDMEkTnDxCaQkzeP8Ubspbt4z/
oAx41XWzyEsDZRAQ3k32PBcdkfBKqIbBIqCraGK2w7YXlY+r1Wg5xPQeZeQBmmAvXIj2oL2Fm3Ex
0oCW6bYh1GNbRWOc+y7d5wczQF0sq51V9ZDDDgcEpB5QDgGMIKEuja6+h8h8EswujKnkzz6GodAu
1NbCN1dxgKC9C3K6pB5vANIzmhPtnIRgVz6AJ8SNq6KS+aiTHQAJ2wuyWgkR6IPtDBmmyH/IGUPU
LgDeQqvb5LzOXinrQZuKrp4q3Zjv8YbSmnoaSx+L+ZuvjK2ayza39UoNWvK4dd/4Z2Zr/gPq9Iy7
Khu2e6lfR/IXrGnCqnsTD26gsuOpPYtW+p5XMGZw2QAA+XSfg21TCiZU54414S0hUltY9XCGmStv
I1FAhw+5kuZxGBkwrD6NF50ivQEgrHw7IE2jPr2N3rQgnkp9Ex0wjIzdxY7mADejIc84C44J2XNg
YKhKXaHKSy1y0OrxOfwIhmhl17zjLCrEnz9KY5PVLbdzWP+uZmfk8SI45taATAbF/t+uS6xu7WTd
QgBg2ysQmSqAMWz9Mnxr13u1wAzhgq19jgvqq0m9f0NhgNAfbr/MWOfbARFu5lo/tQEM0UjDTi4c
QRhNC/rItSbc+cL0uVFtne6KA7vfO++cpTOJDAOvRvDekCy8MtjEj/aXnzzoSoAWr2ni1z4HimCg
6vdv+hzQwwRAeUBzKPE7Hn3+oljFPnGl0WQs53+OJLihnSN1Y7NclnyES4VdVrKBqqgpZIaYWZAy
zBo1Uva+YGuRrTDIeOUPFYNMPrr3eJ+0h08zhFJuFauOJWFMwxjjpdmWVBM4P1BBBdAWkX37ooQj
weZSMzWrsxFaytnlYivehsEEZaG5S3Aw2naoq0cNyuNBBx7bXJy/4172jDb2gHYhUXW5t7CdD8+Z
BwMyPig/ohgiR0BidRDxQb4bmMy/05k3w9KL7LHSYTxuhs6YiERMT5T7ZQjhQiaBV4U/stkgzT0Q
WWddRyWumH8ns7ma4anZgfIFtITC0AbAmMV8im8FSCYbTbgcuK5TxMFX3YNrDxASpp6YF6iO89zW
DylE2DsSU9T4iIHSN20dSZL/CNNVYMVick/0IJFnzSs+mBWcWS/Y+fr9eZIOl5GQI49GroKJa1J4
mWxSU6s5gLSKZfIiMzlvOkiBgWwyWuz7Zwwhj9iNDRY8E3EBGEAkE0JjD7V/IqFI2qq2axQ69M9Q
ddxbE2SioqTvsGhyiJflvSxDZMjY8ESFME96xhN9vAk5NryA+v8aS7ZsGPCiQYI7hEcghAejicjR
p+1Ra2GOoEh87YMJWWGaUaOaWGvB5htbkC7AkzV7Yt7zmrz5nwwtq0VSb9c78msGQKeQEOVCq0Of
tJe0ZToCPeAYLMB6n/c8TME6UIn6/RrBctCqkucjauRIhM2KdqRqw6BO2938IpOD9LV0cERW2N7b
/zZvMnzaEIkly4wL3UW6ZHIz+Ae75DMNgaUslElYIhLa/dWsAYMBzhldQrwu1sS2YLMuUtC3gHrz
dUL2L6WMXKkVsf5NTAbtdzz/mJt1dHJVfbRkFRN3VOMTk3rtN0IfVauT6S0mzRBhFvBBsK/U8hPA
h3hjE3Pm2uhS3q11cSkpcL3RXnGJEiumCZYlF8TdHWdbwrl5KfjidVzAZCbtnM0l0jxn9ARSauHq
ljK5uhDlnACtEIG01cEBPt6yVMw/+IwwjbeOdZjP8MiRlSDbnI417F5Tk2wqiWPdJF5a8Oak+sZS
vY9M9Ugx0OxEJ6tSV4+xoCn//zpKThm23EsJvLrGpDiEtk9wd6tDEFZRhhB/ggMsJFJqO1ngjC2Z
aim+FBXbxcSc164epzLx9keXwcSKJvp6nYNRdNUKQXcE/iE2UVby2Q3a1rbvt4Pdo0hYQE0fPq39
N/TEwNvBB9ZV2cf6E6ZwBpPspGfHqFlU/DacMUy5w5ajxS17Ad56huzLo1MckKaQzH4SjJYNvtrA
oOuLIhdFoP5cl/XPsiXZZubQ3Q2YYNprCM/NUVRkK0gTI8f/KYluEBE19wRh8omtKfZyNWost2hi
BhBRVx2JL4BSCwXjBE/D14RV+Xd8OcI38oD1rHak991fqttKiE4UpgRJoljOe3rskrAyJYrt/T53
lYeEv1aHHjh3Tdw5/ufoP9Mf1dHm8zLp2/FB6T1QvQMaBOgrVUwXz93CNnnsydIPOTr7GAEa9YJ/
ZhQ+Vn65g+WLksx5Tglv7J3Xhy+48jsfkFytAvuWj6kQbJuPS32nn3r6A0NV21LVWjwNSoecIvy7
8/zDcbqrEHrPmjvfz+LtMedsDYBor8B8iZnF0B1lWn+GtHcZs6rWHrZEX9dCvK6hDa9kJy5aFWtc
/gSZ5r3p0GayqGPNdjH2GuJbrtXxCNhjIUegD1X7ANn/sPwVmmmnxAQCaAP9kJ3cWMBuQ1AHJxiC
3CyTN2Eq0q5MBnaHYwxjbSzek/CTHXRffspdyqmXAKpmLGgWOeb7mXd4enTQOXWAMQV5UOf0Deoy
Otblzon6ZXRM65skJKYR00YIH2DEV+irWh83ZKA81dObelsKpwI7eIubJnnepS2YMvXPFXNMuLjJ
4mlTkaRtzU581pTn0/HEvRzScbwuSSDHKdboV9Tt2RoQmSl5kB6rdPo+vFheMYNK16+j/NyGuVCk
PLCINt0d7GNrMYcudtjU0t01wTj9zawb+V7CWetXh8rrA7FhARVEhujGiKLg5DMlo60n3KYpKFJp
bcWFduNjg2zJt0FmyK8o6LLfzzU4EFFlAOK3fyFMKgj+Sl31g1ywd62qZj1AtsaUyMTb4dVV6ytw
DMHP/9pavVm3jcRz58BygFPejSD07Wj9pEzDIYq6hncPjd6dnwQ2NkwYsYNmWdGIIIcp+b9msXrI
Jw8uq7aDRDbrgpQRrsqHhiN6Us+U9/jSr9AG8uyS35a8KPajau2zK0VDpFqhRa2Qi93nDhhnqKNe
NHrBWvWuReKAdkha/7Oow8BuqYUunxPRabyxeSvkhriph2sy36UUuhkEpHSjT+xcTZeE//n27QuX
26010L8leYLWveyspdPc9+CdM1JbIZ8CgFTF/7YDrpxqy4XlgFnooiaxnzJsA+Lc2tPZSBA04xXG
NhZyv33Rx3PkPjrmDqSH9uY6Sz3DguJTI0nwiebDnkFrnXftWV1ol4nWVUMJ+KU82bEsBi4iTw01
ZbpFS2tjh5vICXeCU4MJvbIQwbvAg3+dmPpl8roL/SubdfgbGcDKlzz0YPQ4+4xnuxp8xPguniD0
f2FZwo62VUCX/qhOUbiebenvDlk8X8YOp+Sm7wlt8M1+w2niZuVV8sq54L5qnlaniaE3e3SUpMAp
gO+sonNBGqjLGpiWD98FlwUrusqkCKlAdg3bzt4FO4nUxEsoK5GQB1exWPquYMEeezLr+EIWK3L+
bMUOcLEIeP+8W8SyOfJbAE/jy4iTrHSrnEzp7K82gD4ED7j+sGRKzlStPoA7ZPp3iCONibV95h0N
VjkSdKauS+e/Vzj+oAvI6q0gyX/fzYeuWn5HlrmT+tIt5nAHG2qy1FZ9gmNoSXorLqbImY4Cbsam
lpq8JMSrRc75P+kXuETcVcCLYpE1iMhqdv1HRHpRfyR2HMj3Ukk0kCyNla5WjLK4SV2XDR8dDCKH
tfqos7m47f/OgBL/0ezgEfCUeWXY2mlbOfUpp2z61cjxFTwc/F1gdVD4njKiFPSAOceB3LHrD5Cc
cQos3spDcqfdup24jXpReKPB/cZP9nU+QmJEip6Qa3NhFdz4kJoGO5zXoQ6ELGvARVp0koq5kRKI
jOyrwRk72/2khIe6JJ00f1IOOETydW2ofXLY8536XJyr0o8spPvNeM13myye/2PTJIzNtGnq3zmf
UzER5iGi6KS8nChr4KVZ4lHaRna5UGzAL2RtH6tCS3Ths+taWcSn7jbAX4rinkwcn9iJHV+cK4Zm
ZtD5TJtzmX3LM9uek5Mpr9d8fvmka4WycUY5k4qnvq0MiYs8elgS187pmkLqnFMjfS8LQDdLTCmT
a2vcuJcTAfb7ucQACq+QeF1AcQVdeVSunCBENXf8hktEtzFCk3NeuxHUH4OrgGHyIKiDCI/PQAmV
9H6wC9QrdAeL0lNiP2OaowRt+VzaSz5CoHfamGliAO5b77ZdDhGJQnKtuEICbbVuwdJeEIHSIjnR
+hIrxBpAuXlNozCBfG4dR6bSzdi6Oh6QLRPa3fp9v7kpiBy1Jmh4sJszI8nRoYzTymWsB2LLjT9v
y8WJtcN1my3xmelee8oYvdLY2VwsRNXFWPl1jE7lj1z1GZQdwL6LmNIqhfxMZzdT0vbRFac1WjD7
2gC1IMwFURRJjfR0l76arigh8whZAtPHNwV4SuNCenXnXmsvnZMAj+lMI4XY8ARsfldchYz6QpWg
7aMnBcwpDc7UGxKwieZ7E+AHrBGlo8R1DJN12WsV1dth2mGkCCvtoUrMhowGGQR7KZjDd2sm+wEd
4/Y6f1ql9NSaqQ4vliROVFdIZ0ZUhsXy5qgeyECpaoyjQ/c5PNzoeOqhe4zGNKeqHdQZrB5zbFnZ
qoWbSP6bYucL0ngONc952ryBlxWhAWej2SJY5xKrg91TCCAuh5lfTwcxzSRFdVQW95piBm4cpF+f
nRvICPQvvBSlG63e4HVY04oJoa+G+XWDoXzqf9nU1vm9/lIM6OWRsigYMnrSZN5ZIAQlqcu78QFb
Ph2MycMtl7n6pjAGo6UKGiuiQ7VO69sRTp2GL+jwA8gEEaqtbCnr51iTovAys/uOIkZCzXgD0trv
gVxoePrSbQaiTD6s2wg4CeksRNftgSBwZeqQGaZhm6MfE9cYiDgwngO7pQg5sy+LozGy4U2UY1iD
VCVCzP7ChfBk9K/MNM+qRavX6H3BStd2xx3QicsoDIpf2JxNAeh0EC5BNOqGAugRCj5C7IlBuYxQ
SVcCu8L5EGaPIJ9rILahIyRX9PI/qnfQCTFP6KrLsw4xzSUu+LUswtMIIPc5jOrjo5af+Lyrcj9J
6Z6N0N3djt17eCw7ugtljpw+d4xYvviwGwhOd3J+ALflr8BMh9TnSRVdlgX3NX+erqQVoWwrbVfu
elY8dIOQlOR36W1xfuhUswAkIdOPFgoaS5YCGBsTZSeoXbuITOPJssT6+N0qXCR0LaRXjgyU2TEt
BSPu7bhBC6JZghDq+I8dPPdhzG1z/B9jDVdD6CB2PJcCLPZedkh9o7msc5PQksCRbwCqIbgQzMMm
kBbzjX+W1a5xARKk5CrjTfFzpzRWRpa/Gsp2+I6Rg69//5DwKyCPxTs5Df9yQftbVM5myntHFD01
w7S/xSpFBx20g2h9vgzq343U1cnCw1Z0zf7jX0FugcVpSou+AzRNa3cV4rMRbuhavE19QWuolwJh
EYKq3hN9TykxdhXT3dp6Fmo2kvfDHb9zPpFJiJcOvc7vYG6qdsYbSvaKCH/KlgXzHiXlJ+KP0KrJ
LJqPu3WcA8rRRTEbHFAolVqkZYf8M5JYXvSRDPCgPCcJ5iHeQshxmX0lleegOz3P6njmm5Te30pF
7LhuEhanFN2LdqtvRwL95z/TjzS8tKhL58WG6QildSTebZ/CPn+MQinxrbBmEojABmKgIeHZaRTB
KSGe/sL91w5ZOfyDGk1B6GwRWQPfstDJ93wujgn3LMuK7IHX9bG/MjwsSaEhD4+Mlm5P++kvzhOi
L9cEmXwWdm4r1EyIXBqA/MlaWtkfmz6Qz6mxTtzWejQA6p95Spb+8YZ7iYzvM02t13XrimjOMBU3
yJJcIQZzgNsRlWmqx5LFcWvShjviekhIyN1EOYSy1cA8TnFMbcLB52qJu+k9aoaKAON9KS+4S9k/
NSOnmZCUXIycQdbYe6I9a+CRuAgJyOWiuxXGPe497io49BZaFWzO1ziu/khUZKFZY3zu2qVH9/wE
m4RWYiwcxnpVikd76c9vpjdtiqUDTB/13mtC5GHxWcM456j17u3kKih/+pX9d82c7EjckMzU35d2
WSHPPGq7GX4vkED/vU9eg/Vc3v60TPL5IX3vbiogyTYVmco1BvV13ZWbCWwdn5BrpLeSV4Zx6DY7
HP+1hhe9/mUZWiFV6XrJ0CDy010nYLbaEmZX9F27EjB4zpqK4AiNrZ8KFdm2ayQ4aJ+tmosHuXHH
qMnN06X9II3NT0HrJYW4/UiLuA0ns5B3PO6MtJlukviymBna4B8N2gRCWe5nWpRw371DhDKGiYfZ
2N1Ah7Gr8sAigPHFVZF6bNrLKR+gQcXP0mVawn72kGNVoeyzWSyL/WsRSK68fKHOGG2Igap/BE7Y
tIAI1KDzFNPZ3JBDzyraWCa99gdh6HrGEhMM5zQYIMqu6Wy8Ae3Zmag4ncFSV0j5IlX/eo4hmChz
tMO9yDWTAp5EOPMmpA3t7QmsTtbqMYar+/2t5JITey+KNezpq9xI3xz4zDG/1Nyo0H/4eZg/63fg
q+Re4vZ0IYLl86Noq0W3EMCZlAdWGjVieBnF0/IdL3lYRFw7/1A+/xF+0r3aJajCDJ3Ty5W0S8na
8W4ggqJX1a7yH3phvruGX5PtDkGnBlzctxRuQkHbE3lG6hfO0draKAKWtp4u40ljD07qvCqqp6l7
53wX7rNLzaby82YjUrBB5+KmUTvu0jrXhpTLZ2wzNE8Kf/b6sKRhlo+SCqqENWybIiPCBjhrrgaB
hsx7hehuETqXcvxfb56LNgEO3KEl8kcLBRSZoLrLmZ5VQqorZ8lloNXsw8+170iAGZaefHh6FWTf
P0r45J6/qdEGvLzAqvTikhNG+1itYR1OZnaMGNuUbaLiA/iTwRlnGUsW0P4iz/uwknRk0eBKMs0H
vxwILoygYfPOKiYunDtz75f2C+g0JT+6uJAC9zL92vSvWvx4buaWGooRjTby2MzYH6wgIWWBAPZb
+Pzf9uemAb5H54VxNC+F8IcdnYxMkeaAd3yNifxBdUs19LGKZI133Aqv89vgzpr9fX5szsjcr+FO
ok8o265xkSiCxXd2tqqclR+yN3BiRKKGS8EKZWT59Vi6KnS3TeSvjSEEg1lDy+3yyMcDYx4FSYbG
roq0M084T8jqhSRtVtF2bwaGE72bfe44bT/RBM7Zljs7q0xI3s/T+c78+7B9KpdTI1ggmEwZJVAc
C2I9ud1qKgeqD8w1/5KQ/vVWWGhGjAIA4Dun/OEGTsYCtZOS7vqQRSb8ACOiEH/ZiPH8Ylk8M7n4
xGS9hxfODnhrT17I8/vFhOBZjZ2IG1SHJ2ceZmkoDTTDkZPg+eDjy3/GVt+Fr5pF+bX7La0hoJek
fZJPYKDOk0BnQwIifb//kw+fF+iEdmnRQ2wP6cUvfyePxHP3Q2NHSZ4gF3WQoEeUfYl+FHOzkeKm
8CJrxNrNRRTO4LGJWkTWn00DxMps+Zb7KVeIcWvFYoS81LIv3vImxoLAz7/9SfUJ/DjOzmCr225T
js+Ddaq2mKYuNLfcmHOBkITGJ7eeMgSCIiEOEfW63y6YmO5KYkUN/srYBV4nLjy0NgCWTFbqV5mg
J4VpAWTk46g9rxFgv8JPLpRp7nEneHHgCkAALT59kNgFOQyr4+ocYGn2mUGuz3PR1NLnzJPhvJ/B
WFW9LMuzY6Y2AtOYtVUj1lTYyQFnofFeNUizc0iG05m8jA+cypDGP5pOK9UsSwT4A0QhozmnjggA
cWFZyGc3uU2GESPpws1CaKKu81Yt4T3oPPiFt+bZCIHWYzq2tTkh/Mn5xkRtafDzz2c3X+EORJej
GTPB9wAth0LKRFFs4r3X7qMamqelhZd4e3RdGkv2TDXkcBTELgZQ4JK4zWZNr8bng1rru0iPfqs4
seBTxq/FVbFzYEJdfTVoO3g2/ePD40WT5Iask3be9vLoI3YlqzRkjtC0CPP5wW8mK/7KBFKiRrUs
OBWcF31YaqwquHDHbli1MQZH0qCZnpLkyDMzYLCd7PZL1/MMjojR6GtMIBIt649EdyUE3KDuUEYm
O530CpUopaMx5jAHjLMLzTA8P72Jo4cP9c+L/05a2C714SNm3MAH7tEgk+R6TLUGXN4i93uxbz/v
sNTPJOmFuxGak35LKZKwjPnMEjKu+sqt30t7ZLrHzvRV8iTtZAvh8Y7I1dEUE60g4f4GDuMhDGXD
AODcgh1ZLQMOfQcyyfNXKRILz1qtrcC5lULuvQvGFEKrtbyn7luTuDWQHeYDVqik9j+TMhN8BmI8
obcwgWHIpdQX7ZvOa7nA/aAVymNyuaw4AKAAgG4q63YINQ6lhYCUeDfdofWjyhx7iyDqDPbOiCMh
XZ3lxt7xizrP+R+UAKX8RtGd2uGYgGwctI6pammXWEme5tgE0FRbP1poSkT6ZAoUSPlPnEGpwXvE
pAmclVh3cExjG7hrCh1xHlIRUhqWjdYKeT2pZKsBfPBVs/qMsaVicX9+fk1Z1u/bHjbup585emN+
/hHap254yLt0EDfID/f6uCoNV86o3dvCVGrkzYX3OIctX7OqBDHx+EuNMua91gPg/Xs6qzi4ZboG
Pa2Ajdv1Y//3QTVeetY/x+D/XJJtftghoSdbz8F+IENBFSf3qBRmG9I6xG6/Svj+HdJlXiB9phNI
vHQES11jbiAfhrjkjozdmSLmhV5prnGmSgGfvvBim/6DxXMQwlXuZOGcuNKPgIDU3+8spToCdOCW
C+tjRDmAKdHN2r9jyQAVMoy5dYhw/auglG71i9xbj1e0xdREIYdp2JX2TMYogp5wZxxhiFY3GoMM
gAIuag6fQJl6NaYMuLkGv+QgHEww8n3/+LU+n0LIuZDV7T6a6cFFBBPoVQwdaWvXcsKGU8UmEs51
adJY/JAS5QED7eCxdDheYGYfwpaldizErJeroJOwtxu3qKsc2EE8E0O0ordAltRLmYox3LKT7WAx
OKP3YqKufzsbsFArFSS9E49IUonfL/XKiiJZgoGlwXdIGh12oKkY11ygEevDl873uPDXUlb91Y3e
28+odSqhj7Eoalg90Hjl2JQqFapO130BuOaLX4eRK7Tkpe+puuP1chV1I6JBL9RaEdurra2mgGqr
xXi3Kz6+I5DPMtQ/Gnc8Mi3I2Ib3JSo6UmfHYxP94zF8p0yFES5tDepzPXW4lHkSL+cNx4AU8Trs
gQ7USkCTFEZOAXic2/orqFTatUtwgulB9HjuWH3Z5ntDDh4UaNQ5AHvrw20fDUU3whVZ1sgE1wVy
/T2cIkb7IRi6/LIB/Pg9jEusgbdz5IQhdtwt1vN9GBXiD2GmrpDRlu7W4H8bVFxX68ujU53+C0Hz
8e2s9G9hj2Vc1iP7MjIY9WyAZ3TWH6h5lAVL3YAEBKZAG6jtGoaBHRA1Ew08+dGFmGqctPkU4I5G
/ycab+vI4N9SzQLVuzbrOsjoajH+8aZanOa5NzQXK1N48BbZDDHWnu2HWG7/J1pmEXkWLXAq4XAe
9isLzM3sYEliLyEaWfXKf9A0v56y8lQP9a+o7vahAWudZ8UBnSAfGeuMcVFGnuAraQTZNveHIV/n
e4zpZotv3agHQ/lavBFE8D+knSSONzNPdfK8E7fKlgMC3szuTD74WKgLS9dngnTrwmg01Ew/ZETv
cHiuCu0spAU7YH+ip+1IeERotcJC8b3wSTl8nAGA5gIrcYYEL7hPF55H1K5JGc8sV2fTjvIkCwml
N2qMWQ6O20eUSlyEsm3q8uJYnLAq8IV2+B93yinUTHFftNSPl8zV5FE3BbU/kKS6P7pW2yKpzvFi
Iirq6P43aneYvBQA87g7qg/zQFt3QxgTJOxDFThto80xSsLZVhoSAisFnkUuaqUmaXpvPt3fBWSq
E1Sfdag4yzPAa1N5MviULV0ojTPaJgZTKaLdGi0r3K7qoB2zQHiW6DQtv/oWYbFNsmEH9r5kBw5q
Y/a7fBDgAUZ10w9YCGr4Mj5dRoe3MEAgHwsn21Y1r8GF+sqrTqMCkAXj1xN5D8qXjpQHrclp9Wgr
nujmjrZggs4LZ0TteWrXv6W4bftSS+1Ymmcs0EX46bE0/mqHUMKeXM4k636Cg3aLFs9+fd/IXPCJ
Cy+u5QraalRiTNRXSB136tODeQT+ZrI6Z133UrqG0vlDpIjqmklysKWqyuy4jpbWkT6gIMmKSMSq
/i21+Ws1vpeOX7yuCND05sM4i5RP/G25rPpo8V/UpV4gzkotG4eOYZVc0MRy7gsPcLUVBcvDAQkR
BSOJcA+cxOeBN4QrnVOBfYEW1TNJ6S0EzQEex2lO289g+8wZDgUZe+6+klfYNAu4EXDqrOxJp6kW
41kdxrn3fzKsnqaMeFr1pS0MC+GEMyIXc2Kop1u67wnC61XBLu8HvPgy3nmBFTEXhqyvh1rikhdc
czBwcUHcxQGo3r0I0cVIh8ewLain7/9pxrmT0hY0pfx/GHgUzsi4PKS5q4/t1htDpWeufwxZO6Ln
epRJIYjMC283iQ8pxdTl5wLIoWiFUIGxxYZqJY9Gqe8BARY6J83HQuf51QQthcpNEhZaaF1dfLNz
vk8TZtJ/HHJe0+JWRZfGRPs5SlkK7jso+rGQkWmggfVadweTbFcirrCi32s6Zs/BDoNE5XvCUgYX
qzK2G7Jy2DKYoTFhWTLmpUl9aDjsyf3Vku64k7NdbDOnBlDH1VTsjKDnRLsrfGY++sgd2F/xq+YR
zu/HDCjMzNkOMm8lxIBwJ8aioj/kAanyy4QXcnLg5JsDHKA05KyUTuihSknWF7MlvlP7N7lSD2BT
2y9qCqfX+NNFn64Zpt1U+eQFmK5AS+1GpuOcS8y1+UE19nNJn1QL/KYMA6JY3FmKREns9ADDSK82
ZchlNsROXIjIWoPdgMaI2pNkd4Hb/fCQvs2gF0+PIYoAsGRzfRXKPLeoqdArHFpCQn+Npholc7rA
/cZNNctlz0deOtXtk3EYaohw/SvXjYoadYG30oQye+NVYezr+NLKhkzzFMC5E3Gc0KjRUN4JR2Zv
Qg/OEwuLg88Csrv9EzylravCAZeSuUOio9m8Zno0BxS/SteSQz8cWbB9O40Q35siDplHQZWbAvLc
f6HMdfXoUpu6UyHhtuzDeHBwReT5YRADpUWwvqN68jFNSKbaTeywFQrfhgt76GBVR1O8AneHZDVH
Dq390001Ng/UQTmFPvART7IpDw6OT0c0yOnEYm4UMVXRoB5M3+U7gujloC25S9yHOAMqeze1OZDm
2LQMRMMIGO7QA+1mJ4uOty9D3UDegIoiTk99dhmHLCiCFwovSiFAEFzACxlJrpjkAXJztcNKdPoG
Ly5Qy094f79ihTGe1tl63KzRY1w3cj9IPX7ufgyw5NzUURYOZJ0CxlGuNCPCxJYVazs9dX9lwu0Q
9wSmw3MzhySK9NKk/o9I5Tdutaapr6HP1VRIcGlu+R3rt72idxalxFJjL8e5toWFvqfb3pdIF9rr
OmIogEIByp2y6d9SLxQYNl0evTQKDjrYNqJSBjgbObVThPtu7V2feey4vN9V3F7pQ/I8/fAefkyN
9xEuXCxQYMs1iJ7+dkIAhTKw2AJwvRlv6ObL4WHegP0p/hmn2gk0DnQhIPfto8Xwx53vh4JLcyad
BLWJyqGb6GfVLsO9rPtTW45WcWwlDZYCi2V5DjKMVBRMKX6zeUR+CKd4dr6+1M1n0QaO+EgITjSM
tm4YNyN62WioQeVg0q66KldTtrcW0awSlqYc+Xunup4CNyCAH7JV9ZjtGDftyXCj481Rmf2rWXrt
kOnLcEJP6S0wuKLu45uY9QaVA1rhlpi58y85BtmolMWGbJXtgZMhSik1v0DKRqhDrGoiD0XY5LJB
NdLHug41dTZFheJkKIu9FNe/wDnwpU4OyvxIDpzu1tzSiRE9WXeQWqZPaK1vYOyatQ49c81grGhr
SZGrRyjb4UUiYIhgPR4x/4l0fGN4bo/chcA0Mwf2FsUAmWNLpdV+q/rkqv0IKsHxigSpQY9LQZuD
vwXmOSG1qy9pd3/IvbFfJxg38Zvvk2S3y7aL+o236nGnX0h3zT7s2GSY/B9pze74Al7dAiGXCbJ2
xJdhKttkK79O3c39wNyCpj6F0hEVQWzPR3/b5VTum6lSujgNzuitrMxYUYJ7FrNYRsTkSRE2dj4n
4mnWF970lzmAt5qKFIJ2BW4oONtUkiazuXYs4BGdeTMNrklhrTVUlTaLizaxMznvuR1tFJ7Zahee
J7RHBpo1ocFHh6HfagC8YS3niKBFDgbG8Kit+2kMRSFUYehuaITYLnbDhlu7mqx61lCxUfxiMvps
iQbuWXn02yyzr/n4n7jVE/jmAd49LonM+ZOnlte25AKbA6Dg65+0yfDFSg20XUELuTTS5N2lS4o9
74Gg/xaeFXK5g5AJLbGTMJHxII6O2A192/yIi0/0eAajvkHP2BQ1HmohxT8U9QtZjCqhOZnLY/Lk
lXLSs1lewBcBsOa7nr32vPnq1J4Ttq+XUciHm4qOl91PBpmS68QwLNQrMhSu13cEErK/nQ8iN91m
2rkTzsJqidbKR5qoeLWdbtjBTx9npT2y6+IkyOZ9tX4YK7+UMkaUwQTdcK13ZVaI177bOUt7SXyI
5nl7RnsxJfmDzDkWSk/uwL0qXDZKjeX4q6h+QDPVuuqV1x0tq/RtFtvBdvIdkTj0KgU+PL1Kxs8b
nnTMRqMc+kWwrwxDw9Iicxvu2VzOYi6RQnoyfokFOid2v/xn0rE5TPenGZeS80FKNnfNyCkLm4Gu
R29xPysT9n+BiooQ19kD6xi9urogXXn6z025uoyciTu4POKnMw68mSYDS6F2o4+s6gJknJsls4Ia
l/PcQlRsCugaazqHAiQNEf65Q6aX9KW0rW1T+KhF5qGce8Qx1mmsXzoSAi3OWJYbnyaFHpoEVRDp
zmsvfBP1TuR47XIiiKUGyuvly5x44zCKpdUSo8OF3cCa37CsC0bHE1amon7CJYoJmU+pJ6PiPSj+
L9xVH8aneuwMAKdmvNcxYCdNXXLxmD8XakKeoIRfe4VHb4YBV7/IgqgIEcDXYJLUuAV/DPxEH5Kr
ZzCTtLqbXpSUYmnXAvKqt5L6hpNR57z07xchW5VJx3X115dO8k3AWqelNqpN88J/M+H/sF8uEvD3
84w2Hf+NF1pPLA8nr8P7Nos4gVCDUL9zS5E9FKsu4+ZvyTgeDbDxpoO1GpuDsZPYoqgML9O+N6pR
y+yfcHYX2y87hDox8jp3RTadgd/hFqF3Wz0ZQ9sd+6EdbPWYcs0MB/05Qd7iEUhUM6KfYWOfTv4+
mV+O8eBlW7ndnSkEvvZTpAFAbCMD0kmkYMESpON/+I+7KBCVPDYxYsBWzhMJY1xHFYnob+TZQ57q
3xz0jPwj8UeSVOR3T4HEv9oF9aUFqO6eVX3lW3yHRKYinNT9zEKLWHtRca+Z5EIx89NbMkAGpVSH
eWnDt262qxn6uHUdklYb4o2w0BSmBPNlsA7jFm1MigZO3Gtx2rKaLH2wkBoKC8Ue9Ysi7RuYcwSx
Ohi07jC2N1NtySSFWYQClo+UjFkNRZpQL3O0gfb2vdAfXvgEqYGA8w8zYpyNB9jGbW0lrw8M/Pog
vudRUCHFmSW+swXND83mf9SyJjWFUR1XtUb0l7VhgH+fStAAmwGiNw3JSOYHfl+TQxyGUfi6WJEu
T3Jf1bxt2LqaFo8yIpY4z+NqvlNlSoAvowlWkdxV71F2SjeduDtAIDXuXF1iymj9BJ5kg2PhIxZb
0Z86UUhO16mXecvl03Oq4dRwOzKX59Vn/SxPrHatObqHUf4ntBUjVSw8gmJMx7E63Q0uGNlYfg+l
ksmDeOP3AVsjDLFToA2aogypbzcyDZsfjxpMxQNZ4hHo5DNMmbKOY+E5idzMxmW+5UzSf2lQvwbR
Uelbazc9WrjR3H3/RlZkXH6nn1Bd3eAFGOs24PdJI/RIEDbyvBD3xzWc8F0Yc9ttKXDWXFNnp+a1
rxl6vP1517Zfa2kXxEBTNTV2OfaoQpB8lXYGtfrhoAGnRqd6mSXnw9prWNwJDu2d+HFo6b2zGoV/
kW8pSFbgVhgjooHlU8AueQKzLaUwALpaQV3CQtNPRTuG9uwcvgPxqFRo8eP0zFS8oe1Rzo7ODq/Y
iqmE/0q3Ksh4XPzHmQqDiAdp2t4EXbpjhic7gODyX/HepwrSAw59jXOOc8xBLICERLsr9BxPd/vl
8374IJtwUihI5ZgHIoz+spBAESF9/Nh3obGWqRMpM0d9F/4fD7LZtMoeOmAJgThy/i0CQjOHF7pp
MccwMqHsPlMscIf4CPw/eXUdcCNyaxlYYSWUO15eZjVxW2LCcehDVutsuOmmpHWH9kWgxlCSJ1ra
bTGYqRjLcTzOB4Jf1cvvyMoIMpcwMHFNYcrbMXIeZvSnPO15KeC9HgVZFxoSSZiF2B2o2hSJY3GV
Gx1x3HTsLrYqD7aeXqwpsHrDXyuITz3cWHLTuzPA7wV1fHyET8KzkPvGJWKkQtaJ0/n9MxQnWOX4
8Vpgt4Gxl/mKJQBQyLKr5aQiBugYxMoPUy4T2mBR1ePzvQJ6XOANOHAGsZNmIhEuYDwckFU+64hI
CG4bMHf13LvCpRiDIDt9bg7AQI2pgCX2ays8W0/+yI5OJtAcDLtSIaNdciiulpwoEy4r0Cy0mmxF
HXbI1kLFetRTtZwRy6jkEj13tOg6u+a9ihlk67AtXRwqK60/YDonT/0KwJW53Vwl/fQFX1pWTCll
plSKcm2P14I0ulxc0mohMWTkfk3WOJF9QThUUuF5j3Del6n3a3pCCvpL2+20nhSyt+TLyBdwMG4J
11y4oc+ZZ66kzv7nSIj/Zq1NpyMKeqGdr4hDy33eL9f8qkWzmExQp6dlwsa1duUSHVH61u39/U8+
uUI710EBFKExTghXzhAJBRJ1B/DGKw3jggoBsGuqPck8v6PEA5IS85QBT/COqKC9uql/v3OYHWyz
0l3JffvzCt6oaq0FhRIfmlC4s+2CkvA/qmajCxS2yc7/rVLrP8JUEJyq9F4rNNO6rMsMcjGAg+oR
65U2gdjYrexGV044bjtF9UPqviG35/MFnzMpNVFaZ1mJx3vytVa89oIScHBanzIGupmMqxSShdzy
d6jbbuaz+8xe+VUYql6k8fcQOVI8dJrFK+qZdUWj1p/jPoJ0ozbzsIuTks2376qkm9SODNyHW+1r
KK9uUdr2Un/e83rJCxBaUvUylNQmAtpqPFkVY/kTndnG6fTF7kAZGN7nStQug/Aw8PKusUugE8Q1
vpHoyc9YUz3QvIXUG2jbw6Df3tF5pD435IDwKp0nnLbthmo21bk38tSPb7jyuy8dy4rCOGxTM1X5
XTzzhGy8SKV7P+aZpXwHutF73sn7mPl+jmjsl9CPWoMgU7WMNm3Gdhwjnk5x+V71h1RRKgPV4tkO
+zEXvzCdWY4Xeb6b2STfCFpuVheO5Z+4RnWZOy2qSeQEsJX3itTUzR0/kSif+IH/x0PzmQ/d04tP
viunrnpCX7pT1d/SQoHptY7MzJkeCMW4qyYbQrwkNgO7ZFVTxbx0jEvgZDWwiqJnpjPEya/TtxQ5
zW9u48QWb0Mlw270hv1WNaJPxjO3ccYsNUKsSqdVBYvUmsGBv+uPe5tjCylGFGs53LXb4hXuLr7v
D/dxUvsKTZF8P+5awEOD88uCO4a9tGtmRW3fVXUjuWIIdjrnaTyTPWuNlepTX/Nj2jj4klIRDK1h
ILS65mULwfbVZLDpyiBZwOg1bDVNG7d+a3PDr8MTAGOqB6j3VpCY5kM7yB3jxj5bffoIjd7VmXfG
4fGKqKAlLpD6+8dR94+jGyY0VgdgJ5wlxHLDIt6ye75SsxWg5Rfq9gGo0WHnHfNiATdURvCnu5J1
rd0rJoc7bMDUCze14cn8B8lYITPY98oMZUXdayINzpPiy5NQ6FKBITNraMA/KUotI2jjweC+0FF+
ifvtWw2Bhmt1gdMJXfupi59BsWFn0xgloUC2zUg35hCywLyRyR5c7ti6gMVRr5yX+/wwhcZu9Ymk
baNQ72K6ZhrsCvjXczmUXwsNdvqnZEpP7T+FF0Zb/Z+qcS2XLLJxlj556bo3TRDrkIC9979VoP/d
zfzdvnZXT7MpWTbfviJsD7kooQBPvoJWYHCjsbvAIJPO/nxQtKHKHlb2xtIO65+I9nEuenSpJH10
LvoNSPrT/5HS1LhLsFphiuIoV6/IfDCGZRj2PFnjUWN998HqfdOYf64faCHfGpJN9hdmlwDWwcYd
ub9DhncikcgGDFvJ6EGnOJ69PbBIIliJ3KAVi/5+7NDcLXsjDM24EpNo0G5FQ4X1TAxTHEWrpjRL
vndC1OmPMKXEvJT3U00m9+cJ6EiGUiZB/ijqcED+O7UjOqGcinUE6GqHDM8C79SPH9towqXPFiJL
2iBizaOwXC0Xjhuj3x3m6LmxxUz4B3DawSja7+Nhm3aSCFS8t+uHdKq9E7k5lrugolZkVkVsfMSL
M44vAkKWmE5d3QgqNOqR+AIxSB5NUR80+aFobYLzH8f1sgYturl1Ac8DWGNRUrcL8ZvVx39DMT0u
46L7gcVTY82LoO+KFo1496DILFtIGMEeYG6q2mAzCmFTwmvrXeLz0a//mpycbslMneiCCnaszSC3
2KR7qnSMU8tO3BCbVFvG9R+ZtyQ004+6Qbw33SODdwzU8hbGQMWDnpD5nPDfAQMY+aTb93X3kqTK
VBsSA93gTAz5WLUA5cZ7OfUEE7WhrY7yQh464v6UdgHEJwhg19TOng25LhGnRi9vsZGcvOma3dec
eGft8hwlJrDPgyFC4vokv7nG8xea71yPquPEUXUpmlJtCJnneOsnpUhOt+rkxJU4BGX5xrD6ElgL
PSIcX92bGrRBEl8n+6836GYBxViWTXU9+Z+78DW7z7+H1hYcKRK3ZB1uLJ2wmPospPXjgKkQAYmS
isfJp3ql8uvi32y/TGJfMkHqg/04v6I6H1KOfV315utPolJuwniR/gRpLDxCul97zwjeeWNXQa08
yRV7NtaRrB/08KbF4viCPZXmmSmcBak5obz1fNf6B2AeiG1Rf6GpEJQdcQOFI1EZ+6ryivT3ef6x
nAPwTNkCZk8bQoUxrcfa9a9cF98BeArBIvg+Yj6sSF2XdfHxX+f9i3Cg+iJU/nHiu1WlR8UeP95+
cyTr01Vo1Uir8XUIHrNuLFWFchv8agILg+fK55jroytW49tUrJKZ79mP9MC+LU1XUkEKF1sOjMla
pi5IVvXE8WxfvFLbVkAtIs5c/zbSx3+odfj7OYEEbS+I4uxVTowsqtELWnwq4LWCCkjyQ/ODApyH
tT9oGvP0CnQdSaDOtw0xBzPNG9r+YL7MuAOkLMNIFRRRyynJYkmQRzzMbjIljLqrDq2liPOy9k/H
LNhcC5mwfdXNyihGFrPUVpNJC099u7IR5UBeCurMhJ0BV7QIVyjKgcnSHz/KVTWvj0hWt3iT91WT
USgqZ2wVXOjWsYr08bhWZbIaHE9BxydQoWmlimi58x0sc62jhgc9JPkjL0/DIhxfjxYJJAVNqUlh
WwgSxWSKGWWr5OuZgn/PZ+yUQagmyfa8dZsOVI6Esp5J6Y2LGJRFWUcVAg0GwT9gdfOSjr5g+VHp
Z0i5hvl8HraEm/yP5LI8u5rEZzeyjU1lcJtZiLOszVRNjsn/NXjFQigyuiGTrpPe06jkPiRx6tFD
EdMtidEfc6KYaAik2/F+yOY+d/ow5UEH8yTQ0J0kWpOKhQRfPgPNvaTsNZbK0CgW1U3QqNNoMLBM
M3b7FgPgYPgDkaniqqYiROODUseL1bZVDyform5CZ9f41ax1LYuHU7DjtZ11ttCL08F4nHj2q1zb
/2muZLRkCcXei9xeDwkRX8rBx/yHwnX+MKyuwyklNj8KGnEs7qMe0Cr71HgcNE+0w2m/8jR0IMTE
Fg/x1nSp2cq2YD/FJTZhqj0H68TZBYxX4gkVtsU6Dt3WcYySmmXS3Hv1vg/4kjxqTh12IRzC6aDq
VUpE9esM+nUYq4pB+GaW4ob+fj/PhJpbuQ94SZAf4tqO1CPrb8gezMRb7SDHMfBfzu9R+A49PurD
Z55KKeOmG6BOVfWEDkMHHi0qyYbGj+go3Thy7VYcscH9nukc0dPwEJrZ7VbAjM7OT9bf1Kl7oUSa
XNp2FinNPjHo6wnUaBBD0w/S+bjdEGviRS7dAZ6v0hgxqGgbjHjFoG16/O5cAkKuOAkGsuHLiGOl
eRtYnPz6e5deN7WNPPzFVRI+WU9+OOW6YdHjezMemUj2VJH0M3/RZufRjZyd9numahPuC28fo3q5
/C6ToiEZBpTN9jdB4hzwOMnELdiewQAZlI8gGtYoR6dkzet5MlAZw5AYNqEgLeip9JyY5AxHt0ro
JwkUV8Vvoyeay+cLZWEHade5DlvEiv6gLiEzW8uZdQ4N9Z71dX2Sicsvjps7xrvUl9czRzVcRVjL
z+HluCHUr2qssb15hHD3ZdY0IoG8TQibu1k8hBgWDNRO9NLXhhrOMh/6E0rRrcYZX8zAErvvCrDm
0XgjI85UiT5uP4i3p0QiRuHnuq9kWEw+eloA7k2rc4w4bDc9zA+7lhZhsDSz01ZdHOd//ReG8sK7
jsJuif03NvDV/foPvTAef+am3xEppUnM+WsW6PIwoViXi9sRg5kAdLFuT3vPEjRBzcAmaP4CRPvG
/bUTYVg2DksUh4+LAKvNvRR1qfVDnwJFvSdRIR+otH+oql0m/xpyT9VzpAJq2ECSUe0/w/OgYTS1
f5F5RTQH06AHTLajrj0aUb211HC9ubPff1dS+lSXXve60HrgW50hrS5XJLJHtBCxJpEfZM06/Lqt
CBBpYxCC4kwl/ncPZe+/4l1NZQkVPVGfzn3NRWH5pMElZCEAFTrxKRjGejiqDwkNvhHUTwkjWTan
B4sdPkReVPgQgjzxdk8IVwd/9bOj9JFIAa1kMB0/bfmNbHNcgeMQ07nkvfSs2vXkQleUGKb097R0
rSgxlAqiGJ9V7NTjHFfMv8j0azLtHlLmNOm1znMkpoL6wzkmNRyYhJWHkvmyFjdG0zw+f50ZapxS
Ml7RcXJgQlS/rMhFvqki9obPT+j3YB+/4DodPuvt5A9IcuSzXk8VJzLTL+olvXCG5xZrOxGaLlp0
N0+OIIloFKQWZQsboWWYoxH9dfp01a5Ov+fq13vsBpdnttY++NDP0Jio6LUQZ+sUpko5juruyOHQ
ZvVRXueAgQJUNLJQwYD1lrprYtWCx95l/O2g5XC1cx5leYDwHnE5oxNHLDdoyGjHI/Za5mk2Wa2Z
9M0CkkU1YaDrsjEuWc9Z4b6JQmDVwXSE5NcbiGbOMlnkoDgaUMDBHTfnDXVucj7QC0hzaLKzJvCy
kWwUkqFyx07cz0cvsyJAcQUAqxIwRryEL5Qtb4C/FqbxS9qOItdVPKod9p2y3YP7DKlpnajcTV0m
+lFDwbWnQ8buILzXEjFpm09WIeU35nt2M9QGghRNZkbp41rvj3f/0wAQI1uNfRShB96ZWxZ8m70p
nqV1KSK76hWoEaq9hvr73y2GYtZLcB9WE9W4AtLNaH1N89RjhHqtfXZ9K+2idV6e5yw1JOcuBZ3R
zPjYDbi2r3BjYxPIWGwN5WCK+kkIYTgmeczGNWPFmPVSmUWTfxoNVRVrM74L0ALnt/PJ7TGiMVIE
arIObEtDLnHfEYuT+vKewra7i+USCSBvP/gKB2DpPWvKvLf+opPF6r0AyZBSP1395Yi2fGlG/soF
NsdqxYmmo1f+dPxC2dCY7Pjo6FSMSjBDerV3r4eaa0SK/VqP7sLXF56oXA2eF8uER2TinG1iRQJo
5z6r+/qUUbp4CoqMddwMJ3dbGk0ztyjMjfpDi15oxJlLHgR3RairYJzVnPox0Ne8hF5q6QgRw06s
A8FlqsapxBzLuIhfRXlO/E/UvBRijn1goxoZ75HVuizQRKiAW/Ku4UM0ZfknipUlQfavlClSr+C7
2MRvrhwMrXyCf1qVewd2f7Ai49NVdixXmyAn84uWjT00rn7Kfl4+trroV032PQZySU1tdOeIui+R
2jx+T7BJ/G3ZT26yeeQBZ3wV5sqrvYl0pwvLBAv1Ljxj9H0iXcF6eb+7kht3f+0o5swVlZvvAz8W
7BJmOF43eSG1irLGAQbczx9TVzFQo3UjX/TXStSzA0R1zbTZt3LmRjzwRuIhObLO13ld5RjeIYLU
5vhf6iTAKM1gZx5wjEtB8QyTdRY8sB5sznerCT5qt7eFJkw1rdY3WRJHOGlmRF4e9KRzBFYEMJ9n
gKnKd8aMkC0WX292CTw4WNk9bhg0AvKIuYOEzOAQaC5cej/f/nG3/Z0VWU1S2OVC1PR3T6KZVyfg
1S3plbEjOTztuOalm1ppU9qq9iMLUGPF3H2xsc++RUMTMX+FPtzhxa+u4JaS3qv8dYwyzcykbJa1
cH+tfrMEjQjZAHI+WLmVFUNyxuJ19Bi9QV4ydxHFW+bRzuqfP3zqByp9//M5ptfSf3XtUZn9dDxS
KDi21xxIBJJ0OBgajtGlvKsdZqWaGaQpuMpAJxxPLL/sbh64mE1dKHgnK4nDSXBKez6L5+UjIE27
KQpdhBoTHWcZx77jDAar3DOxp+a7l0ljbsSKxrGSSjXQPlHuVjzFABMjq9WAacmBESf8RUjR1Hgv
6/5i7LnXrjdruSu8Zb4dSpXWZ7H//nEyvjlxBrw9nRdY5QAUb7rftDd0U+AwIQB2rhmhfOaDaJrp
PSczYQDH4QJYC3f+DnUVs3xdG27G9FqnhHDGvHcoflStZ/DhCyIEqDy4GOmEFvjrweiDAjoA3VAK
UMHKcxMfbHMHzAGlhXmeDOPwVcLfGq8F4gnLEFCLbfHlCOXOMwmpDb807x/e24PVSVzUeO2vASz/
dtF8ntNgc/93czwkkxRWy3wypQhz4oV5a9UeQA/SfbLCeuQxwgRSOAH/VVR05p5BK/G6jAGPWC/7
d+XOgsbJxJBFNiug03xWAJCAetLHHZgdogwXZNR1dnviCo9hicMaxD6F2smn/+QcnZkwJDNVGUbe
9PvTzmhMYkfD7YCJU6DepVy1szBU5ragW9elY+UgzJBW7l/3qM2Ycvv53CedYUbnghONIdUdNAKj
eMUrRuqa1P9wsBWdD43fLlvW82lWUzWwKnSIh2yhDbdU80OAwnXtlPCt2ZafFpi6AtgKd5ek1WYr
vSgAkkure36jkyt/4wHBNhzB8Vca7SkL6QKVlEz8Df1v2YP/RvV072qCW8/t+fQmO88wjBCWBLBU
DEY6gPBp7+6ydnXjL1Vy/FSNWiCBrGHrc2WdzKnzx1bOH2TcaE9IbGXAJfGfV67MiNt8X82x0s+q
leRgTGaom9Auo8kow3MBTAJLfCM0Q38AmW+Npz+zwDtVwC+2JmHaAm90Mb+eLMiflHpIok3JBCpy
/+uNu06uS4e4CwPoy4uSVYZf+qfmNsmbSmVDr97NUsyr0k+wh/3ZwsdF+0NvVZxfdVmjY4D3hg35
X/gXhyP7rywhoqUKsp31aQIlqVkYrb5rkkiOPNDmO4GgPQt7t8f9W4UUh8MAPmhX3GccJ4wFLsif
A8QqUMbqjaKT+EMP9y3ZIGxejtJ/Zv60xX9RW9HAoG1nhKkBntJxcpB6S9oJWI6dCXTDTeUf+BjM
EO6mm2HEqzbiIwccWNznbCpHI50xIkS87S0W35lpwJn8BDyuOT8Ka4HwIkMLT03vwZJC6/z6mpqK
b/5vUagpgsJvGL2A8AZ/HvGHlwC/ck0/q1fvkJA1+miHE80NukVgnDSXFVlRSaH0H3hgvh42zptc
9e7bjf9fROZzUHUZu1wdCmqGG2ynCGrT/xDyTxCZEY+gJN88Ouc8lj7d2NQ7eEVeALe1r7Snhp+e
01CUTrUQrp+TCJpli9RcurByMwu50xUR/mbrp0PpEljU1b1/XT+ov4uPR7Oz5qKJ1B/Woapxnw/X
ASlp/Xel2WC2PZ6zvaVnFF5wcOYSEnYCuhi8v1sihtEkGyXGyr1q1W4yw2ff8I5nV5FzucDDvWjg
QS1TqkbFwPlvS5KBba/1FKmUbtz9kEfzG1Uay9IzHKslAmsoHp8IL8ld2BDK62G/MzMfYoLiiqmu
iRn7q9LiWtI1gytJkRIcAvt1KkPm9/4X3oq7JfXZ0YYWtUsQicpJFr8o2NLH/3NHrG1Rto5gDm5Y
GYiqT7fthKC17PxUtQQQKRpubpV8jggiCPcsY1YNV22RyS+DI1JU7I4+Qy+6pUKyPcJQKo/YnCCU
8VnIOqTVTUkpN/JtSJmvqQLqsbItW3Nj6ollbhBNARHwLkrr5k9tO/2xa4YakRepaXuYJfcgex4H
bOFDQyQdkbZkCxx5LLV9AeS7FHSw+BT879g0EinblcZJkXM6a2OqWO/b/RE8Asubr4LZm6h9IZ9n
vpSlKIK0f+gaGPkR7gSahKw85Ipx5Z6QYnOhHmJvLK6gk7uM3pOQIzbSQBCQC4G/NYJRUTJe8VSR
fam7D7HwiIWpAIdZYpyExB7FkfSiJCe+B8+aQXsxtQwLfB/vb69Ab5zTaBTSxlsdzW/pk/+8FZDS
fbPLyvGs/EZsD9IKUkzRohJa9eu15Yb8sSWubUelGOkG0JqfH5RTFWoWxKWEWkWSIdJHmf5XNaAQ
thmz7XHUg1nJ/HSpCyMrWLn+4RP0otd9U5YDeQnDfni6eS8tV6r9d/FYWHfZNULJY17Ilwzdw9LI
1CaPTnSTptOvLyMTNdRYSOchLsDZivKAzlwAZOGfKgDCUBvayfEEM/590A9LGWL3YEpxllwpk5O3
w9uZiUw/cJfKbnQzhdcMFM1izQcBGQnoW1sCf4fgFQ9K2gsHduss7AduafKPwTkp/C5RuLDu+u1V
Hd7TnQedEsjPRog23yfS2PenjkuhwoxwqidOVjRyM2XXcjZ8jDRKXbfNFkiDR7jebF/rsEis5xf5
OM59M/pjlHVwZ0eIg/kxi+HrbPgjUxzKX21rnwaVbOc5ieUIAgH24VbYwRIfZkd6JSakOypFPlUF
bKTBgSQ6UU9FZuPeZDJ8zm52ZvmbMeORv3H3Xsx1C+yP1WgRuqxiZ9lRg6YtksIRDyJR9heuSiqF
5F2J3CoheENg6SbUiTrLPEFus1lgRrHta2aQARvGicS3W5RZ6F3NNi9uzFfMecvR38z9unipGQhG
Gh81TvdBMiNw48p1tpdWaUPARYrcmKoo9AkJHRl1XwsiJ+C6UsS0H9fuSeW8O4MozrJY9XDdEoMH
5/TNLnY3Onc6cXs7g/7ehQDux2d1QUvs+0OSyrkRQ0pTev7DDPrtB5Kv303Rj1HoQhbLJMLSj/oS
PNxxrRnYD6sV6a/1yPzUfXTkcLtpSSWFssPTM/sA/6VHgpqqSoNxkLzWzvhoYOFlTjohhzLrVBvx
RcOJ+oWo9PbEYjvM3UwO0VexSmaWNWHUUoMCdGzV1NYonkNpXYwWy83i6/mFtjDC+y/RSQmM6C8Z
XUJBvB2Dzlrg8cxCT5GZIPhTWLq4GJ6b+CBxXieAf7/LJE2TB14+52DSHYfecvo9D6rQx7ZL8SEr
Abzi+YImjfS5/v9SfmipphYPXafR+7AebIGlR8KWB00LosK5c1Qp5HYyXp9HTBaQDCt/I9VjsbPr
3XeI43q7s25Bsi8hAuhF0laZ03EwHndRJw42B5bHMjOsesFX26d1cTCyDVxcuUAb6C+ZK95qR9/0
MYpSjctenZj+3SHTh9JniEiEKMt7sYzouqt44Ir/Ok3dYevMT/qRJxxfU6xOoXTyewoRhyoYcKAm
oLnofe2G35z2b+aVB+98dAcmg0ZhuynFjmtasCL+RsbEbEMpKaOBmgJPqjvxr8GNiSBFcuBHvqRr
5T3d/x4FhzQ7HW2lpnQU9BrzY0Gi1RikSTRjW3aJ5qep6trGhLdRx/3raPxLCKF70nZxG0MsyF03
KWv6rvN7jPnTZPluND3qOAyoFNsYOF9BX8Clime6R7y9KsmQGY9j1sIQXelwNYYeuYbGLNOOz9kF
T2phzNJG6Mwz5773Aj6h5w48in8CofVndN3jehvdp2Q7+lBUr8VeTdyzFFEu5TzVymz+S6i1VMn/
EdWdd4FkQ3jvdcLKx15+Ck6+UXuGfiShz4NDBCcjSCeHInyF4P4PmxZ3Lvyh23aar7PdCC+gszO+
vooHivGTy3QFmN75hYMYMF42i0POFzWIPfJr/BNN0FPbsiAASiQuoxbdJEqR68sb4TRBEWSS4YTT
5gvGesk9puuMnvyTMo+oxKimIoI7sQS7Gj4CBQ8AOK7Zc0FiFsDbBsR627JWXE0G+UzAPN8PxIT2
QdBHqKhP5S0AkbFhkuMmF2aeDWu3CtSAR+C3KvCvxTEY8DaXE0h8efRduiY5Jaj6czcdHkC+7qkw
Fu2eitw1jUB3MUG6u4+EaN46F8MOyhuKq3VFP9QlId3JghNpHmtNsd/tL/Zst4sfAi+idLkUqQA6
YMsDy1f6hH2AOEt7vVCqmatespJi9+VfrSBGy4bfSTV5dwkTXXvVfMRDIOgQ9/WaK8o0FYWIEE+y
1RaMaoBMxA1r/dJL5grnk8kNs0zXAz2HNd+3hRMasHZH2ZiOcrAuKK995zGhKXJT3RQQbMR0Pk4f
cwpH7aSKozGfNBaTlQtfSWMPRiOBRbDnmeobMXX1Kz9QTOcsYiXPWy65Lla4S91ch5zcikHtCx7U
GIBks5+A2SLqhiBGtXmWWfN15pN7uOGOq+iMBLMxcS9JikWrbU99jtua4fk1RGdRHkFhDkKSgVDE
J3EDyFz5DsIhLcbKvIvgHawIj05vZ/j3bG/CLC5MaGwNWUgm8B/G1RG869acFSE0A0dpNuIpcujM
e8qvVIZCWQ6FjTCzepDuc4LG7UoBvDMrLVJNGYR5cP+4V/poteuP5VdXqht6Hq4dEK3n5jiz5pXj
gsz3Oy44m0uCjDBV1zTkhhxVyT/fHLgp94zR18hLWxdpIntUJf166M32YMkILiyY1Kzvac8j3MPL
MKzjuqSyZuHJ2RuFvfcjIq3u5IAJ0GuYGlrMTgZVXQcYO4m2BZCAw5ZwZ5vXFSxJi239U9BbmmYj
IlKOV9wDMEMNMhQzQbYzt0Y7OK45CG+A4C8oupAwrX6KOr/JafLTxJnURUU4LCXRAlq1Syk2chue
8IstcWM2jprrxQpIf3dkVLBfSeuFnCHNfaU8AaF0pI+OpR4BTYKfx34ktSOLYRNV25iB4qx7daGa
X5FOMC9rJ87CMABGGEjZKsBW8CB38fO2xTTwAZeS3RzgnzqmuKJxdKZ7MnJAklVMAnmOX/D9s4BG
UFu7/wP7+rob4StKzZLQmFRLNwRw/zlLaTqmVqctzxft3uGAwcsUqmx0jWqXBw7E5biEXojy5yOO
R1XCbway9FioRXSyYYDvCQtNe0xx8lRc9GOGn+hfC6rJlfSFzqtOJz23OWp+UN07kzh85rwHhxbn
n797CVH2QlfdGNqzVm7Q6wNdqUb+k96zxQV0CL1r9CxuviymPBGlF9DBy4iG52KXtOc+JCNG6CuY
Kv21Rv5KgqC1sNCFoj221UYMKzMVhzFZftcnXN0rGj0EZzGgVIaapH+zmDXIr4nTX6Cw1E8KuYSx
9n8mZygNs5eGoCc9CEupzANPnNo0E9tKgd03PIVW0a9yTr1OfrHwsMKOdE6O3LXVcuZs4/NYQIoS
PpoQzVrLHtcT1GNNwdLcScOi/Hp1XDZnGrF1IK5gZU7k6LxGQs0DdF5n31S9N3IR6LkkRRYfWUTO
XBDyykN65+VevMLm8TwaRieUYeMhdoJMKrXXwtAmaJkXG2iTfmCncCGI/L0Hv0LjmQKLT0YlxhO+
ecOO6brEpmEVKweDnO/gQHIGsGdj0X/LSjQrDcmXIxK0zojgVjUABHhGSNGeu8rkNG7CTusmIUr2
+GoYYSsa1uMJsWti3mq0OAWy1oZqvk93TRoexv6ddphYq+/6xwKqaIX/ggWE/tX/BxtxLyc9l8eb
4UbUHTfeaQa3GIY7wSIoGAA4H6sH2icYM3HxM8UjQrrdI0KvPFutUTFzxfcGL8RgXU1/GEhE5z39
1hD7kzqdiZKjtm5PyKDP/rgg2Pc8Z8q70oNxvJnnSape30udlDOC+WIZ6bCH24EWsAkMS/YrBBne
lUiFiY6W4JrkMPUsmxKEdPK5UKmk/4rSYPQ/fe3hzaOpMkSIW8k6Iky+sEj/4Sf4Q47GhVLNwJ0t
y6PEIGUNBy+ALcW+nmjfeG8rdpeWOjfj997dhcuS+QL8XgGYNny7nVEJcuSVL5qFeX9FYv1nJrlI
fYXaIl7Usb7Kv5/IAxb1t8Z8vU242Dgxwez2V9IeNo7TCbAEmeo204YwaJdRdiv5RXw3A0G3nZjE
OHanE7PWkKSiu1N+n4Dw5mrmmzi6RJm4EpPUlEYNhOIjSRaIG59cIv5Ue8Ylh6Npt5Y6kR2PFpKn
mESrdd2Ciwqkz6rvSo9W93RSiqMZ68Sq47O+qSJlXFNhmfzZmbNtMqNCmoRUy+ZIVVjPnMPsYjJf
pVkqa3HAIBkooyAltCRWiGrmq0QC4MX7eHmuqbYpDIRX7DPwzNB23n+yvKQcfYyVQ0zcM9vmyq3A
bMvN/xCIYLYOIExP8dw3nx+Uweh6PXQeRCTJlRons1iSoMGfH6qJivHgnuRbXR1KxVUPeAPJmcGk
dOdj9/K79DDQYk5mrnKmD+ZNaYbFl6fnssJYaFXcz42NbckEOkyHsO1TWM76sT8Ge8iXnQlbuSFR
8X6is264YbWcscmSwoJ3f0i+mmnmb6ock3zR7huKYD/f+tvdjgVGAhhBIbwxhzEDtXqZmA5+n5Jd
vhpTV+ioYAVHGwXZZDREVfDSDRlCYefepqF7YlJpTPCqMr7tCot8w/oihV3/6meYj9/nGCjL5ihf
JdjXNHKdQmKdp4jP1umX2rJ2If7XN3rIYJHrCLgqNzg5y4RNYx4Bm2VPYETq1rFQ8IEWnVrC5sKq
vCaKjfnHHBOAJ6MODVTNu2yjtcO1/L70Nd0DEcZVp2aBkwiqC2YR7JOD+GwHbh+m8oOtyyWvONMZ
s7eBnorQO0aUbhSVzgQiZ8Mlz5j/V8WQe989xTehnS9m/ssiHHDr4q3rJCGmVuJLGV0yq4QkMpTn
go9318fu62Gl4ezz8mskBkhS3gvdeEQHQJPZBB70xY04rrbqG0SCocCXeZOFQeLN1HRiHOmcO1dv
JE9nNLrIv68DPPPvfQBr85to4VLASP+IS74avjc5yi5ncu07nIo9GwQiE1TrnQjjRhCRFF7XvIkC
IzmR16YcXRSAKsWMo+N8w/cNRy6p7C2hMY2878foFAEHGJc7gGp2a4Sp8bkpzy/1SnE8T+QTTwky
ACJTcuVBp0B2a/TSUerICUtn5jjTeeC5lj6XHR3I6u5NxXUwdOv0xC3Tt+lZLm7JOiNZ+ybaCzik
moactVstWju7Tx4GoZW35YpVHZzpSWk5zweYGi8QDUmd0yu6S0zsK0hjbIFbHI2XUVgPfEkSU3Fx
gMd0XcPcpci4U/NtSpvCjMoMCYxb9NTzyVF9fvvccusydkZHNzox7LY7CxEWwL0OQqDbe5/frdtp
3EybkWZgvCICxdb0+9aUEl16me5jdiTAzmFHVD8sV+kSXw8KSnTr4yw0rwtRZSy8k014BEPH8zDz
U6JNMCKusPlEFmrNfwXaYN8tDLGpJlOWF1mi8f0q0K5K6ut/Ycn6hpa+Zm/aOEmqNw0BdtUb4BX6
Raq4Ga3u/jXTo4tyJL68iKs52gw+tvSuryowzyn2qfOC/goy7Q7+Onnx1M8b7eagLcXqlSjqi28Z
lbdBRa84kh5HpVdc51FzaTwbHXmpONRlyNVh5U8z96xyfqwmOmku6+1xHIjpmJDYipp6LN7ql1fn
kfbHJ3uQvMoFTZsWTbaxgAbuT1F2FEjf8J6mSUDQGDLD9SNy5/CIfi9EUcZfog/83kWWv6D5YpOd
MvxPmRU+bQlD/lwKucQzmxWr8Jiq7EU7eQjObNBq/BR0jAf6IUREk/PE9O84smHmyMagIgLNKj23
FHErumFG2fCYwWl3PpcgbpGxGWuorbxTGrcuaSVe55mJy6Qrj6t8ROh45YAaM3E4Vu3Zs25ueofw
mwRk9loo53sbA3tFSmUMcDf+sRYBlP9ifXvfH7a4X9glkudfIq8mysC/0XwsRLIviIGskThtbffB
gY9GpvQPg8PEq5J23M/26d03iJD3R6Y4Mu2BUKAoeQxgfqJUcROdIufnRgxBJgqOwCDO5uOskGNv
GN4Pn/Rm107kQ6QPzUi0u/OGyOqjY2MqQMKURDu9lxA9cQzLVbtSa54Vq84ojfMJpW+P6+yyJA9I
/mmCmyafPHqTM3I42CVZYBhBBmrjM3A1GbVUJ5N2QoZYawzTfJXjceUMx5ZZbmEaB2qsV2dbMtPv
i4oIeM66vy3qe9o3Y90pwGX4mtZu0wEC9ZMbYtaJ4KYhHlabFwPvUXwj/P5LVdiH3bVSXAod5epW
HR61t0P6Bn+9vVgyhxYTGMrqlDIaGNy5Al0XTACeGbQZATi280uJGt1IgTjtC+xkl9VXoZOG6EZF
0BN0QiVqdTd6V8WvmxfUI2tCY/Sf0g5aY4GcIro8CLiEFaBZoISRA6aarOR72SbFwoihtvtCkGke
qWNECY5JcTDhQgTO73lSeqdLWmPDxJot/GxIr79TY4FUqnBji/qi+xaq4o5PfkUNglkjGhE8IUUJ
N4gx5BJ47R5Wl+W+fq6wJysRA0GC0h3QzPDgyT/88PJitmGV6AcxPTc2AAfyYjA0i39tEX6YYjdP
n13UT+sRb2erJzSpB2bdi5QIkmf2zAWEe9FS0IBxtoKN5IbJIKO5/n1oY4gVSeftuzrwt6UalZFJ
N5ob22MLa2zr7naoErIFEjG3KPVabvtjpSEKoryilZK/myv4zj60p3ZQwa4/VDCFoQb9v/NTVKHJ
rYdmZYIcTvp0Sos10L3lo2V0GFlP2SX6IKulcZWK1pgvYyAoDYPJQR4U9wRbVU0zvyhrD4VQuGEj
GzLKoXo4wySfeBnYPyCsoDMyGEFtZnosZOtVEvW6GFvN6t+l9Eh8SwsEms5Nc8c4klJ/cs2hHNZV
tl60SQNYW/EXuKb0qigTQibkcFaHAyP0mgOGck3t5fGD17dX/yxGLdLHs9sXCSHHVWlNTbsZtSt3
ZQEr6CE3RXHWtWyw/IrgvH5jv8qVYiHqpjEZ4uYJkziV34rMMtBnuRR0hSBpQ+vFHn+Aw6+WK+th
ZH7+wnzFjmpoIi/JGnhqex9pWAbHRTxHdOkNonvhkuFNMaGCfEksaorKyUVVJ+yHiQJqMdHVj0f4
Aee/7D2YS5AXWgV5BErJ9EcUKUV3Bz0R/AOPIrKDrNnBxilVOA9TzjlzjjrwNh8Dw3MBmWv49iY7
vkHuzBfxDeQZGxlSj18QGiQBMjfJlWSEfqnVsnX/7M8QONTU2eIhhGilyGZNhtDp8GG8W/N7R4e0
Wp8oAQjjJD8CIY0ylMIFfd8L60mLTvSE/nYsGG5luSR4yQXPejzOyC3D3DyG7r+4JDhvXURNlGD8
yg/WX8i1Bx144aA9xWOhUnCWN1e3SC6mlwiLEF+QSV9p1aLi9Ax78/513e4G9Q1hRRQ5mHZHJDcY
eBao/WKZpCwkrWQ2bXPSrSJGKAvTC9spXz09F7q8R7caqoIA6M0SuKcZR9AiO26lojjjfuEbEi1R
yI3wTZJSKms/d7xwTEh2iF4A9PfhG7SzCjr/Dlxw+/8MIblqS1X6h90we5/r9oDueT3CYlWr2Gni
+RbcwrQSr4aTOd96vDPlshZoUHKenc5HyTnfCB4MOY013N7sTOVH3aBm5+1arxODOLXUENcMVWwm
Fq6hSSQgZLeVfOAUV2eyj+OsBM6F4rPQo9r8rzWj0a9HW/cjzSEnJ0820DntuLqskooveVhELWLF
Z+X38Wy/FiUNHCjIiX+rYBAPSA7IrgjFVQyYudczPnC2+hnPBOSoxPbAr0+D1UkxpL+A3UD63pL5
7L6AzuUqlyqoc7TZNt9cBGeKiEer/uBqpgkqsu1SgetdL0/2xI2O+8bP6qEQH2aZrA6IsQrtCZA+
Hr8NjwGg0i74c5fY0VXyJ0hJ8L1sOynW4Dq8mY1f8Ya62mFFzgvW+Dr6llwcOllkBmoxld3BTj22
ut+HzUEvrCKSWFE3NHTCMX3p4VCUPJpX/PJJL/g2LxpUsqBy+1FTJosLWBXeudLFcujQ3ULFmETF
erT40239vAi+lTb0x4Fg5LChC/DqRZHhCWqAEXvGZ8A0JNSa3NTUCYTosZ8bIR0Hel/pHPNaOXgg
+DP3ge+gwt4oGXEGQd0a2apws4XQWkxUerMzeterTREV3z8tx29PXWE5967kmtUWdGoTpsmlK0SH
VT5Xm0d1zaXfPEgRPNyX11HojyxGfR9Z/R1KP1DYKjwJ+rmXf24uYgREd1eF899d3YK7B7Y6CmS3
1yjqACQhY5T54PruXDRtf96dYHk7aGVYQahWcCEjRZMxYORNNUmMvAYwTliz32DqqASIhZJTvAMg
FXCFAvOB9RW3l2/V7wftefUueX4PaZiMGj1fpvGsqB/raVO4J1oM4iy4UjtIMdgKEw2T1Re2xj0l
2usS3JiGUVQzmAhmhRVVYFhJgOuJKFlBVR62oC/d48e4HpWvkpWkH+XLscvQoqBXDYJba54bcP/e
F7IbWS+tR7FcYV2RTiJM8YVWtPnW/NjZwBEPnaaDB+I9EenTLfHegGEbE3AQv6/9pdnXCa2WwLIE
x2FnQGS/7V5nMnTa7Mn6T88mSs/nA+CxC8Op4D7V619L/Ere02MozS/sm5rNc9WayCjjVmwu180k
8vtpnDQr4gCp38pZ8fca3ONgx/D54m12D8INvpVEcVSHab07aT5HbEAdTD8K/ka9yQXr/mphm0+I
nB5s3mQ7xD6gPPVwi5b+ox7c07kTEDgm8ZsVZFr67LDl7iUYRWaPsn5NpKHhOJmm2fUZQCkhbC/b
Pkjsi7nhapAW5Bcs0aoLLI4L+GPHucMFGCygnnPFBMSN5v/UGvY8RWyzmLPufb1DISe5WqCCV+Cx
wIbq2S6xAz2Qa0KCppZfntIi/qgMbMxr4d+jendMEdeaGo5Bj0bB/NXn+k7Fe5Jzya+Tflo0Q5Ez
cBglG8li91F7xhprSxWqcQjQ7bet/j2ugKG/Al9P7T/AwHqoZEq+wxlQgVKn14yXVJ76FB0V2Ljo
7Ha/KQAqf9ld7DLQxLySkSbTA4jc17sCxRtwQB1Cp1xqLIABoVJieT9KGNBeg8TFCdnxm1ZNIByf
SdIt9fgZQ0r1mAXo4KUfyR6OsJnmkiot/Z+Y+dFTGOv40fpGtRvN31EQxe9rUhJ37ucEDnpqzxwO
dv0N72xCInyxVmYU8YHq59NcdJ9TuDHowgmIsy5nfpMQzlR6sOjduMN5AOnpw6mULw0oBQNgpPQe
btGlarT46bjgxevQEnvsarNXpFxspQwt5w0KaDETKUJe8+iZM3NENMPJ6X8lISXHMd+M2GKh4W5P
H22ud5lJVaJfNDlgwl+AkUJLw4QaOSV5j9ZBiUDcRtfi6p3OkGorkx4l+vcoFxTqfwNAQtN+zx5d
drEobj4enLC0NEd6s5mlUhcr2ibcK8t/Iq7Agel+6czbx8BMcA+Shv3lW5gezqqfGZJe8/7aVYYx
oZ6fF8pIT4+BOCbhEaIuhwN36xUkW12YU32S6SYN93Fv4OyJ0BXoDd30NLUiiKGtbhG7sjIyudCn
E54Y5UPuaXZMS6OAAm9MUfgmBP5mG3+x4e6CNU9HJbqWNAOpdDZNcFxbTpbudKMzAcxdpyz3lbjc
Sb1HFmp+Jqyztx8pEZ05bAwggbswrVJXbOCYsLv/yEf3b/GdRxGoemupTYAS+xkg2lkSwF5ZlzdC
I4KjJhir9qgPKgUjCEqc6V9n+7KRzs3I9H8MDZlbjNMvxJEgOmY9lRHsIQqJC4KFeZ53Md28I72k
/WxSp1MEmBcVLYjo3UFdcyns/uuFjj7sEWHhMf+lGIcCFnxMGla3QYF4EjwrLYAdVp5ehIzBrlLb
36U845OlVtDXdYaZIAyzwqUOwWNumL+u9b7AjQsnSnbkUqFH0HGG7fGRuaB4ZJIemEp5qMl4NM0u
EPP/PPD5+lC/97oLLmbuPfFDanasrH74Z+VmgBGJon1dmre4gjcJZHmgJ6inPrrDSAKQUSPYVEoo
YXtEDNnRNu07wXjZzLE2Gphs3Ms6EjrtT7ui40b5gfS3hIatW06K3dSd+KE1EUnG6Z8lVwfMhXVB
Z217yuU39rW0npAY1mUGUhjVZKhTOqb18pUPfV7XNHWb79fgeFfKX2zRbNZ+s/WbXEnYl3dyTHoC
HAzBYM7GrQZJ+qKhOcC2kd8EXCpE0S+txQqokmVUNeF7dB94WXf/PYyKm6NzUGJ4pvUSzgjPkrPV
WWTCc6KGDZeFkOZnY2EWGFpcUEjhuqAkwaJ7z/GNYJ74iNz0Cf6mR6D0Gv6+8IpTLlCP5K/adLcS
R6kZ+INrPWazefhCgG3yKDwuISJQygoXZURfT0qjwDzQxmdmaaWAoE8L+dD1b3BbOo0y0PUTiZOa
JZy09ousvuBUyr0WvixHmcq4QMhzIqN/i1+PjN0dbr+xDllEPovQKPMlXHx+u5uN/zL8ykWtZggl
X0GCA17uttFCAAORdvJsx3m1elUx26GW+6d5AoPfuCclyspVtGyFbeNujLcSRVE6tDAzcvSxWHE2
ytsQmHTirDccEz4OFCl9gZGMDxd3PhAvGjVEj7NMeKKUYsgnYNeU6MExR1jN0i6m0DeTrri1zTQn
jCsO+tZ2dn8bvvE/PAPRQSo1u8IfIlk+Ur2H28OphvT2PDGqnaS0QQqgGpzBzgp+Ibf9fOptC0t3
RcyRo+aStdnQZ11on9AngVqqgf6IbALiV0vUkfxIvHSMag8ElUwZRliJSbh2c0YyYnNdoLeQLfnp
sKJvI4sn/p34A4Dxv1CTM22i5c6/YsLVRjT7p4MGJerXzKNOM1I0XpnBVhuxQtxvoAIfKnbVAS1P
4jai8RIUc5j6A4SPEaPU7iDOBGQ4CGufdCRHLm2WAXR+zifQn0ruSUo2cJKAbhRx/YkHE9Oo9C+U
+4UZp8NgVhkrroLILv0bOZ6LzrzlrJrQTIXtfvN0atQ1DpOlURR1I32zWi0LzxTJeeBvwzzKtZY2
h7HmFghEBMC0orMYBRc4LfQVyYM56G2yEoAjRgY/NiAtWrcR253clZcnzOyPMUx8K+3/gVm40Fxx
4OCCr5aTvnmvOE6ydouR6YCoR1R3IyMSpmq17FM41Lwhl+86qfv12nDSyULuIk6BmcL12wODHUqF
QKMD5YAXiAvaVF+atBwmg7QoE9J6d41ltTrRW2or98k+Mpr9ROzjE0m9wLAGCmmTDsgO/mnGqAjJ
NB6wLiORE/3TKs9LKVPPeUCfB4oOojQa0rXkXyUX1EUUFKVfcWzJBBM2vaW75eKW9I5L7K1zz/No
lFIP0SEWViQ+XvDzBemKB5kyBmNP1f2gnx7mrRwNeKS3kEqwW1HuTYI9q/4Gmhpa1IeX71Z2+JxB
v8SoE9ZXONNNDyM/weTGeyOannlssGxFTRkG2Pd5X4LtRf0Rgsqp4h7ZplFIgUSV6frdG7Oajy8c
u1PmDQOGZcbjvfXZVhRZJ7iYEBaFABVC99tUJlAVxBZmG2ufZMk7ocTw3dXMlbf6lbRY1SIwXT2D
uq5rwKZ4B2LAa3d6/zac3epy451aLmNExlpsU2fuK5Tf9SVerxwmRS5SNW96Vu8o7MaxunDDqF4i
n1r+a1Dhw3EQy0Rr2CAgR0nGeLyg99PWHy9zmHCCHXfedgeUtKrJjC4L17HOHLWNyA/1Ex6rU6lu
XYaLP/Id+1OTEvu6lFNM8XqlXrk8oIQbThO6qqQQpLndOMpgDNZ1+R3SAI82DmCxXFkSp2h3yT+c
OvnK+ReYCRdf6ZN7y7O5qAfl5qosXcII53dCo/an1aRswNNN9U7gUNnw+rRGbfevXevjsHHTSkVK
2mATwyyYiuXlgbAu2KGQ6KTh0X4MHfBjH09OSkAq0zfNgokYvW/BIuZm8376c8Y3b+bpU/rtfPAO
uo6VJa2k7PIfP9SmGPiN90zLR4C8AL6iNOqazD0SMWi7t60VJPOwoWHRI0DHCsqV+Rnxsxn4147c
Ed0AcynGLGjVcZRbGv+U8PYDSeW1XVDtnIO6CuaUFvnVUWxxWgCaAb6DSjQPDEK6J/vVIV9Q1ni4
sNYDzu3qGIIuRc2mje5GsVapMVz2SAwU6Isoa1A8dybK7ZTmoTo606Etor4L0EPdPG4qUYPkX+N2
FmScEUbyyazISD21s5/rRG9Dk/z9nvivh/0VSbiDgbPYsoeffCk+FeokgnJ0RgmmXPylPMJsQTi0
NJ6SUXktx4R615Ek8CCIsIs9rL45eo8NBHS93Gws/8bEWa826YAOTf50bRjEJqkyGl8IDITsPdHC
zcdRCILk/nprbOO+/FdYnLb8Ug/V2LXIopQ5AYs31FoCduzGnivXlIEVrBWou/U4YRFbtuRKSZfJ
ryX0JssoZA0ufyXb/UW7YmRNZ85jUjp0pQd1DMx9KfnxARxZZf0h9JFWV+dYVy+xe5AhZDZtn06M
+cvo7RgtVjLTOWiYpZL/cX3xLMnQVFCVW27bJGCh6ZvGu8VUVl5F6tgHjEEl9/vSQj9nHn4wFd5h
W8oYpM/xIf0Xg//5q0VssFpEENR1Rh1BqO+1J8cRVxlLt7/4TJQqF8VhQ6h2UaRy5hfDrvE7D/hh
OptqwFebmN1alLA08uBCllcy6G3jWKyAUItWW7B0+YG1tl9oBdawc6k2haFIULslC3eFo1fiZvC2
Q9R85NRZDX4bR1Rs5Z2nh1CdqmZyEQl8p8cdJp1p5T+887GSbciUvRgfXG16ZXgt/Q7xI2w5aNhX
McYXn5qWArrhHZIEB4g4mvzZYp8lyBxpw7JhK15SYmbL72XNsMsg8zKd9sxA7p1PKfbAZ8EbeDE2
H+xtHK9cf8y+JfzTmeB9K7aU/QpbfT8bDlWbpNX7zRjZyVNoPNHn/Ggb45uvyKlHW3zajnGz9u6X
59+oBd867RXISCemHZWucIX5rXeOufXpBFvDtZZ07rBAxLVTif+r/+BMg3rB7wnLbT5RboRbzcum
+7p/1Q6pobF/2Jnbe4eYAlSTLPYEXJeYde1tRachFYlgepbf7j8E0IWDRk+MzLax23mr1xsatloI
qVfEAxpM3Qsf0rBAD/85KqjXgk/AXio4mgxGQL5M9D7Vk/MfhfUwxqwSupMFHRWqASKy1UhqeF7U
zutzxOjCUwYh3bRMSgUZesQ1DWPyDy5PLXXLb1ddHjFIXN1xgQOCC4uzuhsPZZMXewj3KVw0YZ6g
8LB4gaKynoqGiPdBvlsahZ7ZeuLgfxtYssOrvyJKX+IjIHGKoFEURdznTzd7spqfUSHUON/S7Sz3
Jdomk4qqGkfztru11i4/yRh9AXomldDMmvixG12DgM/M2D8epVexTcvZX9RPahD+1JaV+/fGX74/
a7vlSF4AYH4wRUlDDTKaGi/Vh0K7ulijT2H2y6B27FXdxg0NjWfGRDoQo4tKFV9vzwb/wHHV5Cl5
T8aIEyNeL2Tcac7iADnGv9iEBEO8n+96CrvcjXb7DTEXGet33FltSboAXVLyNTG0STFGngVCmha4
LcDBsTfcn6MtQRftCgEsURT2tQlkmvuDOj5Jw79/CxIrfwNcSLaPfPK6J35aokxkomhwEdnXkoP2
idoAQM7z5jiBhTRaB6gEkkL6t5mKndEsUMKuAZJVjBphqWG5ockKrjgUN/xNgEgKyO/iwEERVbdv
VTH+q2cdgJ7lu7GXDwPj13oVu3OojMvZ+3XvKiCKS46x2b05ShvvyuDMmQXS5x2eZOtm2uSgFHAP
xJ4dog8JS6GxtYdGo7+sYHpHO+izxsMdMyK7kRrsrpurQ/wenizOUlpUGgZtJ0fqgj9ZvLusChYd
hB8C+Sp55DLt3oAyNxwpg30ucgPWS15skmGj65IKaPb0weAfw+L2jZBnNDZ/m+P1XnhWMo/mk8dJ
5/wHs4hdRTyv2uSc4Eqcw1+OO12OC4HdopNZEBISVJ6AYxr5ocVucIQPTBQvxl0uM6DVjQskFyAP
pLThScPsC/tL1fDnXvo1urBz+MLeYju9lUB/A3olNtQWhgfUF0pgq1h6aYVcx7Q69d5Y1OuAKOq8
KATzWwxc2rax0SbOFIGdYA5vdbcmnifvUHOxthbods+gADiWIArrn9BTBTfqCfbMUFFB71cSBYQ6
9KcLWgF8TnBZk2OBUQXZNHKq+uOw/rLau5Ow1mHmwauS9CZHbv1K0oqR088Fsoe+ol5RiKJimXz1
5kfFcAKlvVpwW+2xesenP7tuJXJmYkOo6NCaG0BHkAAVKypG8PK/e/rN5AsUsam3D+O6TB5sUr0q
F/7pL0fnZV8W1b0KKpBd74BhinvRxwSEybbnMurEAhx/72b1r3uxVazLddC5cT3cNc5AM1Erav4M
HFxn6p8i4W7GxnC6klYrXFqO9aOOJoPmPGBr+al7/L+Jd7JuJLUdcRVAY1tNJc3WObOdVZ2Rvwy4
ZQ179KNi8vDfXt24W9D/Sf/mzWaM592n9vDEANgI4g8tqD5GoY9SZaxp7IBqFjSbjBdIv4u8mqwg
t6h2ApPYUF8jEc/PB8DVuekjBnmsVikDqgD6SYP1fI+buE3xd7M+xc2zFuEGcAmcEhN09XapwWQs
YbVkP+L5n0mIm6eTbwMZJA7DcnXFIuDkxsagNaYN46RgmyjwguBN5hBG4oxuAIUbt1MLknJidkK3
Cyfj3hCGcI82G5pLTmzzJGBOL4Du+4ToLKp2RwMTAqKqskENO6gu3prOG8TlHxwn8xBQ0pgCIxln
hHO48AbncC+G3rErVU12G92V2kM/o3cd57Gf1atJQZVm2lY/7dsAdi/fhqg62DqojrtQPE5cEHzh
Gdj05xLsLQUH18L6w4gfr+QOKBcu5fjCxEMHPTaYRgqL6mk/kYt6zb1ELUVcbHbuqYdkPmdSjsxV
lmJCdTHEeQL0HFFdm2sYR7GB5GvBx5nlG8VXgyBNA15564782Zo2BIhYJU4vmneKbug/HwGgRRPZ
wGgGI3ygisMCUY81h2nIKRMwN2AW7aO7ueHdqeUtcvPQ/YLi7utw+9WfuAzy/YeqyMIjVQ+LQWBo
pocPiBgTV1kuWjo6qSvWhTzK3mk+kOzCcRqC8X3YhwcjsGAIqnfGECUxH+75R3Ekeu+Nn0e3WQSM
Cqcmipx+6FSRlWZLfYKWy/P5mRH4nXIwKpKKYBedJk5qfWJxA1QmUycwimSpuh1AlttTvtmcoLWo
zD5QWMrmv8zSxihQivGylAePhMKcmtHNjkFWUxK89Pfr+nU55UwQmOQUjQPDbBmRFylzgi/jP6d+
FuUV/4VqI/PNRF9DlF49Ii448NOGSaFX9Q+nDwSwivRa3sRlOwdLp6NTyJgw6jEa1hbmS3zl2hbH
s0g3A3jlSrtLRfbaveZsYsTXLnOtd/dQFoNCAu82JYEMez8BN4KEu7QiNCieAHQ/MdPkLbwHk8AB
q2lwHKzbSEq2pklSacCUIKIv4fqae0OEAhdFKjSNLnstWSkQMrgoDU0yVmpqIU6VWMIyKdwfBrrE
MbWgJ5NsgXx/CMH/CKBPkOHo4FqskGXhqnFqbXzilTlDyLDElm6TpoAvKec2ortwwfRPeUWfU7BF
Mz8Dj31iRd1V/ExSCdaECs26Xg3WrJMBudPLPMRXnzGm+92HhtMWqnPfKLc0mTGMRkfatmcDrw1K
gCmfM9DkKHNyy2+0GNlJDeFSXX5L54LdGUvls+VixajAv/3zPJpOlwja7DhI5XkKN71iH5n+Qj4e
pjuqke022smNc1NUsyVQ5yK1Kzcou7L6qRuYG4s6eVl0ZPurq7vtEKV/hV66LlJby5DO+vJhyv/o
7hpA+DV78dBIIHAF3WIh1+X5Wb95Fs8AmHFhNXxMrUhXlboUkVGFYo5uD8aDWNGoe7PixjVoyBta
5FeoVJq/EJsPGROAM1/w0FHA0IQ0FdiBbQbBZmbgMQWW1nHwQm4M3mhAyAVI+PQjKdSfSLlIjCcz
z30vQdDGd6prGq1pMbIDx6Av3sYVSQSUfOd8Re1cz+3U9M8QHSmiwbCSOzsV11TwAradhgwGCk+k
GpsW3/ZIlCfIeCuSD6ntzTEAzd+NrX1vskFDElpgazq9h5O4NxDaDUfZWbaIpX83YxnVUAmwDfHO
KPYk6dv9dh3aFPBujwcjqEKmPwoPP9IJNzX2JhREIE+oH7QFt+sFQH+77T490gNLJ7S03LYlGflI
qGwfY2UbNhojSaR4JbxNbaYk74iuKEgnhHm2wgRp4SHjd/3E0FsLSvggHqd0KdPke6evona/GZf0
HuPGCPmYEZVQmHiKGytqOB3T1KABXtuHLtH5k86erV7jOQzcQgtkqTq3p/mg/eiWiD4NWWJSkViM
1GRll3YAdu20yWjjH+zz2SLlYCzToJs4dT6h6F2n0OtumxDxOskaxJUcQGdi2V7XK7KaTXUWlYt6
Wn/GYchA0FeGeTfZIm2AAwFG6I5EreuRfb29SAega/czoZDiIzz5kpeHvMMDe+0W9Ls8qYLt9x5x
KRPvyTCRl8hZTdgAG4NB3Tsj5PxPjw6XfnsyUlUuVD/r23hHSug7u1t8Tx7YSi0qpv6FMKbPiFk9
FDx+zTDRHfjFrx0A+E9fstQmPe7rO5h6C1FYFPdcNhN3TdErCERtRcSnnCS8G6euDwQkqYag9pYp
TFn72wbnHL8e5wsoC3nD4Kp9ncgCWlp+ZFYMj+vz+IlhqreymIkwGGx5SyR2Lijeioau8dOwxuy8
FywGqxmU7YQqJS+91GjE37BAtThqBeB0kn91yQQC+CKslcpf1PG8GdctiwRwBH0NrZFdlMrKS7Eb
92AwlfsX2uYT65d+MVvtECz6eUHu9nbDtHbjPCwuTJUsXHcNbGwNq6EZzlafRE0Dsch+aJQjTTYd
R81oV+TM6+mSNr94fWsLQidvPGs33XJ3pTL+iuk9udPuzym6xy/vHQyUmRyn9/6LxuRvi9jH8Ssz
5AQ5Espldzzcp5qYJdVRjb8VhOWcm3cRh8RxJ1c0pb7DqPIS6rS+o79VjlY5AGnhwGCgj8IAJsTM
8mkNBxDGRLo5cK5rmXwVThaoHHtDGFa9Eoycs98fInKYqiVAguJpAh8vAqZxgu8X3Q/bQ/77usuW
M/swnkuPK9N9LsbUC1HKQi1jO3nEQcB0zkmwzt065mQ4QN/ltXCX94xPf88PsrE6grwAp7dHwK2a
jVyqr9SepcfehlExQ+Y8L2s2Misp10SOc2BF+Mpb0y5Lvo9s9IeiUx0Usq04B3Ljr3DOlJbxIEP2
n8n4ixzyf5A7RiT98XfXBr83bkHGsGwFRnoPXRD9dRHPdVvFKqfwRxZC1ueXokdfYci16s1yHtAZ
L4PxzhzpCodiX2V1zHD6aWPamTNw34EOZa+pfxah34RBvPWaXC9hrv2ojOSGCLwWU6F9R+YpIUuo
eq6zwYbBEC02+mO708lNvjxP4NhoBd2hx6FEqSCWFZeU2WUkF7kRQdfqS0on0X3UF95/AqZpOj+X
jSeYmCihCOvY4mvZvc7eu+9y4AS+GcXCOKTF88RucNU4a8id+dzz/L2yASL9PshttUVIRB/PwFL6
Z2xjgpr8PAJbuqmplaexQNS5E0/kFKaHHI47AoEi/mPOv/zHcYm+TVcGHk9UaRIhM1dT4q2KFC3Q
ib9ErHQSaSVQWasSsQWLmN3FP7EI7zVPZXcv7W3jWFIAI4/O1E1Ay99mNyUGSDeLIzvsRn16Cs/l
tjbFtJle5G4jtj8vQZamQAUhVtaTLkfvBBQg8WceuEkmSeNfs2c1KTvKR5llU3IfKFNh+OAYwpFc
L6WX/SMXmwmurRnHnQSqimDZYpT8HPL4j6NhZNTVAth0JRgPycresNd2AYtk1iiH6wvBuaV2QdqW
IicQ78TAV14xUYTuxKxDJDD/NCN+d5ZEIhmHNR4+Hn8nFNmSJPRmhvotkvdGKfNlyuw6rIHlpTmP
VKawhIta24laiLWFeG7/5G6YKwDIm6ZrpP+o6UY/Ia3Edo/l/E/bylPRYeQCKnwP1Wm+feHsokJw
TUJHwNObwXWw8YS3645NK6Qsa/24AIgfjwAaoOZWbvluexXbWtefCYi5QuEefPEioqj4+9wCDhTr
RwsoW9spCKaMIpVF76ChihnVOAu4D0c8iWNDwJZMA0f2S81e2yH6iKsE7pRtweiDBhB3r7j+48A5
9EA9ktcPOW4aRpSSCu75hhrFhFWIMGgSefgmWvpsOKdc11irTZKxNZMhYrk+lBdl/T4EKDc4CnrP
gaXS5yBgqWhXlt4AjD4YbDHt8I1/PmpJ2+10OVcs48N+os8cVgME58GyFKq3sN/oJTzSI2zma0Sq
/e+6GQiJsOjFOp5BbcWGdHEC955EyBwo2efjLPc4C1RBCIL8Qbvc7/6OfxOLcWW1Br5NU63NuVMZ
dYO1M4AgwJ6sSh9RgSPCZhRvd2xvcgOqVFMEBWop2GRhuqUxUtyBJi8aLBFX3QwnBPLLZYGAwqxF
+camyVxbUf6wY7cyX6uCdf8rquovkyK/cF/Q5ROtQuUGcP17sa2rqkUTFgPsiCBBlX9YUxRzxH5C
BOHUkoSdM81z3W7g2Gx0z/e1sLWw/GWhusluid4sx9At2QXfKAehHPVjhwA+FpgcmL0Ef8jio+Tt
CU5KT7e4ICHiB6LOkgNCInegWjR3JQ9ahaSxdWs4UQQWST+s48Dxs7SHO8Og8nuNIPbSjHwtQJCJ
HYwfy3FCIrhEmHNjYKWGnyUomprcvm7ap6lwt8Y2Q1NKxRZSu+FM/Gzw219u9m2a2Q8EAFwPhtdP
ev55U/mK2pTLQvogjEnipgOVEBecAu9a2xoS+hr8AdRm4xruj/phNbQcDppmW3MnYoBs085JIX5O
qHfk0U4+0J7tMRe0zWcdDsiBhJFld0SVbLDhHsuAmjbuoBgK4GkTHhidMLqNw6VbSt1swU8Txuvk
cFTYWYttK4oFfmCG0WM7Jm3V3DdOHtEE2M9dCJ1mmmM01Vd1kN4eJddl661AK+a1kvzBrTLHT1uR
R8475YMZW8F6YwIUu6g32sZAgl5tSHUEgAGfqnopt+uW0mTC3wwjC1/TJiTCQV/8D0WigHwQyfoI
10sHVPZEN1Db5xUsICbThp5Wh6F6rQmQQa687PuUKEiP4BB/dNKNWE0A82VxsEbLMPoLz7xaNjUc
qU94IsylUbUo6LZSDLLHcUBv7ANEZpqLYyEdMvgIaL4IGlMnc6mNOV0YpSNjtEQwQKv36Qo/37ju
+cQu29r2NdKFEEjbl1kHzb2B1twaJGf3NSSqgFD+LDgNfT0lSbWQes140MWpy6W5q9syDxro7JYY
QfPDL9Yr3FQIDKsgEMvHt/jhTtEHQSPEsK33/YVsqAKUTgxciXeCIrdnYWnHmLVKto9fLLyJqZaP
mNMl6Vlx8daK2M1JRXF+l2ZaiHKt7n2B8sug2N4eV2J2/AGYoRhCF06lvHfoKCD+6enc+TdoKegG
m2PLReAoOKweILZ5RcVLGGAsg3opLVI+S7Fg8KwcGG/L8Rr0eeqFPLwuxC0SndggrRwsk3u38u9B
vmq1u2P4t/c4JNr3/1HCVUBBQgVpLdjeCyusHBvJhzm890PQL1ctrzXoalBtIvwTVUaAY1SCgyYi
C92iYtoixQeOokS2bfQeuQrhOGw0OHQ/yAeI32gaPRk7vYEI/H5mh+Rx2rsZPNuoSUeFaJGdpGg9
M8zWV0RyMsYsLUsgYDiqorQW2PyEi55jhzAw/uNz/nPgZxfWSWook0tX1dEIdIj0h3ThJPRksv3k
K0ah8Cmcy1llId39OdH9YP81oNflH2keaMdRHS63EDea447RDOmxRcJC7dmXf70XxFZNub8+ZEYj
IzvxXzsHc7AtThommRDQoAZmKQWbAsm/EIjjZ1TvSaNC/1vgBLWec4ncfnW4z91GejwcOdCVjcqt
CDNZrq3MfxJmfICsB+xnplmZLkiRGWcRK6WhsWLPWltuo73Toxr8LgNWrl6JHCEtzYa1LPQctmHo
X3HEq7tgPXxMURAOxDuaWv0nnr5bofpPnCCcWExZcpjTinSBzjp0qh+0yqI6DDY5QKOxXwICCiCM
b5Uvu7E1CtztackflnqqTgViRFlHlAbCKdBR9FpXcJ09izeki/Eh2u4Qs+brP3Guyiusp1Tjf9Zq
VlignPKNap9ASuC0mtiiMUeP3d6MrmKSYFxxUIIVBcV6LgCwTqjUXDcPhvVj2z8fsOkwh0X5fxdG
OmiHJeCzsL/PTzCqLRkbhEmP8d+k8O+Ee7AYIBbGSYhzpHnIo/nNOMu/kk10SnqS31TcjRZNKole
4v9tkKhEkJewP58GnY1h+GlvddiS+noiiaKuX5KidEtwsD9Sxci3xvKeWGdcpEwbr8p1mlBqd3ad
3YEaNZQGFhTvg0C+XT+i5c0Up5HLb56yDZq7MAX/AnWDnIM3PpkeMlx6LUVod9w/Av9tS9gPJZG5
jDTSeFOqreKX1kw8OHgDDI0f/311bT7gRDJgB8KTkcXryPfqgH8rtWc00/SAHSG5b75hGUYDHZGE
cLDDUKPNSxZEUsqqdqiN8Q+XGyK3cEURwALoytLt2Etq/omn8+HGJLzAsLFQ3lOljUH/2mYYOIB8
Nq+1fZxEhr4385/XhRirEuboT+MN92xUNNzS8Zf/P2rONYRlio/1cKf2EMtr8fiiBfmwO7kZL4bb
KqXv6hfo2xGqrtrOQS1wniweKzZhVmJ852Wz0L+EU9nbBh+BObed1/yNJjg/RJ6ZPlVkHVbanzrp
xTZmTWhCi/eAChXLmpxK6Mnxg45q+xrgDfEhJ1U6lTk3NQIY3+V2KoQTp9uiKnMoZ2CkBbWpNODq
azapqyg+FmijPrcUQ3qrQGDnaSqTBrhh0ByZfSpEdUbY1CemH0NIzGOES6Xe55RcZ3GDstcGh/KO
T7aQTXMd5UdK5R4dGJJLQAAZXi9qzWkU7XqBQ/4gV48Q29mZNrsvk9AWbt53H88pfkYBX5AZeq6D
1BLXPCnRiBEQGDM9ZBYi0q2eHqxAtVC7RC4Tj15jXSyMIPUzv1U7ceStkTBJlFZZJ1WERT3wbUPM
hc2kzgdX20CWJXLpw/0Kr2GgwxiQ9n2KGAoR56Bz7lghfFA37XyBjnGH+yO8dHqUiwyweqQzDoex
osK6u99XSGdXoAZyEx4MoU2VqPSANWsPTyMaiGXve7mM4m/lmfHLZYInUyVJFe68Ti2vvEbEK+M9
qdPbpck+MpNF4XKsVo4AHwD3OpYFd/OvfjHJK/uD6US425kBuTcT+yHEc26r2T4ypXLChV6qJlR7
gKCQIt/OV+6UnkSC6xSXmm9ijY+YsQ1+fyifTC0qskOg+EcqWJN4/PERl4LO9ALu7fTAduaaiLcU
izTqDu5JpohFTIjqK7DFaaJy1weqRTv4mlzHhg+Kf+7OiKCeadAftl4592b3IXiPicgfZDnX1LXc
Ykq/TIDsWoQDe3iX0HeDKbqpMdydnu9oP3n7ROe7yf26PkvqEAXiuQslrh8RXs3hjfaO3T3EzTpg
ByXtZ60MmX97X0sNDisHVKjtUoEusqu5ZfdVfchkN9o6FN4mR1izh1DrPsidoTCR4U6fNuDyHd4r
lRe/M+x0bS8Y4CxOSf6mu3R4+KJAy+ifTyl+UZUvhYBCTV8wpfhWlHYn3cTKWihmuAaKjS4LC2e7
XphgnUM/qDc55t+0pWSN9IwYMHIQucjaHDYhm6YevSJwyaBJoRGy45nl5efxLyMgZ6ACMC7YpIHE
XCffxbkxd7D97rK/dNdC2um5/00bzeqUzT4214pJSHCbtiAteGQE5KMkwJulXMgp1s+NYDqX/YdM
Rm+Om5XgJopeIYITVr/AhGZwTVrpLDH1WDXjhvtFmU294RoPPzQzQNaB8Qh1NcTKaieuWhlpC+80
P1vpibV3uznCNI1mn2K1gvhvsspTApm4P/PXrkOJKyslr6Qvm/KGuc0jxT3SmLwwvio1ND9MkKh6
R07Wlf7SXeX5LYO1kgPuFZM6KJBc2sCR10LwOEL42YPlLQECGcJABZKrj2LhTnB93HML5ZOI8oZo
VuBzmEK3AlIemfU4/1Ow3DRVVGKm0L4rdBEyjb9NxA1AOxrf+WRz/wgoHsXaawTx38x+M5PZZ2FR
MlS2mOD9/a3/r3L+on4WzM+VcZuasRa6/iJyUIV2A/4jeS9E+9GgwjpBzDpiSrlCxLnM+PAQQMwO
ysqdQnWhivC2sQqcX4I6ErAXhC4tYDqZyrIeLY4kDC+YqeQtnL82T2RBotzqHgWZ7S2uaJQO7pOi
SgfGi2ZXFhOT5v7egYHg0dgFUSkCW0vE8VK+3sGF3jWpC/4V1ylFWTS5nyzHSELDVi2SpO19D+eV
3DmYHPjutoWp6r390uQg3Y2h/3s7x2WDqjo1vXEepQJiE5BAxHwMYn1GgECV2qD1xJ6/Wb7rJd33
ANbJP5fb3zshCSSVdZSZRyYfLFQ9utFpp7akGUcPOI5ZLf8X4x60/fe96Cm+42l4Fm8r24bxSrQ/
LMjbkq5RxwLO3M+mMaW/qgT9m6Jncpa5kNk37fqCYNK+Qqr7X2McO3KEYSNxw8+3Mcll0+ZRJRKw
sGAAxIAO+eG1YoBxJKr2Pi+sW9q0B9jRDqne3+ZyVoSnaN8l1Az1gAwGCVEQaDXChB1fExuPlNbE
Ee8zJoVHyzGYe5YOsXczGYu+6b5GHXXDoMnqKB8m4HFICfHrkKcYa+27LwpezEyfaaOnbnllZnA1
HLIYYS5zE5XbUVz1MdyZNJb/vhobV4MCopEr+XRwyLA8u3SfyXIHo1pQnfFRqC8SSf0VMO+Y6NX+
xImaR5hdB1QiQIfq4UpZrJXBxc+itswxAOI6Ko0U2xnm6LM9GDrKZPsycUObfkj5TlycjEyrVBUV
AdVhvN5QSZSULECZY9Q1aXzZ/DSk1XsY3KTTTak2vTBDZEN0FGBVviazmTeAFawLOWdvtYWpIp36
QxMx9doQzvLZ5NLVShl+mWfwMYrscwGgb0GO9bJHAYdsyyG/AhNiDVIMFx8mXci1CzToKx80Z08q
ZH7gjQOxweA4QNjGTkVEBth+nGRmP/pAxXNoDmHgkJIfXGpO1YRY9MEg3hhagOR13EJNmkxAdhWE
xlBh5PJS/GKO9VyJida41UU6CXfx1Y3LTkE2oQUKN+sGmaYdqB0dxWCXOKT+dpHReA6yUe8LE94S
1SgqOBG1X4DJRZxV544Fz0p9epyr5Ow71RANGXobuJpvZ5ZPj7Eiujc1WD4ONuFXgja87mcvkKsS
lgD/Mqi+ti72/fYj/Pz81b2PKCpVjyN+xETGAFMkA9QCEaIb9TrHVncs4cPHveoqOd9OqgUES2e+
9ID+fpLF/UKtGSJbQbLTm0EobMx69X6ouOcDDsAFpxhrc+UZsuVbXCJauT2koBzpBdjGU317/0xM
2f6J2d4eagGBmBk+juVgylzIRhD/hJyySDxbEJRheEsVhYWXeC/y4DSXH+IYaXyb7EAI3QcXbXnp
i5RzdGHuZVoNSviDr/BTKTeKHf3hqnW2oEkuk6F30At1y/DBwwb1dBCUxRWq0huurWAtX20zAu1L
OAD4xA7G4KELjMm4c+Lwu0M11m1E7juI7yrZc9QZksudQJbsq1mwIQanSCqfN4RX4LBniQfR1Zw3
2U6Jh8e2YH2aI84NOrS8u/Ojpv/lTeTFJD1PWkqQGCnmLld4aH63A/FEoUbAlCRluWQM3zZ5rNre
OC8q3JD35y1+Cj+BOVyhunAv7ryUwwCK1zGfvj8qRCyfQE4pxvmnpy7kGmnzXJkn+6eOPl+Fe783
SQBraqY0nCO4ac5p8HMsGCI/VSpPTnx8Y/9TpF7OaZKNXqkpnpDyMKfGzK7ZGEpfZY+FI0XzReT4
mQDm0BLoq9JhPFZfdQZemS5v0fTYTod/lGwedu7mzrTAREgBK6QOgqqCDeCxrjSBMeekVwf6VYwx
x8wMO7yWkiMgSfzXE/3IOW1l9S7JbT+S81cFwD0tBtN7rc15mv6yrwZovTguvlIqhrx5qKpQs63v
/2Y3OLEglIOjGKWdGnvZ4aUP97OIHFVL8rNvRlLsmgTvzdhigAWKJeewv8kUvzfv7FZbyA2rJqzQ
t/awTrAuAZhE4Oxr/U8jY4z+sbT0UOSXMLwQWzudLrlHhTNkm51Rg/eG8UZ8QCZZ0q18uChEIlDs
anMQU5EaZ1KSKpn7fOUGtywVL8KuPrU3SuaA9t4L1cebQvERTD5D67puWmycec8QhTMvSzexfrZF
hH3rt/znphXmmSvhuUeB577RZE4Sril9vc3sxjhP1fOHhYnw2vKtpYRPUfzum/xLWWFVKx7bYEBw
WXVidnu1lCHpiwLY9kCylZHwIlcUD1DRxgZBhjpNcXCN9+uFAzf8H9Q6HRs0uIEWsGFuO1Wt/XS5
eD/5EhDToU+YFczbU1H+bsW6ARLYd0JXcwG61oa/HqdVFgFU2nxSrVGwKZsYb6Vb/jTZyn9OZdTC
QTK0Vhk5BRwjD/T52kUBsy8iSlC3n6Q9UiFQqNmjed9+nj2FL86/KuExnYjkicgYX4MW4Q3ZEr0r
dZnjdieumEYWWpe+bKWf7owrqqwVtMxgYespAwj4gUW1HyfOzk1yegvkcTapkwK6TrcL9u0Cn4ly
KJDF1ShcZm9SMrRC512pWVU0eAA6TELGJoUaLw8PDdKeZpsoojDn+yjrH1pUS0A6IwwADMxDiEp+
tpS74XqZmLqdJR/Id/sJyj90hoX/wrwurlEELgt6hRtLTAQHyFUWkhzEAcSbmdbZVCNaUG62hHno
pEF9W92rVe2Bg3FaFd/aC7xDv2XdDVdr+w4qNDLzKlaKX/kFSG2vdMFjngSXZdkwfoTSCnwZeCJe
WNzG7wbUxG06yYt/Lw+VE0iIihadaRNUlNUSlwAvKewIieFzPXc1Zwqac6Wb5z3Y5xsPNw2q+utD
PoNvx5SQKOMBvcuSE/f0JSLL5Q2LnolLc37yx7EyWqgKJ+QKk9aD3qsJ74TlAGKPUCYGb9EHWqdR
+7afiz2bQQa6vNvnKbOf3Cjq4kPaHtF8odDQfcrgfi+BpVdz0sG8pnjFScI3jsSnWsTKJrFsFIn+
wPXQt50dLjjqE3YJpgc4hpUxZL1Ulme6ZTsV259L0EjzMTR2VEWeYYn9rqRbqJlSSX7cuEYNOI7L
Njf2P3/mF8eoKTxfbg2eRSRQFFPyer2X5sCNP619y8LExgYIJbahfgqcIXXAFwSSNkWMHZ0w3eco
Le7rHYUsPTuemegjk5Kvb5hwgB0ZjMy/gZV0lpCG3oEOkxRgshxN68Gw9ai/Q5L/2JFEfc96K/Er
rCuXlPWb8wnQVLo5CIHnVeU6Ks2Cck7VZE2p/Wee1pURAD+ATCOBS15zTCqC4SjFPak5tDccr70s
KhUyNXBfVzylamG74h6xMl1vvxw/D7axVn/mWknIZThrcCyVCr/W7Ar52lZ0GIQeafqyF1uB2m/y
DhvCOVVSRnRWFOO/cLEm5pQD9GMO0i9LDoOCXR8pamn+LN1jKAERPNNSmombQSh5RkbmGloCISHn
S1+MDGNdtB/axpCxMRtFNlWumT2lTlvy5OQRSTKp6okig/Z9xwU3Ahee4pvWLv4AJCzXoqsrGR1i
9Lgp/4i9E4O+VqMY+kQUG1fMlC3ZkXlAggACdwJIpnpxe2rWO5AF/EpysqBFi1RhUTN1IyXoO4hi
X+zUzGIEgn21nsJ1GAHmsaYqLHRT7dUkZsurSVHjkkucBW0yUeP6qFIPc6sJ1+Wfh2uF3sHO7KiB
Su1HtBLmaSSeOSuYLKQ7S3L+BTjmSNwSn6tz+trtThzjClVSrwkFJsdYSJtLJ24McCJ+t7Iq17xv
ZCAwLe6gLHMXl0chOqzRD0zLuCHM5Qc638htzAo8WEndiIw21p3Kq/mqIpZ/7A5sFigEghUF31FD
bdpRJHaK2o+7j61jD6xB27A36j41EHSM9Aan7lmh+mtvVOvmHR0p+jSyKUcFumtK0iYfACX0OJtY
a9CyO5ZCazxrNgGhyNJx2GoV6dDd0pTXTQEQWk3QzUM+7yIuWdKbMHez6FiPnYHi5dQ+lbvs/Hx6
+LJw2b4v1phymGIK1AO2el/RllcIYhuxaeynOT/7k2Qh6dMVyhWnZFyIRd+GEuvfdMyA/SZD3Mpj
CMrDwF7/kVTtTec4s4u/pJCWMBn97JEEGifITjHHl56bzcqwduHflN5PQV/AVwSrEOy6Ls8JBZhT
zr6nDktrS18kYAl/zh892EgYPw1F8azARRqcz9U5d3yehdORzkqAYN7Wh1vWMSfds7TIT38Me4nx
wYA28o3QyYGDmMEHImgms0FPOUPoOzFRgujbnOPNXoCZwsa1DVI5d0TgPsctGulKZoH4ds+PngvQ
PiNTfcIPFh2nm0y6vvvT25bzZ+kUf/BwZE2V/Pge4i0qWW9sR7Jj/R/dvcklctvRCYn1gobiUwvA
ESKHjOphdc2b4gV20Rsc19tA3abuabJLGYkEiyJPj1Of/rExGahx7MTotAvib/l80c4ywUE7TJmS
GkvS/p2SQpqybDMSlBsF4E6e+vZHQSIM4BBVEjn2I8aA+sbVGNut0UBfoWpYeAggyDcn2Yje/5rY
QzX9U9jz2WG4eGFRcUobNMt3bgVX3WMxe2anInv5yZEtT9/4LBjY5FjuBjeyqlZKisQXu67XIlfo
YE4vpcXG4Dcpg2Tb6Wcsc9M/29GduasNMvdE/rREN8DAv74uaaZAPX5tCn7dsYC1fSp44Z6c0ooX
p7We1vIYn4jMj05cYhMKxo+l4GMwL+qxgL3viwcZK1KSzfoBcw+EiLLx30Ouv6Ysxl5GrRv5qKFX
3GOJuBu66VmpHd6XReuEnf2VLqml97UIOByCB8Ouc8CuNMy2rJWiX9WvO8bkUSN7hukMsnS72X+k
0JK0bTVPCY2MEwmmFjoTqNtTSSHOxzvOCZK/56zee6koga1fgvZ25OIlykRVxZ/h4GmHo5QWuW7s
nR+aWpeGdPKdtZtPhW6mk2w2K5DjOozMJZHBfotVbLIq6UiUeeyEd6q5F0U4dV7ooOV6k0S/PCoG
Afo4hRYLIkZyUANYInPL+Cgbrw1wJd/bjhXJLr1AgrR4qD4wXJyYxcPSJjUQAefj4Kp4Sd7mRHA+
F21F4YknxLfH3mlacJuzm5IUDc4k2oKj2qnI/2YuuOvDz0LWsIvOLLrzDmS7uSQKz/LEnyq+vbNr
2U30hJ+3zjcgAwPQEYfhoMP28twDCO6tzEpyYzH3n8hl1rWNTiWBBCProOj0g8VNuKZQsxJsSKBV
z8loLnAd7BMketnRvOWuVnxBRX8vBOdsuFqqMcHrOqc9flScjlVl+i1AyqF6Zed1hKBEGiuukgK4
W8k628yUBreGc9RukxKaf4bYlyOinckAxL2J/t9gzxe9n5u2MrDjrazvNJiv0mphSYUg6pypFaai
EApl0EL7TcVpWWXlcwD6cV7d4jOXnUSF7w9cRpHf7vGNPDeqgW401Z8nNEJnQ+2L7nglB4qWNRNx
YnAuV44Zq/HCCMU0+stkilFBoX8tCli/lciIY/G4OfT2nD54EkDYZ0rw/0WLnypwwD6hshqppGgi
VYet0dqDd3Kx/S+dXJWku7V9AZJNQqko9QK53ifDtRAROKXB625NXuybdaJr5CkXu0KHlee+rvg6
0BWFoVk+8Ld91TdRy+NT7iatR8xuxg92dpaf7W4bNmM3+p+qy2sjubXlaONYdJhyRyoX11Y2VMB1
VJ+ztETpd0cXaD5jFZARgF7lKH+Z6eSwK51AnwvjpJ5fsl2wPLB6zk9avErLXhm3oHou3OQbNnE2
zr3EaoWtOq5hXco0Yuu4cWNVD+SHvhl1C9NC87rnNiVUWpgvIRCM+sZ8dMeZiquD4mYbEsM8hLWT
AInexmCrYtvPx8x7NTTGNvXZG4IHpe5l37y5lIx8jY6s2UQk6+ur3BT1tfMrgbSWxcbWz9ozEWCK
H6qVGy/0vWOgB2RMl2DSDwhxNf8p2p1FrG3muLugDZRIKQ5W22eeRVIFmLLHjWvIstF8cLnJN657
D+7hqUwG7HQ9DNfFbaJU2vM9yZGxabBgi8QsQ5Gvg8zxoGClIBY+hH9ZtKOz2Rw7LRuIYPxyBwKz
IZ+ZoApjbRT/FvCM+YtMaqEMf+C+8E/5NGJrSNq4cJg+mEFENmNcvReMzOUvzHIY1Mr997ILbC2w
LGnLe+dZKgU5UH0XRwAGLefGUePTppyHzLS+cLMd/oEjSy3qCHu55AoWf+0Oj4hYjsT9RNVTwAjB
CWAnaA6/u2Ma50UqEIq9YSgYJPFeUSAoxHp7PkXTn8HS4JfbOYFtc2+xBDE1uArev7er0JrsSDU/
fvONyVzwqHpmXJi0eZduipo8PerR/Xe8FuBD3qJ+clBGSMbTDhI130ZNkviFNHmdP+NLSAXxITbs
UMcZavoiIy021SPG8M/Wi0Ck5KgATjr3a3gSPTIefL666vUvuh5ieAHk811IGXzyI3c06UEyNaAP
xz9IcDIKvCejSRC8KNwFq8CWR5Jf76KfGPHKA58aGQV8pKKBExMnXdl2rbksYcQMj7JaNNfgd/HJ
u6DXJY7L5vbMETDXoXkArUpLy+kUnVmgL6Gl4HmTEmpUoqqvW7YU4azsOe6LRif6E3+GI7EXCRu9
0qQ779XpxwwyjqUY68uVJ3eN7s8Q+bDovEicVPaFKQjhNzQL4BQxk9Tcl3ZwWsd2IGVWIlgqgoJP
jVYAwVHuxHTr1CoQ5Rk9KMKjvmUfvMogikkrWiZHub9Q1LDoS4Ptp/HFP4BT5cJrs1iOPn3NM8aI
IQVcZvycJRpamCJaxCt0UTsICBips99AB44tb7syilKwbZyxIWBJ/nx5e+WaAjTqcKusGT6NS+X/
aJ7nC+Ppolfs7rDhERld7DtVKadwJ9GQd/guchkZX5BDdQ0tzsY7KZv3jB8xx2QFvVh5UL/Tcpmb
3pC1l/6nGu5phaRFfkpXe05HRp5vUKCw4P6NHxvCkWGDubeogZZiTyrTgCxhOp9TKCj7m6WA/svu
IIB7MZFE0F04e4cnkTpFEbqeD7XHkIuWByvOOrE0K/m/lBO6Zg1aDBK1airxxeM/S8TYOu7w9Zpk
6zxZUkWcKzht4DaRSBhGWzAwm2yEBAXBXK53lNwSjM3HiJiFfxv+p5RHfBDXYucuVh3ARedL8EBj
KxwChGyDDNmMYVuniXLUbnj/qNCUWBY+1cqJDekGffSJmZNnye49vjLFQd2R0Bm/mRa9ztBNGSvS
BzsV5eltNqiXilwaRvfDYp5rpxNZDO3n3T4cgF568SPupnb+NouVyW52Bj65rqzfacOSfAy7Y8fa
0nshiYLG1Diux0EmVew9eH7P+RT/jkMlQj/t2BMz4KG5UQpCLAuDcHTWWRzUrXDYAkdk8slki8du
7fkFtpSWkSvHGHXekSM9gqSONGfdoeTrf4bWoaUs+WvDim0Qt7s2E1V7EYtfOBxYY2oSs1MUtaeo
olE1Qcsrwl/NE9j46iAOE1we2IrQf2CO1EpCwD6gjrGVdadcQeXaGEd6ptlDJR0N/an40eCM35Qr
ZZzu9TL/RFQZ/tGmsdJXqRiCCje8aemZhSqD4Cih/9MXP09ociEU3ITDoP/kNo4Pq6MsYsSA0cqs
0AEw0J6wwSJGcFkOU60nJqGeNGNsiFDph9vEJAHYhT50l15FXZfvIZC+CuwEI+2Z6Vir9R+VUka7
3pD2l8hGZJI/wWuFP3vivXNcuLFIdU3jR415fQQNc1p/eMS+Ec4av0dN/HviiJYg61RbmFIeYkcU
zfo123LWO1GdQC9YHQigxHrroY5Yx/bXxgdzqNGXu/0dVVHosl2TjeXyBkDo12FQEBc2tC9P9o4H
F4U+1jMx99XGCjhUhd7oMJUSgD6MUChK0XpnNFEbp/hVZ8OtzxVTGklMDnGDGB2XxSbSCsgFYpdC
YN14X4qvmUJyFTMuMmrVnVaURvZqVqNtSHE+j5jlHHlchW/02G+LjFLfuO3xlPF8eV3RvN+nDGTe
ekYvGAVfjewY1hGlD5xVIGKSVNlqExlfykDXKBmFJi0ZWwi0oTcykfsx1ceOvEGnlZRKtHgMXyFq
Y2FZ07SYv8VEu6GKEe2Tpi0HYLRaSF7Phfz24BlrW53aN+3bYMYJ0cP0Jt18cINIC9qyIoMDFIWC
nCymMV545Mnqsn1cOiqPhUS+LJDG/eTRLCJb9wY8e9Nl0ymZmrSdOEhK4I8CSV/Jem5p2pn52gpT
O8/+bcAd5B275n0WhHF7NYB0wpT0OkbFeQBD1QAjODdjGGYEMkrQMQDpzu862kHJq6F2mNedq8Rq
l6MY3QkOYlXdh3mHrlmvBzX9NS/MVcqyoZxBbfz0wFITclltoVQuf63gSb+QDU3PPdRYn5KHcGVx
jHg4XZZbXwdoCfikKpc3R42Fd6TnTXk6C+vs7y67tsbPt86VaiEDfbTVQw9t6pX/xyRgnDbAOCnM
yt+u8wKMwCMpdPgNKZf5SZ2parch/yynovN9ZXuKF6pD3BHxvjaEyi6zHqt3Xm0xw6vHClJ24zrm
JtapXVFNk/a/EsjEUJw4klTPFigMybZ/sGP21PVUzj1R/DbwtuH6RDM5oAq1G+Coo8UcyIW2YGKG
toC0Gr1o+tj87ZbGpU4yl1SA4fCTetNAdGBhkJ4gHjdyRRPTVAu9qQne+WgLtR/WIP7bYySPj0H3
DqHdaW/gGehK1hyx8WU4nc+IRG8HXS1rR9wVAGKAUwngJxY+Eb5gLVvUhfmFMQMJV5hWNRMUgt+y
F2STqtDDpLZhne0YHeo7PXXpibmF+xdMeew3lgkAlBF9jEl8J182bQsALT5iM3GQDw9nEujIPI2f
jMiCokl6G+O8KbIDZUfIR/caSaF5ksc/uQ6XoYmmEDginUJpeLe5KaLpf8PT26KQTyHwVx6XBJtW
EP2nF9pXigpKoZC2IXmePURtSM+o0TakJzk1k/pHeCtWahD54vHgDZFxxhemKDa7pOiqqSZMFnmS
Y0Z3x3OwrHXVs1tCQQE3tmEoN9/+ar2hHCU+Ns0FJBSVVe6tWG5Y5jXbTKDrKrXyXDlx7q4nJsT4
qCCm/py8WQI7qbtqxckZJck/9l0drgBVVyF2B0V5CTOwubAhVuLltQdB6pNxDmfNdUqChbSS+8CI
dh+wqWlWkiYDSWWVDjd/73sFhw4z6IoBNDI7ehRZxjoOlmzTU07fN48cedDl9Q2QHcpmZnBjqcFg
X4MHQFZuCzenpWcgf7PDg5TTGDE/lwLrPDyXsmvw33zeYnXj1tmOEvS0eGKToMnSClgfTmyKSkvu
EtMUqskX4F0DgtWMEWmZaEBWWwec9YpcgAdMFc5VRBC3/1Na2nuRk0mh8UOAdj7QBRw96ciHmtP+
obIchgLUtZ83hysIZWZfikOJH48QBnY7Cdt4XLriGP2/Ya+C8WpiImuihBSmoQXn8zk43y58rmrI
28j0i85SRAwdOspz3R82tMvXyrlD7yMIKailMw6mFnLMggKmQeDE8Ges8k1wq/iqNhoHnHQvHge1
jFmWAHfBCQlzRg/yBd29NZle5HRtQnzqRPgSxyqAvwgJS/mGrH2F2UV5CK8d3DOsW80JlRLA6GTj
1E8yVUJn5gkPCGT5PIY4oUgHpw1rBbhQYgUOUxdOEDfc6jEwVD++VEBOKrbtGLC0yyvwLxqfERsn
+0bmDGUbC3t1/vVtYfbW6Pmie3nye/MhitxLm4eL5pIyaAEtzWEV3j+EwckzeoSORIqdQmPb1SMQ
Zsn5cKkJsq4Rl7M/F6TUJpaKNdCSzYdcpOssmuy21jGhoP3jJeaPmnnLDj6Nqlmu/gaVZReajQ9F
HFElXoYzZg7B9ZSNmAITmRESOxNC1mDyEMraocY+EUYtjqWZU04KvW8ULEa13GcFpysOH+LVXN3a
5dKx7MdsyK0Ub9c66VtI3helZRWbVRmL8CRNilm0OB6cNHOL4iNFBsgJQeyBMIDcn74kwzMNjShH
g2ZLtZ+HnBPI+PgySlnBQSdFmaoZg3j70GL+z1qWDZxD9CyV90WMLMsRdNRBlcjx3Mdc8N3cXvz5
ykYrEouJXUGjNB9ZXk0HxIMpZDatyPIL6GzXF5fvOl0MdZs3oRtLAqWUg6jt9eeAhS0tw1Jm1QZN
Yozh90vEuKIdXIrAqHNbb3IGr/UYF4KMpL7Y02BPfkonzwh3BGP/xTnDebk2FIj5Iue7qANXTzex
6gv7dmpTl7YeRq0hYjHi6obiqrUGupwgXCpqQ92ENdtELexTkrMMgxzVw2zZS0UgH48Z3OrK/AM5
ecxMBDcqn/Wdi2Yuwo/+7SWrccaOWaAy5LIzBMzHZ5H+Hs021wgG8YVCgPXq67dgj51Mz0HnHx3q
szUieOCIJbqkpj2YSMN997/+pf0qW+oa65zrhkaO2rWEKq0Rypt/fw1QGk8B0xma9L5daSw/04FR
Psxn5fqW0rjebTSHpMfTNYCFJbD/CaE5mZgHSm7cP7QxGq+LSuJNSw6xTZBcI+/TpGH+qsTuHxnP
EtPQkYBCxjJqrwcMEvkMv/W9z0LS8Hs6F3KYTdpywCgwxst9T0u2VsBIdDjJh2s5j5qSCcf1Y9AH
2o4Z9ocfsuZxygHxr3ha1iI3CqpgbUb2qfoxiaQSBuNZA0SHMJCCEi1HnPROA95Pndm0JENmeci4
5e3i6C4lbD2qcHSnC1Jc5/DoPFkDsDtVHbNp4VZaQzhXVzUCCiStgFYrgQjXTr44ZJ7/f4uIl5f9
0EYh749jmtAiJiHfx0V4b+AxmvhlVYUXOm+6OKgeAEj5hBPTiazU465HjY4hHCJT0D747SeWOks/
B+Vdwy6qfYbnUtGWHU1Ix7SkCbi/kfmIRDZsgnhtNOqkDGKdZGOjhkp2B914g1Tdpo7W2r5rXZ3u
dF+YW6IfKQNC20rSB7r9iwGYOjAlPfAhFKhyfzYHns/p01dHJRrYO+nRI9kjuCWf+SMWLBhSMLuI
23EY8xgUlrIkEPwowinM+XL9vKz9DehCB+8/oKmt3+Hq0u+qJo1af9xS3YeshmbEbzbA/UMP1ujp
lOSANsGZ7qJmOUC6MaaXkN/L+ag8/L4JTmBCzplTBclVuiMApteukU7W1oRPZe0UtK5eImwvsm+/
Pt0MngB8XAbsRpEfSu5CMsZKw54xYhF9zgYEBnIiLetqfZ16HNqxhS9p+7Oz0MhnyonbAVi9rSv6
KhoMFykGGCPjuK0l6WpIPo9GXdHP0ipfoWCFypPeGthIMFSvheN5EZ6HX8t3e01uyzFvl61ZqY4s
QFVpdZ8uHojjh3vUXjZkJY4jbhATTKTmSDdyQgGJT22gbaeNBj6IzUDNYd2sRRZF2VMeuZoSc99+
Nk2TgLRYzGRE7WXYp/t5E8Z0ENcZpG7nrMfa2W+Wr/7gC/HXZGbZJbPY2M6svjBC6TxnkwDfuzPy
OcDVei93yInUVxQfx1gOLTkQN9BO/ZnT9aF5w+k9XTJZqt72x/jZ+2jwQTNhMEtj9jFLxKuJphXx
nAM1lWtQOGAWxYbOXgWkyfxwwqG6932g7Mi9NXeJH4//p0vKBgM111z+SUB5j0qztOWqtSVqj4pL
gL0F/HQjLT/ege5sFF8r913UubHCzW/RKENuAwKePt8vs99fNy9yYhByf+wEmmT8eZ23nvbD8WHZ
DLw1k+7t6oARxE0gdaDra+0dQsmjb8nBH1u0J823ADvUhkEMf14KV/pMuvNdkWVs1/1eVnyRGCeg
pugZYtYcnS+BXm6Nyo/yD9indPXj+LNR6TPiG9VEHWX0A7peWeLxVjPeyeMvQIA/PoFmqzfhT7RP
p0IiCWb8zF6X17YYG7JdLg6RUelQoUngU1DI+YwKM6bcBaQwqdU2ib/6eLWN4bLAPBtP/37TTQXt
lgRZwgSYHU5mPuqWsDf6RfSgPv7La32MrmeWXGi5T3UoP9oIKjWFSoaXSwwldy5EuJPzalTRZptX
r2EnmYobOv8CBv/9sqWeR8pHSqEErXOjbNf8RuohAlApFyTNAUGiGBTksGuwc3kraVImxUxevheh
W7xtMA9H2OZtceC0uka6fi3kneM6H6RqaEe2prdh10svOAQJm5yoomQBe5j9Hl8xjg0MhZx8xmv6
IALmk7dBptaeu3lrQeVsd7/Q5xnhMv1vWnNsqrl6HaHR+10nNpfrVXNiI420slthYGJdffALJ4Xj
faBqjazBp60NIP4sBC/HK72dr30/hNGiYjN4yV0WTnwaLBCchTFFndCgjPZ0ztoVMtllxXQDRXRE
TEZQO4USXzUy8g+KVYJDKiaufrODIAgzz2oDuKhPAslty7A42h/ncJhg1eK+dmLz6haWsCrVZQgE
IzbNZnCTMTf3VS+jFKiw7jpvdtq+QuZd8X4qVagNtHZrZUVUkCic/ZWziLe/YBWFpFojINfOVH1L
KKmURVkDnpaSRJgdKn2k90cIvo8bS0KFyMgzCPK2QSS3769Uvc14OXIAHLhm8dKEFBeb8aES1TML
qB+oI1PJ28HSXgNJaou+Ygf/4H+NkFls9zwKAiQ2TOtpSPtfQqeTYJkoc+ip41ga/Ljk0TuJBD5d
oOwNltsh2dRuLOfFqJbVr/ruaPAMw8+Y2t4adb2YG9w5AutAt46ocsGmmeqV+JSHyFJVS08o1kjY
1IkilPS3pHBPom+pNujsfdgCxSQWAVcb5nGlUALPF5NnCDZDJm+u+p/ZqoWbP+bQkwa+zc8sYKX3
ZTFCFh9/yIvMxIhqEDlOKGR6ArFwnW0Ob8euV16ql8SvQOl9jdv0pSX0QG/XYgQ9Q41pXVf5jgvW
1LrQlIsfk6euHjYZ1KQsNxiM97f2+bX0QEQiB8h+WYFl64TOz8LDfws6lQ0VWNl1xSqRgUfrYEhg
Ek0Dbd6ufIl/kT4Pxp1s7Kb9nXkBgKXqiAB7DY1xGk/hJKiGDj2wY4sPGlGxbE9qYKteysWvIBgU
34yFjx97qZBfS9Pas8nu3yqzD7d3lf7XgJisXhx1Digy5+fSjn8qRcg+t2D7WvBwrcd2Qtlpaq0f
xZTNjsenZXlXEi0XW8tBFIPzVrX8iPVxXAp0Deh+ObNe2IoAa3B1syMYZcmenewz5ucUj8CNl8iS
uhNbnKMOtyAs5D5pJm/FDZenIcE0T+52HpldKogvrZHrwPYS3T0rTo04FQvGb7fT1orfivPrVmDL
pEdO80v20N9KTU78m20OO9skLkiGddhlG8SVqbM5ppPKb8phDrJRIDUVuvxZE+hJR7iQkAab2irx
JpKqBPIgABNdAcFqo48jQj+u0oTJOrpWaWDiYRUR3mr78uVXIAKym70jDCj8K7LQKjzVUfWaR7l1
3TzPZz3qr9keq+dwwTgIFlhcHU447uH0L8yJDV8eDlZIzj7lXQYuK1iSvF6PJPj4q+HYwdAFV6Vx
Y3oHFRFznF0KwgucaZ0tepOxruc5TwdJycReU5jZpkjgvyoJEBvx248BO9liVB0fm3uAC0BLWzjp
DQBPdZLWtWTj+mK42/Fg7IfpAzcw5XR+LSXm/B/jMXQx0WzI5jUB8j+gUdQBCemQKBUp4o2U3MOc
bomNioQkOcRTYbiW8YpSG4TVkNqoO8PJFrokmTA+eY8FHr/aaODiCp7yosFuNEsWixmitBvnmOvf
aQqi/QqZnN9nh2ZzLoHkSSPB3ze6KuJxExakGn8ifJWS5IjN3HCPsagBhm1vr7P0YvJHswJxMhEd
vq8+ditoiTkwXVPl0667RnX1kLYyG9dbfRltQjTM+SULkNjFWHCcL2wSoUKPyZNT09H8mxc3a1O1
KGUtjqezmT72ZbIpCbN8eMbhPpvw7m1OeTQwm68MTQ8hSsbre9UvTS9eFVHlQRFB0QPv7HbqkXN1
z7t4kDyIB/wWdhZ6qtfDvZ+o81NitQpzuH7nELnGsxCE3jF/x7iRztB5OQ9FwBsHrnDZ4uhtHOiZ
9LOcA52huRIlXns94kzNOlDwdq5G2xrjl7kvzI1zOqkqtAu8uZxeP40RNV8R3q+6+ft+AFVJ4zoP
Gb2oDgMeDv0SW7OUJZOEiM1NpeFFjfvVM2tIP9Y49jBiCRfViD7j+DNy6AC4lhdnXuAr9kWPApj5
ymv5kXySxVnCsXjJz9nyBDg/zFu2pXJrrfREfN3jdwXqZ5EuG5AYTmnMygulz6RSvEvoco72VodR
QV2U3QnBQG9fR2rswat+C6rMHDbRHF/YvqCbCd2IrG323aqviwpaHUymJBvYGEZtKfJGiYiVbAwA
+ne8xjfCcA1dJtG5g1KpwH2VUPt0oIXvHqsIWK+hn3qHmEyUplDzBrNizZaqELBJyBGj0ilIc1Vj
8frbZlW8wAjUZSh9jKLshXq+yEQy/gVVkhDZlq9eJCXFX27QP0nLf8Lw43gCwEafYlAN9fJ3KQQx
qSHxF3DdT4x+sRNms7qIQVd2opdG3paQHzaMdq+ZOwvMAw/IQnA/VItagptRIXMaip6ZX/CjE+Yc
kbfc3uVLg2dMEv6211dyRL+p0L7oyKlCF5+z10itIJ/tGP9lQ9DTGsOIIn+0dBEllvOIdNJMoauw
4wzU/BSa/Wmf/qXDM703+IcMB9Tpiw8bjSMXre5ZTDRpyOSIIlynv84L/ZK7mnlARJyMmRe+QPhM
pG1mODCoae9Hdgypt6jA1wv2gIEdtZN9O/4QHiuqnKngD7wgmdREyE99F1n04Up2GIL02D819gvO
Ayn1ctzOnRHxDLmE0mX/tY85e2/RHNg+UpgvcgY+lvOA57I4HEAGJKXYd8iMsn0WsFH7j+6RbVJx
bvENxX6Oi1osuyp+HMdKvDeVuACNxm55lGZZ5/AjnF4vYtQCi/lDNDp6KJejTgh/sSIvXqXDII2p
VWxns80nQhiGAVIODoMPqGpa9ElzSKrxUQ4N30KRdGovWIsLwcrOa7z3TQFgQsVThl124ZGkuI4p
Rr0nIZPHk43iF/Mg3CrG0P7ZXkoj2iP5Cm0FKEdZJU8YFLaNHfSEU0UBofQreswwDUtvDxVWU9ME
rcnJBDB4eZuXbceiYZPYNKv2T8Nb38DJRqh2aZmh6OZcGNpNz+BPfyTJAu7tYxQov1MFrZc0HiK7
Vg/g9AmdWSUXgjGKoswH/goaqHppNcxSGYKARLu1YwMS6Zvv4Ik2/1HnHOGppzaPuHHNvbI5eAXB
e7MOiZNcWWf92bPRFXqIaKgSdpvpX/ivmXL47gUq8eYEqU+5HjsZVPX3wrlU8jsKZ+C15GwIQHuB
SwkjKYu73fFdeaenqksVD3gtNJeKQHSDC2fv6fyALYyxo/UFEOuo+2hgvoi3M02gEqJvwj0OPxMJ
n5qRRpNIstCipDoWJ30GToVeKOEyvd4zUEoaX2rueyTtDjoea6YLZRPC9hU4J7wj778CjWYpWg+v
CpQf8CwQNRGH7fMuLPmiB/79Z236rcO+zy4z1VcU6RrpO8dfd39TeLfJFkCGnwsQf2GridFPK7P5
n2uKKVE/4AoDJdpJKpPl826SLg2vL3WrBsiJC/b2eQP/uBh6zXkwZjVGnZ9Q7rxCp2Syeyhcb4da
8VnvaKu0i3aAXAnIKViSCf0Wgd+qYh3ABq+Iwp+2utHPJVDaHm67AE4o4M//9c7N2FIKWUranpoC
egTjSOGaow2APa+Ut+hxN0xkR7H7NSqer1CUWSLycOQWU62Y0ii6b/23TlOVzxPjOel5X7Mnqqfw
xaY7RZtlRhQl6RiF+2LLWIsK5sys+kbJJ4y9EZZKgWxn0rKz4ooLSyWuOQx9lJoGqgMa5Pyl5ghw
uX8aDIhPI1mDGzcbnQL1uDKwmktp12CLoOs6psHptDZrA0HvxSx6HTwPd1DZdy8BrQuy2t2c5xBi
0wbA7ckbLrQ00up58nkjHGRudIsvEUwaIvsvabEvoOMi+8/Ri38Q9tgiI0Lld0tLAim3yWZwmKd+
G16p6XlUxbX6ybAyRu/+FKkXbxEToZ03fU7VoBICuKjoq6TSlDlm+0iWhqaw1yyasgMCMN97PA2i
tz0eSGmjr+vy4eZm/W3gQ+7qdc7IYbtcphKVfkdiwzPe+sLwK2ik5IkEBVaP+V0TqvTSeUt7Ud55
YmsyzT1/mdnXvbMjKgKICtu3UZD/HhoOlD1QL368ecQSuP1ZpwVFO4UvZzxhxFo2Le0l7z6gidn/
3A4os0FmpLsmewxTjTdoG5cpMnhnznXhisrZh0xmStfJVyY8v9kA6IXvNiBEYdFw3EY+cVDG2dwd
L8UuU7HfrAPDmxMkgT0cR5Bn2M3w4P7OdhDxV2rsWBuFD0F4hx1+CIbNqQ3bNlJ2BY9Rard3zShw
TwZPd/Nb6w5kD/Dj+tx+1mnBZnqgrttbVBsb1IG41KoPPPIG8Jg4btjj02XdNLTOFxicVr8i8kVd
yQICAkqX5qA+Q+EoQZw9BrnyaNUz/rYSvE3zuiJ0imPVL6tBA65d3aGCHy98VAKEnwab8eze6oxn
MYCjb3EqQipf7vzBRZXYSvHhQGz8ACdNsBlhHKFTv3fBFY3c9PjiFD/AuVzt+0Y7Km+YNGSY/i7n
EvDi3j1QN4BwOIY8OHHkciv7SECUP0yC8pRTJt+V9lzyxydPiX079syJ0R0uy8VSnT5i2iYO2BZB
WtOErxkRsX/RZ7pEGTUVHWsVzpayu0QeR5udzEoAQEktZkLQqTW8MGfWPETYf4HtqrqI38VWy/ES
x/lyVHzKJgAgvDwHlk4Ns2N+UBtm+h+JQvZEaH8EqbYntQ3ZeFSC141xeRy1y+WIEn5dtXOFniLB
gJtV7wUF9rNgaHfERJcfl5wGJv2unYmpxqlRG7il8nKbmfQWd3W5hD/sZAnqjJukrnTnaY8AWaQs
GK9hdcjo4fK1QhTkqmBkaDAy84kIVV78EVQ/ikdewfx9izlUvFMSPe/IEpBBlPXSEo8ei5sex9jP
yzJTmtrE0A6ttgiHvye5vUPwylL5SWi/+HxEft2+Va9pdDftDJhsJMFNPMaGnqJQCblIuDUATvJw
V3rD+0dA/PsmQ2P2wy2DMARM/tho3Yddh0oG2MU+R7h2NrccWmSn8yyQkL7xL3HB6g1aJ+Xyax4l
Ku9FtHevSQ5jiFsaILMXj0kIfy7lUsTYN1SS/CCHuT4m8i0PnTrRnntDJ8L9HFV7T/xmkQvo1GXZ
qN/hCkS98+e6e2wZ1NXbCkLrWspIkOYSktUO4VUHTfOQ8wXLEae20XdtfnynQgtpjgfOevDHvLhX
xZ/DD/sd9G92wHRrv51FAJ/8/Sw9aNbChr2IeAWwSdPxj2amBz0ykO2vmiIO4ddEUNCWGAT+6vOb
pZNi8ZlffgCtRYyL2SPUI5mbkl6v9lCBnLYD6ip/YbyoT8OqUgRDWKWBUHZ5O1Y8WAAhrZVDtp4y
8jojUGmE8n1ap5aM1RX3aKV2h44r1gkD5dMkXsiYZrGlur60bgtjfFYnZu/ooCYkrAs6cnJ8/XhO
lMCXySGVd636R65CG348xx5fbheEfgc1S1lRUhZfdgBGlrNRJY3ZSzlbtYeXWU6JbF+n++OkCgRI
5aw5KhgMaCz85SgK181oEExpEjbKqL3zlcHVvUqD+Kio9ZXwgwMSBmfSyg8SAq2YVFe2APIrdFXH
fwSh8c3rbgCOEFzQ7LBKZ2u/MkbBkSE2omM35JB+dcvOJPhLjlZsnvoFLddRnoPBQL17H5ioeweT
J+Q8jTGEbvgqleibFf7KpawxsUv6ZD2I0NV6+Q00DSVSq1EyCSLWv7owS0uDiHSUBK7x5IKOThIL
l6pYevddYjvrgN0leE/TsgoO4RkdXqk4ovFR73bIAnAIVUBpoz7R5/Nls3HMjSim1e/GudxKq4Su
kvxub3opobGLC498iP8/Sf713HcT/szrEXK7gHWcn8oIl+QHoxCZqtkJNG11kcekQgHtwwrrIvd5
7xablpufy0B/CZEGfvBJgM8fsUmlmp9LHq4CN6O+OG/4+s3UGdRe3Z1UHXA8hDsA9MP6zIbG0qRH
Q6P1ZgkuZ8VYXYz4MPk5nDq14E3i7ctj4iu+Vc4SILd5B9tm3HXW7l9S661MjtCmZpDeVcR0s2wK
NonKdbGApAk0cGEClTwbQOAuLMWFUM9jj2PGjo2PFGFdxlJMRBUhp8oHse1LbaYQDhTGHm1y6D6c
/pDgh3acndUjIRnMDUNRnNtljJpkuzFz8hvAmBf286Ft14qDzkVxyr961ARp8ophIYfqY4RV3LKX
GLFavDE23Ei4DMbLYqEyn5emqNBN+hFQXcgOWftBf/YpIuNTuiaN1bbXeC86gm2UdHZDE/MsTUhR
X4PCt6BVyIaUwoPyCs2WU+bJfwbuwjviQrpc9Rq8mtf6QEmUcbXnFWmcoLLuheemehxdopGscjRq
w5aLWiCAFiNBVNFmdKx2VYQlKey9moDLu0Iz00SQGOssbnm3+fQLAh5XPp1UFaOEcIOkpOvDnOF3
KirDxQsaH64dFKiKHTQBYHVXDfWwm/olxymy2ForzWmk4cVR262r4atjlkO1KgVSEY22B/iLK2is
imIl+4Uwo0sI8zJuxYtQiA+dK5YNW5Buv6VUU8wLbDargEMPH/yM9CwNJI09cye3OESHK4kO/7MX
lVKc9mPXB/wiGzGCPm8Iwy8s5WDiLwGYDqF2WbD/KDY5l8a3APJDcQentr2WnHEiQCxtd7fmv0Bq
D2boFsSHi8eLH8wlkHKegtLUiBnk9EBNc2mQZRBrgUm4QfH2C6AjEhEQI6YnTgvW035ZANZeZvB6
CooeDd5LZHwKoMHupJjbs6uQUweg7v/wHXrv1TAmveUzVcs3NWdI7VMw007lKJbvChyq6vrZz/6p
rQDtbyy9s53vlxKdR5JFlHV0Q3G82hX/nsOZ5j1PZqc/If+dyWPSTm9ntEJB6aYuyGpL/xm6kaT+
vxDK/owtls4t4u/XQTqpUj7ZB3RfXnpNjvhZCkFHYNrD8obRDqXecjlLe6xV0+taRpw287mRYHIm
LpfxqXPv50BokNYfT3OWyP1Cxtt7HrJW0PPsikgSTqWuMA7ojtiMdqbeMufPLv6ppJfredPwu4k5
G9Nq8vhibrT7j8DJmlP79uTIlgI0VqjU57D+KasaX8iuEmUyweYZoy26xHB9E3gU5f+ZoQKkZHhD
VSTid6FZkkq75Hy1pclo1wDRNdaFF2GzFYs9HlglXTMZmF2rei5CO5srVDQ8R335ewpyy6957BR4
eWyx2QxQlNZu7BV/E8pyeakX/XaodNc6FaG1DVE5vOjJVbzvSEJPn1xiXLvYll2MKqKUS1pb3Zzb
5WxwVY+YENq5UhiiTfy932cuwoJuLOdYcLZ3q6ixm/gc58+7raxvpmx2oYfQ11xNFPxDTTOU92/v
4w2eW6is9Zv3opy4Ptoxjidd7NlvMFwJuyZcxNVDjF/ESph9ojWZU4v/CIMW/09HnPMu0mCbbpLq
lZH6/eDgZeRelTOL6OPiElqQJVXf2ck8s16rbj35y2O9gRlzUmmjN3WBTQX3slwoPCWcHd5s2Nto
oCiWWsXEhOsJrh88f2f5A8fDclpAJh2Cz3qx9KNN0oW8evoNyO/xb7ztlQ3aoIBjvwUXM212a3cP
iH/ybOxOpfXPMy4lGsXfcaVxsZdOW6R65O9cm2d64PXi8hcypCqphHEgBOr0Vk/Cf8zwTUSzLx2r
Ys0GxlY2VIi8jqoAnWOXNFP4BYTaSEhYt2tfRvcZRApCXbuggR+rKkbmwNkuoa+Rr6EcVBYBAP2/
kP+KdLO1WNQxbyjyCBINnWeEk0SCKkz+0fFmgc5ImV8QmNC6n2ZQtjf7DG1x4rjgsfa1HPmsTxqJ
HjvHIpnqIL4E64fblLGiaafOVWmicsvnBbIL8h8x72URT3uyzHszYdZ92e2L1BqCXHUK8eIdFCE2
UQh2qPtSttMN2uwM6zQhjYlKHr+Lgap3R77lXRtuc+CHvUSJgo1vHssHn/tMKlDU+p8aL76q3Bst
eioU5QCsaQNfprX4qEtO01vp0QxeabR12UAo9xDCkNfw0/6nAKAcbLAp+g6OPlo4shnsvDwDRwOi
59Iy2TL/Q5dDJX0rXW3+ie7UPTF9wZXCwFnm+SbdHR9mSWpAR52FEl677/9sNFHrxU5oaZej69y5
C/5jk5Vnb1c1gdlaFtoBspGdOIRr+L2w5kD1sEhsiZN9zLgH7qjjibb/2XQ8aIJGOTegylceFUJx
HpESnOmitnrid0crbJsy5rhwAk0MRyRY60ww1t5BFJ1I/ol7k8q4T9yuPHJdOqMykX52xzSoi0g9
7z8ItSMA2/b7IdVgmYpKGYK2tOXsprdiYcar84pK7fp0tZ4jMOgjx8B10c6XUtOWHnaQuLfAxl7c
pw4aP9GmXkdBFsjSNl97PI6SLjyerrTyHDgEjpX9vfYYQotZbHKFhgSNU7YYmpGwwzNGJndQkBEj
ceQzTyzvXZQks7KYjIraD5GbTPeQzgpIE7jJxppXYStpti9eQ35zObDGxYMLg2pukSklx9OmpNkM
rbZ+V+N7oAU/hI/GOMrgplP2+NvVchblAcbfIx2LIsDT57a3rVmT6xPvTq6EYxJ5hIwjPQBVdAeU
4j2S5IelzYa+B+xNsu7nzpQ000ddQpPq5DkyP0WolZ+vqEGDRLFBns4qxq8YIamG1zMex2M7SHbj
34UY/Vmu58QSzFKZMuoFX4M9KjJJEA3cWbpafWMs4nqvqzJ9tJxfT/UeoTk7lhE9UoY0R7Bs6iod
efKiwNpxP/WRLIsWyDl/ds/EPDZrUvUitRlWq1jWqZ0l/XtaUfoDg8pyy6mtMMGn4cmHVZNjfAEE
LWuk18BfxqSVCV6V9uIKy9CaQDD0dpLyiiJTWPykkP5PewhVbzc1q7U2GxgoVGkn9R4VrpKky2zI
EBFFdzPzwZoDewCwAIVGMqE0PEEKXK+0Hk97qc3CYZrN8QjCp1rKcnq3vohelN1erBgu1z0btEjC
T3Qpl9RFXry7ocPdT3+sX3Pk5tTi53Wd1YstNHW6QuchqZTSBzAwYU5dhnRQrvot4AORdjuSpSyr
KZrmCS2yqiNYWJNYMbEtXe4anO8kV0XDBeXww6DXscO4SerUM6LeYJCW0SfrF6mCLSBY+Ye9r0nc
eMEOSPWkiQoVahuv2oZwMaC65sWr9v0/wYpItwIgq6YASgAEVgB0cxYwpkvyJqp+MO4ENXbGdyIr
Od0i0q08yzhcKL+ppnHhNhJYew+z+c0AC3SvsokOKWLyMuWliIKZgCbrw3cFShwGUpWDQqB3XJ27
FoM07WR2mIQe1h74IPwViiFNjzczZ0OnAyD8kdsAcxL4t7AWte55+fHdNsS8kFFOtAfuwcwXUqu4
TpBO95UJMMO5kSoD+KxJEiuDH9lcdvJAA3t+UYGOK9zaKU3yL5eHSk5FcbayH3a2E7BTC9krK+Ud
MIdKiRapEIVnsrsZilZRUUu3TOgWOQgNEcdd+r8+SqyvK6MZgI4VIP3dEIthJIAmChrT2hqSOIt3
5oSFpq5Q3honZwvhmE9bNUttjK+JrVTUJdeLD5dRJa3FHrob0wrECRV/9tlfad1MjG9ef6pD4951
seN+Wn20pBqQsJHYEcyqRjSuVdW//znZyLmL1KHokqRpm4gS4mMbTq9jU3hZ7ZopHz0vug+fMhyg
6hsc/QBk/JvUk5vSZPt6PoqgIc/ybcKfG0rh2eRP/K31BGl6zOV4WXx4KOBjWH/x5ViLJid6uGGV
ak3oAmKorP+Sp6nuBSW6U6CvQfmi8AD5JcDstggBGiZcHdN5X98uJGowGXwtw/oHZeE0k/FzyfVE
MNB4eI6E+Xmxwec2IziTuEYu/dknaRERqWi7999ecYCR+HmOSiuK7v6TCdjvs8EN7WEK4s9WAHCw
UKwK2MFwBIbhXRtOt+BKo/c539xaADAIV+2qyt5dPoeQCXexFqRqsGZHRi6vYRExJhOGQTosIXdv
tCJt+zmW03iLAptcydgv5/mgNwJ/k9lLcg523ZFlVjowBSdV+ljJk/Tegael646jKJmf78gGY1gI
yrPhNKvsVvjTNksQU/WBCF9Tpv/028ZeObAgHVTSAktCikEr9jphAxLrROgDxuwRyDnbxSM9dOf4
JAGMrHxVIhNq88mGJpvPhsqwtwWeD+pd1Ri91hfqsfhXb9eJfbHRAp4KecxyTVV4P6LR8fbC6Uyu
UDfx0R/FZZUf+spaa5MKd7qp33QyMCxYrc0Fg+hfWJHofXjSZvHczz2wRvGjbtBXUb4mASs/eN6M
EvJ87idKBKL8FTuhenHTMJD1xFIpMeQQRtT4IWPfw7V2nlJohgdr1UGnAUXarvIz/C0npKTXHuw6
s1eP2lsTUKt8YQCXP4rcKfES4UHXp2ZZdiiosn76sg/S7RcmEOQAmJ9PqH4onivYpAB8eEbvuc54
0HvemCc8p00+EzkVD1GCRIZcdaPVy4byxT2UrVAYukn/ZjZHzeyQ+UvHrcsIfugeZF3FdFHRJNWl
nRLQc/1gGFZG2k/r5BfHKqmqFE2tkyCNHC3GHYJ8UjFuumq1XfvsL5U+7hHeqWM17f31W5RBUF3S
+ohQo2d6OjzlCE7q6pdNjEi0aKKl6NUfdC5t4uABhM0kzIEfknZCdC3dc40GM7zMiDIVc4u6TdJ8
8qER2QIjOS21A0Hsu0j3Uodn9WG/bKHi0jaFzJf1o6pEbLDEMkuj+JsGbQZ7B+Fy/EiX5uotN3if
sV4VVab8cRfuFiVId5qAGCiND9zLLwNhFNxoOWhin4VLNGdlTqTDFnKnVJYPHO+IOKa9xDZgDUjq
c4HpC4hl7DI/SAbNbwjWOWFViaE6S+vbEZloKtTuqidu0WINM06+Sn4Nu83SpCDQp2s+MCg3SNTG
wsCwRtzO6vsYBXT7/cbyXTWOcQKb5/q8wXJZ2D9U/MrDToMtR6OCs1qpWZco12LKkvKCaMQu+WAx
kTEhW/LjcOX1nhk+lxEqXCzeDA89HKluct9TDGoLdw68d3JvarXBPVVqY9D2WaMMnvyiY0B3nvAe
7/LyOfDTdd+6rNZyDHZORUezau/IDwEdaTCm08otqJQh/bNFNWpUMrDGIk3eA30mFP9MVNPwEGN9
UCg0/Isba0OqayZlBYGm5lvaF4hVeA+1uYluYP3MXz52rXZcVxM7DPZlPpAOgL/AXB0RKq3a/3KG
Ag5CfM081Ix7IREyRMGaFuuxZdstO6m656HCPz0yErM8+BvDgYi1kcnPXxq9M5Oy5ZJCVBGHKemQ
vtZCYGOlOxkwjGODMnsKHC2+UmxTKAER/YNeo0lowDS6U56m+mHKddwKpbIgD/E2PWROa1mQ/HF2
ZIwb/A0rdq1pjYYFVVkfFy8YgA8puVClN0y3LmGvaSIU4Etr0D1F7P4oXKeeYUMl35+Ap3maG3Fu
1DToYTgvtdKfQO//RCZuaIXbC2dFIh0aeTgISH/KZgs9IgPhiCoLTZgnn+u3mNChjJcu9EVgMMNu
Wo6IPemJYze+JVwPPzHSb1OaVkgMYu4FinrzFGQL2nHFTCnYI0l/CpbIv3YCdJJ70llareyfK2zG
eMljnrdmMoLXvneqfPcYdpp+z7WWtEK7LfLZpj0PwkcsG971Du0IoygBZsDCKoKY7TfmQjRONiPD
1ISKz5nRDX4kANstvoKgyF3wu7TW6cZznnpLrfsH7N4SbaMomjMgETDVpvd2q8uxv0vs+EMPE773
4gcQiN9Ot/f5m3cNgjMkQ2UtvbOmGVmnD7DcA5OLYgQXgUYMJA2TqA1j+Ctvr5nkVyLV2KTIe+n+
ENSmtONmBLcAa6oLE+Cp74Fz61t/D0+N77Rj7oDt6epgxeY1D4ps+5mGjouQ2xgYasiT1gT/KvzG
NXuGWBav/MuTuWQvefx8EgHkuszF7Pq2V5OpQJNuYlQTfzRKhGbDF4QnPpQnQ2X0hGdx8b7WBTEg
yUOgmmrd7pdLQb5pxa4lumOG13upYKmbM+9tmUHwqUPrtqc8jqDgE30W9yJR5ZXgA+bx4e0uXvMw
BRhwPEJYz4obiCtc956xtWidzvxVfWFwrBIs8Zfjn20uSMzSNWGk3jwrVfbEIQcDGdl9f4YYNl8r
WQMOLo8vyWF7vydIGDoAxGhnr4Krr3WwLGvfnXJQvRw1tU+4Mx0os04A1G8RdPMsmPy4MvMfTBMh
PqoAaSidvvwOywze8xPtUYAgCQ6tyNIXLxEc7ey+zmxNIeP9YTpJZ68mybhxIRVrG0uPaH8heAi1
L+pQuZOnXEM8i4soNstea81bI0ZijKG7f+nCvcQEmCc+/zj3ozuhDE6Xaxgnh1+NsXp14umKCFUw
lT38Ys9kDMslqHCQ+XStYdOv+eZk1KpfVM9UX7wHU3o9j69beuh3zgSpK0v+Ol6CmdDODvfJDMTG
c9g9PSlB9Fg0x61gxR6LGqHs/fxm4aEudndu47p4BkUXV5D5qr4rGmHU7Lq/0rmxdJxfmkuzHJLj
+4p8xv/zcKSQdXmUOSGLX27phTpEQeUo/oxmLmo4T6uP+4zLCXjXg9Y83PQOT/s7vmPPh4o6BU92
O7Ab6PP0eeibYFp6LOUFQtv5hMIpxhn12ZlXxhbhrvbA0U47LcsgMhqpi8sfPH23OaPtfJahUkUc
0L5N/beVKllOdaccjEGtypCR6SSV281gdBGNs75RKzsnChg73PRabLJ+gJ2BLp362y70GXnKrUly
BrK4IVvMS5VeMDxHTw+SWhXWVqB+dyUZ4CLkBapw7kxMu3A9U5EhePUa0hCkXLetRZDKSdlOEWzp
GQrUjdiRmZ4oO/6slK1pc1z3P9HP+EOD+QekfujP+4a5Ok/PCUvpUgjcMut+ZBq8NY8BbhqYLNLX
MIz5m/E/+ZfW6zJMhKBl2KrzHgC6yf6vI28ovt1z/FnVx87iGFD5nYL6TCOvoQGTioqj4wH+eaFg
pZChkWMnZ8E4kc0xTQf0e4dLfbdCz+XT/IQzwc62hnCRACL8kU0J5F84g21MUpHIkoWKoQn813Yb
WrNTVfrVyfaKSC8x1wjz2hDe42mSYJ5G0/M6BcX5oM9lF0M0LKy746zC3PCNC5TxNk7jKQTZmat8
cZom7Gt/pGO//vgrp2g29M7zKaa2vhlHhNtq0tkYbMDgEK7JTeSdcncsLLJAOXsSfcHWXdSyrfwM
GaRZL4gUWEZvNwhxdeJzIAGXPQteEqmgxVwCKflWwEh1FJnqaLE3zk7EWNGb88vMEJQA0GR1bhJb
+7qGuhDR6Ot0PyBUDRGgNxe+PzRrvJGdP12yn6u8CTQ7FiUwLEQlQ5civXU4OMUL8h4ClVgDfFom
8dHL2yfySpp4T2JoviydHkzGP7d0BdCxZqkHtMJhAPUk+Eyh64R6Y6ufbhWiZHXXb7Pwc5lW1f48
IVTP7AsTUd4maFE0rQoIHffQ4A2+Bg3hF4e4OJKISj1Lr3u6QnFK9GtvZwN6fAJNPpZLNrB50YT6
qVfTPifwgMPwWSYXt0IsUzU64Idmpz7FZ3M68u0LIWe7G/HrVnfkLVMDwnoIVVXV1iZIrjTs0xK4
EvXHUti1l/KyNeeqMIugrL2WgAaK4erml28vMzCPvtHkU0rUOarT8CXwNedkTr2uzrWMASUm8t20
7lbIWTBSkb49fM68eBC2KNURWMw2mJaH0fVYArMTyBWKeBJ12Gopaq2ykoKy4HHN6LynMhyivJS+
RN/15cBTWWDk+U6BrDawyS4MW2KigDlgt4Bv29mMfK+sEEWCH9JmqTQLBGsrQzfJ5WzQFTHxyStE
7RSJ6b9kv0i1cF6Pzm/1u8PqOw+UDPAR7DGuPM+nROA3RNePlun+cwjoFnez/VXl85KFhabzN5YB
oOOlC8Rrve3XwEuqAqXIVqUNki3gXMQiPQ3fbnpmLSqxD4NwhzOnE9ynwLCPExaUTmr2+FsUHtlR
ebAtUcBdJW0wrXpJpJZ7C2uBGvCDbv9/JB3+X8nFw3iQ9wOBAw5WM2c0mcFxQGHqs5t/7Xdpq+yL
TM0TuBH+1CTfexOBwTG0Er96b0HoH6GgEQplvJiZcyaVdRHDno+0bZ2JSYt2zBJUQwwYd9TjKOm3
LjPNTKzndoBS6d/6vDaxzTODIaqqGUs5y8GcmOxWktz+wvE3n/Q8OZs5PELhtMQMoRyEz1Qt5Uxc
Kq8arV+nKlmixHxDVJP0x3axoOOXDKHz3cvvxnOvpQP+eCfJg5mRiub7+3wUZnXhD23OA+D4/OMd
EGJuv1YYV47tCZ0HZFjXUpz4lz+Vmo8zra1V0RHu4+ngBVSFpNhge+kB2Y2mIg8Hbd6YMQwCzs/j
9eChoX5kLcJZR627FFBcvgf/KKJzWvTqq9RabWnanZDJZe/EnB8DSlWQwE9UPtHp9F8bk1j3OCw2
4A08OotOyl+dgGndvwj3c+GDdtFCX6iVCWucWoOuofWNMThLT3HEnhVU1S0AxyIDzNXI8MyKxMzS
ZzHX4q3mpAO09NF+wuBSizK1cSh1EILwTbYa3ZgrkJSXiGkSapeXSqoNyKqewVZFiv9Zo4C3qyYX
Tk6RhTOx1tmyR14INxfm6cyhzogzNQXnDFZT7JyT6B/Kn/mBYREuy/f80vjwACjQYB/F3am0eXZd
vCUJHTq7b2FSvrron3qgxtQLkqLytp0JlTPeSkmWPyTkqvCU4saTCFhF0+Aa1pJvpiYoBiN4jrU/
ad1ebONGO67NZ/igyBSArDovS8/ajzHsPG+yv0sOCVvzCQ9bpelS7alKkkq1HhljYdB2XpjD1pmV
LsyZR7ePHidAP0Y/1Y5IL+2y6wt2LyfN2mW3r+eR8mmbkHXAdckPhRDBs41y3pynX+aIAgmxG00q
G1GEzEwjIvptgcVd4JUB3Hm/1QK7Z3xoPZ374y8u7ZBald5gW6tMeTcvGPa+adoKMY3zYDnttEy2
3rQj32eJQ9kFJS5YEET/hi1cSLIEWJTjkfPN1jmwJRap4WFnxgSFhPC/c8gOm8u3h384S+NVLP7A
l6MdhNnijGHnbz3/kcevy4baacPNV2UZ/+aIRDrUogFEmn4RuhXsJ1+bn//nJ7OZga0wqoyLenft
ApbmG62BuiyhsZBjqltXdUfg8c8Q/XsEJ4I21qQ+OMx5coQuxAHootg/iHIBHbYY9PN+EmHLU7MK
H/4x4bYvygiXFmPLV+rJ2L1ZQkEabegKyhGa5XyK5GmHxk0AG5ph8Q8tNr3qYdKwQC0m7kJAQ5mi
GPHgxZobz/d/IYvNduzAPsse3fKP+mn2WEDwY4EcIzS7oAFVoPD+ygWGSl2WxmczBjfZQo6p75Rk
VbaSiAfuIEA0wbw4cYFYL8BN/27PGuan8g3/JdkK4enQhjBwB3SHnU8NO6nEcS1H9unFkp+PA876
vR2LxMALxziSWySkuxaXw3v8aBxzCU28OT/OOa8RGbD0MzksFR6D/12pSItuIQ3+WRNsOi2FkJOp
iNAfnCqly6Sjeqv0IduzzcbnsFaSDKya7wvTdHPFSR8eoa4WFML6PtU/pq5Pr5G0SaEvpE2cLHEN
HPJ314FMqLTwY5e560SjnrYLDi5dJ1Qbpv3ZA5Iw1/060YpMYBd5za0unLe+1oy/sNoriKHOw9QL
DJdz3aov/YIlvmGWALQtj1nhqfsjwTl1k2NJY1PyAEIu0vo2sbKjDNt9E5FAizRZzuqd/qEqflmI
BE1oCqFZC0XlFwb96eR9AmIypFwwUPBtLkNR20YmQxDZKqnXULpF+fAfy+MJ/PPv2toIIXjVuE1X
XqQAie76WsedpDpB8iMOaL2TQTz/oM0j1rZTPhDYde240BI4/qnUkq4lABt+hRICbBBrbuzjkeAi
PcEJD3Yx1ugvvfguxNVAq2tH9o7nq2cddQ9gwj836vlXcBM9MjuNwiupRBh+aH6J/KQ6xG3HqaNF
L2kA/4ZFelEIi4zDuc7QR4rNiJVpJkFNd1Wy9TcJNoRCEMAVDUo7FEu30MV48m18V6V2owXkXfSp
wmLTBsooWx6H2q9nKvXsKdLO6Y9lf/7okOK5ELMk69m14XH9g/tmAHKUMHCObBxFhv3a702lIner
aaSX43OOyab9R4bTNpbRfdHB80MquTPDEH1UIVaeasAhd4NRFAigELzPYPIPbliFevuWgxRGHaDH
+wxjXrILFMKRSywdzTsoKuPtFy3rnDLxfQ6KvNrcpg74/8hEDe1dMSnKELrfbxHVHcvN/jA1NPWp
ozkOplj+X4vG9nbKi5bzDWl4NUtKYTUMko2FVj4fwtp4zb4o4b5Tm8vRcoU13ZjEZa7boiHc3bc5
F5CVJdfePbjhA0EUPlYFCkJGNTj2Bnlg2CQ101mzV3EPzRW8nw1GlhLWPRf4HoH+fQuIUMpKvGNB
mv2tgshUJARwvi6seR8CKxnUX4aawsVgLCuRIUKecRtjdcTegXQAhQ0nDzFtdpjYikcvXmVyCWZK
312GzLWgYh6+6oHU+l1DmTbxSqNxOckvVLNLfGVSy5B7L7znW18XtSaebw11m0bMERq2nQ7Z3dpG
6x20I0JpDAGVqjiy9HydjDj5L0LfaYSyNTYAsakuNTQQUQY6UKaw+C8bMEHwCXaCQjgdSca1Ly2z
QngtyjOiG6TTn3NiMKQTYmcwGuuF/y3aAv7OnxTu7nEUT9nw4KsXWMuQSA0/UHLsJKfDSQZYCagf
4tB1GyC41U5q5KSAPjp1l4gn5ds2i/XYV4wcXIzTKfIxntvYWFGB+UnsXgsfsJHbrScaJgH5i1pH
VUddt0oH4YN/RrVFLuyii1Sb4fFc+XYEMFJFq6AexviHEAAcdgM9IXTEn+q328U4N1iMtEz1IdzW
Fvcg22vUTO0U+6/21UsBcq+OnYLglFo0uch9aNbCZWOLvxH622RGTdFtwYNCsUxy4gn2y2iJhzcw
QJJyqafgoQz/M+rhErA4PqFQOgZiWXuI3yd3AnWzwTsUY2tKJW7ojYcfGRDgbxSXRoDqvIqnSgFJ
Jh/3nH3EshT5QLIHdQhNUI73Zn24xdKac1V3hVwV6yjgj9EuLhDTP7yuzfUqmltHeVBJI+HfgiOF
EEX91pfGLFL4z5LyXMKk2v42WbbDgIV2ZbiuimbX2/HJm047yoCxa0MegbUDKeukljJr3joWwHlQ
g8xl2aU4ToJYT0vIBLdQ5QF4ukP6IjMjaaN2gXUS8A8x5sE/meA77i6IhUWxR+8Hag2UlnPu4J0u
vYWAPbx7rxbzUmCRHPzGNoLFDbYIBq/4Sp/YEOk2wJ9rDLPZxElK6dnJe1u3dMfmnblpCrVXNcf9
vkAJqntK5AlrhHL1sspeNtNoWX3lowyjYl8cx4g6Tc+WHIMJOoYQiZnts94c+Pek+W37Xr0AHPym
bzfjPRCNkR/HhaNATZzodMO1whkxP21uMnRMfL79rdJlZXJtX/j9/KYzwlmYWqXhLrwmmdZ5rgUD
HvBHHDg4NaybePAGgDmOvYZ6IG1YtUoysPl3KqLs9pLLH+4nt4JjI8eWP7gTAk9Fo0NWFjoNxPcj
BB42OKJzfTRcLDOyfnKVGviEf3/Yzvc54J6DFpcvw2ZHKfnFsI7kNuKdH/TSYUFgzD2WzpiBZzzo
nH4hp+BbxVIcCo1IfczB6Gl3uBm4PocJEMvKvkA7en7anRBagDo7f+wJPmBJBQXopmIrkoZ1wurs
aG1kpL4K2x0BbQM7WZx4Zw+sVroa6HMvu7aN/yPVLOqs18tFVGtqPMkE/SywaY9BF8u1kjXg1QfG
JvvB+pmpNe0rGXN2ZG9xhdMi/e5FjBuNAlLkVUwdz8tJIzslBPkBxPno0UT4ZHiqwzq2IbKAKZoz
2kbbdG6uuWnGLxJhRqqqSZUxRKrj7xqKZdfx4DSpdl38bVwCLd8ch9IMXZIqgwH+9Tadw+B2WTBo
Uz5nSJt5Ft9CDSolYA567DwFUQaV8WaFeytY5aTGkB16y3JBoMwoA5n7UqYx4gQ7aC9HM8lTTi+6
rMcWzY5TtXrvdvatyAhYB3TC7xOuIz5GJt3tCX64YTxoWTXopKhJ3GqoNF4f9LwX9xyKmNmC17kg
sZRX5iTDNk2xcJrpGoZEWvFZHTCJZcTURmtRWORh5suDpM6ktNwfVNnayg44z9dLWU6Vrne9ba/X
QOD2ZHd8P+G9hyF0lCkSQOhrrC1jva73CJKGUYuwGHs+ofy1FqL2BSf2ejIiGwp7qmclOMtvm2FS
72BpOpsEyOoA8BBWbLHI30/WiUJLDi8PSGnyKpoU7fkCmPIxUZnfX9L2mtqJnRdokMKejyMpxbuQ
EMWj3ZTXaOydxXBweAnLWj7BcjlkMCbkvk2pQRg1tGz0ZuQQfm1awMOraUkrwEpLaS2wyirC0q0v
ZWvwodP1x2IcW9m0dGOpJiW1boCYGc3kt/w/Rg7w8lKwm6N37rCBjFJ2guhN3TljaVBSUGIxZQpx
KSMCB/GscE8VcFBDaEJgp2qTiweYxiJ0SVAlWGSCH8ZAJr1nnE4GmDVqpCK2UddXW2Tky24cnsGe
N4t5q0x2GxKn0h/2lCeTdU4P7dyUyaqVpdiKS0HP2+Crubu9jd6OcjWD18/PEoWuzFoGoTAn0aoV
qwI67en9PQCvUqR/zb4MY6gtXcENS/c+o2tBYqlxrHBERi34Kghdb760mDrOOjOShA+JJXmaJ6gK
AY8Haa4E61Qo6MRFLl+Upk+OQADtkY+Fa696Z7dy47bW1aMh7HMzIUtQYBO8228eVpDbQhDA6ydu
0mMlJV8ExQoEHawgoaWOXyrqkgup1MfDWAK5jPdW3KPhALQSQHv7KrBUBIsxDqZLWqHM88UfNl3X
irapxKILiQXYWGOcjLGQtFW7Uzo5qQau/0J080tYTPqlI59L/cT9hiR3PfCuqG80dY7uJhe8TDMy
Abz0HRmJWlrlImQzQTX8YjEz6gNL8+yeIshJhW9vyRT9GV7qr2oTeG1+SExBVeIDeIyVPKBio/bt
TKHB496xEu9vJMmvM7PslOfRHMLV38jKHM8l5TBYi1HObNKvpu4K8ENmbbcmH3yypa+3DNtpZ0am
x3XZJgqUTsuQ75BIrzl242NGBbXrvPpLjtRL1hvUvZL0TF2sAOid8cLpWkiOEbRx/piETu/R7SZT
oBZY+SrcEuvCx2ML1ZUAHPeASl0dNKG4hfTcW6HKtXnBAmevX2rXgLMy26KXzG8pF+nHrKvBRf7Z
79psVK6Y3UabBlk2SKq+4AkVYZdYc4xTPHNl9enaOSM4WnCriwLL99FKeUnVO5LgNwlc5NiIVM66
nXJPG+akVFk/vIW4tsKVZrMCa13o2mWuYf3Yu/X765dEYqcMPo6iZz6U/dQmnItB7z1mMtlQOWuD
EXKCM45rAsFdZShNG9YgumdLVXqJy52CQe4jhK/bjBz3fmj1Oie1hMPGjRaxtwbrmPBSZVAHSK11
Jo12PffVII7pgIrpoHN0EmzR8jWU018eiS7YAc90D9lYHqN/vZFCh1/jeW+3Z00FtnCGL26vDFNL
LWohf3+YlKya3C7j2rKe0BudgzdieYmA2OEOKXoVdH3hJvObeEIzv3mb+OcB34DcaHhzz6CGnMDD
5Pz+b8gGoHyS2+mEakMyGwpb+rKUL6m5JvhNlIaQStXAZ1H4LV4E069cWJ0mayvc1SV4krrmezAL
6ty8P35V2ZqM3grr9OoxZaQf/sexZ8jt2adLPf8QJktHKArQXoXIf9Z1f4LEmKJ/r5+viRiRuuio
o9EPNFo1o6zMhcLh9+Unfc59MK7GI1W2VYYHWHN8FesSrAWEoBe6UsdO9+/rXh1gibPw8NN5bRDi
ONCqlo9zQKgJHmIxPY3asTZ6T1/W+a+ZYkD8uzx50i9BJQTaVb6E8to3vxiOiA11NCOhNuILi8FZ
PiHnWC42PGzGlMU4OfMfLYIMWgIDUdbK3t3MF5UzJSLDyvoq2g5lGc++D0mZZ+9lyXAYEPsCKQI3
0rO+PMcEVNo/g4+wkjsHUm2iuTDxPBbJzdPqF9Xe3rDekufGKIhbNkGqOQxiEs5qdHeVqRJJqo1A
b1X8Afdsr5XkLPz6TaDBlrHUPW0+i7nvbl/clusaiIo8xPj4Dzz5qwOY3kMEhyHvCDJE3+31qpXc
efxLSXEf/+LfwY1TZ6pE6fre5WNZn9fTt24GWRMeacx0jJXEeKzoe5iDLAg/igQx3toGcKc7JM2c
YqGgLuae0L2YpnDOrXLKluCSzpAxavr0RzY1YS+pveRa6cfMSMIovAbJ5KW1AlgY/2+7WxnFwaLm
beZsGHAq+2FlzCYbAJ1g4XDvu58aQbNEhTYpAwEFhUX7eZgthR2pYdDLlQGXmiCJB1PyjlBYRtzO
/pyEm4nEe/qCI6pxunUtAuYkHN5AZ1u5CH8ClAtdHrLErVmKKT3DZt0wdw+vUzJSrdT2X0XqfMAu
wQCxAgR6SwVKJIy3leHafK20GN4Ys4zFBbt7JlZbRcvLcbJvSkfAeTcMoCyOKb4a00IH858woVO3
YkrSjBbuT7HLxJhDfSa3CFdgQSwYijfKtOmbaTvbbtXfXYmYQXoTXbRZFB1gXfVoUYAc2vuQHHSD
G+RRRliNIqLDRFmWt6r1resJaXQKoNYZqzs9rvhNQle8YDa7WHJZRyvXgCeB9JhUts8KPTNc2uoP
facRGMIfy+24E7Rf88D3SKwWj4YOAhpLwSnBpU3Evb6O6ZvbQZIPSJxTjfckzibz/BiFGBJL1J/k
zu7iOGw3JMpsEiHf1gfVy3Pp5ZNk87lBbBkI9MlXwFbMaXX/e875gsSFQJI29abuIx3m+c2x+fN2
JHrsFsBLSZg2eFazoSKPQ/rWa6BDy7T5de/FNEHm74ujT9rwGg55AZE5oNwPkFkjMboPqnnia7Ek
lDtcaSXNAVNk1dxhGlc80UvtVkXJl6EEP8DeuGK7UYzfSrOWmPGq2XDOSoxJkVUzeE2YHkk59EqZ
VDo6s8RO27d5lSCqTlsjbiavO+cpkS/JbFlxixHxyIig02iwDtmfFvIzEcgu6zi4tPTs5p+TWs0J
2Eaj5MgO+8J8rYEWIBrppzM6/nhsbz6uyNPr79BbycPVoqZ3xp6NQ4sOT4WqXpDcOp2J0xCNz/1I
SIrIFdf0deCBcW+YlwE1P61qG/oTS1QHZWme+vJcmoIR5jnc3v3mws9FN3bjGRLJCwMqQDp/rc54
Kp4cNfq+Zt+HdCSXrZM7LP2gJb8VH4NMfkWSGhyJmxAQ07mxDfbc3Bkuzfxp1Xi67Wbv8XO1S1jC
nkvVOr2YBr50mCPtoFU/q8qusjpvU+waZc+xiWiUkyb1KObK5piGkEOmdY/ChgD4DsTJvewH8Q/L
2m5GFS1G8thKtyt6kK/w2aCNhfPToinjcQ+NCzTjm61Z8HdyOVgVqFjuVV7W9KFB4BLXH7Mo+Iix
+bFgJpeH6zJTnqa0FQpeB7MH7kgJh/V79cEmvezqBciiyIfrVCK5Tl0HeOQpDzwW2dya+7JUJhtk
moLph5vvcdJDYQP8S6vZyXQCUG+uOpguC8+6iaVmOkm3k9bVhnTm0tbvk4DGMtcUv1NdnS4TWzLA
OFRUMUG0PUUf8utTnZkyvHagEbRC5GB3MyKFOdcAKMZ1IE79s46sHuJwqu29Y8B//BC/1UxqnUfE
snham/LOZQyvAhFZWLpTDtqCIhuLIqxSxNsUUxMu+eRk+Obt3Cd8w3kTWXBKkAcRaXYnjACskxED
WUKpRmmjrks7H1Xu07/BxzVOQzjeISl6kKgeG6ZD77bn/GKuttn2B/Z4AQTrsppjbucc+HvuGopH
zPvoMhhsyjREVa2e8eN8LgBDkubXhO5hA7VQ8YtyJp7K4b3pzIlnrybgRs+x3YBAhXxcC4+0j6at
UuLFFeqlnJPpavOW+HWPlR0YDOxGveePGABwTRdIQX7YOAr7snOReQe489T6iVGK9nW7Q4uHE7fi
klE7nCJeOOQ+PnuDZOvjBx9HakYSoMfFCMzoJu2bdGYSN5YkjhS1XkMWGQcQHLQpdb1V1UdIjbly
WcLJjkmMCOBzyR/AhBVGUR2RuEnjEgVGRZ6R4K6imbnO0K/xLfa3pRP3zoyVZg4fMqshbpuPbzkb
S3s4oEpmZKjN4CYyM+KqW4YTgMqs22Vm7UkkOBeVfQCKfEeqpLjySOeKc3nhBgW24Ly7bjLJ2Bae
vrcVnZZtXyHiZXxDGK5Em1/0DcxoPMXoXDRh7pckkjGcgZQrPuL5Ke2RcagajZwBbbhgt6kIBqIe
aAAJRpNvxkkjki0tMMJSE6wZFZoG4IWNuBa837h0B+iVyfNkT8kRpJNtcJJBvnlN7oGJgoSfEmC5
rE2Xu1UFcXnNXIDJYa7GLlrOeTLFCetR8JctbZXjLhWDFI7aPDUy5jIk+jKDmMwo+rnHAZNH5Hg/
zkEb3HHWqT9sdo93Nw1rNawIAWJGsaWx3L8Os62bqAiqORsAuGqX/xOEDFO27Xipo0E3VvYntLjm
Y3R3Ch1TfUIUXX4wFZ4Fcfwln7ohtWoi2cu6CgwzYPPCuVWs2hr4O1a0bMjT06iV3Bpke7xIxgfj
/rRl3iWOana5OYSILlCXDS+XRH9K/NMq8HgJfiPylom1gHJcbzZKZTY97DLsa3jFMrThmWad2vC7
q5GRXe5SuDM9BmQUMiDxOH1Iyd2etJ40JP+vjxDMDhO+N9AzPOPhi56USs0x8QlrHMdP11Fsi3nn
Oe1SUV3yj6pQ4sN+FR7NDm2n8vlUZXm86kzEsnhhWbGdLrGs83T94pOYoDc4wBtf5DJIq3SCDaTZ
hpEwJwpJGuu5Kht5yO8vu156bCJ5aoIP8Xj6nRLyxCsvO7NhiUau3opeUbOkxDeGxLlIAdDUzllT
wfkDtPe95p9OrlRxQNTV7DUVjPSq1cTrOla2DmCme78WAcokFO5IlFM2SidIOtjpDykUfm4Y+JLr
NLb9g6gY/tCqOo9lmRSOom7r6HY1zPk1DLVqya3UlNuXnHNN/iXD97OtmjUN3GRfcS4yB7af+p1l
eWpkNAqEKrlQ/UVDNiwltKPbHm5S7+Nx6YP5aDBKF8qIKaX/2QY5WefGnM+4E1IYNIaVdWA6rdzU
+i12xR7x9JiXsA3qWDy0ElGX36eK/zJ3jW8ZtHzg9lZYotKQDYCWsyu/uwMSNCM0gJcImGIkS5ZN
QD6LSsBmqm+blM8dQAphtLoMUVHflHWxbkbso4r4Nf6+iD7Lw9CjRRpQSYNcxzK7oF20OxZUufIp
uqXj4Zd3yn91HAWglUoUdasSIsVfXg5r1K2LUkhwGroW2yzTYqphDEc6+bahDI9Hlo2qWehD9I/L
IzdKzdZJTzJtstAnPYm6UtLgVafXFPHKqMq1WIDG843pnuvxt7rulhCjM6hxEaEYOTia2f1OmpDg
HtxTGwa71qag3FyVQ8I4b2bMT8EjHojT/dz3j6SDWIuwf2pZjsteHq0cPQ2JMMMvT54IhRdUwciD
gJSUdwlvHWesITc416MT3gIm2Bj4uE8BJF3INEMKW9NxhYUkzHp3tM86TYH8k22UMdnzD06cQD1W
LUWKec8hTewhvj2/mkisTQBKDX7VTRnTRx3IFOTQM9bWWE3hFl041eM2mPo9nnhHiUVHEHnF1MYf
0jw/Y409E2Fc4v/HA5vhOXeNgs1mpww8a9532sHUEPiynMGLSq1T4QHeuTuaa0kgDnljJ6sn6ZEX
mM0K/01aM0LFO/SlXuTBcWBigtBu9WBIMZr5LCUjepW3WIy8t0V2wS0gRcupMvs1vm5x9pBgv3mF
s5pfltBOXHP7lLz3ZJz2fa4nfLqu4EQq5HG0EnXyDEeOSCRf455WHyKuomT57GfE3qyrOgWu7Uwb
U4PlSHMGcOM+2t1wI9LKs/RKlwXwz3eYyyWYewhiU8CpH4omx/7TinpAfMn8N6aGb9kWMWA0DHGc
61KAX0nqOskeIT2s01wAkZTdPaKX0Nb9OvjxtTS8h1ZJ22bUWgP2RcJKlSAwbz2slfpyKZNHlPnX
Gfr77xqP5Vl4I0gagtUrWkXnC2OOF3b7CWuZAvbYHnDCPjacfgp+Uc3jd3r8bx2kGylmxC3qclxE
8R50RBz6Vaen5vbTmGV4g+E97rloBSExMlUvImIQ6eOBVAiCbsUA69rneyiLqD2l8Yfprgfy081e
t02w1BMqryJwmXa7o7A08FBMsipD5SPqyBsqIP3YG0V0BkpknkWHb5GO7mJQMfqPlvgSNDvsV7HM
Lu80gswJnSUjnASfrzU5Bk/J3b7uqCGjdZv/FyXJGsuADE8rLGkQc4Q4ZkZDspSiAxyih3DUUErn
7kzNOKA+7SqszkI4ttU/GUGHz3z+AhRHdKnTCUKJpMr1TXmMX3cdOx7wVfMHk0nY1xu6rFRUjddy
36Eh+ImDRztVeA3kJ1jhUPkoVq8eynvL5K7mTls6Xr0dQUo0e1TWMpB2+Kfe3/QPxqdCZ7fievh6
9lQ+rZSJkoQ8q8vcP8FwvCj8cL+GZAkvUqiMw/hc7DhWBR639Xe6gKl2OFU1p9pz7AJ0C0f5I+Y/
3c0LFE5FYq3y8Uz39599VHRiccL/snJOgnfHBdujZdPAlrcFPE6toFj18k4ZlSwSG0Pl4yxxHWEn
mEZmG8WZqmZc/Oi/7M828gowWMvOzdh/jmE/oa/YEW8GqXdESsFHohq1AzU6kQb8fltEX2bKgu/E
RtLHWn51loeX5nA8XBd8W3Gw6GCn2C+8I1FhhIEbP9TrEQpcRkuC50oKPGSydaV4r267RJJhGk0+
chPuFXQVOGzh15Ut4bHj+zqG5+C64+Lb8PzpPymKKQI4XIVfINvCgOEJLhUl8FZa1yDP8OUX8Hbw
4VCU0uT4y051ZyJAfxiLkj1PKixE7S9bKjYgtn0s2okG4x5P5dpfVkVctzAX97n5ZA3cO8Sc3NJC
3Tb2W5HsH0KmLttGyY10GbFY4PVcHgu4TZfbZzWdZAzaeJm2e1jpszjOgICVA9GaeMu/2IOz+wBs
zuUvWtEKGHns48T9XsrBsiPj5la/173YMToAcelLbxkwFCXdQQLM9Tkh6eqCZPivkcDPw4bRZNr0
3Bx01A9gjGybN+2fApsX9lYHmmQs+FpYd9ulCJL5yidg2U1A4+i0IypDKWX/qiyrDKCiPnDmzHUI
OJdu1e8GjKBPGODAZqHn00s/4ixuhtyLZM05moL2TQ7qsiFXknSxdKNbMUF7kw374jOAjhclKesX
0lrZWXVx44a8blIdlnZzCwddXRcRCuI96N6ba3P54ZP4mLmJVD05sVluhFDDjbAlVeeA9UgG5CjB
xWJC3aDq3xdexh15js+LRDWbhrfsjLMxBODMf8tSKNh5IbrOpitQzzDvHPm3F7h7oxueww3Tx9ZY
X5PtMRmCFlbx365Pwqa4Wj321LDFIe/cZj3iFmP3iHcUBuUxznBRNhwo3lXd4AK0F01MHlyoUwkF
ZtAXXhalUW3/4dkdwJhw+9go6DOvXBSeNgMkL1ScOkFxdeOnrT2D1f1unNsv3FC63OG/vtXllFK6
EzNmSFjk+xgbB4X36fjzbkX0OrAGIppv7eBIp9yP4opeB7dcw/DMCebMcfikvhwDpyphXjdYrPCp
hCPshxQPBIlXjSyz1FQibasVlZ3cciIEwGfzv12wQ/QMdMGdg+W9PppvdaaROLRPlBy/fxSzHeYh
GX40qGU/VILjlraT+0bdp2JGroClT+jRjMoHZXYe8OxFG24qSfy2RQWHtbzckd8TkdXywByXT+nB
E37U9o4qlu9lVej64JNvN4gWWhNk7PcJ9nj5JowisJBvRzCJSAG5QiIW8uM/p17DqIjhItq3PWj3
0K05sqW69dhAjwIcjQIH5PxroFCmGY2qGZcYaCsQgPWZ0TWcXMmVVABS/0zC2lYgXJkLCmXFBWxc
OXAo7GGkrgtT9Yc9HzBiEJfi8Xf4sTKsmIfMd7KMXkBefMVOQGBMbeODfpMFtsRnb6y6qXI3q7ux
6bXNCglX9BIzcRj5m4p4WLZ6GqFnPI682I7Z4IsKT4rs9FfXB2mtAb1L2PKrA90d9Uw5bCxfMR1Y
0Fz8Dky2HPKpeR1EN1Vij7NPCFBWjpiz+cymK4cjdw13fLhyVgYgiejmZWo3gVjww9lrkpAFFIRZ
vGE281KdfJfCdTfmYZbkaXnQjrAp77LoFyZ7ZW50q0W4MKbr6cmm+dBXuRVvZig+Ku4+nBFX5/lg
o3mAaWaI+D8XlSJjam41QHXapZu7AVSOniTJaw8XhVqGXxCdGRX2cInYWkkrO6q77efNfD7yDblr
j3aTOkedFHydItem4zfUZFD689KrDZ/RmQohSH4eYUNXsGSNmb9Cyfp1SD21wWl29s8Qf7uHbfco
SQrYerVXQBV4YYt15qf+/+8KLkcKHoyY5A+2PAJGYk4BxrRTvdL1eYabhOoUqbVZKzkx5PxXy0LZ
LaQswGona70nHTf42z0oYSVw6Pm/73Sb/bfcmCLj3I873HnCsomcj/eupoG8idyQn7IU900I8AK3
VpavXF9PTtVe1nETZHnJ+oQu1wQTSUV815bQe2gS56hUWyG4l0SE1luUisBkvfYKxmCg6V1sDHSN
rJ3h5zc7ZNmvxTMcUQ5OwPYamHnYBKL3Q529/wis6joQPP896Q1V66gtYWJWk1vhGFtjkcJmZXoH
X8f4fCJszKZOBTRkQ3JSLIwu3BOg8Q7hfSkrXz3T84UwRTUOr8bVS9BoM4MMDcW4VzAXPbevA+T9
kPQNl8Qh6qItnRBP70D3gThDqcmZ9Mu9FLotmhJoiSn9bDNoeuYZBjX3/wPA/RPGf2WuEsIuGfw6
t1D64hIvakEU5dYpfj8oMmzir3x3sxvIIOn9DoyOEjoH381HjTlljPPgdeQdHY5bIwKfhnhhzrMQ
yi4D9qeXBd5Xc462OaXx1CivRrSOfm2wSBIt6s7q27xxh0ifqNjHEZKuRzxoSGXoMCwSD7wiLel9
74kYBi0JmHt+Raw0jXIrOjdLmxYTK54hAUMKBv0HSRsIo0VrKs1qDxRYpNqO59DPR7PS0eIhASnG
8MEARdI1+kdTseiyUN7QXV0u1EIcBaGmNUQr3RMFPYkWZDJMENA4TT2+2q6n6JeWj+95QBMqeE31
Y6D+GGwbJj894F9APTtINmfd/upeHPWYL43JGR5ls9SUOIvJcoJefupUXIScGzsF2DECikjYmckq
zI3IZ2z0+Nx19ojbuCAftiQYJQSos5xE6nDaIzlWZQMDwnGA6RiTBIm5ygQt5RqeMQzOOfmidy13
lhuTf3WKM0GYuHaHU7A7fQt97h33EnZRZBY/KYU2JLOWNOWvk24y/zFAdXvRuAzMdjjva6kjOma4
EWjO9Yw+wsv4jG1KUskr7TKsDGbQhWxUoPKzitlIath/ntUZti2c5mPqpZeWBiGiWObdvYh4MxsE
aiSAibLyk1Zl6cr5NSEFv1XkJxg6GKmC1CZ7iiRE/a75GCUeYlum/2Q4iSrpswBeDldykqnQNFVe
q46bQksVLsdSwL+gggWT6FY2Vyn+2QfMV0HHmvvqHlVflaidQu8xtdQsmI8TGh48I+n9XY88zGet
KDABJJ2HmskMXwubx5A61LYUXIF9Prp3kvlPo4j8uwSmR1gyMPoWZiTlb0LVFRjw77hfeupchg8Z
5V0sQHHx+ddgFJBM9yN0/9Rq1zqfvPgi5r7Jv/eHNPsa6HS2FMcAj34TmMBiBH82jIrwak219M+M
LeXmHbmE1TsLOjjZ+PikFpwbFhrWi8wjuGIV9DvlcukSuyEMryjoKM5JHWBBo9gZ7+7rv36iVJOI
AJB3eIb0smAZ5L5ayUUNL8MnbYGSyvhBI/RfLznOM2M5WYCZKE/i3hVvikNwGhjHrg9fRSw26K3b
D1l7EGuVtVhB6/U+iHeZcpI2/x+S7/f8Ch7hBKHeVQGGYJLRK12it/mUM3NHK0Ann7e4xQrZBrwO
F+NbeQlWtimLwHqZGdBlDyKXvudDXF17wF/5chwECpodYizL6d7M5MAScwgtHgs8vod6lPeJUYP6
SCwXYoQNGFk1fiyFyzT8RaYT2ntQlzm1ar0ENR9rLl9QTBEf9ketEHf3yqE1XfeTYWIiL5THISor
2FM9xCEsH/dB9TAAXA9174KrwD+r8KtI1rvyOe8D48FwnRXcFJGh5+3etITlnw4YbpS5YpqlCyVu
aZEdHssCxI6jfDOnoSUBLpP8o3brigr2V6d7lQZHweZmMGlRWcsQvrZxjhw4Uh3x3jZKe5tOeG5o
tpwX/zS3MVVrUM+iOtok6JrOEYZdv3EkKs7cBlDBrA7GDuIhoh38l3Waf5W0R9QqDi1mFbY8z325
/1nF/6dPs5EOpmFAkNIK5Fc+UzXofj+XitHlewJUczq/v3aDn2bSjArQom9Mbo4o542pxSoKKRr/
dGi0uhMwYl35EDgQ+/1VHCtD21joCsnFPpa5yphjv1OFBIJzPE57ecUpKb5OSyH3tzgUA4wmMjiy
4MY9v8XSdqmAKysn9WSYSdfmMB4IpPyvGK5aP3RmHhDfBe3+5OY8DJHc80BCYVFlgSwd314rNmw7
Y0iUIcxFODd5nUTVg7PITC3pwz4VsiBjlqpCo5ZfwSB+TGubkLV/8BYmAuDmJiqmsyCYm90Pgfcn
U94l5+iWs2Fv5BPtvEgaZYRmyX65CNTWyCFEXX6tGz4Uu7O/D052dfaU5mOnaWRps/JyCrnyrcA/
ymei/Rrj44LIinqopfufYJY4aBEqYztZzbDi+GHQA5DS8kb50XxxQpMfj70L6nz3z668+UrTNPQ7
gI1503oVS24gn3Am4DuFC5pcFzGa3jS9k1rT6bUUUgTJnTOqrjDk/e2/VSBcwWpsM40d2BPlOaEe
SmdVtpnvOBsQeLgjf0us55hx1DZm5Eck0yJka4CgthnB+e4ls5qy/a5ZHstxdgrhltNP0BPkovPX
GrvbTYHq7xR0xGWupbVtttze6DQweITfFyy0qrAynDHDZbquBBNbqXvGL1k/GZghrZ6onk4Ow8Mc
E/M3wuhnKGnuzZ3lzVuNGpmmDptIi4Vg5lfTRgVSn1M0GsdU4JqksGrPZREJiLKLXg0C/wqiY+sr
Gu8nluMdxiLcL9XEicrSE+LtDN6fWXF2+A7JZrQKNeIEI8QQgg4NN0Fdcny72sUEzZ81uI2FBzTV
W1emLzFcxtRbvCH7ok3ou7qUTv/Kh4F8lxnT1wnE3Z99l92Fh2q65LRkZYiN5HdwL2s1IbDdT77m
k3OnxD9tI/cPKbXu8EBphzr6P6cPn0L4tw3kOkc+TAkimEPCjR4kYRxrWJhOG338YpjgdfqRDAbn
xAqLO5kq9MpPUj64oI4qoGJPjEqngmwY1WZUSfvBqaqm59IFICNhEnKarFqXBVZ4JlCMY6J35bLa
eS5gk7DPkwQOO3b4tDiJ2uiZMUbDL+gxnRsOqTcOy5DIsZ7Pjh3C+mQQGzdNlXZqv1kK5eIhJ80/
f4sMDcBUh1GTx90k13oy3JvHXFVLeoM32AUAevlo3ExNbk7jQeC/HhigjQqJnE51tvsfddmU8GMN
Owc8f3NQEI2GEwkGj/l/s7fLeQmOOQINp7Lm2GcreFgR7G3Dvvl+VMuT6cfPRg1nbMC8NwMsLaih
sDHi3IZOKY/eTWhr127BlE29tMM0GRYoJOo7sHmeyuDDNGlHXBvMObrb7tLmtcfVfNPbdS4FX96q
tVt6ERZf1eEiIZfQ5UO18J4vP033hSz+h0gabpBFfucun9n+XFoL2zIioM2XzQQmHZSXjl4B+9KN
lhkS/A/U1KfCG8PIsB5O4A4mwoXE+H8bhYmZz4p3xdQORgd+fvHZu/GlQmVlI9cPKLkBAyfsyfty
LpKn1k7zDinsOsNHmLOjcKbEPCFhG6A4z10svMcwT1JCG1C2CfsqnEK7mA8hRztaWMhVV2EjKQsN
J8zEj9d2/QxUcbC7CtvW+diVdS1s2f74FSDgYB1kKdRU21ELlNc6MV7s/1Qlz5LaipTWQf5R+EBF
bc5s6TJXYRJSidWTGUxptkKqWctKPp2RX+nDR97xfbtzd3tU+1XeTCiWUsfifRKO7gm4uEqBacG6
mRR9+bYu8dyW9pkA02tp1X3UOlyGBuXvOB0y7yceitoV7j/wbbwDPu9vjeXpH68ngIJx82G0jj3L
XMqaV++hazFMdHK88CZRZdPB/ULChhJCsTiW2ovQ6WwDvbs8l4DhL0ITyVnVzeFfLSUNUCarAOuo
60L444V/TAZK4X4QABk63mH4qoK3HWVYZHlRyi9diIww3ckw2Sd7UZ8mgezb6RaIvcjlLLYfnuqR
C/PuoG4TF7VbqBa4BJF0M5B+wUzj7JL9k1QX5kCl+nYLlBKZSzx+rldnMp3hWpxIXFZqBenPLT3k
PmKWaCjB1z5BYxuHylO5NYq/QGIPss5BAjZnisncJGKZLehCTsHqyWFpFlJVo3/O34SFVuWaG1KX
yjAxr0xT35iHMqbtFkOfb3/PRSrfFkq/kK1OWyhm+HL0klGLBigbYybAHbgyUS6ftZYt0ZoX5fiT
5n22heDWCqiXhj2fv0HvENrfnouT5c81iV+9KYYzaHkXi/P0o9Whtgt5KHeNIko9+OQWrTN1LW+H
KeDIAGWz8Dw6zsq1bJyRPfIwZtssMENXtilmtWeIStnb/Nyk5eWgKP0mYmUPVEP4FqB19Uv0Kh8j
/PoSbtbGiv5X9x8rzZ529bTdjuGYWNqQ/3xI2Zgk1ag9MaGdcS4ooFk1dagQDcqM+Tacoju6qXab
bA+sfvb11fAgcgNMTTg8aDeeLh1LTgqYkK2AgF2jysSTmK8/q22dQMMqYdhaoEpGjVeglUOC080t
oGWcKTKK+WPEkGfGkNZiTultOv/jpRhpBaAXSQzQBsvyeN1eq1xZ02JEDhHtwwoJDr2vFYDVUxKU
qOZsverxm+j2t9uM2WE1oTDAeVEDlCBdyRZfiG1EqmYaxUBQCJPcQaqHQbEPg3gV91irS4LrnXVa
eJ+5EiuLzYfWKVpHiRZhR4SKJ+pdLkFMkhYDU8/B2T2FP3rYaqdQexuWa7FW9dL8yTHZxDiiiUdF
VexhsZ+9wkkfQdNGxBDPwhXP8tAMHTiDM3DwsVxDu944x2X3pFNa72HytIewc6fchRAMODwvlsYO
wwA6slH2YseQa4VewvdvKfegSg94hUtQ63s6EElBsXBpsep62mV2ndRgfMCbQe6/vVOxa+s22JBN
j8VPckyiqtsne/kpckMuivJFCb1QPjxLqHOGkb7Gce1y37joP7L0seRoZl52JEvetjoO9NZAbCvQ
iP62MDw3GgfDkWSViiH5tUyr+ZLb1JkMniuE0mZ/FHXxZNV2Y0CVog4H7FnvLf27ZqbAKeyR2yLA
Zi8YmrCxNfw6/lEHKv/rK8K3uixQiqB/m//DNz3TelByOyxaSQHCJVeZdseNnKoZHPphna5OvDNW
WXM6cX95/KaOtzx2Gycuzi/V97C6BABUerkgWrb7iFSoKlQCwefvegDC+ZFeoRKtYURJEjdN3td2
8F3HhSjv7V5ZrlSmgHK7YDfzCbfsFpJQArm8/fTsCc3wf4ztJyttXpx4gvXBRl5Wy2lMFAR4jj1+
KiYoh4m5Rbnrli2R61EY5ieNM+oEIofu5Kuk/xmxWDF0XnqEnCp5NXTKRHLFoamUbDeUwfKiTcZw
0LdeGOJpbMNqunZn4+FWKiYW0ob1yGAhAhAwUUSRbR6OYgPmLh59i3mDs/lm4l5rgrr3nKwJlr1p
NobFkXXSe0UAoURJRNma+ibEn/f/QZJCCb0CYcFBbWCJlyCYNL30rr04nox0ZMe4k5TRAUStMlIS
NSIYV9mh59vHH769TboQu+8Sq67avDX/PurpYpuEu4OT+Hu1AQySrV+EZce0gYTk7C0Wakn0ctLL
l2hSJnNZsmsj03K3JdMgiGI9XLet+I0aE5qWhy8objlcaKhlB7AmawS11A8hE9hgp7KZdozejYOX
4MaYePRYBv9jj8TRHo0eWt2z70TMj8upJtZZAL6Fa34lKNZXCdWPxbXnQ+H8cCbi4dXCSAiM7/Wf
Jxdo24ULu9IH6evnIt9m8uZw4Dk3/7LKSbt8fOLqnMADhWK8bxxnbRW/Kor3qRAv5lhdfJoHoJXU
5KL7QB8NoRy49zWx7VfjdPAmpVFF6EnHGb0SPBr1cN8/pBCLCHNZcjIWQhu70CjK1cxlvTWhr4+c
G1aoWuSiGNE9BlZ6QDwiZTvJOoA1g6gzFEYyF3Fy/zALeCiy3wvF6sF+x8FlX7uHSvOYMtPCPlHK
HPQ/Fsse1fuiDY1jF9YMvsMKtKfCZ0PbKybUc23VdCUm9CpY4NS1qONpTUHcskx5oX84VyzgDien
mW9hHBoGajAeeJYFn9i+SoLP7G3sTJ/0M2z2RHvJOzuAfvJUZRzl7tqSWm8kR+3+v6CxMqpd+UGS
HFXzdcz8gEauhX4L1CHqxmKO+lQkWoXGknhLYr1vlCIAwkMx9WIanhYOFsmr4/deXwVe12kCTC4H
z1pB1W2ndwemzRRHFq9j6DCDqdAq+gFTfyhYWemZM4OuDiRwp9cQpayK0ASjej59xxBdqpRmG1ae
vteVdT39wlyRLg0CAfE3tSR11dBUeCUJnOEasuR2/07ROh/fW2Tp0uRLnibcU+3fglr9SPAFKuY3
GS9j3+eVYE+zo8SeK2mQEdXxrF5/E5hMw9Slup8Zh+F+CLKbpSdPIVk+9Ukmadty1R+kAPBho5iP
3bDeIF0clCq0P94q9vqfy1ZCD3nc1hMaKvEJNAEgIO1HSExFLgjYGbDeMpPU9gPCiaHW7VteHMrj
POXqJQHNjsFPdrB3yF02PxgXvattWa3M+rWIiGPNKQ7ufbckIq1luLDLV/gqRF+uubyFpQoqA/2+
6WXklP8DUM/6KR7z5omKeTd5n0REJuGHgFMDJ+caBmstkfBhNiHGXHaXXMCaftCq9rYLnffTSm47
ErYM0JWr7OKggSIoZ3Fo21Vx5ogrgnh9qvD/YHmYf8iqvN04Zx1lj0XcxSlmPjyD/0duPRCbPVMR
AX4HBRpF3mHm6W1kTGyWNoHFL3/WGlICFEkGvlCOWvt0FCCZA2ZyU6I4zi5U48x8jtCPRmzjDMqX
D9MaWgynR84KQX5ZSemqgBlWg5Hm8OVM2ivT5rRlRxl/3S5vYYGVnH4uJLGrKw6vxlbmAYu0PC/p
ML7wnyoMsOWtiLuM1snnjjCeczWJL+FsOTFhLy/ps/SkLpvIBbLCK90DD17GoKx6KM/PID9Fy3xS
8wA9G8zM5BkhU4BeBUUkq3E6nDsazPfstxL+xBspk+AG1kr51ctarOLzCXsCIMpCThBkk4ugRSFb
PtnueX9ZL+Eoh9vDNOrUIRObid8QeA3nPBx9qaYADNIluPrZPk9HK4QYVpun0kS/4cmCRQVMUKRK
1YB3LIQAH2Wg8+qoZ5dS0AboH7/uebp0DXK3OarWeQNoQpDat/BzcrdjlRLo4hv2GCbuTShBMeOU
hd1q4JXUh2+cFHrW6MP1xyHZKWDiRzSRQUn7ACqWomA9QfOPKX7mptf/74w+FfXH4TE4dTbIM4zV
EiwlzsY9kOPEgIOGzVPE+XMHnoaDc25ANUSBnztBNHOU+ZHi0L9CMdRBvsG32OVLBLAZztOspEmG
uDf5s14VM5d4eHI2G8KwmeRv4JY3jyM7DS56icWwYvcDgAzUHv/BcJ3+e5IIpE74L4PRg16ZLQpn
XVR3nXX8IM7G99ZdRwZym6gr9Vh3DWh8utxgiCeHh1Lv3QvzFDspVo+jMXph0dcFGwWPsjUXK4o1
eOyUF1OORjUW2V1yEh81Rl5oZhupdzOES/6ees9iYUvOGt77z+SVD15jnBDmAewRChtY/3tE6Fwp
cu8VhF6cF7UleAz8Bg9rpW99Mj/KhA2hvmTz7isuLd8cUMDzXNCM7fmDPS/l4byYhRKS58ToLgW9
YtLSn/YSg7D6jU0M2Z05Co9a8PvPu7f0MPlgMlFwa50ZfnibSOEd8/IbtbNA6EcfmQdqkuuvb5uD
c5PN3sUyfvlLIRZ3R3+r4E9/BRZetDdT9aX89B1HydKwLiHa2W2/ItIGT2r/8b5xfvAlU2c/uvc1
QYAmtMn5iYUsM0+JCcOyKYFTbwq7sOQX15MqOlmSNk+voGJg2ujFlaPxgcGLQmh/0dOCkJ7sYk4k
6690mtBkIqyGpmOWyaSEPWh5B8uFk+KP5elqH2mIZAU71X3VlxwG4JO5Rr0ps5hxO0KSnjuLphs1
m6kK3gv7hXvxCPTvjVwDCUTu3PwWltusiSRa6cJ5oHUA/emicD+Z+2bjFRd9mfYNZ1XtrVsM4WjP
0HTxCzfvEiavogjKsoogI9OwSseGrGkdP/8ejixClt3pPOLOfAOgLy6RTv7vSM/NBKDoDUuxI68A
crYkPkfcFaoJRMEv8nwxLfemygsKyn07uN1t3XSN/UqBUmgsGkXbKTKxDUHiNgcN7+PAcDInlUMr
eL3hRDL1uQts/O10MMWIE8KYoZu72GvEI3b8VYMAzxrJ5hPjhUZvcjieMt+qnE3KPUPslqkJbAvc
jPAXOL7ur+F1tFezEETqz1AKXx8ktHTHsFf6cIZnQhLwsy4cobYDQfkpvFYgTevsVDlXFPUBHbXu
1EUyxolgVQtoqPstTSY7ncSS5H/N1nXECLP5KLLxUFFjnrYbXjZyUbG9CzVtNm1rBYGDloHFBCe9
0YblqTwYiYGV7VvO3IZ0Xju5Ug0Ze2u5zcF1mmdgmtYSWxr7BoFXnum0UDU+13kr4L1+QCoOdUmY
xZLRe4Lryjjeo9haafFp2DBpKEbDbbm8PPA2dLCs5JyK9bruTJRUY+u4v1x2QTtvug1ilNGMrQu2
zUG2Kxvyh8AcTL3Q3AnGFIVgkXJsiWF0tW69r5v9e8tGufcMDPVQUoKUypPxDY8+e2QgSD2xjU1U
Vpn5pBkZCGm1ooY5Hjd+e0IiSCDON404NBVv+ceGYb0RZohsI+tnmZv834RzJ646jUPCt+uzWBNt
+klg/50XR4STzaDvgBICxTJ0OyhXTjKC8fsUXFMwE21bjLVim47UElNwWbdIc6BPiJLDQwLMOlUD
zHgLrJ5cVsqBEIFzhlT97Xukzt+K7DMX8z0aUudo8IyU0YdpGKXfQAfPNnOoVm5ameBJPVrPYTnZ
rQFbVtlY59s+LXlJrSuuWAgoagbq6ubyxHfZFCTbilsghftA4RDi3AnH1UJMA3Svai+0gimBYVKJ
6OIxTZ/vR5zsiYtKRbISA+qHmadiqyOFYFk+jKl9HqbL4JGHKAKtUN94SInuN3s01fsop05MO9YW
j21xl2KjDsOIfi+s0DJurhro4yWFw7+mCdyAKUUFPDN8ZzPJzH99HRXMf4YVgP2znPelRpO2iTWT
RKgwscQ87U/71fpqR5x4Xfje+MgmD1VudwqZUnwNGjdvcNtqkV6/aFuQalePYfh92rasw9Rb2L38
a374xf2kM2Svc4eNGopQy77nZv6akgTPD+op8KTfivjyYhBF8Cm4k3S0Lg0bd36ihhhCRE9Dxz58
r5Gkh23GNtwXOwYFDFNRSIz1D13xpDCRAbMKfD9N5qA/R3v72JYGDf49Ibs8PD/6JemH9vjYR1Un
VdzBFsTqs3cHiQ3QLIjJJtxVNxWiOZ5IAcUuG8LPAuqYUUTvjc0TuCPe2Y9CYcIJgEHebvOLFP+z
ZTuEdwVdk6wNSQAgsahK0shjTzjJ5rupNxc9gh2D0ImDYaPlL5p/36NeQ+JgSlyTvoLEtM8zLTL9
3kfQAYVahOccJyyR+yPBtdByTb6SWYEwdpkC2kiqfZ/QeL9EgcUhVpHUkh1sPK7rmsNqbTmCPedd
m7/Q34/XVHwamtHKMt8+rhyjx42Y9wd3RCoDcDR2pg7sbIyWCiJ9zgTLTIb90LEZpTr0CHFYlmnP
QSqdWt15LUmSYKx6US95qa+EcU7nQAbN5TbBfzhRDe122iJqViOOXPTIjsz6GHLpHBuj8lcyhC5T
Cyd1O50EWTcOGD1HDsFzdn5YTicgEsnlGrr5gWbpiyFCoclmZl9ZhFbOYRqkr0/gEqvdeRWe5rHV
HA0DNcaGrgObuq+VKEOYMIve3Jdkhg3wsREWxj19EbhXfG3bfL13t9u/4MGy2h0wnkFSL9zEy38W
7d59IP/sc1Uj/mxU/l4qVNS2mYQ6stMxrxK1etT1GqGS037G/rAtCYIz+DYiud0Moaubk3XDfkuU
KtJC+VduN2FHPpMtsnP480fwvCFNduh6juYA9fE1ugXACBjT5feMNjmgVdgSM0YAe+ZMaVjwixgt
T/UOxCogxcSBGNuPSivO7AtGrsNeeiB5Sar74Kk1FeQs+pwZb1lEbSraeJnanMCOg4uQjrSGuuln
GZh+hvGtAkm/z09T2/XDemNNr637O5c5OdTKNL9AnWmuE5FzjfZ1XUWlsTApqnJIvM6/K/HmvlNu
qGEnCRNB0r6fKEpozzYON1duED15lZROPYdh6xpex14tNAhQUI7WlyyKt1ETXD6JVDlSiNOoT54S
4/Y727SSHqYPBCGxVPF09J+QA8EqUBY7NETsh45sdJZCNpBkCjSQrG9v3ty1zWBmJUAS4vbnp3ex
GEjeUeRy+ZaYQqU+jY8iPLsc/xfFspvC5TgPHbF62tgXVeETRi4JwuHrQK77FB1U66JRt7Y7dqNC
IvrZk5SpLlNppNrhFhm7+kMJNEJAnGpga8kUUXHZKkA/JKPp19Qo3mvBJS6o8aUY4CrNuXgWdayv
Rnvepb/jSw4F+bx3no4updJ3mF8IEUYaqVhNS/7AN5+JAAWzSlm+V5/9/yxY3WuGQHlTZLc5VhKL
WnuaYoaAZ/UV9RZaLDFDaECXAJ2kmxBz30jitkNpLzW5V9sxPWurlhYfhpPCQQ5DTM9qZ50a+fZY
295gtnzDYkp+YtpdqyCYHhLNEJabn1m0KlP5mGhDkTG5DqEuEvYtYnUqmQqSkNpIBMExIkXBD1v1
u17DmhiKQErnNnFVKcU20BHdcznx36OHcMRKiwa2WJBuoHfYSN+pmmgBFw1zchEs7SoYyyeVBJEH
nipeU/GXLNdPbf5cEauNEU+KYknEMRqR+XcuIqWyBFgLQZd6r5kb2ovjVNMFg/Pn//xk0EIa9h/i
u0LYDE3oVTNVqzEPspb9SAiHybxet6i6UyNfWcENu56OyLPf/2nD85/N0bCBH7lpnhuX5GYDEE5U
YFNNaKQmeYmJQ2/fxNSBvhFXB2nfS1fuOhBYPPTPwB3qYnr0Q8Wntq0BErChuINkvDuruF2HVvDu
H7KIS50pPQUDUHw6metXbij8eyhU5o3Si8ShjK4yhoVGdx98/KkA1iQotvz/hlxycGaXk7ARWOYM
sFxGA1/9Uxe6Bdjm6CWXzfnGb4TpEvX9XmjbMwStR12TiW1fYHjm8Ag4r6e7WB6niHdzOc7GMaNZ
uKXlk8kthZDI9E53/s8gIn2ztvFP4Eno/tr+6CdvNd9qkro1x1CwQSOo6P3mv99F1cHdX2iFxruI
NAHtm4JnJAGAGbKvvII87ersdWb+4uvye9/P8B4hnQjyFNzkvI4pyQTPRst00/dy011jGhoOgtS1
NzKE6w3RPpQOeBIemoadRJ8nu9o652/KhIpSettGF4NPO3RaNCk6C8v9owe1Ru9o08Nlv+yuijLb
5P7C7XHXAxQmIHLbYh/K18oMUbXp/wpdLKqP9uBS21khyZ2dwQQaQlU0L5MJ5N2fVBdj/oFfqNXI
YvwfX30wQ6Pz+XSd7fg4PhshaXSMS2s+gzVvuYOIMX4XUsiXUXemH9qS6ry+dPSyHDOiEmZqUs9L
xbw9Mu4mPH5CZ5epwyym9h+kaACgtZB0kS1xtcJ3tZQ4IKuFZAOULYjmPxEM0uvORFikN3iCOXk3
kEQdrMoVwbmgol3q7lX0tjZWzPfm7ZbBUxOUbfM1Ha6tXkW8dUNJROmBy/Vp46MwAxJvA4+gJlOT
ondxgbbwY+I0WOheIj/Z9vwrVluxfdy/Bqe9sLuRV/qVVMoAatx5ETo7PFPoxszTfppMEGlStjwS
mzeB8p2pkE7vu5xhVH7Eey4W/aztp6reoNG6GnGzqFTR1w/pIK3el3w11zG76QsarhuFFKq/Nwep
G9SRGWXXPiCUVpEZ/0/Ba0d2JTj00fFa9tqE94yDlcgRBN85vHWQ5QQsJ927DWt/8b2KOaOchEId
gnGJSYG58pyyAQ+WaolqQdPWfn2HVhm+iO+T1EOjP3ZFdgeueaCAcLL8GeX049EMCxCU3lWoQnwA
nxsggv3G4GG0rF7OnJeivmJbS2Wzy7NA6x4d3HD/8dXaSBskf79aIZLviSPReykIHmzSNsShu1AJ
e7r1ksgyFZRDo4B76dRHpNztH7jGKhZbpz+KmlxbtgpZnmQsGcnmtHIrv90AzEwT3Y6UqRpZycnW
s6cOG2hsxdLsbUunjkimX4DVa227Tu0+ynFSvraF98MNuS8rlzo4Vi0UO1a9r7UbEwGZgc/WhdmA
A+mpm5BT0HN66FxqsuLWU4hPc82eqo9isHySHINWPi5O46V0o+cQG4ugzRIBuYdJJOZ5p7iJ9DRU
f+SW6ASVpTs+jq8njlfUV5A+jWYJNo5hrFDCv6v3OWh9yVbohCmuaHhDdq7wrzaLE8REhGKMLFfh
YP95wu0O1VAG4xeMbSQ+hywhpNSppexCPvIKr+jNRgCOPB4VaEKLMYac03p2pwNxR/PRUhAhykML
Nnddhmx136SkICZ+JJNP20Kh7RtimEKLEj7kmxgfMFgJKTzDd0NtOETU4EcV/qVjNwJURhXH9dxw
xmzenO7dtgHIhC+uFdnc1EDObaFA5nABOSapKn/j9HAc8RIzmDhbDvjUNxSVLtQRRvRoR9X5+3T4
Pa4M7zVOwoYdxzgl1pTj0keRfqt8tq+BhRaEJKnxInFUISMJgfNfLjp0NhzEKL/90jxIF+bDGHnK
uiXxSi15znyyXfUcOcEJtplKcoZhrsM8JAtPGlERIjnJYBab9eXSuPSs4VGijepj37OPP8PkgkwA
A+UbY80pDwxqryZv+qjsn/gLd/v42opUxwFhTfO3DzTZGlEauCjDmZJzaUhpyxiU4FJAMOfL25PE
NLqjgWjPHsCVKij/aMABAy54DrCfhyVqMIJA3aRDquyFm3XLajPNd1tgAwM0JCM5TapVWng2x9sJ
gXKHgYlBYXjhIkCTX7UlmsneWSvdmqoGLLGvyaHqf/q5yYng+3dEW/IV2neUtIt+DOKqm3zSIyXU
JIDFUr+9np02f4dU71S1CyAd9TIfz47skgqx8SckO/TY96oQVogHB/TgXQCH3M0+ShLlQNCbNXJi
JjVhea53x84jkHmHb0rRw5T9Bui1lIA1hTWGPcmEYvbIMAiOHZoR9VRpW6Fzso0oXy+q3du+F1EF
yR7/gJf8lgEFvo7nY2l9sdi+Acp93q176zsNJuHY8v9bMuUGANCSd+PeE6dA9+gNW6GEhW2IDCaH
+Mf86ZMEiKfJP3/e2A5Huqw5hMMVgQB4+7P8Gi5XJNPY5SYiApfXUn8lvKdFHSbOi4z4awBU8pBY
jKJtLYoNmMcSsTCMbR9Wx/qc6SK9Y4zkeDRCmgugtsFlH3D738rZemCA1wQ+Kj6v1qRqS5TRhsja
C/LA6Bex6BBxviVcBIiQaEzES4DdUzSIQcdk4/Zb3eLDh7tQwAFQbLvFXEoVgUGh6axfSU6YGbNB
lS+u+ksFior+HhwDtXyX4klnBCnzWWCl23B+szWu25cOtf5QiySQPhx9myuRdiwrDmwXcPoJKJ4q
zKXZemhXtINyh4gZQP/7lb1OYWuWLaOrB1RGwlmnCbvyUfP5i1MbYnpzgfj02/QO6Xfbyn53kuni
ydtvOKcQu2cP0Iy4h2Y1vmqSlsX1Y34lp3iusvTd7FqwIru3jiTXV+24YxmFVcdRbX7D8vz12P1x
PCHqeGdcVpFpIHFlqi115TZMyeBmeYoDFQhoSRB6xT+C2yqXALTUVNU29s5QcEIWllXH3QGy3a/n
mO75aSWDKsw5uuR3TeGE6y3mMzuU4PN+rORrbbmpqvXkLGlSsVc7vVUrcb1tGFTJ/oYTuepk3AJS
3fw3Mr8uawMVZxmjsvYeh4qaZzdcd22aTee+G/50nhAsjeXhlW8a4WxrF7gMVNjWrfZckpTaVYQ/
1+eEgR80Gc0lUlIVxpZEeETwKQI0DdYbmpkRFNBdAZ9zNGINWeHW/jbgNiul46QnP3F5gXYPZ1Yc
iQYBpkS5MBWMfT0h+vG7Wfx8fKnER3SxnG6AXGJwNzn07pvP9Etqt24Ex3I4lw4W3u10VpjJHKua
ge6mSKVpvOy7qXv3rl30QLyPWbM3YNsHlTSAvGKQtzMgCI1BU8iFe/3+BxYg5pulm3lmDH74ZAXu
tAlQfLvmiX1wuBhjmD3VUdluzY6VIeCNXHhAScAks7fkSqpSHzIVJYIkPOJczGoN3YDlYKOUQLDA
g9QCEohuC5IBmnOq/G5ScMvDAIxKnFYUpEk8qqHZs5FNgL+zj5sUnWbx1KB4GhLfRZoZKQ8dplwW
auclO3h84UaKgW5cfzE2bHIzT501ObQzNmETJNMoL+ttcMMApkcQRyMqpNhPgbjb1/JtVj4ubtwD
ENxc8Dd5o1Cq+QwSocsLXCE66CrfmW88Iutkt5BJsINc/PeR4k17075S43PSeutLcv9zAF5aUycK
gsjtyg3PGqn0qmXyghGn60xXdHVIpGtBE6p1zJ1fu3LqZXUwm+fNZdNseb2Cskg24AxvbG27T6EJ
ihUZ6j039uKip1pVgl9zOhmP/YNVX8LV1MnjsyhS2jko33ReICDA8zIwSojKmGjuWhX1l3/5yjXt
3O+R/kam2VoSdJkX3NCIetofCDHWTq1Cy/8zlb1vvWyjKh3N+SN9FqgDqbziMyiIiaCDNqDUagkx
9nHbS+Xhg1m4PzsJvejKIRGuRVNkORFGp//lLQjxJf6WETODquUv2cEhLrEDPOqUJjuEvYyYvzhz
Pptg8c0OHYKh5OdPa2/bME/ycHNUcpJbu2w37T3Hm7TI0b9/GLlU/1N+hqXOLjNWxq8e2dC6Zvig
Ca5Bln1DwHsXUNFLVkAW9UgZbTglFb/x2mslH8v7opY5tvFJsPXHsMUOCHMsCMqC1hPeUCTl6W53
lEiH1D6Rrbpq7vqLGROyv5lfthHwx7z4jhfypyVntxYQGMNIYgUq8dHKsLSUNgFx3UVEg0x842I0
tujHw0LXK3bdepSe1kp/wJ6jmmrZ1sBb13z81Fluo2Sj64obcarujOje6C3DTUSx9UsuX4WoTO0Y
5fTqUUSquOiKQp9xwZy+3KYH8Kud0aNOLFKbW0j0ooWRkkJBOf92F3LId8lpw0k49ByQu6gnOMUt
GA8oEJ5+GEquSradty43qxfaeJSp0+mNVO5Bstjlzr7gkQps2umc/HvCgomQ0CdS2UAb6qLeJCqG
q5XPJzt78uiwvReLrRKGNPexycEMGHPbZaKSNRYbFTdnz+4XI3hcFw0+1WiGfciDkVyoFn06Nor/
DFywzXZtapwvodEkupdvyO7rRez9R8lL2tYcHXIHm5JWDl7PVW90Sm2V8/w0qgOks4uggMyy5BTx
q36349LZi2xi9wxfxIoDtiiXfsRTxf+mcEfgVdnhmLY/YSu9A9fEuIVRd3umM0mXEMOxOndh1FL7
YRwQ0pxrizlGTu9Fj34FmJV9fYsOp0/pJUg/s3LyfTqeAkhxPyEPt0CGVgfIhY6o98JO2vNvmaae
HA31A0KkqIwV5lsTqNVU61JYN3IJOWv3ns78OvI4OQLjcB9fPyGFNxsWVqUrQZhuq3CIiRSqVBVn
WvwhjuQislL3Yus/25UPrzghxuSi46K+QL6HHKX+2GW4uy6JrfrmYZiPMz1AHIzxIZ5Zsn9us9s1
QINtmfIWWbAIj4bH7KQ7TM+OBsOArNmWLyJFFtUhQNevykh/GsHLjAe3acaoWho5HIXX8HMwCMtB
HVP61K6MvNc+CG/c8KPDlP5eOZnUZfB4IAImbnXdro56EbYwbmEjzG36o+qcnJ0+GFnqiwAch8qM
LEoawZN1sJ5/6YadjcH1GB6v3K0ECwCctfLm3ezXi4pOML9FSHgQlP4BbbytAeNzdIDY8XpslhT5
gAHmYZhaACrv6th8BkVwuFdq1DC11lIjjlmnbvN0/2ziDBjNxdr13GvNRPhrqHbt5EyrKFa+Jplf
ov9mMfqcjZv1ehS3L6BnReQ4S7Cq7UuSOwHEsH+I/Ti88UQ4Z9rpMHrHV7BC6xGKKkvyB4N8QTKX
bxqg3TGRl2jJgb7pftFikOTczgcm9Zi/ELEWQff2XL1lLOQL7eAsdfBcxO8IF7i8Sdx2O1KQ7rm/
9ZdSwYsWqq7RAxPcPaCbHFUDDI/RzBF5ErCL11CsAytvQXYWwkqljXJJ2jXmGf8SUQJvXzVFvCOL
s3s4SpD9BaSAEDjj62gR2yNfLb345slptV1apJYJavnVWhk6eAmmBTV50qR4JoYmuWqnxKPM5xYx
1+wUPCVfTgYurs9cCCSbki/bBajFWErKOV68nKTk1CFMxxzMxbuzQsnfHmBjw9enjioEabMNiSpy
0eGVBRp8ZyBcCnr+TGXJ5prMAWiYSxj7EVhoJhpdGjLHIHuOXPaSI9tut6f3sqMyzHcB1VvFc88s
EppAyMf3veggdLGvBP7Axyju9TUW8wUytNeEp0pKSpTNoU2WhbFaLrd5fcRdLqynKm/UI+ZvRGgr
mqDPs0cbfFC+qbtzebBbpOTJa9B0CGkRAsQJdDkRHleR7O7GFmD49lAEwtk2D0d3sU3B6VPOh6GI
64K9ATcPHum50Elf2eot0zuAKaWoM2VJ2f+QplDgfwCqDooJQRGMo7h1gZZx0z8mJ2WL1B9ztz6f
o6FTwHeIY+pImA0bY45oONIlOOHjC0mdjHFH0l5WP0vKVZTn91oNp8wIHM5ytOdTra4/JLDcLuzI
snPrf/uD6vFzILszGldVPM7kXNjcqKWh5JS4Q1L+Kg11BFao80Xj+iKZDlM8rLrfCm4FxDZnoK9Z
jqISO/CXqECFz17nEAc+8iW03/5AxkOkYjESOATd1nBz/zyVeYyUyM8yev8MypwrhNzi2CFeQGRM
gPz2Y5vsD8i/PQMEZ98J4OYdL5eb6kKW0e+/QlwklPBypfTMVAS9uBX+Y9YCKlyZGQDDoGes42mA
DadoGtW6OkRoD/JjVk1n6yB8AFU5hEtSGVeTszChs9lElXORmhloL5vB4ki2VqwHBqOpg5ewxyXc
PlLTI6mao4Y4YIor+zu5VbacFPPdeWc3PUgkprvYHxLISZHNEyjTQhEWh5F2+7dSpAq2gWr+velD
pxTPfMIqUVJlH9nS7CvSHMWWxAalbFzADtOjZBoItud07MBz+XWIxmQqA+F8LFHuu/VJniSHqOAI
1HTHdIm2dZY85gMl+gsZOWkVS/gwdKSavYhhcogHOUUaZ+5qjHqli1jbu+vpyrQ2qEtX1kxPUMyL
e8fTQ+wslPx9B1bbrxxOqMOswhjvSxEcRWrrX55tAiPNxRPuYfXdVsz/UMJtn55a6XptAWC4l4yl
9WrIkhRQ06BrB/Qvw7naTjXRQgPBeWjK28BYo6LpCcqjbYOpuKtfaM4QAeSOCGerrTPWkeA/VYMy
lJyKMwFHSNoGbvP5S7tAWoc2Nm0etkTpU8Hxd6v0/kcTrH8aOhuwtOBYqNy3oGbdqnjo2TTizElU
emH8iZ4a2LnyOuG42DNhikudpqjhP+vgK1uos3myH2Sp5U7xIMNG1keIWuClTcw6mwxvsw0NN5wl
LD+z8d+e2u7bDR0APM2TRPsKl0IqHH7vwEW4mq8iosu4oFz60c65vq7DH0X2YfoY/WmvfxwjJ5Jw
cUaJGpp10mGj6wEMtaP3ADcUypW+d6lHSVIZWpC0b25pLGjNvGupO0QepMBth+8FyIObsX1Gd6JP
Xa2AhKSuuwdKc3Meg8ZjJx+i22SM5m+SHmHpLrRTBpPDTWo2+u/7kR74uW9fjqu9bEJIJdUKSBuz
XHCtlv2qglXhPYYcH+baNK8FCYzZsCcvrboSpjR7Zf1Ya92Pzm23h4YUgeHWtpVaZ5GBm3P0+Gam
2TryW0+rMNyUwus+EAhKPMMtASWG3xFM39IoW7jgyUjgD8jdKWGXNNXwb6+5lvIcHEEvZs9ClRGX
eUHkRo1HB/dMlEqs3/GJ3Ex5IVeOm9Qs0HVWmI6RAzMTiMrpS/qd2TqcKCDRExmUJvohqaRPsePZ
dxqqZCvU6AFtrADZtvQRVQyRhSER3OmyB0XC80PdeewcQbSDCTdzCmXBPnq+UchM/wxTR75N7qLJ
Lhu/Y3GDYpi7cN3fbUXx2LuFeOSzoj9heADn2R/ONYdryj77+le0rsB0tJokq8YePFZ2H8iObqMY
mznmecNDtvFAhVF/hBE9p+nFRXXxLGB3R4Lh1d1X0SEgpeaBg+LXl3yxdlADoqCLHOSWDotELY6Z
2KNA4XvWcYPyESOE6h9ZTUTM1orJvN6OsQQ+3Idp/82C5LqU4ajkZbZ5l0Vajv8ck+v6ZWzg8PDJ
iCXfM/G1UMwGKIhj7B+NfCirMb4MtMXWkUoSLDk7QQnd6/yVjLjEoFNxzc5cfr2FK96ERMKuqlS3
1n8w6cY4jPIEf9odJL0M6WZZBnarL6xQjcORDgSLrdZ7xqfJTWiKrdFOomoEzHedA7sG3sVk2uNz
ZVUCBS9m5q+Y8qFauzYe+oIC0NaUJECUttGON52geOX4oFYTLu4mG5/zc8Ufqxzp5BzQmoj+hEpI
r8lgSUYy5ocD8KZB386NLw1KZpVL8ZvXGvy07yologNZwF9a3QevkJkpqp4ALjT64LWfO8Tjo5FY
WCH1xmOn78nO+tLIgxQ3C1rMulb9pnMi7fis2GesYyjcrB2SZb5A45RcmmhtTBbeNxIiXtWF9WOu
2aB3XXWbiB4GtxUuOPgU76H53Zqta0JvZA0kW+rit0TqqONlKvV/z+SDPJ8Snnh7Cs8EMURyFOl6
FtSRbJr+MmIlq6Lh1Uu4oXM+YNnRMZnhpCN0G5ppF1qfSZQo5TvDC7rs4p4G+85G8sBY09UgMzct
aOURnENj4Jw/EzsHc9o3gpmhSTBMhdtqNQKk6PYPGA1Ip8KpSxNUvgrjKF2l2FA5bm4MnQemJFEo
cgYJssuPFRx4e2tu60HjMHMjojzzn/pMuxZsc9t80cNy5ri22HsJriqSskoLFpn3TkVvBgzTpddl
lCIRb/yGLpHf5xYPpDcMwByp0zwIGSLT4BHagJV74PcZAmVYsHI2inL55C9VXh2YNmCvHbYaCs7V
zbuZszg4wrJ0p/UnR4nJKL6qmsoUnKsA8BFVkuiULrE1PBDStKZCqtydKqmF3R/O3qgSiPgH5ptb
YjzO9ahH/TxQ7jSubzCRFeJh7RIxJSx+RMo1/wcViA3uLIMk1QDa5QzCoxxe14JvhLgZDgbEeHrn
pzuswP9YM5+92KCJqMQLJ0cUmTqRiCblaKAk70nZhiRM1EBk5P9roJparkPAilHZrVorJ31F/uMr
fHGhZgXc78N6/Uvu+wcPJhKCOxhp1EBAMH+kCCd2ugA5Oac0F9DHDz/HYef+SqRp+AlRu7secgqM
M6pEK/FviCeMV0y3LKxyleMjtGBXXIMKxjNOsJ0IR1tjh0qRt85wcp0fulqHotAt1NIvYFZD9XZn
hYUPe1beV/Nm2+iadD1E9uGBPXKhDrr64j1L4UYXveV4N5doCJU4ZnJ+ldG790jzNUauMlHzfRFK
rpChQYpEeNY3TLwxRviUIUEsQrqwFgRHKTJlctPC3Isa4DY3gJpDm8RUZ3rTChSJFtR14XVzS6bB
lpoUk6CthbWVOVufRNVfAV+svkAHUcKGHOwtmVOupPi3T1ZfRlnvpWFu097VduoEG8qgXJXR7VtH
BV59hylqLQdfN8PEQv78VcmepjGDfW1M+6aMg+DR5/U3aVYJ8HLhpuK0uP1SiKg0f1uY32aR+BPx
jMURSdXzYMccfso245LFHCRIw7cDWrTK34uzu8MY0w38jHjNOD6ssx7aiufPayTwET4oGTRoGCk8
9uPHpX4iZYn/SNcpsEkKQ5S3E8IOfn0k2H0T7oriCURhbIsPtsnAXH57tH60lNcOKiMbumA0Gh/M
V1U72ytblfZxo8TPcxLKf/CJX/pucWTBNpb9lLWWw+VjbCqDz5Qzg29A137FtEsowpG71oUPSFWF
R1DhlNQq3yI4xSwDEWjoUuvkupswseTnFTCvG+U3xcZ7AAYmxfjw0UcmOavteGtjo8cGqkwKhK1E
skUpbEPuOVT+t6w58KbnFO692228sRqH+7fzbt89bTw8u118V32kgY3jyHASK/vZhDqY6onVMXYd
amr9R8sxq1qDrbC9xVJ5dEGP/3wqy1FnW8SXw6EUEUBIg/K1wvthhYrnRSaXYLEy3WgE6L2ailb2
p0AwjGU6pEz9LRjIiRSiHCtQ5qHO0aV6enzlggV2EgEhifM9Z/ms48BtLQQxcp6ZJlMeVkh1q9Mn
VVWHI3JcSgKhXf8QdOBYz+59O08o00UoNxcBxFCxlRvuRiyAlfyRJdMqdAQFPUKwXFnDARfWxGcd
I6/a/D1di6hcQwGF21HOhrMzrzO0iEI4eRi4C+uRenQeBu6S12yncsGxvF4uMe5gPRw19oaRX4Hk
/K/6CNGnB9DlFQy4icaFr54QTpGpbMTRnRDLoNRrp6uAW6LPN+OONujFLrCUntwi7lzDKMUgwQtO
mpR2G8IJlpu2eZ1v6sgjkGyvo2p5+DWVXwJjyX+Lo7EDnHtzeYnXbmhokJRyQIlXnSpOBDKooOsl
OtEVtlRsOFydW3kYNBBxHbHxpouFn7rAPreenR4bdZbmjdEI0Q1Q+iK9oup2O9G6jtrx4a4lR1lO
2vhF6l1pyETtq2tOkT2z4FkqYCW34v96n0EbklKYFP23zbJa2QpXrqKYUuq/BamxRPxinxb5E8uY
XEdHetNwxf2p+GOKDp8yNSZYKDO6vCl/wuiaRRz7ykd1zyVBH0jpwcmAIi83smbSaO4UKe0xgUrp
lCBmPvUWdOVpDShNe7o9pY05Lt9EO+Mv8L6CKtLWKhxH80JHV7/Ub94UB0cTEzfgaLeJU4SszJkY
fWHM17Qwq2lpUaIOZ3TLPiAvZqwj3Rf3UirrgsWfaGDHKbPxBiywUXXuHp0Z2k+GNzuFJ1Km2vNX
YRfOLx3Rpzw3LRTTVgQH/R9GqORZX0Duda9OeR2ERhJz9B/k9IK+rKrtI/U2VPGuGryEUS6fW5pA
b4k8ZJk5uxtIjwPwN6QaocO830rAN0pR+SknZb4B9tvNuLrV2VdNIHoPFmwOFMbLNqN2hNsYvymn
Jt6AL+FG4+pSfBWT68XyRMCB/W/udrvSFCGwpYp0MF0S84qkgX34FG6E7QuNvshjmFUJBd4a/3Bf
eUT48Dc0pymtOx8+0+/j5jDFWflNaZASAu8sk+iekzmg7i3gzTNb+or4QQfFuwfM+RbDbpMH93pu
YmFwCnXSCuVQTPQNhlqcH9FcOXF3JzZhOMB6iLTLzkV9YZ+R5vbBQ5DuO/uBF3eOMb5+VUBbbMgB
a544SFt1et3KsnEQbV5prT5DrzUytNKF7J9899/2HjkUSwDRqHe++Aof5jUVIURoMomqaicy5Avu
ztJUKWBo5jYJA9M3yehCvnV9oIWd71Ms0qdAoZNqXdUXXYrlBfjKO8qyjJcZOW9LIH8PRHdC2Kpo
3ns2NNNPI7oCmylhawNNviDQ0dvvp8fVrGTu6h5o0NfYIv4GHk92lE+VpAUu+anFfI0fiIuWx55L
IwqGn15P74JEIHGHSwQsvAu8PSwh1AJik6Dz8MhEoZwcgdCe0NtBUy3C5ggu0v3TflzcWs1S93qs
6U8wei680m09FTpd5PBNxOL2PJlJq/fviyYUpMps/MF2BTyDRfE/XWg1QyR1rXiyLbW6Hi2y10yO
IXh1oJ0uuLZFxOpuoV6pczHoRfzCGnwJUWZ2nqhYclsxEOhUfpawTAQDVwEW3DrbxnSiH5/Oh6WQ
LNO0XZ/MeQ9LaDNq7mPHhyqU+u2HCPR6p2nsZ+oYCb4j9MgmlqP/YetH6ziAkh8HFmsfrY7CcWNh
d0VLLcWVm6wIbrKshiu4q+mXxK2aixa/H8onLoVSQDB6MjgfFPu64cMbViYmeAGzxeZtYF3BBtPi
T2VzFTy+8Kg+4fqJb5MF0ToFfWuMYiA8fDOzq6UdmQaMOlLIRUUmP+h+Ee1Mi4k0+ofHTJZf3UdA
AQfIDHXvQfbbWDECdyVzk9vK/4E/aYEPjECjzDYkkVlhDqpMwokYwqHC0OCpWtjnyeggFA7AsBOW
Igs/gCQ/qtS9LwVdZSHGfxJG8HGtFaMzfdaqkg8ZRpNoXXxoz3s0Fyg1IhZCy5Z++O7uIw97YWhv
8j+gEs6jpBRoMh8Qti6mZI4Q4seQpl1YLFBIG7U9QPwgUkw14/h9IWOMKnORgaueQDpi9MuCoZDL
UtrM7Ta7YSq9z2yB2OHRNbbCermKvQeCuZOPPETOGpWS9nAj4uRAuLIgHcLjkjdUhGdOvyspiEf5
dU97AQ6SSilhtrlRkW+dARN2ONaaLC7MtBYYuSt1uozfh4YuqSHnBmxSOqQbX5T8nALmf21JlUyi
gwmUa5ZPEMxRnPEF55nW+ugKgmflrUe2rRpqnXLa/HYFjO3L9DWFBiMSU66q5KMrLZxIWGNe2Nje
Bb1+yOuCmLWjJMdXqtJZqM0ZkzI4XLrJcXh3iwh4pm3mUfAcy4HrKg3Hm+8IsJARTF1gY6+YbPtQ
GxIgYixnIUAwsTvsSw1jEOHaGhQTjlBCQJBoZcdLIoUYqS0yIVrho3BCbI7efXNq97UHxop4O41B
NWjB5BVpBK6/mLoKU0yuedYBXfhCqLhSo8w1PlcdTN7d5BSMd+UX7CT3P6xq9YWfw6iFRbMByzCC
qY0svIFzeBRSI9PaGZ+itjg6xDss6nK+GHY6h8uTx5RMm9XgAttguFfvzLXWWRSWQgAX1DtRzcBN
r4E2Pjlh9qTI6CjBjK2kmMxUwExGOZykgGMvKn6qni9cQXosGlVGQAbpZM72MeqGZa9gJX93VR7/
DwiPeh1biYCStnnCPElwrW8o2SGU/HfjJeink//nDjUdWWId3BoCW9hVWcnC6JsEW7rFHwsI736a
Y2phjcb+uTrPg480ZxmBu0AnXOlTP0AoNurqb6LBjnRO2KQRXuMiIpq76A+CTI7cBoazS7/AUjVn
/NPc6e0nTL448ydeuln33rMia+yPlAAaX8FgmCRqH0y3VSrqcGy1xDaOROs/ezsj9CxhA4xCSIQd
tXvbAfb23eN7290Pu5/rHE+0fDX7sprZNsACtJcRojwvB+lchsO8JZRQqfOizOkxMx/iNo1URFFO
kWFqzbbcikmBGYF2usn+Ob2JudngE9PYt21utiH/lQ6HoF/wfCpnXuUj8Jjk9eynCUmGkDvOB+ve
pk7WzycB77Mv6krktHkFVKqE+xwcsx94+KffAH9woqR52BwSmV+Bfh/evvvPY7hJMkXso5sVcArL
C3VNV2p3saS2MgAEE1vjQzMWJP2tnh8xa1KpSoQo0C3RS9zRFKSB1G3pkx4unBALupa8ZtmoBksk
/PhgVv8pE2/uHLqpca3HGa2IJPajIpcty8YmfezRpt/cy/7XJUr3qEFnpnW4hoqJqpPFlPDfyDsN
+Mb/Iir4wwTKGinz9UdY04umHH7RBVr9kNvPFnO7VOuUJZ93LVJ7bgdNUPJPvl9Deqt3hg3nVLVE
sQEz8sNpel7lpF5e/LDk25BIgs8+qzmh5uEmafaDF0Ia5vh6SsK+jFZhvuc12kOEXn/wDWfwXH1S
7JNA/qw8HrmWUYmZPSrb1rA9j5hTxl91l9IlkuJiHqytkeVt1ZGwXlRsryjA9OsJ4OHVnz0gezHU
mgWMnQwQJK26GoG5nLIDaQM9oBLNIZVtoxn95mwmdnj5YZobeUNqOLh2gIJ1X61DZd8+FZvF5HdM
auE37Lk1De9dhp13AhGd1wtJwnvhqLYvVCHpN64kSMQ3MKFe42E3hEHgQw3AYX+LjWWJeAEmahP3
xgQL9uXOTdWfFoHWvUNikf47dCy5GbWA8r6cadwwMgg6ODHNFvKfhELL3GNiOXRIgwCPX9wPLgHw
OCxRoiXWy+S03SXkLos5ta90BeX25LqBTMCpdNFvFXn0G4t+yxjy+AEByzg6LTiq+REBxY33amLs
HOjKoSHS6OMqj7nwN/rJOxTxtnc4pRHqSDNa2ibf9Jwv3iXjeqNjl3N1Q6E3Vt7/4oHEIOWyRnEc
HrfBwKuoUNzHZzd438mbGHNtQArstaFiv9ZbSXgnIxKELEy7j17Gj2JebdIzP+dpjlSUCEr4QKU5
VTHBVwsg81TgL61dHYMlwN+KlCr4ctV6s/b6IJb9SF74Jg7JozH3ZAJJlqDPPndwQ/bSS2KtdJAi
5g8lLVdfy+bnCWXBM41avIN3ZV+JQTrWyZFmx38ULPjFYABqHyuH1Ap28P0f/lE2LcmhE2YFpKxL
Kh/HtpozbfpQYf9hz0QQXSJOljFq6FPHoX4YoNsIdS6+I7AstmgQDJC0io3EfoBF/YBaW9MCfdT1
HUYbtD7maHvRJE6i15BZAUvT5hTsM+eGkhWBzG9Lg1jKdExtutXX98kDOX8ZQWffAYfE+nq2pjco
UFAJKXIybc0WtQdeLw8JcmqUqjsdQu0JlL4nJeQFhbdJw82loQoyc7fx5mzKF062HjTyC5pjVEZQ
uiwVrpFSj9Ww2eY424lTTli6jy18HmF+5ijHAHMhsOm3V8jDV61vcYmI9kaj1eX/jo5ZCVxxfhO5
h62tn/JURYrbvBzG/dURxegOeIUcw/UpueYbmr4+FNW7QHcEr3/t9Q6rul/sekoFmHbSvXB6+JuU
phWA47ciwWNMRcBQOw6G9+YhsuzZLt6cAg8RtzgBrYin93+jPE93mFyc15jaUlrXM3dJnVwz+Egq
uBzDQJ8Zqga97yHpYxIk20NY+w7lusS1nUT1ox6aePFqjA8YFlGE0OSW2g30vlYqgmaJO499POs4
8iCuo6M1YuyTGufsOTjEZfMIVjgkiVwW0brF8oUNpUEmr0miApUf1m2e2rYx2iOaSVz5SBv0b+Hj
3JEcZ8VvU4XOftr/UNQhU1PVMp/e940uR+5aJYm/TzwXQZF0r1AZH1HQk+kMcsFQVQRZK4Y7PCaB
ptSPhq/BBbiZV0O4RIc0BMvtnMaUjn6tx1uXF/TnjVu7OKKeWCIBDcVuVaQ2EFx5yaLibvuNtywu
T9+PCGsLe4FugBQpf3EU7rH0tiUty3vk1GMQ8Edm+LPSwwNXnZaKvc27Gm1kg0OCFErc5oxnWmqt
3s9bScMSJKJpKr9uL+mepls3mEzseWeIr5x4tPYOmL95aQXtZI5taDPtVSdnxfU2tr18y/GQidqD
MBy39ZHWoXm6hDj9UE6uCEyzPWupSHRin/asht6EjKb4g5TA+s0tAfkM27IkAYuP+XKNZjareB+Y
kyGNa+SxbNAMHd9ifK6CIZxzp3tFSbUfmoEe+x7rCwErVI8JwbWJkg3m/IpBP3thSg54SXc17eTH
I8iwjD3+zvy9VTQyeQKejHeWjKyFGoyIdUiYyCs9MSOMOGvP4h48eye7uA1POkv8EulQCKKD92Pl
dB6pMpeitTUg5Rc8DMklZtyeLuqT44lNkHlRAvf83PJ45o+RCxBRP+VFuFxH86qYdo7vR/Cs8s2n
0aYUHpgM6fCc7bDJj3kBhrdamdxyP16B9+vMQhYjbgJoFwIuFL8JRmXNjSMEZek93oH9/iS0b79f
bEdh6I1avdmdoVBYH1AGHv8u7TmL4/9cmKpKZhuaRcCan/KoZJ7rYSSt9aq0ChMGM4u9obCRmUaA
BhncFbAk9xiV2YsAJt0hjiw29T0DP1ZRdYK9IusUXkscS+sV9T+IUqXhv2uGc6Tov3nnYp3qO0gU
BXG2fInIxcbORL1bdA3zATUohhB8YH5YhScicTABIMQTPrUBezAz263p9IDamUFLiVqxu8SOifMZ
caq8MaFiR+MLEgEKufO1GpEgaY6lSoMzmjccYtf2gZB79AFsZTFrZ0P/ENSoytBRJdJ51cmSVDPV
Nr2Vw7Pw1gImyO/doHLnmwt3eeUE6h56Up+DdcnuZmgbx+0Sor56aYkSbtEFEU8O5PwBID97noRM
jnh992DLUfXbtnxIa3hqjnqAzScuX+OFyxupc4M2aVEfUSch6cB2bVRrblvl0dfc1GV/qw1PIDuM
gunlGebLeOZxDfCoMcagYhjK8eLoYyn8hbITgU2c5i3b1v8vsmKbGxZWYcfaqnj7JP6zp35nSumY
jdSKfvhmotodA7uOkbh49LEoN+fOM6rSKC75Q6szs78s2iosB/odsNYoNZpNgq3Cp/eztiWUD/Yc
9SrQMm4dGk2oUr003WL8wq4wNb3lz5BTt5212hoBgCwyGHo13hIvz2oBpxiNQCBBavuvJivTsDnb
qEXVvimanC6zrDQngQQzOnihuCOtcvXSdoa3QEb2wj8uO6ZsIc1BckYO3lvcZRZMKnVGxjh1f/cv
91VXIYY+3YKJ86dhn9PcA6NncgePPByPNptREQ1Ez89ga2BslLWD0OwWPWEnFgAKLNBAqwsInLkZ
Z/3g2TXil3mNsRS0rjpG6f4fVYyj4PvS9YeaM5OEGto0xMZds3dYcojzXUprs02Gv1RZDfSs0Z8C
Ud0EqLymSbTFOkjHdSEcfmmNId78jqyg9ut42wtVJ5E38fNzs4kDxj9G0CsgZAlDFCNiNu9BDqdg
icD8YqEIeQIqU7fPrAmv0P6ISv5eOKTEGfZkgiafgh/foaPDPgpIAqhCY/UuHYwakZy4tZoPf7h5
856d0OWZRRTua1tBo01NLlx20Q8zGHn7NZh0KmDkTHSknE91zo3JH++jBln+nHUDbNjf9ODknIEw
Hjtob/GrhBeOhY91oWtB9zLk80/ybNS0Hw0USBX5vm2Ng62gC8ZlG5PwIqIk1cSbbeHMJH2iCwDg
0eNlPiJCl3uxn4OPkFeTCCsPr5a9/mVCwd3yuKIKPdNFOYsj7VEbKkVNlfettoxYlooL9wjyTtBJ
Z1uUiwEoOR3OWZWjRL9T73bZE9FkaqRiWDx4VOvUb35PcadW+LIgtWA/Fuao61zlhnajPgzjPQHh
ULLOW5o4epwr7lljuE5HEpkEC7NYG0A99wNHbJkELEvrI9R9QYvs6p3fMsWy/ymBD11jNvO89VUS
RiPwLx4HMI6mNQ7Bl7fEnYBkj5do3lIylMReqN1xs3yqEMlTdzc/bTYPpNhTIdoOHpt4oFj0JMTE
zx/cVSSHh5YY0hTDj9Xa4xlS/0U71Uwdq0zOF+tC9o12NNv+fUXy9P39zCkh5hddtgQrUdL4m6k+
+ZQfPKc8WT5XcY+lonw1nJkNlNkWrTvzjbKd7LmVVA3QJ4OJdTTojdLbE4AK3wCP/p8c9YHTCvkR
XQ7DkuNpFbeSyOKbqTfZi00ulgyZCzgkB7Cval7XHG7D6ZKZlG3kUAK4AIntEJTduL2Yv3lNvGmb
eQo4HCnyJegFy4WepAoTQapPd9jDrp6oKO+pFvOPGlT555bQ2wHw8EmxWBBVeirMW5SwnaKBTYMR
wxi/+vbGfIW+LOWHOR7Zlhvg96CL0qvrzK+GoSPYTHMhuyYHnZPz5u9wcOLGRaX9iG7z90a1TYMV
EGdTFbeUYBzVH1pwU85FPHU+e3rLy5ePy4AbrhsKOefACydPa1Tg1GirVcPphe77qzlW1/Vtr437
3SQNPmtIg3cd+71WIZIrp2vGY6fmyXCcttXBC5oG6Nm5rU31KrFusBfOvBeN07OLC4VhLh4D/4uC
CDyxuwtgITjmWH4v81SMre+qzsPpZoBH6RQ4+dKPJ6xkR+wNH/s873dtZwpJoa0SlfeuTywhOZzh
pyy2dF4jYJnr9M/59uJo2eilGS6M2Rc1ppbzIoOaB50AgYvuUKZQu2SXuryGK7HoW/9M5tUsXLmB
6tmldtDQsnq6aSN26gpQ/QE05Hndi7UTZlK6mknktqgJVAaqJ2XYSEeuau/8b0IfCYC9oN5KtTdq
GHb4WLOi5ndVa6BumZ8yFr3VtrQWqb07HXczzaN3A6E0U9vdeKg39CkO2dHMVbcW66ZOAZWJYMDA
yTsDE1u8H6dBRaWdo1C6H2gikZTDWy4cTRka3FSQY8HWqMP/ANwp/7X21/Q+DApDooVTTlafkGvw
OMVWJQaCKS4WLe7rcMAMyD16oFxoLAEGESSfBW9dJHDCIxdiI0x5/Jj/QScjvMIllvqwV4dhGkI0
Wbprcg/0cj0/35Bdmf7hLi11AIUFBp7ta2T5EqdDoiW27f6cLPaVDkDgtqOlMdyhZ2NuU6kJCg9k
Qjc1lZ62SihOPCP1aCDJ/mkD/jWjWM41Nv4HqYx7taGOz43UhF6FBZn/Ytja96W0x2Ktnn1I8/HJ
jpBT2HAMOKDWoYOLL/rQCxQgpz8c9+R26zzp2Y7cinnjUTYeVV9P2VTkhKC/CYSgr7+A/YpMD8tO
cs3sayLdXpr6mEcF9PouQGb+hhW93cEEbp+ggSpmDxP8jCMzgXYzjQ6KbUNw45W4XqxKp6q2YIac
mSF/KoWZnelk6bMtJi5inYzdBHCFRau/N7Y2y1yVxIqeevcAR35/T78PoVGCToBvbditnvw3PHgB
0+gueYDoISmiyUqNZCj/EwBCcs6f63Mb100seFqXtCrXHtfOLBUU0naKlVvHRqST9aGmnqWtcR6U
5t5DM5HAuA3XkegcIqP9H5U//ITVa/Pnvp4e6gUDoNqoFddxldqgyuBgUQMrptktpum4UmqR22od
1RZbSzBYRQh364RTGRPj0iZb13PGIVdDvFad8JV64mfJIQQDME+eA82D+xiHnu7RtCrNJ286XxbJ
NomJ9iS7hyOi1tmTs9V0fQkJ7FawcDQmoWYX038Tc263C9myeRgRs67NOIE5mkE/xvmxVKpRR0sM
fr0jcN6d9rUQIjsa+gmb9syhPtDcCUXG5clzQnGHOV85VCR4p6uF5Cl6KHqMfpUBE7bye6/u6qRd
eGMKLVxWGK1t0BS0OD7sAtCOMCasEZ5F4nU+TEr5F9FXt8AiWMw12WCmlVysJlJmPxZRn1FSuysJ
WOcxsmxXQTOynoU6MKKh+JBo3kU4HRLmgRaqNc4NilKlEC59jaz5P7vQ2/N1SnryzRfBNW+n5h/6
QQZQMeSzAQyqRH0OeonIta9JtDuwAFLaKpEiWDk5rdhbPAGKtVloKQQGt2k8KcYSP89IXO7nB67f
1WocbEzu9XdXhPidXuseNKsX50n93UKXdP6nY2roK69e92b8J3eqqr4BkTlUIv+7C79b9+3iO2fZ
SaEJ60D6qfJETz75wungzu+PD1dm4qji6u3wx5hNm+jTIxlldLnEFK3KXH/h7mElbFPnrincGgUv
eHp6nNtgqP5l6XXek5HTZo+uXhLucT8glQj+y/oV5AGCi3asuKjTDGzs767K6LTNG1ftwLR4EJh3
VZsOwGrDpb4Jlss1B+pyg/9ml1IQhz/BTHm/FdR/fHuCDnmNExaUASCaXN2fPMK7I8dLRLOp9mLL
sGoJ2aZgA+pthYbbjf13JbvkzH5wd2Ws06KxrdvgFZgK1w7PIc0EGXtijhM///M3f6JTns/F8FY4
A0tmiTIG4mj13oRqTiFBQyxEsFNJz1T66s8G2WndaELKwE4vSOuFYuev3nDpqxt6rTK8vDssWBk8
nbI4+LPTDg9CRdQPATblUlEagIWQtyvgua803/wkclY6PR4Hhf8GiHyl+NKJYWZFExQXVdla7vzj
+ekgAeL4jY/olEqIRu1iSe6lHvvZEmzEx7ZfF+6wyU0PNQ/6WW1smYKxpZdiyLyeP5CDdiGhJ7ky
OVdnLrqoYt65vMXyzvcfvgl7ufp8sfrr8xztA8b4MVvh0+Ou3d9F/YvCypa6J+1L4SVAsX1PST1O
4TEzTCCqzgvwg3+THh1TfU+I2fyEK47ggAMIqMdx5A61iivBbdYk9kbAWD60nlHH1XheiJ80QRK9
c9E3+F7818tDQzO9vNUUTt2AZhTEQNYJY0kihVfWa7/7PYKbHhlSs7Jkto4z31plh9Rrdl9ChvZH
5+X7VwBrEAgn8vIqYo7Vfhz7df+0DYHczTchvaWsLwfayp9J89JMXbkmI8t0VL464+ucgzdTk95J
nnuGl0WdXZ+/NREg1HySlbeE6wX84Ro1UdYsyyV9Fw87Xlz1YXTZET0oQD8vqOeaugcUdWfYmTFt
ngjNxh3ctvOj9ckfXur8/nayV1hHYW4xsdTjU8S1bRo44cyqPdym4PywiF/7H4vZpcoSPdpPU8zl
N7DbUPuxiQHKHiEov1JrPbyD5rBvMK4S2oCyToh5L8mLJg6fqpT7YGM195iycHyk7RO3UxrH+GSi
Gc8rJ5NIz4g2HWAc+zG1VVI28MgM4+HIgxQT9wJrhLR9tKSh7Tfm3SLrRmT8sebOTRmz0EpJwcg5
y/YUXE2FPDDVqxf/T2caj6PjRknd7kl/nIVk/N2UbWWYXcq423yFXo4VMpp5xcXSpbIw17kqzhs4
fgrEqWON2n242tLhP7zt2YFhLuf3BZE4V6GtsjkWj26rp1OAOduT9eRwGpOJSm2vAw+tgQO0v5Ds
jWsbjkYpQ9o5UQ1KefagGvPx0FjYKiY47dh57n+WrefVoT68Xua4USW4txBMVuKz2PH83BAknyYQ
fbfLFHUoITYgyakHpfiBHqonAH1g9L0xchy62OuujSA1mqlCDPqtxJBz8oZ/nz2ZiSC6VnpHhPGO
QMhK4KeWaEB9zcyHnGVJY5MQeQrGe9AJsjHFJmfAVg0o9dcUZpOcGZUFwIDWd0kCKu+YEJvARbhU
+0qijNZVyrw/6Z1gUkwgJDirdGd2ECtZgZteXxSZthRzBHzLeq1xs/AnC/UaT4ExCT64fD4Riw69
MywnAufnBGgQa00Y/OG445pJQSzkEDSshgxCMGmIy4diy3qnwCTfGE+Mwr2DTCIDPJe/5h0Ns02y
Angd/rt9YeGut0CEZ7bJXBI5N1dE/at2GMtEypSDekJVMEyERSjsp7tdUuVTZaO6ETpqAYMEcqEK
LGJ6atCTukfu5BLEEXhOtQh/geNEvob5RpVZ+xior4oC7VkvYpfAig6yqWYS29YfL6UKXQyzG3Ae
MYHPspr9pXaZm0MZucv03pifBlArr7uK15b5BMK323bwQ0kIIEnUD+ZpTTTr87JMJST+IESXj2ua
oTcVbw1bjbarscLQX/Ci17GJJCivEib0Pg4jvqw+J371j1utpzPbX2bsgKTRip3iE4sMiEU0BulO
6i/0gjlsH3Brb9xwMNy+axnZ+73Lgi2c6X/IzdQbXASg5lynLZUAwkZzkpdCH+Sjd07r9QPud4sJ
tgULqfOyCjOq+LU6rG1XfnlUvy4rSYN5unxe1+kdlCdXj+roqDns0DlWP+I9C/QEy0P33aomwLQq
NRRoXfJJFWY8YoDTWLQpuLPdJXm3VvuxGJZDGyydtMC4zMuAbrQyugwpj5LgYNgy6uWZ99En9rUC
czRnTa77IwAZ4GXQLn81a+1TdW/vt/i0b7KftjfmZh+igeROxl++15u0cpo/vdFoNTvmbhSC8h8K
eiP1mGEd+ZT1ygzLnszHOCtp8sXbiAsm59/qihs0yxWdpX39lW3mvQWbs92niUmSsxrT0yUV1s+n
NMkeY5R3NCM5c5mm2maUIj5uRc1ViCzoD08xSo9rAs26GlOGoUhwKYNjEvG1ly2a+q/FIeF7zRD0
dOx4OVwa64+XXRJ0gSxlLNBo2pfZ5SrfoQcdFq/EHnLXIyZvL/dyF51MUg7L15o1oTnGBlZdsu4G
fRwce/DW1cKGVrzBZkAwYDHOa8H9jFqIgpnkgNeeRfIxCttKw1WW5Q82fAgfJ5FZpVLIUn38/Ftb
lzzU6U2GGP6/GIcCOBnDiuHnkDQsemhrsl8BLLqd0oOQfohZ/K1AO3g04htI6SLhuPOgiyx70qos
uq9guzPnsDEQgD6ksenQtE/mFRliwKW6UCZ2k78VYJB7X0bMJSxBF94d5R5kCw8YJJTTRjOG2Y+S
45RWfNZLHFv1WEkvV/JViww8g9Ec0xj3yrswu8wFrd+QcCRzib9OTc/bHnBoaR64Fi/ecfw4vrgH
v4lZz1504RBNK/G1BC/Y1MSRX7GJAanKjmg1KuXtLnfk3kMfQ5eNLi1rxeeIEIDNf03drJPLTIOJ
pM5cV/SBjOBnbROkcm9TpwG1qUWk5JcbXQTsNhbY3YaeGzDv556fJwnoBe+1vDPMqVBjODvAl5VE
T3EpYe1jvn86w4PaEkFqhF18al34zPH8rI1Fko6qeqbhZZ/55Yi3YrAqprrs8bkRZXjOtpayX0dC
ZmHmsR6+Xv7TDblPIBJ+ZX9o+j05hQBfJSaNDTyK1BGrfQNtZX6PR2aWtvDxqf8CJ09qb7zsCCF9
I/HimcllPfZBxzBqtuCSOzAyOyoT3BTALTRN+PFcBF2FH+GdFontqK25P12GpxLP5h71TQEmdtdd
VIeP9ZiERQKrjn5Q3ilek199BVShUKuyFGKHF4QdbYVCrVdiP5aHbFhwsWb3XPIQtjvwfDn7cNbx
t1QPqLNo4VmiNlyHKdF3pntq2MUc2k91EeTjAKxX2G4gQuZcP9cBiYqV5lLnCFIR7YeAXmFqUhAz
hmiWK+yUmFxs1a2CegZmHG+/36YUi0mcGFcNpkV0/DrcrdwDdhyAp2FWWV8MbtnvyoXQPi67BBk2
xaJp4MqCGXho1OdIfEq8enGaTMvQ1Mhl2p1WwbqBH0tmWVEfCJyYZ6LNfJGVhtYMepfYSvXDSNAF
f/LPaJ+8xf8xoa6ffl6HjtodPPIGT9MuKXjcRP18HFOqsaRc68M13M5x4TVo0T5VzWqMHEUGEWG8
ShJLEs8QcFZwroGPcRjX8ZH9yRLW3kP7eFsmcOT489prqdnYi858q4nP9N2F+/QAap8g0ZUfIWpi
lrhBk6jmUie1Tjz546FaocxTllAylKCTnpjD2ZGeEhTRyCFl0OsfYU3c+oQxRxt4uCttyjgMEn3Z
4J6IMm0GYeWbfDHIhUNHUDgeHfwhp9PF1RCbX5SU2pmPlhV5GHuHssA5Va105bXtYqeLqnZ0Tbs8
gnJz2NmQL0Deg1Io6NX+ukvg2ciN0a21OwEXouaytVo6tmeieANFc7gW3cpj9fFrTZLCgZCjiglk
XWaH5gyl1ze5mtxldtqriwkZT/zU3h+IOcGQEzFwNTa4n1qOzD0lWc1bfx8dMHQFn6GLit4DLSCa
wzErG89GJvtaUuoWoczSUIhSbj1G/mpxLuycKPMuP1okFJtNKfOU9lWfAPS4kdLyQGX1+Pw6iOiW
KSxO9VtGBYT6ONiQa2piAu9DZI1AxWfZOta0uX3EF1DFx+eX6xc24UsCRO8Z3RjKI1Bkp0J3KZVw
6Slc7yT+G6AY8K8jhdZVNejdOgQcvjkjvZ+IVsHxxdycfUeYG1Ns8coUPka8bQseD5JghNE3rAyk
zpRw9BZ4LQolrZfYzkeBucShCeOA4XVyGj/eaGy45PymXnVqfXdVIjxJ0R4Cbjr8SH5KXEDppJ5g
YeoVqvmpmSVB3ozmOOwuJyEVQNiEJq8qsODggZw/Po7PIFFUVa/fiIOB8CB9XG9RydtBYz9VXxCJ
eoe4Pv/1eSfo/aO6NO/+IrdqTatUE7DlLtv+imzKXwF+CoCNb7syfsIpSaD8CbpnhMOsWETtzntQ
YCrNMqnxkEI53OD71SVLNeGHM65xRsqVUDFEHKvFWY1xQqNYX1PlPqRpianv7xdgPnG53YUskZy/
EHV0JlSWrWkQKh0BXQunC5gtWxSFD0BKwPngXT1ja2oDyALB4ZGKeQjVUm+6BVzoLSknby4c3vO6
oF+zhU1U2L/1fUhBWe5K3REYBcz7pRr+qvdwv7xWtt+uM4mbgWGnHiBtadk+LPbc7kjzVKnwEydK
syPFzusWz1GtXVagLpgQUNWFpHDXxdeV12Y3/CFIeuNmg9zojKbNjOhamrv1kLugVAH48ou+hTdz
9/GKK9UkPf/E4x8/n4HHBubnMFMX8o68msENtVc6aZB7t8aA80lWeCjV6AEFOb6szcT63s+Jzvfm
u7E80Rn1QoWAjpJ3p5kL+jdkZHRB2TNwW/DHeLCHnsbyd+OvIxrtFHuPVh9F2UbPpDVsF0rIuNxz
76nbr2eBGLR7f3DXiNc7Pc5pDH0EEokph6W+mCR3e5cEq077p2rRnRlQXLe490G324x8NIYqxXql
wmhf1pLKx6Dgo+Kv4LmR+OrcFcDaPTZ2FQDJAmNM45nmG2CNvv4zlSKXanhCEvXQrSAyc3oe8YpS
F1rWiQzJTFVUTi/oSqSvrgY+4ktEwrYctkmq/jdGcaeSDjSqj/p0MQ9LlRUniV2SnBnYZkN8jLJs
L2e8dIs4eON0PDUTOjTxRi43q6I8FZ/F5Ec6RCkKmcjcmQAImiX55Hy5fxDe0YzIeY0wvHM3kX88
Gedxd0MUnUkW48Rj5w83CBQBgq7q1KqBzBMP3vqxlE+kH/kUkY39IXyvG6n+pDSqgikV2ndW2wTR
dEsnS2VoCF/Qcy0Z207FzchI7XGhU2fG4D+T7MrcHEw7K9S+Mn8fLJiePvnnkAjTGp6ggfll23WP
PGTBrQAsl/b7jIBGjS+rD8FSvzQuMzL3rR00a903mQEKHzkI7x82ydEoFuoBtqKo54SXNYxLRqke
QB7RpwStWitoN+l2meEkHWXl8no3NoAma6No1sb5aFfsx1w0xCesXDGfmryNeUpencM+erW4wjNE
5xLy5pfgcje48TxshRhiEWIVTSNMwDxEgQQaMLNzIuYg6lJuBAIgNxzfKGHtKYAcrkQ1jGe58yr+
ULB5jyjLC0+oLVJKfLVO9x0tdt89ItHsuRl4bUuzwbM6meyIAVxu/FyJuqn9lJ5w3O/lWEe1pNl1
WXFg4GicxiWSTRccmkwyh0XveX4lCRG5+4c/l6OXunqgne0yk7VqZG8XQ/G+EmicYsIg13iy56gS
ArseYImYZxTbGpYbf6mUESsAdEe3YIA+r1YwaVUzSANOPbhtK/lztMP8s9vcsNs/fcACXylWp3TX
L7pce2Avwi/mmbJNXbUS6sDGJl67r6vkqjNp/noAgrnFLlp6l6jWX1ADMTNlo5ePkCwEwT6tVolY
YrGuFyhQWYOPwZ56kr37PuWhSBQl+oVeYkKA2IvlXut8xE5CRUGzyazHooVkGtKtm9S8HAfAKhkG
/L5+sFFv+8Ds14f+DPhpE07bcF669Eo2I9V+Rtmnc6NZPdaQBKawmEogNRuEaJ9v/gvjVf/dgcQs
HNh1hny3TH3Zn3gn6NKwr0zrziDAc8UQZq/kgS09U/DIgl0+PjNoLz4MwECE0svycZkwFmZXIoKY
2bIV2Q4OGa1Xn0TUMmLmI7QS9z2W7Npqwe+yPEbW1g2NLO3NY4OA+vz84KdLgdJJ6a77h5YhAvhh
8Wf1q9+0E/n5roOVvWFwbDIeTReZd+BcrRnc+p08IcB5dNXJpaTR6+20TwnttNzon3yd9LQny160
oPBVAmY0xK72UM2xFiby9D17opi+VGE1jwJJgXaOAeU5VBhRt+aay95n05LS3srGcDvROOZ/qM+m
J0niC/ik46L4UxwP1BL9dMPaULkhRVr9NR1OEln5I8mpRP/jUJIf1c44Q1lu3BvuAslbhi8yhXDg
TDst5i5qiYtXesg1JdepAwtIQWExF+YpcEpIC951dsgq5941Al7rItRVaZ8LA9dJmRaJC/4TjOs8
72b3P2wiyYU3NiSUnxsu+SA8leBUYm/hj6Hia+KiWkYVPM2RWJBWqsw6pVJiByWrlHsOJBxBIFcb
aqBplY55Ga7vM+YaI4CknxOHIMQA/eiTYvOyJ/6lsh5PvfN1zyud9lqGSFE88JuNWpCLshKWRG8P
PDgN7cHayTp7QEdnHRo6pW8Zw0n7SnvuSjk7LydpZChTLXxaCBc5AeEklLdR1wSP4YTa7vGO+Mkm
pTwIUPB4ljV5BMbFXp2GdJBENLXNIJ78tOQM6+CKQP/Di/RoNF7cJ/Co6CNw5w8xNHarB1fgqi8F
Dj1EHzNK0rrnZs7xKo65jga+3/o1ILpbC4zGuqCgOQGZ1ttMOc68DkqIhL5KCsXwcVqDBV3MccrZ
ZGdRBo3wES6h9Fi/SNQ8isvrw8VlxjopStyBZulx4fU1qLr6l+Gmfs1p3NxYCFUEHuMon+Qji+1s
2FVvqLAPNo33FSpCt/DnjNjuHWcJ0Wk5+O0q+OE6Xgs7fy/Z3+8grPUSEj/Vq2iy/0nkMYkFDpSO
unLeT/qZqDnFNVwOrWqoq0TZYlkKgigmpKBritgqW62jTEL6KuIiV9oXJERIsqM6UqneuZeq4VuY
ta/KvglPTGixPHeHzaEUbnPJ1pjplcuIcdHniC2suu+bDsWUw8N0jdiZqpIo0emM2cJU5vqnzom+
rcIwCYUXn64Nxg9fqWNIvDUCHA7g2Q5rGdeSvoWjK1KY2nAGLt5T1dbfzN2WgLTB5NKUrtKd2g9q
DiDUrAjYVXa7gLwVq9kiTaiAAdU5cIFGPUXGRDFGVaQUOo92YZepCxIZdHZKRZCNcrc5DqR5aiwG
M8ZaZbugM4cUxZU9VmYKRKXF/0+Sxg54q43IDLqYe6Xpw04t0DSm/Tjn/vDk8Gv5VtN41RV2KnLq
Mgc6MXDL6IhEN/yUvt+6Y3KUONdffeQQGTmrd7NbFTZaTs72byfcIpJ00TwIpDlhmrasBMS8q+9B
IeVrgb8HXUJbioh8NNXK9tDfhD+iCjK0JBy9HpedoZeQoYFYQ6ulVrUUstGkX27wC3MXsAqfzctS
DDDcRs3XVH72JEEHk2h9zqpPpzDtv3OpCMh8fpBhGNyv2OO5o23E6N1EUbVBD+ri4K88JYf5eAbQ
h29gjWBRbD2ROEGnPcu2HoX16fq9BXjopmV7us6jQMAWDZhY6CKWm8kOvFli1eY05OquCb2xHxjC
4A5UoT4DNFHX/4IupuGaiL5sTcWI74moVBfljPfC9d+XGJTrQEPvSjwqZI6OKYXlMMe63NgnXA74
qZH4MybsMAgYaowkRR1gMbR7voBOtTX6DqlgJYlDfEJagFRTR0ycyBiujWq0O4w1d5jK5ew/gUs/
8ksTirQDomBIU6UyS5GjVWCsJkDjRdnDF1qLr4WQJSqTm2ax3Ok7hii1PM/u3iH2LOJkXQEnl3Ee
wxPrR0zv1GKKNGZqMhby91Pd0GjgOstIGnsnKKl8n/2ZoC7+KDlDnjIKba2tIqlVYt6TfmGDNg1t
RGyrhK3cVGx3+MJBH1wu5FknNpz/xQJJvh6a5iLiGPJZvFCYYNcJwHupuszdcdihPS+XL6T/xoBQ
SdVOw/hXLrhq4LqxxJsKrXymVIs0WEbdiTKbJcrpag5SteZ1x72KSeixG7ouU0TWkRoDAIyqsRQ3
2bVMOzqJro/7Nb+uok/WRt7Of9jzMIaUvDs4466J2tEq7YAzWb1TvzdU2brIIBCDe3be22CTtLq9
Kxii6R8ndWaZcumxlpzUKQYhDruXvRuwCYLuGOAIsyMN2qPx5Mpuc1+YzpZG4bv7m76p2bJyD9r+
/4u/b064wFCmc7a+U08CW3OKU+wf0zYOlIciM8DlnPlW6ZB2JM/WCf5e/5n+FoitSp2LmB33WoGw
/JCsLC1IHeZlfS6ibM0w3NnJrydTVoyYXwNhkzBnIMYg3vbEv7kw+cBmpFko0lxQ03z3nscutPq5
LwjwE23gd8wzVPxtEqWqpq69w8nn0w7A5Aqci/lEryGkehCbSaw6stwKndo0SoaSfvpF1QPKVi6I
6CrBSaHYDOJfx1hzkIC2n2og9aEuMEqZ/WHTQfc1vqtkaFv5Hg5DyxkI8AbVfMWZQSqfVXInV+WU
DjsD/2LZKzT4It5OI8MDjrLdbcS2867l/H2ubWiX5IXgbdQWNbh8mJBUu5ooVC+o96yPEO9Ju9O5
+x7HH5T6cQ67OMiw7g7rFly62utAxfZKvzkmFIlJ6ckjrBnlr1OC0QwnqxeTnQApMjgXTMJZSPA0
Nm+XpAt/bdqb1K+DNaM2HCycc6cR2fKstgUlgDEc8ydknoa5KpI0ObapS3iZq8WnV7HYE4O2oEwk
3IA29rE5rTdCTUeyFeJjH/MoaG0oe+7N7VyAj8xBfnj2vgmIMLsw3/LGWoFtQ5xLYTC7pCRn+LjA
Y3ZZ+h25JHmhDJYUi+IM1NUbp/TtjfGZRAfLiFBBR5y3fBr73AdlMPRLwUROqNbmRH8/gDQwfADl
9dx/l1jOCdFY3bbD8ipYigBhMJAOvROJL7bP9zxZShck2JZwChAi7AesE/F3g5XWUasf54Xfnm2P
DlThuouVf53VObBcuVwzPlIqSYlYRs7bw5L5u49XfyhyuuR8T5j7Uih+T4Zhc0frdZIdrbfFxGhc
fu+eOW2rroTy856z3AwDgCc7c4UT4GiQr3AxMLZ/bZDfa6L0LkKf/ulk+TJPIPz3NDMEQV1EbkSc
tEH/1E3CYjUt8O11H6PZ2qBB3Ax8tKL82pZhScHRFaqnk9/lxNVhyl/Bu32gpmYiCFd1EgJBGONk
k9Qoj8sCjpcr8ntitWO+DFE+2A//Vo3Vrq+G83ZkJHKTmDZYzGXhp7zN1KAbcc859cvXRPqdxepi
zh+RERlDl3zK/BPIXFPUhfm9w+f9uwE8cS7S8g5qttzhbxF7JNld3YX7BMusBbQw7qwposN7huzW
cQt8NEJOuaBnCfT1jdIuByxRTzTslDY/u8DMSW4m0RKvMP/+GA0AjsOT+R1vS1jvlYFzsyOqQ0d3
ubRUJ82PT/aLNxM14XQeqDnl9fLnmKTj+R873CVUlr4B+gOSe+KV2Kr58CMA4uqtWnM+DzWzvLS5
5sPMkRgg7d1s7ZYUTUtlBpbqBoFO/k9m7pDTcOpkXWviF6BuXBDLnR24IIfDLxC2ZjjCeGU4d9A0
b2LZjTgYU3iGnnV1dneCx0LejkzgWatk6WpGl+yeigoHm0U4z+W7lreHWfNB24eNG1gqYxMifw3C
UOCODCI3wtYeprtYqDZ9WdD9CQ0Gr9trUjdQgtHryqZmL4nO+A8Fu/UxNvHvn6smOJa2ZeuxaNzd
XSC2CIzZ9u/NmRt002DWW/xInlbzr9LUx90XPnlEm1A0aZQcPxprU3LeSWHbNgcWvJaN5aaj1de3
jP5GfksljTZVeFOFjfGr/C9ZhKSNWq5lHKp4JC2UzMbw0uAQDXm6ERnqCdp57KtwBFDfOnaDW1mU
JKSWeQf0YhT2aF2l2BoHNy5bJnW8t6pr639sa2oVr0Ib260bRaolpX2OfRKy07nK9i7+tkpL6zZj
IfkyUNHc/iXgnHh0/YzdZK1wkxeRb3C4hTtCh2P232R2XuscqUadZLgOspNpA3SeAgsHjFFYWDY0
ONPX3+VGoqlKs5MIwd3ViygGcJxlkE0F/jKPodYYNpDFSx1xHLFtDAfusSygIVClHgDtivOfve4P
bkNXRWLOh9J5TTX/oFdEvF4Ih1ApauX7bcDuTBHN7RWDnYEe7rlXVyNUouJeeoT09oF3DA/zDu7G
cigDkGAhjyO7OxfcfZ06qkKVP9/tiIVUI5sObS6YxVOC10ebUPTfKKGtd1o+T9Cw3c/HC4KxdBXU
EmXyiu/lrkaeHpibL2VJnjzHS8KpSNyUFnoy+SA08DPF/zVNTVvOSppr9S5gbm7sTgMWCMIdaOVb
98hkRE5XfnQJ20mEYKdnyRtWwnfCcPXMPuHJSqNMwr9nKSYlMSM9WDaYekGSuAXng0e7KBn2QkUy
wb9hf4k0+UFGIEuC63wSJR9vMLAznjl9lYr+D3eSKyatHfLUu8V30ILAhjt8pIwB/WV9I/2eU70X
gIeiKExa7gHAXidwuKxNjtFNZF1IEGDw/bNjttJ3sEg5/rXjO2DVPYNHg1kHl1L57CVxsLIIenxm
YlizVi1WuCsxQjoXA+ASYGMnwjA/uAZWHTjfMVz0lee8DxUNUFgt44CmGT9EYrUjwaG2IRe0ifMS
nXfJZxPH948raiXMnThWtOI+b+hBiev52QmLIqsWFr8uJ+4i+48Kzh8+6Qccw38czaNxWFLHTHmM
SD75RIVzSltA+B4JX0WIT792uykpmxk990L8mGMPAx3zm1zUMN66RoDTl3jo4AUN/unNUEhF7S/w
8zYAkdD1gWM2FNXW0vRetf+JTjRGZEOh2SlC0vjTy4T3K60pxz4Rb95mGdFRnIIdLRMVAVrQltSH
NykvMoJZ72iVPmoSuhm1eA8PnmYllGtWqcpQw5Vxn02Qa46xE3a6dxxXeufKjjvSMsZC60wBmwIy
HlBY8+5TBEGBQi3WLSwrgcPgAth3q4FpjkjCA1e8lJP9W4mO49IACtw/UxkXTRHrMh+AwejWPbNk
4/f+ajVUGWMGP8HG5Dau+ArzSPUyAJGPXznRB1TFNMKjnCUrOxxxK5ae9qFPeaRkXUx41mw7a7ds
XHmRj00g3P83MmsuephQg8mO/RY/EswuHRyYYsYL+pg2gzGFKolu7xVyUdVpK683HbB4ec4IMrje
8ubJlG0qPEXPuOqXXeEeDdtyMCY2Ys5Zk7etldWMQAgft+fWOPUV07BCWKR4n30Z4h0W/iqUpZf3
SfxAClinIa95bvW23FsYIug8sM3z7B3qWQCtwHUNQiRmiPbx0yKRGE8BbKYzY/FAdhO+RlHMW2xG
t7PJJZ4V0KD4jlaCvakoevEzi1Db5lBqQCZVrTbmstOharrmVF1vrXUc1gy+LLrtmJOyX0HPO5cX
7wWYYY4Y00Ju8wWeA9+80b3Jbr++GZSZVV46M3R0y5mokPDXTNxD39vJwbExK6cbSoGUE0jTIAEw
ff5lkn43EwLi2btafD0c1U+6FbdafnWwH5Wf8LAooOWH5eATONeZ3VigmJD/owEBHRBGGW6g8VN9
d6owr6RRtW5GYFTcUftkYWO/WA8gGfj/64op0vUdTB3pKKYRxS93qmNi1K9go+MjrxoOWNyTwvzI
/zHYovdOCpxpBNlofSqotS9v3a7gyQBrAyIhnPFqKwfIsxGHkM7Ddlz9fokMvrQdRyB4k50+m4/T
XGWpCLpZRTdPI8Qkh+XYEu3onDslsF9ajDC04KgqF7Hyvay0inzFpTTaAEpn7RYb1QxhaxKk/KYY
SoBmnb9zuqSuRvRE6rzrXPL8GQpR0jv1n7r+mr993Hd4PNeW6gv3nuRzfZ82J4hVZ3QW5pwaZeq5
/nd3ZhGfAfFhaUU6jiqaI1J0nkT1rxzk3sXo/9hwtkwcVMKYhb2aFF5hNEoaI9u4fxCwEFBqyyX4
j7wAZLugewfI92vWsN687p18gqiRtQoIn0ZwbnRWGD2FSj1IMDkqLDmOIZAJ4Pygs9bs5j/vR3tB
qrZGp0enIsMqPAwsL+k+1817dD5fVu+feSZW60dJZVtNtquXxIK1DWVERSMl1J28VMWFCQvg7Tac
GdIRjbwgSHI5o8qYD6FQ3hnhetJ4gVlgxcyea5RFd7Ulu53LO7iw7793RsKB6/gGvX/635MqMIgX
5IRRRiIwe2eWiMg+MU1xdEtSWMQwr/gMLL1PeBshp6L+CMXDTg2Xcg8tkssYob2/jyD8BLQpBeV4
bKHfO8mDssTmDcG260lQblqUMOlHGtTJK7df5mYiQOxrlVP81ZuckyAho1rF3outrs164WPjZ9ni
0MejwHSs6FrAIa94y9w8zl3awcnI5aYD03TjZ/ji4gDjf6WS9eXPHYZjHoGkidNGLndgMfIuZvqv
+Str0ltjHebO/opcv1Aqk8wGzQ6xMBDVs5blelcXkm0eK5NI3RAUC8WP3BP0Qux+RFVaSyagiS8b
2GbwadqtpI8ABlj/fMj+LMsUOxadTrqbu54/F2w9YwSAabOrHUuWyN/Ze2ONIrmSvzmApOIBMW3p
TdLGj2WeJCVJH7OiHESoSspKJ0QTNkW+UNouVzovFIAjceQhx9Pb1fv8aypuOFNmizzG8y+AjHcb
lGh56RAECAD9z6tgGGSm5MTGfhTk2Kz0UXujzdqQYXUfwtWILddMO14e2SeanpENglVktSgAsdpH
5EC8ZDJOaPSUUP9I23o4VqaocyOogBxLAHffMehXcBaDWEIwQjHBi3T5TQu8h9CltFFbvWRRfLvs
jhO90wWxM0CmEefg7jlGGH/XiJQxXeBVhQz37MulNj+CUhwXwND5FgKzyZeglBcgjCO6fSUX4YXa
UthMUEkLTNzvSPkZzq1bIrgKX+F11x6jQH/PyBybWPFzSLOW2nXvXybqrC/J9UgjqJucC0kEEbKf
6DL0dyAjCCoGQx/2g1yJHuiYO6iwcbCEhllQUO+n6fUbWkqaXl6yv466hpXKGvace1CjtAKz42dF
9JeJqgoHF0Z0gQBxlRQf3bevBzwxPkO4tD5N71rqg3WHMV4vT6pbaiB0l2wjxw2BOp+Eoqxg3cXZ
aLGixuEBvYmnjtG38XXPY5qs5WxrrQ2uY9j20Ek0eukuI93esTW6/NOz4UW/zpIrxEVf/69z8pmX
MRUKyjV/Ks1fMqhhfjFe0jMepfOQdh+Rjr1bNBQyTwddDYxxR0d5Zreigh4aztHHUTHOlvHkqM1W
yvwlgvMh0cQ4YhmLV60WwPY+iaxrXf+mMAum7q9ifCM6ElI8OtYoSWo+UsoWfMMpSP9TOwazIHTH
sBFu5wZfrVqh0EglvzBzXBlAop2Tcvt1c3Cwe9Z1EiBj42lLXOABVgphVA7wWGaH5MUIy9GpgWvp
ZDEgYlx6NBKJUD6fNtIikB2QnVHTD/YOG/rTFMYJ/3dE05tOD5mdv+D4omyAPqi2XBscviTgLX7R
wUxFB0eRS5n1ANYhReTzv18/h02UWIuuZLgPKURlSCgupvYgs7f54P71JH5Dhiqb4HiiIOzQ0fAc
Nb2BXF6TKCZPPZpf7vhvzcENomOYNh/lX2lRmNhYUKwwgwkSLcA24OvHALnIayicx+DdC62CXWra
sBjc2AIMlvUn3StJoR5sAqMaFS8vwu7lCZ0LdhHRROYjOS4KH/vHEJuXeC/zG4bZtB6SCq1T6CdR
R9hNxYKH/4SVObLqgR7LKoJ79Ivff1nRkOTDI4ihHwCEB/FJAaIUvE598rO2i1GQzfU2Z3NT//ZV
Q/w7JrX0yNBlvNjBOWE7mNor0qfHnAggcc3GhWK395WGi+jKyJUSAP1JXI+BtY6X2hyMzEB9622h
Mo0QPeJe3nSO2+MmJX+mczeCykz6JwyGeL7UjgWCbNY55CBgJ922G8N57GyepX0e/RjLP6DC5cUL
CwaizuTBO8wYpiRg6456aVQSaTZ/DELT2g+O/6UIZKC69IQZbptLEuVJJmIhwls4QnDn7BoQTM0+
Fpi6kjJ47eWXEpolk/P9SCrrOnc6muAJdKYssY0X6JUwgqNWffuC5i11jhjOLWIysqHoPUBtA2lC
rdDHossh2yzgMzvHxIkiBkoYp1n7NzQlTEDloB6f5dqlBomh28PWh3sJm86wxq3Yx5bn6zZG5SgO
DESB2vH17fg5b7V2i6wpk7lsTraE8AbMVNkXoaONBCHYcP+8XUbUf0oUENJ0vQnuoSBw1SQeRSz8
+JqbLouLC/jxE0/2h4NSb9LgnzPCm7UTwmKRiAengONVIqLERjbqBSK9lKieWPSaJFtqT75KpI/i
oUmpP6UxFeQGNou0DidhODHe46FaoxLkwfjMSZcA0CAiJt1MM6ROrOSQ+N/tKrzy/YcWgXrqmpji
SYRm+feUwipzCy4c04pEDh9ol7j5BiHxivton4k7QY0NFQS7vHPJMCwqFmJFpMp5dlcjrTw15KOm
dPo5/0K6/bxrKgHErpusDA7AQ5j5hp3elEMzpsIuKl6TfBbNear7lEKR+l+lhNViO2xoY4GbkPKo
OEbo9sbX2zoiUNG/CMRUYm2EmQi7iF1pVHtKuvQAiBuAHI8/ObpazVED7XWPZ1UXNjtaMTkU0jyO
YqKY3zqAAzQE/3xIbrf9ZNwiPGSzjV8qmTBBdjZ/57M0o+7NX1L9mmYRsMCTKN7E2e9GJDySfC/r
CXuipuaaE29WkIiU+SlpnqiTiUJhrvM+uoRCs9W9zXlMOP8ISEE0bq55X0XZZ2k0KvdBf9+0ZFh8
TC5nXm1KQOkwJd+jYL47OH/sm0VKSE84/+94wRpPfd7Rc1kovi0YuU/DqsAsVLx1mjTQPchv2Aqa
HY8uHAnAvSmJVFLRw4EIj4gba0WStTrFKrCMaIf9K1bCwQcMTpx5d6kNAW03Y67A8lOElcjgJeUb
Wd0rY4O0cSmR35nATXMJat7TYSyiYSBh0lJrBoFyq0iJMeBUU2cwnq+MdLRlneAeq7+DPTx/UjOh
yGDKfHgeVtVp8BWHATujMkh2ILh5ZYIBo0Krfm6P0PnaWmbtt6VA2xHAUb7HDCi+Dvt5s+updp/v
3j7UdKudsv7X+sFkVF6VY8XrRDJdjxQgcRN/P7Lx9qa3zlbjQotD8WxsmcPVpC/fjfzDcKfMXqN2
7BjUx893atM3AMiTYX7GSBM84nxraTXhxfqMP9T2QaSwamZWFTBfvBSN+ElNXl8THYedELFJQnOI
VUq2xobIDF9Ag2bnXg8x4Xa9+E8ypdXkJiudw/cggsSzTnoN+jQPiSAwXA4q5wf7Q03heZxBdvME
j2VfdlYg26eMFGtRwwWqtaUoE9R8EzVVr6eJsYN7VHLDhNPbh4DPyPwqZ6OxEJvln7GawseqS5RR
23VxKd/r61kObEc+lulfDlDF6A0oRd1jxT1cTjq9jKEhuiNLM9y119+vaYbSa4u0XoP7mUj6KQpE
+EIP3nfeCjBOmh9y1XbBfillWPo6BJayoLdXmFe44wkI4kOiH62kNZuKmHQ7xMqQP7KlV3vFg/lN
AYwFsvok8I+vZHwK+1fw6mzG9xjYQ5TectocrrcR3tbGjcsvi0hdd6vv1KGlNalidLLyBuy2jHw2
mib3Xu1CbOi1Ask9HZdHMDbUov5J8C/fs7kt7CKi6L4yfibqxJuZPANPNTbgPUJQyeJzmL0A3Pk1
K11lPshj0xvQkhIC5hPM33ncGyojl49Ii/VO097X8W6fyQ97jmLc0eLK3gHpu0otEsCeyH2p+AKf
efeYor8uVbLOTFZxSWAPsWBk/UpQsaA8fvnmqVJCW7crbduwZziknKI2WoSCtgmfaIr2/cLt6ssM
Gql7YwYTTRsnyZldQAgc8A1QM54vlOt1bijClzajAjWb/oL6R1ZkV5ff6qgAjA7vq/yfJXTN0DZO
RCxlDX8XVVvQCRmbQNPsqJF+3mETEZSqSguI9jmPSp6Eqag4U60BtWTnHn2uyf96u1vwis9m//DH
BL6grjTCza1CHDCIUvQJSq12ZxGgMxfNfPDeFlEDxT8lTOFTV/2Yh1T37ybxZwlxWc8zJUQGoRUc
n1xu26jduqUV5KMV/61cJr6G10o0XHy2hiFbrGQt1MAvMMyQ40ti16YfpuBI4EP6fJUsfS/U0AYG
K+u+Rf94sHkK5xEeh3LsJR1wspv11a6dTuT0s2zNzjz5019Jkpn4TSmccOkvCvErOfdNGO005B1u
YpuoJmFTAVLcqsedjbiVAIPwl+cK7Np6BngVCuL9pcEtTYnlp43LgyUWj3bPZ794LgzS8/IMpP3g
aSZWgt+m1sxapZ18AumwxQdy5uCZuPupyfeMC0lIWZTXU2PHM0cw/Usnp1YOup+s/Q1XA2TJgZcK
dHu8gtsAxuThtkWyYQKld+TCdLMK97DVavImneWOcV0EDj6oE0PtPGdKev3oPvKLpXWmVq6phGki
hbjT2K7yubCXc/u5VNtxe/bHWidpwEl7myYZk8shS0vnGK616kzVnDl6vViBNyWt4dKkUJZTy2eM
GvEozEG2RwOjM4pb+iGxjKfVUpPDmO7bmaNVQkryHqAcYSBl1b33ca9bJ0dS8Set25w0O6pzmtyl
NX2SgPyDuJa0/yMZwXGy8WuGL6Bu9tAC/8RfpcG4o6bGIp3MmnDRbjnVa2BLiom2o9aPk1enx8fU
6VM+lyb1FxeMZpYQHWAln5FF1euHJkp1S7Eq02HLjgFsB10NTka5dUHIZDAt6fq4G6jsQEi7geUi
QZY/rp5fs7tKdf/XosbfbH0G4RsrBnkPEvJf1t/3UQ0qUEv3Ten2QtuIYdmckGCjOWbugclCMDZ5
M5XnYuXZd29esiOYgpU2nX+BXdlOHBdkyj+Ry4UMh+2xBB6Fv3wgH2rQ5eMNlV/8/OUX18mpyNlZ
9pC3yfaDHWRyNWUP2fjeGPrxrC59OY5eYcFkzVFVSIio5JcQe0GaxS1q3XADclxyAKsZCqV/zNcy
9YXlv5m1xqHffA2gDiTA0kahQIyN4JGScCvyWO7tkPQz3E6EhbtXPZmZeOPdXIF3gOOlgF2mfNYv
DakAvZXXuY9iZ4QNX17gXxdO7hVOtSP3JzQImtxpp0OhE6GfgEFsouU1vuwkWB3BcnEWIYfEa75z
m3gmA0FsplARV8wevMFgFveIPrvsQoXREvxC0zL80UQzgHdlMfPGjg/P1Y4tJyOKj1VxNdkws9Yi
4d9W9O5Rkgvbc5BR2nuUhEoumc4hkY8zvb87EDY+djRDGguvLdzS5ZS0fmHFvVmnoWqY+2ojZT+e
LxKHCLwcZJr51iOpa6l/XP5BWU6gfSoiwK3lE7LIIp/ePVIesG9vGUXRHJIQ6Wa/iLYSg3d8FESL
0wf+orIfX8lxsDTrzvAigUyMWx0w8S8mlqrZ5FMfq8pg0GtCAnSeEvkn27BPKd+m1J80GYdKVnGt
ebQ/lsiC2GKk2QPbUgk3cE/kPe1/OC7nDnawhLp1NgBZqMWU9CBW/ZLs4ZqEq6DKhOLG8n6g4qF4
jakLZ6sEZRnV7IL9OZLRJ3ZkZ0tEuUL/MRK69QIzlxpjypQ4s2WiTohKLzlnJqz/fpxFIZ2EM0b5
z2wWPiI/ftx1SY7AiipE9XWfJqGEiCXlGtdxd0KRQ4tQ84GMxX1cYihNrHPQSC8/FsQd2WAopZso
bv8DuL2MCNXCRnw8rEj9CDlygSafszfVKuMjsrVD3B18fDfiQpfKhHuoPELC7tIbqjsTO7u+35xp
YsomSqM+Y62tkRfsv4KyN3MMG4B9AYxAEIzviN8yylQq2E0OypQ7bvOjUfaMWiUqLAUwbhXEvi/D
SoRBSNsosIshwaxn5xGNsk2Heu2itdimyROQhi6XN+N2SRrKo7pgqp2uqlRhcIBUi3xTCHGmvanA
cbCqfNiW551aMKF58Zhg0ciC/+ut0i72UXyqbrX6JNoJlLTcwSDZ8krcDf/daONFf2pu+COef/xj
7BhwmF/fzGYIZFak2A5msa0ayHl8TRp6/NzW2D+3wgGebRjF2nl+kEwimkTItX5u0FhzbPbZpw53
kdqN7SW26sHBRqbFPTuu9iY1344m3Bw2Nnz69zzz4xtEvF089l9ZS96xw7ChreJbxfUvrS5XG1Xf
KADCClTXwHDYOhB5neIqN6z0MmBO36B/ktj1PrQsUJr3fZfhJ1TrLPpeEVjU514cGfJnun+sOlMN
TIivRrhHr+EDn+7evgSyCJf1Jq+yNpNyvarxq8ebSYy5SREeohyOVtiaKkm0ckHFWJdhhphVAXrr
vOh5ruKJ2yeE1VCodiNnWfB4iOIvbuumtIsSbZX5jPO5iC17JgEten/Ob7hrmgxYtuhgESLlUZZP
oJX+vmOYfA/GyjCCL24MZXovnS+3h5zS5pINkAoKW4qFA9ZGTK1DwgrKAtW0+CDMXBlLAwa2xMvN
0MWPlEWKjhhJjGEJCkk/sIsbBXYeIFx0Eyn72wcnNBkiWX5tXNjdh1Po6WTrCDEozpXA/94aXM1j
UcTuv2fEC1aWEYnIy4jcjH/oIlSd6RQ06V7baefork/juakbMk71aqa3CGTBHmhU1XGBbqM9xaqp
xFA50m5B4haH7Lg35hBYwLvPtEV3rVS7JaiYjvAQFW9iJ4OQXrhc2+y8G6A5r8xBcsv9hUoMEIIa
HAHQG88KUoi0alSHsa3vgztthA/aNfyBiB5g9LneGuOGDRMLOTP5SKERQfW2wzXwBO02xdj6R6hB
PQuZQwn8+hNq8DK81a2QqjXM5kwFRsVwpwt0SO7gXKG4TZ3vSnV8Vh8tJhCA32llhwZfk5inuqAL
kk8ycO9zwVR5nrJ9yGNFcm+7z/L+a1+tjhS8wB464g8X6IY1b7nY/KM8nrTdfZ+wdCpKC4Yk0L9n
+xc9NLTHT1XipGoJhLbW/lhJUHhnZg1uSp4dhjDOr0f/wISmvfpRhpnHr2u2B4fQlO8BBrEoSOgB
l5wMBQbD5cOiXypSdfGhh3R5RgI+1UgKPMVOAO2UzqTmPRwyyqX4S6gkk5XChVOdEqA/P6SED7yt
K/mk4taWOcfW7mF+nqM09xeQoE1b2unkgEpb68elo7V8KxXmOLXP3M6KKRp6nOAxQ5VrEG/lp2dJ
PsVpCtdWHYadim8kEV58996ARYuV+U1Rt1s5H0p3Je/n/AsD0DYcdAK1uo+/YN5atF58LPSv71Yc
tAlvefzrhL2JcjrNr4YcqD4vBUEgh88oaKXxJrI4mrlYHdgcSSlxuYe9gv6SEHCbP2pZ1YJ4EdBu
ZSbwyhyC6tRGbUgLGQ/NDJx8yXVJHLQUOnrjxS2BZamhLJAVAqI/9qegKbS348wPuawLVap4TR82
4vGJCAgdwze7BG8aH3rWteuC64Yv1lSEFJCR2Upp3vrQmUkcnKfIfjYf9/aDTGEVc49HwZKL5Ddl
UdsrRNPIBr4i3eBNRPOtm2VMEdkRtFznDrETtuNYiOXUpUkKr+A3nS3VHC2bbBUJR9B7dFFqHLA6
Vnzyo/Aq58gzuE1SfmRETuVagiWDOZN2lnvoKMKlmETDjXeHkiYvH2uEb2+nWNgw3WBeNgvJxEIZ
zTBPddMzEUjI6pbME7+tKg9GJawl4m8xFCW9Oc1kbSToYqbvVeP+WAH3ts52XxuAY/BW7yHs9hsE
KcZ1QxnbXaZ3o7/UXUnBe4TJtIDUKJjnFbE80pHfJDFB5bH4jSb5Ak8c9HVMnGNz2x4urv+fF9Sd
HyKvcJznLyafSWtacsZnLL/SCU5/bx12zORHzACtedyrmDHFFYtRb8B3EOHovpSHJ2ELajWuAxWL
3zt6CaUFgo+IAvw8VxLMJzzoQ6rngkG3PrGUaFSrXasEjLAO+EZ+WeBRgEjE0R/Y7XTjPAjCUtlm
NOQYJzfKMjbFfXabCt1Kw9ixXwYNek7NC3OvA7coXfe21A7OvoWV3Ie+1I1AwjLc5RA70A1rZfvW
pFnCaXbWlTYfuIrhpJ5uvNDkfld477rtKE6g59xR2JHHh+lwFjgYf3J0M3IV1NpGzVVFNdA3X1h9
QhDHw0jFOHEEB9yXKeuoxlUJH1nted/WwHQxzcVly7pQpV+3pMXC6rpT+MJYd2DP9+nk2x+LAbAm
0k8Z/GznPsy9EN32s8Thfo+F01rvGmpIvBBjYq5BHBb1CVzDNKIfVBp3SSppviKMkK02Sy+jalPK
Uyl6bLZNIDreyUkSEU9undXmiRlC4l8OSbwUxZgFBaFe+j4R4giU4OKYYpVA163CGN48S/uRSzr+
+btnQRlsPAHrb67/01DgJm9w+09r+bp7d5AEXoswcJXrtrMhKbf3/2vyb7gNRyWoZ7XVIr51rTjk
YpUt1sWwDrHqGXbiSeXVRgppDYDcCitw4Yt4RnxOaN1Nx8lMSwuobfT6Z0jXSzcV/vsH/hnwCLmV
HYblhaEMhLRpry6G/ov64nJnA6gJpBaZwFUT4fFYrX5ExZZ6H1hT9fFiAWoO2FG5eFpGJcywLjN6
bVWEvIZkqAzV8sI7GxTC2QSSdvImaYcMsIm/N4SOwbz8c3SZRpjZ/X+B2Q0rWbRDndaRKS0ivz2J
8DVeWHa1Kx2fQlj3s0DPyRKKNS1/ZCdGRwhmEiFQ6CdSJV0sr9WkAwelTaPbJMXNjXozl2PIyX+x
SUdF6U53uKlMbii0tZDpy8NalGN2H2Mzisagx8FxYalCnpHivCplB+LkwDLjQqJUHS1Q3nW5q3la
yVSImp8U6YZ05M71mnbLVsNpQmvTiriHrGM1UPLFngFydVKLe9Qb/v+RfW/fes14Fnj+jhUYjiQm
WtvYhWzDd/603EV8sRF6lZRkyfU+UrIADsrINiL7sO7p4BqdACNRS8Kdlo+5+cbxRPUyy6XgU2Mz
igJH05619e/E2GLyGUEMq3R5s6ADd6XBJeOAWcT+/65BQtvYTPFMNunsaqvQwZSiyAPNjVNKCZJI
/ELjtkk/rlZVzqnSQZq79CwBRi9G622R6nz8FtBu5oF3Ue5z/ukPNKT2miZmnxWhSNgG5IJ8VUAv
BUJ/dQgJeym/gN6eNdYvwxOVK1jzEEDBQg5wpn5JdTURHY7/aWuJWvjaBaDeKCPaAhWjcD+p3Yxh
xhbXAT6dfYeU8oFvFAGIOtWOZov1/0lotgMm2gCq8suc82ZxNxzM7nJV1w3tKWjp+M8NdIx7jDoF
MEKcBrrAj+gCJivq6Nn5LfJMthMr6AdcLozJRE0N/DwdQagF9OL3PwuQ2qe5eOo24y4oY54lZuAD
NcUGmSIhYRJaJb7YO3KyapvpVFDOivxZ3atQztyYstgAU2xCwriR9GvQzzExu3+SwORcWQjfJ6jn
VuGoSTi4HkVMFF0d7oBUhmPWdoxqym/dX80MiC/m8bh0c6/YM+liJlzNF8M4BNLlrkrz5dzvRIwu
bHO9t5glkZz3v93qlTOEkaOCxk92WDFO3WS5qa0plJaTilcjtjHtEpvpPcQm3ESbE2qoyezM2LJM
2uGRVJSDTUBtRPZsQVVR1csguzht0dc9UFHcxWMLh6eWB7oe1fHx2GBQA+sCpKrvXzIHh4qJPV63
CjdzLzOeH4IYvRcwSub3VKelQlljHpvdyNNsAPPi8pz3qySMcL+LVQHXDYDDWbhDc9QQiPFmbV4f
4ZnViSNcigf7jXC4A5kD4XCiyKbBTFBb062KQxs9SnbSay37DA7IQME3KYFdOmEOvqYZt3YO76xs
BVz2/aJlIzltGw0ZNWfrhfNnRSEMOtcJ5yErpmyYdoIitJQ5e5JKUA0ytrrUQgFVhd5dnXMUtZ0Q
w8a1r82A8Xhb4HSOGsSAlpxQvv+8gyd9NvYvkhFwAJrgdq4+mR3ghcjdsLzEI3ahnV6bYYOBjaMa
XlwIM9JpqpymrrQQ/5unAQy98jKGFPNtq16FgDLiL97UabQ48u0f+fXkxExJYARcRvIRcCtAgG17
szgd/SholASmHA4PPYm2AyKWZRDjijhIR4zq6aAuvq91Z6MjyNosLw6fuPypesaH8vRXazqcwlG5
CiUvbZwlgi+quPYt2u9tXsKf4KjCi+B3kJz5KxGdtEFpukMKKIANi1/mUiLntmV1SqJe2piryzrx
DSoEy0kHcqkfHlb1OG+/u5hq1kk/WJy65Z/GVkhZfUsKrTiWm+ukBvQeAp93Du30Dt8gso2fWl7Y
G4PnKbPvet1LjJFPYIEHuQAnzVgY/e7IgWSsPk2hBbWQnN4pAFViDYcH5D//CFxAhq2eCKEEslVD
zJve02BE2K5xExrYA0Kuz1tU+RuQJco9G9+qw0j+IJGIWdTtEtMoKFYhrMcO+epmmTRUhZuP7DUS
pZwlmvBAzPbpE4qLwG7Mt8LOPOjt994rBxXWKcITGI7GkFtc6/y8FQwghrtC33fjlFOqTou2e9cA
HCj6AzkwvbLjJQnxmPVKLXlccRpW6LjrGwsfEBoJZZwkd5zrj+t9HOlUMDTNRoI4RoREcGHMUY5m
22Pk/aAduCIDNkRlWXK6AyYzDhWYYxhhgxFfXHROqtWLVB5A7EttdIw/l4gdFXmG41TqLjueGGZm
VQmt1p/wM5OMakfX06LHv4yt68OlVTl2mAtObuZyDfysS7syyvqDODD+auweQ2KaCCb/mGF78/AY
+VvCX4eDbYQhZ8IAEEqMUIK2jVMuWZ2GPBWRBRDl5D2oDw8bfPzstNkPkkDvKGCine2jkB8u9ZBY
BgdzkOYezt4lE+LKHiy/1Q7boHs07AZzdYbalChEYLi3LRUFtFBi17/jaAPMijYyEqOMxB5ZJL1D
0YUAFVYlcuXOV/w4Bbi7ybZmRQ59r94biL5N/IcTj4BbLCVQgUgQ8tKVImJAB1ZSbD1p28fw4QAR
r2Ih4vB2NiIOpvjquXu0rfUGQT/MTlQcFKE7I8HYfG6so3NavcoNBJjGQ6VR0OWUdb2Zjki7iDG5
BrAmx7EZvjLMvMKUUz7a4Rx0bX0vSMjhkkcwAaOK35mI5yPg22BUOPaQGeXbBlkDgsXIYiPVLtne
kVcHMlh6xgir1k7TiDZrWWqvLmcZzown+zcErIzRJ8VJ6prKj3pMM3ayQKsb0Kk/7XvIpzSl+w6J
0fmbxXmI3SwOCmwTGn4Gv6SQRaY2hKZ/sRxEKYUDqMZ3//QU1mOU6tUTHnEl3nzhg2OnWDUVRe+Z
zSatay5X8kD8+bgA/z3Qg9KojlAT9vjwXQRhNzAL6sHbeH85K7Xh1uqH/4E62kZz8N8XuVPpQyaz
fZHvFq92idY/Lz/AltHXPE7XDW0o9SMFXoQuQeHFChb+75Xtnim/gCjg31e/LZubPV183H2LhFvi
G3gY9wDE77itKJWmtWy987PFjKruO7SIveDG4PJiWRyi8955H0m+XkNtzWFanRNHELvzMaK6CpCx
MLl9gM8KvK6WzktqBepcCbC9jzoH1leSWG325B7n2Au+UZoqEn7biFnrijnw4N1XWR9CkU5qo2gJ
ReLMoRPhAm6mC/gNSAeN1sz2qRFBRjFpTnHScD4mG3CbtSfqUIhVCrpQOA5Ip8V63VoWQqgD3wyj
JlWwY4QuAIlRHTBv6ufvwB0iZWwFXKTKn0y2V60ZbSgVGE90LwhEDRNN1+cemZZKNHB+LFtbO6Z2
0JSdUVahzUwjvGAmyh9wFBQJLqplAyTVjyp8zEZQGBFJh6EkBzRia9a8hCy6UlerG7VMCIEGOmz5
efkK7/+McJRyg/Bq4hI8NLzLHob43B8CIb9Fht9XCwPfwALwYV0MscaLsm6qW9XT3okT0b5NvWf4
39uPEUO5ULW2stM0XGDR6eXoF+v2ke2V9noY3NzzNwJOEXHvQiFxa7B+MNjIVsj1Dy56+1iYj8kO
In4v7/CQNWSDVfU6Bhoqe5ENoJGzza3eGNaJXydkrrgvhNAVgQraiX50zpKcZ7EZIQqDTWC9YRwS
OGsTf0I9fYmzqnFP3C7KO4LdqH+xpuBjmMOVnOk906XAYGjVQ5Zht4CLNgSgnOKV7hl92RhbVqy8
Cit9QZvP565hgcYfM9I7zd5A4pe+N1jj1juBthVygcMlHGCbUuz+lSiNFUnP3yg61IKc7WDjpNru
lb+s5UkzrjAUnGAPKYZrv7IhKnaFDdCYi0+ctH6Yhguw9ed405I5mCKkKgSBk9ZZqQRIXx3ZHZrK
HC3f8dxIhGBUUBdatuCkcqJrFcg3ndlVQ0gd5nqUnDYRfhwX69liUZnuY+A20zcI3NsOWFIqpzRN
IkvtgHxsnGuppQB/DMAzQaJn0fsAV9uHW7VIlSQ8+/SNcdRpuDUudfAtFQPvU3wiZgPE09q2tfON
u7SAi8tppJeG/cl595yWUE5WmNfKK5CGwvpAhjBSh3Eij1mzwHKQmBvpVadpI+ksMzo1HZkiOTZZ
i4BKpbbZAKFRj9RvYjgtlbBiAV6RbmmeI8CiCs+K4sIJZIri4Dtfu5SXqN5SP5BNuI4tIuJJ8LEG
Q0F2gPEpOk3ohnGHe710t0077dGRYcDukIY6w9pBf1KEET4vuXB1VCKRWYIraq6H2cDzFbM9tta0
XnXt/x9EpFTjRYmDGzJkK+YSRPRr4Gxpb2+BTx3DudOJ6kAdLupdUm0o04aXgPDm5ZpXfb+aFYiT
eE2UXKjJmsyhbhLJZmnM0I+kE5q0H8pKc7mubfuTLEvi9CVnZuswnU8sQgahoPyvOjKmUCc8JvKx
iJRQnwYYUK0Hmd8BYbQI43bI7Rwr9MFypCjxLz4o47mYLDX3k+zyIvYWz0lOq+psdbSUKhFB3Bmn
LRYr7S8bTOc4ZFnEpYqdijmiRuQGR4XBX6DNzsrjKdLgnLhxpH0JaoTu1Wc/RMrzW9/FPu8MXLL8
+cnrY6D/npnzPQD4CGaPWuHjBAD74oIBnCdn+/b7sf60kGOvSS25k051JPfMxgrDbkk3CwVYJK1G
rpVUBBtql7qt3SaNgsUV3XzBl7rTh3QwWjkuRSCGWDmtkShNKS43SawYuxrw8e0HjSq0L1ay4Tup
ldmEGrvvT1tGUvP2cLismhqOYytHrXvEWBNbj1fm2VhMIdThgR/7pWf+QD2x+omk3qgMxeTL1vHB
S0neGBRXg/DmQxpasBpTzL94dJ+cVS0GE9SlYcXkcx2h32ScfxRlFWyCF/4TBhaJjBh9+KfN6mBw
JNLpFiLSXIpfvsEtW1OVLQpxx8i9stSd14GwVEgfxzzGmtl/U/Nhw+w55E+ni/LnpoXiRTFKl8hK
GO3yPEEyXfrUXLaq+BSFUEtCFtGkf/d0PnrGFcZOPd1pVMInoL3N7ezt/4C3XNPtJvDacYbfO0AT
g9Hv9aSon8WdtTvmzuOX80JSVduxB85wlAY3+iolynr5e/8PspC7Wn3GpkW9B7JAK3AtrcZ4V7yV
zkdc7eHjQIBU1O103XXQOjFqXeddwQHdQrgFRopFG+AagzbwdP6JxB8ZOinCNVG8gOvZ4t+5JaRL
/Ql9nrhx/7cNgpe1dpH0g2zIcWKjQMc6qHM+ECxTTz1B5UAM29nZ10lr4r7QROmMknaIjjAN+Il3
VKybxBA4HUML5DxgGC0Jzw/i0Cm9WPuH22/0GxQLZtN7SSa01IX751WIjq4pvY8eUMVE85uOxTw8
DOM/me1CMMmyW38C4rLhIWyrf1HNKZMxLlnDh8fqjO1zn97aeqVi8eknetFL6NKtT28yaVdxesRa
pWXnAjFQWde7soQWPXQXTNJ/SFEOrU8hjyXyYYr2pGzuVa1ijufro4GS8duhvxPQ3xeG2OK/eYHM
AwgxO4EMmW2tq9vc+xkqJZSGE4Lfk2Mcm0Iq7ZtdkpVtx2pB3ZxDEElFu266ZhN/8ykwWT8LeN0a
FfqC5uWlEFfRxD1Ns/pmCxgJ2iehfQQcsEf2qZidgaYGNIorIDk2BU1zsj5iePdV/uHA4BtCi8YX
Kw/S/0orAv/Tf3gjezJg6B4TTIYFu0raOvLFI5dgtCXmhjDnGJqi7uvDLcKXimge0zgx5F/SlwUX
Bt0UGgOOCOuDWuXeFzC9x4jw2HRRaNQU+xw/jxPai3YRvXz+E9HIlHt0rpKsmWp4cU09IwF/GHEA
HdM07xnoxEm0qJFuR4fHX5d4prQ5WZtXhF5+8lmwzCg+2pjIc1QSCr1wqrd+KrEuR4kQTHQkr+Ab
5VWqSgS4MRwF9RkZiEYewpchBv7ad3jL4KeOqlpgm/38hAkep6MIIxROOVWnBv5kmUMz75SoW1e8
ebyvp/4ho6wllSuN1nwnCnAZbZb+pHqUJW3xMhtRYpDccaL9lJfl9jor7YQ612IToDC/O2r16rce
SQeS/20rrVRkQIH71lOAPUBX7Xp1Plgxm7qO17dCvxBe5k9H776lHL0SD76wTiiZeiVrA3lJW0jz
9xMpNUEx0WOYpufgKU5WgPf4jevtIFi0RkUMq5atVGeaYq+nMSY57VsMmLTyl+CHd0lNWp4abJJQ
+1RsWjSsyQ+MDuONAuGrdfhFtx0+OkCvwcMDC3nWrez20V1ISsi/phpzULo4pZG0HzsKaAfDdm/3
fgCZMy8unEm8uipRzW5ddqwAJviQdtmtyebi5BUcZzAYJzndNovCpAlGroelfjBdvRnjmdsdNpVa
7PXG/rfE+phI+gP+l/vUeiNqEAvbtXdSYuHKBD4dzONbBvvC7PcJ7jTW7nkvDE9SkSN+Dh73RMur
1rZ6v80Ca3yy19UZlJP1MGQUdHLqJEdGHTXQ2BtmcQXqw1JuxMtfV0aU5UMrroHWSb2rlvoSLxR6
RXYw/qDpKRjphnQi0U6oqt6eT9FCpfH43ArAeSCy59E54TD27rXBByFjm3A2sAD2e2B48c+K873X
O6dh5iKaBdcMytmLYWmRmk8cnV3f9wLo5wR5a/H95IepweI4TwRZh0gEQaCFGzZTp+Hm3mqO8Gp3
BvCv2hvnYOICmr3Cmy50PwZDG05gEA9VJIgkF6pjMU5ZhNRtCSjn86fuqmHWJ9qbZOze4JybHFtS
+HAMcluNUEpdtwx0ai6JgDuVOD0FmLSTM+ahbf+Q8dfb4Qi1LaoRJKLXpi9qrddtiG0VabgZft7o
h7ePMVOKD+a1w3TmHdwOI7X3SCi3tElIAkPb4UvU/tUMMQNRwKQXqimIoxxzt4myRKWeOSOtaHMX
KE97VUoYVisM0JGCF2YA1tUxNnzhhCpgOfIAQL62RWu1h6EkMn/vIFq70THbSpXPiXnrEdwIjIKW
u8CcU/7IjakFlL8x1dwD/Cn3AvpFF2Agj5N6sDsuqlqMZVf2X5iTmIiVdZWzLk8F5aI7dC9bdAsw
z9xbqxxhQ3fWHScGjKMBDknMdCNZ/zVVFjgn14bQ251Tt7JtHDY60y2ijo0eqGHN3sQtLpgeWcJt
o6DQ76vxORu3PpjDcXPQGgpKA31hwmVbx70zMINMWNSrik6cDmv7TyKG22mt/IKYnN6fRBqyYKe5
BuD8VF3+nFCwDxz5eBipClIFT2VswwtiuBMc7qPx7YFNI5UJcTR9s/JOQN+wgg3r6pNA+ltg9kd1
GLHXT1+xQ7JCXbKJqC/CDUG+wA9Jc3/WNQYeqdfUlpmW2fXwifU0Yz8dIlFn58Yq/arPNCdADSKL
f5iOBOpMLFRxp6ofFJurbAzlep8GE6/nMPwskrXRiIa+zEuU8rMCxDbyKzGcjwek0LHWGl+PamCH
FG2Dge7bkO2HimknLceueT1ms9A07W4ImKmMSV1tI0vRWdx4nY4uXljoWWwLaXxN9A5+LQi0Fini
Wd4W5s8yk5nVXxUcsubPEaHpMQFeRqu/DPVmj4SvdtKEobA7ZuumsbyHbbt/FVO4umOEaWTRlEDD
0iSwbZ7/fqu1qgZEi/Ys5SynGYLcGTK7f71sF5/W/lv4q8hI7vHZFhTRXI5gFCIpW0JuMtJ5El1Y
UY30zHslvYk5xOpQmgmpFiFSC+XRlbhc2gj313EhY5F/ZsHDr0a62mdbgOByX4NwgpzAwqE80Ayp
mCRJYok6WV7MGxxD29dlFbqXqtQIFE1TdV/JG5bGofTh/GZFGpLS5exF+QND+SrHvqF8+MQt9hUY
IzVMtuWTQOEjTJBnYSqS6MSnpUAjVqxGNDx/wbV5uA7k+YpIJc7tjjJ1+btHtIf2A9HdOUw7JbSk
H4njGC9MINAKWr74/KlQBm/3qEgJjbfbNsn72pwa1s4Paqdhoh1r813SleE8C02UEUlIZmlsG83D
rErnU9MBkSYluuIUI7jkpaAFSvFiAX6NL0b6yWodjA/SdORHVLwqjHhaGusrb9TPmZH/YCEP3qX4
KJkEcjAu5Et0v/f2KlhD98OTU7JZodUNCVZRrVncKR3XRnympwpFYg8DnQP8EML5SebxVb7ot3G1
uhUulwgfaNHbSfl/MoDC3Ugzk321iKQm8zU2ywkoNSwYYaogzBAjlO/r3nJZhVeGlFQo89dcTSiJ
h4S0delrBuvz5a2slLPzO/3/CrRhc9Cdi9cXzoMw4kK/3VXnmedJ4EtAW7ox1WuXnjV2xjPaqh6X
9WFz/BTXm7VRH3lbHSRu3p2O+kHlmYCRjpBa1t8m/yaoUs4Sf/AdTiaokRrhJ+ND8/89A/5abhYS
eIslOqL8Fk3mR3rNfd/EB1ifeml70ArSa0mRCQ2aOo4oNzLUEjzEcog5oK+9JcdFo9P0OTYuz1OQ
ODpvS4bASkKa7+PWKXsP9/4WCTE5cCLPwb8LPVI37NUhatYSPVkLGPw4llKhTVjs0gyoEEslBGYo
M3E8cKh5QO9oRFGGvD/lDkPcKq/exs03HV8F/OhSLCxYWzWyYFP0EV3DZKGp2iWPCJ+c/swu+iFi
iMVqhuufCjajDADIiiEKcaZ7IREgUqlDrqjFpktrq0pbmWIuHVd5z4T/YOCRkrC0NCtFUimJArEt
gRQhQEdnOq3O9d7MA10q/5AaXzSH8XZzwPG7yoFQ5Z2QBYxhfxIeVrz15X3HFXBirJZclEFttn5P
uvFIQ0DmMcRgOvnS9FnJ8kZiuQuHgNTX1SmpLE3QJAz17CSZSlkVdXepomGs8zkafyJ+AN2LlG4F
JOmLuSEvAaS869wiQ96xaq9sGlGDg64BK/FwUFp8HNPYnAeKS5bayhIccCYKvD/9rVA/kSpG1ac4
NeIoOXBlc+N/N9xhWY09GMhrn+aTTZOyj4Nt/o7ATVeohG68GdpITL2P0s2Hv6wMu9PXWJfbix4k
fFmo6kJDV8qJSk6A5WgjL12/JHtOoC7bju7nQ6PFYdZVxbxOYXAWFS51BlmJS8Iby7Mxv+uivED5
5PWUob3kMCBNfrCnkROTqTiamJWUjmKLk46o0nf0sDAAWY9qTJwapyroP+v+QFPkChdfWeqkmMSb
iMRFEjCNrMrfs/9tcZauuW3a66nWrI4OAv8nK4xS0pYXglkaCCclPDCW1o9tJCYDuXgODjKpvr89
2COk+vMp8QXvQkkz7fqa4Rc1s7q0W5nP03U05Xng+g4yCe7gQhvsy019nS9rmhEYWTKxo9kpgDSx
du7CI2cXedCpNNi3imasGmwj/yHGHsHlfQ5XD6A7W/x3acWUmvxN9b5OXCpB81Xl3cPvD4oqhgSE
+QHrm3vKSvsFD219koXI/VLU31KDYgx+FBTSWxbywqmJt2CuqgTFyH78s91NJC/Kl9Q4jDNUYLvX
PXnKH739dGLR3Q6fdRbEzbdd6F1ydi03Dk0g8RURTLiOuSGhPLw0MhYNMfRofw6lua0jbTboLpvM
OePAtjW7iuZRFoD0/CfkLOwXtETlKwow4/sF6mH7Nz17UaF9WjazhsEO0Lgvhp2LsF9OSfYhd4jN
BU2XPcrhPefVhqAMdqu2+aGOXvtBNPmreN+Zb349iOSPSL7bwCA9OHcnX/lTt57VcuVxV8K8gaaC
qRK8qIR/sj6bDyqjCEn77aJ1bSmXRXgNXADZcFejSC5tjNuisWGs4wZzkI1Gujnfk5KMWUij8atV
69uLdz+pETB2WdGuv39WYqKmjiRE6XmDhG+Ywc+dyBC9TSNfsNCuP3s48GtMf4XNr5LDZXS2EgjN
Nper5G1D8hjv7LneRZ/BSzFolz8vdG8Cqfl+LOVsebKnwuAI36Miip7pfGdqaPTcpTvigZkHfUPQ
1q9enRAPBGkmzXq0a544gWUUII3hoiWWJb1LIXjqUNsGRBFjyZGYL83PdVG86K1osWJKQJ63JRis
+0LohX71b6gi2rWXxJdJgNDGDmSwGD7+/7UvKuKTCQXW7zrukWqbstZnDhnmMSFaMxcIAgLRbTu9
0fNg4sgxD87UuEqsxglSSA/KcFxGvXUQ+VUqJezu91Od3xf/Cv12nZJr8bJ579ryxyS03LL8khXy
X0TNfTE5bYIcKvDGhBm0MVHDc8J5S5qj999IPzXmk1xnJoHYEnx1KHSldLbv/z7SJIZ8l1QVmCol
2vVB0ZkzbnwuW+3p0AqvCcoc2CeBiqEwwUNjCs62foNflDpAbvZ6mV8b0FAOPDFccK4VmGaTILri
02/Juo4XbaLD7U2f3IhSyYTS4EsOuoKNLaSB/MeL0qmUZg0F4haK1C3PnNGToQ6kRZsecL4LwV1X
mFRjPthhAhJKHLb9YM8pfipubAR9g1ChXGrSMK6xdx+utELdwPqizi0dvcOPpv7b/LcpXOz/8S8W
959XqP+NRmoXyEZ1zfz10tJ2ySQq14xsmfAY8lobbVJErSKzOM6nTLIHUadJRS91JgoEYBBkACV9
5PMJxC99tc0w3dR25fMhxWBuivv/DKU1iM1Zg+YUR4Alm8V/yxc8XPTWEopPnIcYO6Bk1hz56bMY
lmrDsQn8QEkh8/IFlHm9PEXGJZKtD3Hz4aGDqWCQloNmA6ZjDmsgXWFmQsW1YyoETZtD6YF+L7EZ
7XQnlXBgo5vuuT/e9WIM4tFHMv0QbDcH9AG9lnd1nKOuZE8+qkRGnYKqmuKZGgetIo7YF9ROgw74
Tj6iUAzJ27knb5P/frI7bhJvegd0KP74BPr9Kv6h+1WPxo/LFxEnUeT37Z4IQHZjWY8AtYvehxal
ip3oSHjQWP55sbaC1TrnfwGR6i8qoGPBmCG5juDIYbo1pS0wefrSr2dI/0upIKbIVuDYjcyOm0I/
Ag8/FI+TkTZBDGDSfObrH20yzFpxeVbiV1qyPqTYIAvG9rdbd1TKb53C4crQ58eSkgzg72+0CBdI
mw1ktsQ2SUlI+wjsFumH/6jojg7zzMpeRgRxrZOa0jZGM2nvodtaOFQuC43K+KkSqST1ePF139Th
WOcCItN30zjXxFfQH84la1nv+JyNox7cuKMcX0ILWCvy2eSod0NXXawLwq1JL8K767AzNDTbmrT5
N/UVaNPQ/czJDHggnb3sUEpt01E53xIZw0qp/v6OM6S3TsmhoCrkU59whIouuJntjwRCbXdavb+j
vHcx7Kcr+Ot8Wch9O8xOULIAcxNz3d604lmEroj627rMvrR/dqTiUiqPj6mM0j191utZy3ieZnu/
BjhIBkU+TwgiY7KPHH8Ug9Qglt67rO+y/3GSpCqZQrqJCMMYjvlF3+ucyI9Hku30ctsbAzbsFtZs
20mNadxi9Pk39u9W4OpKwoi1ZCY4wd/b9sndQVdq9/aAGxwEcrQ2xF+Q9dIu123/E1Xf//PA1vLl
CosddUXvt3jfGVjAY++erenWA8wJy7e2ldZkgv37sZ5g7kKOt1IQ970RSin7nzlyinqHVPOlfv+z
paesvnE/KjwEhCX8pmCd7QJPwBBbk00DAX0TYe6tcyr/1aHK3VAl54fkewkUCqrvJo6sx3mUWXsO
O2i8htXdZVeqkpodA6Dg+9KZkfePYtIXHsAe2WOXVjHFfmmY8sV2rL7nmsDxIbHVHQMxpABI1BGN
AdxsJBGH9XpS+KkKVTJDqR66pyH1a3bWdcW7ZrujGLLLZrvFgXF9A4vhMmBgELtUFhurD98kxG/b
PqXeYeldPA+LCSA8TKAL8RvZFcOAA+fqAG8poEz0QoFLWiOqzxW5blhj+eo/HLXq3A4+Up9DGLgB
uFnGOMgkYlWH2TEF+oqB6xseUtMuHXXLpiS0ajQJSIxXwqfF98YRHD5U/TlaeixL2jwJm0q4brmB
CUubJUOjX2OkZhZD9oRCV6p4LLGNjlxTMvUVLdvMTW/8LEeiriRtE4+jRpVkyd3h9uH0QKHkZ34t
TJ8gzMgZ5M3zqgaHIxig1i7ggXnXkH98eCRkLM+3NvzJHUje//lw5IfwHkOmC9Y/QSTlRk/GMNn1
osepzaacvElnDlGCh4kfmlM0cJGnhhEQLWTtoNFdH6FrI/bAAv7xBJXretlVyZBXPqOiQAhmyX4D
83xZMfMznxtGfXkzgLIi0/9Gb6buKs9SUSagxdZPs+ODTxd8EGUXoUbNvxzGHYVID9kV18En8vho
wgcwe/RicQPY5/oFSwG3mxbuFPkVuUw+BirV2sHJVXGpBNSK6RqdJ5+whlVo4pIntxC1O7jQXGqI
3hBxtVOjUg7Uj37jWw2mYdPwDR5Lq0FL4gFvzKg2ikvfzvR/LxcGJ/gumwVpr2SgwguZ7h9fCn8P
WUWSte7TQhdzYGEmhXEHVmy9fNHB3TIwenQsshmC1NyV0VQCpHlaNwc+jK9rXqVBltbosygr4iOL
92gA1BZV8J1FCzlaS0qThRwVx816Ymn4jmT7dMBfUc82UmGOsQ9HL918ZMf4UIMQqu4ExWDzPc24
XOXlSGq3oox0nnx+TTvymJ4aAy4efS4b6+iuchoDFmWn50HWHKpJxxBdVqrwpH7WmdcXgiOCojky
HXCT+8+hlAA7GI7s8gZE49lg5K19viY82OJr7TXjH9epN/3SmmaRWMa4t5vcbOXsZhy8HddOslYH
q1yDUsQbxXicHygDYH3OKLSZmj/byP+m/+e7BQP17xmYyTeEiXcwJchp86tO8HgjLB1f+HTGtOg5
UUxeAWYRUCBSyHXbULFtmj+e5XES3rxtZtOZQaFlYjkb3vmvbAmIAONR2lXjEb0B2k5BqcCjU6lE
0tzHYjp4uj3xGHlXe97EeKXaH8hDy7cnSeCbqMwfZOBJg67YR2sN904mJrlqGVU0GkQa389QFt/k
4Ok12q0W71DTpmUyDz0sCGgngsIGOt99CBWH7fJdnxic8FvoFe3fY8W3nAx6x9TqGQi8pHjZmQEF
htZcwq/EJD5MsyUM1lmNjHdrJDCiHxkVL0bejsW8b37Y3AGyUaV5mJV54YKE6Ko8+9YO/oeFV84k
PQgV+YH0Qk6IfqfS3UE/dD2z6tVQEbSM3ti16VvRqPQopVCjkJ8CO79oMJJwibKbnUNlQixHcCHw
Cm19wWLlcxPn39s2duNiV/a66PyAjVECeTu9PYo7keaIVWGkys0aqu1ezwPF/BcJ9CFi4dGxgwSe
cvkKfS49SHMJ5kzbydwYFIGlktJ+jLs85lM/a4Nn6gSEn8ePRPKmwMNR7iy157UPpi0gJ7yz7NuL
o3cfb8C4P6q+ey5ZyAV+V8CFlGtph1EEbbrVf5J+CbEEpAN5JcOSvS3BxyQP4E3YUyeSSrv5AaLm
rDBcz+I/ZdXlfjbEKv3FZbWqe6eAL1KlJro6EJeb3hj/8MCsOKIbtJEt5na/qVPP/1L7kfmOW9ux
2yjpg1UxSbgkaDQDCigEOMcALRt5J2E7nzKTko281bjK3yLak8UUY2Fhlc+zbSMMGMc3GGxIkYZO
DfIqxlGcqKR0VwK6/RUQMxeBoi16/aF/jLA0blVtRInolH868bowyka1nKiYyAt94+bqHrQd5XON
2pQKGkU5JQYDFX6PL0sHJ5JZfsuUGXGj5uWJWqOI98uijViAzY+FDygWihND0J5+R1rMaspsK1Uz
RY8oKnuEvVjfI3CMu+Cj/yMUE/dFCVtlmnwdCnNS5Cw0XYo3iEyg7bLkyDH5MgIzutro1e9itZ5m
Id6H5H9Ph6RPHD031B2aiXEg5zAqnnnwP48Gy23ev+ixs97b5s4fgT/lNaHK1fauQywAiy+TuFMG
fe9FxFvr4NUpy73bpnZyRExOeAL42xtB3ENwV0l9iPYkuuVHLUs5ZxdIES8Bk8XllH0pNNePU6pC
E59fcPz4yR/V7q88HxWMusxd4kPOeyB8Vrt+FxKtwinIaX0iRrMAapvlPfOeOF5bsXmMA021EdhT
+lGV+Hbj4DNtajpEOmw2fMccqEhcj/UYlysKMZrQSmPQS6oibDFa1BnYoXg9XbihnNptDFppy4bU
HtFmJdJ5DCJORCZKkrLqRguPwQifckiW4396gJHNtvgFJNOJ2fBt2FU7O3esVLBt3swqvn8EYehm
r67RBllO6MdWhDUxzCInLFj/rZl4086Rn//7Z6H3p4yoE4Lc7NtClfE55AFfgyXPYRtr/q9Opz0D
lOjfMZijHcHd11nRxJ5KNn8MgFHXyX0vDAuqu/U/azWsFgJzupXik3n8qF4/wfnQwp5U0kTD6cu7
eBGyhj1tsmXTn33YNEyJEmfDQdkfa/lgXPClCh5ayT1W3NLyBtN5mcBg3D2X0pjVT5jjVfuP6KIR
EDfTIZo6sJpHeE04MoLEE3L76pKp3xtfdX2EIQB4fHjuUBXPGCjRbDup7cUSDiNHFzXBQUPMJnua
f07eZmGlMnONsyzvuithsQSxApUGGczEeOYDeqj9kPTmV6LM88IlcwnBrxMq7VKHzsW4VaAnTq1v
MGQbH6fU9oV1aN9OlJ/mVRtOBDx3/slv4mxL60loNbM8aLF3jWet2aJIFEICX3bDiGwuGHc5Hf4z
MiZLF7/apwkQK5n+igOr+PMKmWbftjasFqo7lcY3qO5zVPamO9BNyRi1CRBmAjN8b8eluFwQC6cb
H/XPqjfVnduIrjPCWAzRy0598oBFE6apOtHnQgoIqELLB2UZh9iyAoCCw2+MXc50DX6G/ReMlAGk
ubotGK9Ucz2OvaMSxCCfiZ47AtoQCqBr4nKgt1lUkjmLObibSD/vn8P+0jKYZZ2CkyJXkma6v5lK
IhYd2EWy5dX/tbzTZwoapSLzY0idQ11BKDx8KUlPMzorK2vlA0v48jTd2KgyNMZLLNw/yfAXG5qw
XSloMCwZzk3hcqGzK3d64cYR6Yya3C9BCQMVLAMQVESkk4eLlGbNKt1f0ZqAPQcIdgvnXDwRb9FY
NkZx4CkZUoXE493p094tW/nB+hVCOil2mY1Z36I5Sg4wAvzQ7m1PanaLnT/CkkuDMympqPP3wa2J
BVWjhfec/aiwbeXUcObif/g3h5foKYS0pTYXuGBR4EKjzK15/NEDqQERZXE7OA7REGeNrNH+JgO3
xOKRXnT9p9Rah8zBF01ZNoGXsvBpf5FBC28f4w/NUg8Zf3Nv3KIi1spTpA6iTv6QMdT1diUh0fwv
8YZTAT+zYVTk7yBe8JoA7Iw+oMMiFVhXm3CuW2BH3sdOLUb8QLFcgg9mWsi9wJe59pPjq7LgQBnz
T4T+7jPs94vwqzrLeEdtK76bFlCoQ2222deptWLwEt/qrtOTxtJJoxI6HcLJFKXnxoy/4fdhUjJO
NjxF3jNJjF9UEU5V9E/hUnCyP1Bh2Lx6mzQ7/gWYtEkETaCYAqdgtw16aRhLzx1i8UfFrC962VCl
reM5j0sdDJrnRA3mr+mCIZAiqUhqULULNhUc0zV17R6BpU0n11M3b/3HW08jcDc79zS1p6tEAmR5
0LbCcW+O93YORuzTTqzt1Pyv+6/pN5MUt+p+W//hUslgVOtyKd5USWkCJdMeZq7GGbxVfMt7sKev
Ps7YfQWmQx+1t1RUOXGIpZSVkNd97RLn/JhS+Tgmjl8AoqjfhmzjsArAnEmqJ9AvTnpulyixLT4k
42etlpx+1M1136yDXBGmtBhwWxuuTgMyddCBs+KqDlKKTNtU/PzbwHDfmPMBx9x9P0j2MzYzOi9H
39sLu1QTBXQOKruxWDbeFKDFoUy1kldfmODrrNY/on9gF2jheTCzCFIWbbhKB3Ib6xstbrO7cgL4
NcCr129uJGmBve4MvsXPfKc6sVi6uiF4FhTrDyzWDtmWpvHyXWxiw6ZQ1ccRtqkvCY2F+CBdjFuz
yqfYT9bZzNJgbwQdQA+Hx4PDuFuIQqP0MAlmyGliiKXltyWgEz0lpAG0iN+qpfOOUscsz+sonsJ9
WLsqdFwMf0SYG51kYO7abVjeE3DqBfnD1Ac8AIcH+56wvDff5fTa3ZioyIJFw1cq8OlgAEIXrcEs
ffC/S7YqB3qQ2U34b6zsqqu61Jfik9iPFtLrAiBYdX4V2LLUpZmQ8KwGs2Bq42LRxCpIlKK1s1EH
pyRFpD7m98sXWcwAaVAtgbst2q0fQw76WExaAAmE+PMFMskh87w9xKkkkaf58/7tnhuMg+QzLq3I
RuyE3bHXCHLG3UvZEo1tgJw5u8OZfP2a59xxxaF1w+b1vptPzKen44LgFL4yKCITpwDE/EC2s7lW
8lnw4/0KQBZCcDBjMdiPKdTPw77xQZw1haiU+PftY5eX1NFFSUnPKJPuPR2dplCyHTZCCP1b/CND
yXY1iBUWq06N7u4bJTv2MV+LAwrpIdYBc/LtTnnloAMYcb1/wXTVP461xzKE9K5Ut69n+LyY/l1x
vkw92sNb9TVaDbPQRkcjy0vFhzyEe/miM9L5phhEia9xIJ3hp7enhewvTL58HzFZAZ65sSwVY+5y
bLvJEOrACASV2howcX5Qy6aUFJ217ZqBtp20ya3O+MxrmrgiIrwzNNonhXdFzALM7v8jxVvB5D1i
34T0KTit0kHFrTjOR4VmxzklHC5IPEw8+yG05FVfMefrBboyX947fX/B8OFgsTSJ1yYO4sY24rEU
K4GaaFWTsFkwbuZ8/MUzt8jMlI3625/d9p0/x6+nSGM97Ug0KummO0Rf8pyQw2eqBGwIJ2OMVm5x
4ABDrvEupgpJ/tMPXpSw2z3pwvRIKDE7xTOzsHBegU8Q/otu5/u75Kiq0nEy+oJNNsaCNoOoKAdy
qrT48U+SB41BJrjb01M8T0fI/6v/+jev93PRU8N5bYc2GRKih1wgSeCUjqTHoOQt5irYxCEh2ZBr
d213IXb9hSBJKpWRvPS+FrWTEzzZoE1mIeTJsXQ3HlgeGSn4kWzav9Vw4VgwVfKTFa5troInX8Fo
4GF3nHTK3MSqLG2BNy2d2pIs30D61YEd7IjWVApasFT5aHtOsscuQFzBQuXKhXAeSR1bzeXK7DUM
aOXRNxzjpTsGm+T+8g1bGuHMlXEeFqIDYvqwS8l4MtI/XiYFnwIb7P/Ssc4xPTu+64XKbP/CwxFp
BlMbepg8BpgpMYC/TDHEBYFwK/BG7sUu9rYpUELwni3ofBLhKbvzl7swm2wCz02fD8pntoSylYK0
k/2KPl3XwWve03QV63THywE/hoAhNrbJV9Pu2hKmd5UUpUuuEWEuKZ/9mu6W9f3TvbCBz5C6wPzL
uFEXWAs/uNggTD9ZpmDZ7tPzsaMQ/HGCHcA3sjBCGDajhJdgJk8HXk0CMP15DOTFQIQph5o+gwYq
O+y+XVlY7T8xFCj2b85BwD2FxMugK9uke3UyCxX6z/Py1EV0dSLV41CS+XD3l+4E587ewuFa2OLr
aCqtqTPoj4niHoTjkQX22QqbvOtcx4rOftvbZanl+JrqscB8YZi4yDPls9EXqzos1jSAsTfCwn/e
o07Prffyfi/LAPPSc0+VKbyhrzD6lf+uBkIylmw4s4tK1ILICK87dNDuZkBIMN4saRIuifrLaDRU
kvGqVQ+fT7iZapPGzBaDaw+SztgsHWvWoVgEeMU+DzSKb+GMDKESUkBiVGN2cEpl+Mv0Bjkf/Eeo
CJMCeiyhPA3u1m/xku4GPI7M8v+nJtL34xThF9wUaU0dgQm7L0Cbq6ifRfSF5x5aoXeJZQ/oJDTd
f0Iw1FJ6VR9oPqu2cwOSWnZ6aJ3hvShIjRt8zIS4lfw8Lvh9niwRGg9o0Kd0DJLWjapyn9bQpVOw
S1YYPs8F/ywnmegObG/x8W0Eko4PIJmpTdcUJEJp750ZvR9PmA9SnP2nbvDprnloEn9aZ5iaLkhi
OHxvkzDAH02YW5MUDJOzVwCUwyLZPD8o3DgNcyQaPFwmSLaPKFS6dDoIrRfU+2cqmO+MN6K2VBOm
kWPx7f1P7dwkgDf6jUIvX+9o2DUkqmKFDptBQtrfWU7nyiCNYY1R91UHzGxxm8BOerGKjD0Jx2tL
PJ07kGM2jc1NpFZp/My+B6gh8RpLJQXMLwazmChTO21l5N8ShBFv5MDcxPF5xeskE23743hm9emc
ERpdOyHRBHD83yMRH9T17PJ8FM9TlsRCz9VhQEsTEKvWhEbbMfM9uSRpR2zvWawkEQTGXM4zgGYc
+mOr3urR55R/TxpHvi2oVCe23+Zs10ty4xIqa6259s3iEcppl7/8P+hB/wH6FamtjIP+61gb7akv
18WUHBzi5u6ZuVGwjoC9Hbmeczt8gFRSuv6l2sdm4it348u72ZI2CLnkkmXIiL6ClrwXVsrcWSjH
KwiXuM9sAVGafPyMp7YQyKpoxS4Lv4ONcfj3nnI3YHXBORByZMhTJpZpQx7WyNmqkIBa+Y2V25eb
VzHYAkvYgMryS0ssBEEmWyPIyCwRNsImNdruZE7+2+o8koFsLxWtaJSsed8E2BpONaT0Ip91X8PS
YJlQIr76TXNLBue0MV844gwoDavW+QwInRcw19nf5qOkYpYQJyLMlGP3FtHQhf7YDbRcREdJdoWc
QyixzuFsLxDNM84Jxp7y7eQ5UtjakQt509t5MnZz1D27iywYBQPsUWtOVyHK5c3pPu2xaEdlFXlp
FpksLeiytxcvgI+Ap3rDoa1gfrzEXW0Mo4AeOLJ+z0BlbUAVmag26VxZOgg3n7dXHe/xIqXmkeH0
BUQuYfkhYIYfpwPRG2Fd47yCFRnJMPnWAxgBOWYtjD4eyMNTaIy4dRE8+IxweeM5E1gVaD0d5huI
Nf+slYR8d3d3vAq3z7cfwbC3vuo6TFbjDZbbym1TB2bYEeCBhihtkODhtrZlMw4VFIjVaI2+e4Yd
IsXAoAwjk6HzrlJPqBQMh5gbJi24xrHjtuZFlLoEEeb4EwKPv9wr6CRa95r78HLR9r2f8nnJ+SOb
Q/w2YxEtdIptYB3Gx+q6XPBTPE5yebb6E6u1GT5vRo/R82am53p9MgomXS4GCusMQXjQsnBYTGW4
I/CGZS9m+qZryziLoxcZHMf9JyUglvctVDcgQ06dVbTwiR0mj9rLL29lF99ELfT+B5xLxfkCjtkJ
0/k8LRSVaNoMa3dnV3bCZsZqFa092fPpLc1p9Kykwtu2VzoL0isZ3+q8/deVIg1gWPamBxPiY/AK
F0OQJYt0/VQa5kYEEFHQ7s2/nSSqaQuboFnDhZCfdV8olDtRvNghKhezxQM+8TiTu7Zz2g8eoyeb
4sErya7SqC6mHMsXYb/lSeHbRScH0e3Thtt56V837flpz0LcuMUXuw0FLluUx1JBkboys43kXV28
/tF/XhYPxZ7zshKbiJazGRcmVHOmINCUfsLHaSMayvH+e5wAY55wTHL+vkqkOuyAWL+Mgpq3zUxr
yBHL3VfFQOkhlVKtphsZvww6PsXabkQ3J2NBH9y2mURIsFbJa/YAzkAwG8uvcghNTw4t+Ju0xbRB
dZb0Q03Bo6miNFNibLvVaKrvvRP4lUOYsr8kgVP5Ne5gWrsNnH13PSbORxmp7TxmiyehB1EV+w0c
SIhb1uloHXnmZKY41oQHlZEcU4jnk8aNE7ccTkiIXRDC2higP0QCG563iD/E6BlOtRfUYDdt8kLY
GpxLT4aHQaLTiHtVx8OfrQ+bBpQD9cVv4RO9Lyi2PZGykDTdQCwD/arqjcw0OZDoLapdUojjUCD9
Hj/KhRkEj6OHRu9EYBFUGwfv2RUEQt5eelepYOxGQlxvlOUu8vZ/pSZC3NatMfQD2rq0ceotoOCA
XmHWEaHhmCRzcZvx0FFbdxJDL+saRALpvab3hCAoCC7reJuttJLsM7SPklwK3b+oT6Gw+iCuYds5
fnXCQTbXFYMSXlrCzyEppIG0qJU/7m+7BUQIQS8iNbfKW2cMPKzEodFmotdMSFhXobhP07WcIYXN
+7i3KfgPGnKKELdNXSPBwdVcbiX0LZnJJ7Mokxz+jsVTAHZ/QQoVu/7L1lyws43v8U+1cH6tIjtI
qseGCaKYEskRpbio8k1NfYCj8oS+w/LSN0maUZs5/X9jBifWWyOtfodXob1QTmy3maBWHIwX5okB
d5ZTyE/LHSWvSDhrok7HM3+GWt2yyf/myT3DQKXzr70ZWspFCnqjVQDY+z7CH1aYOdrKC49hbg2q
AcCmizC5uaWm5xiFNkHhkaySyAV8dNfL0dghn9C8dSaAHoOiEoizOHIPs2zDmTrliaERI9IxD/33
c3UDW8k29B9LT++NytU2MpwlEgOJPanG+sNVMgq2IWMbaylBFr5i/0q2zH+ZHzye9dRsHLlt3jFK
twiWqpvBKo27UQAo4NvudGJ1PLXT0Qso34v7yEjHFzBLN3cOua47IG6fls1iYQ05o23nAUH4OlHa
GWgzNLs2GTDlMiPDhphho/kvD2DruHRu8pjzq9aQVn0oghlrGgR1XEMLzIXOSWu5BLFtCt5eQElM
r2DMOSTowSB1L6dxRljgypRvWDOg1u6jvauAB9kMaixs469G3m1pfDK9gv8flW1WF5ssn1jvNlhl
ABV8/dyWS98TUwhj+8JDb2gYTaKHA6OXA51FWhBiDU6gRJLb1VznTeekN9WLdNd/8YQFrkwh9Npj
ECnusVi29QiUEn033kM0kU92htHIbQmRkGVQy0nRW0C4NafeebfPFEp4rTIxtUglqtmhVT6b2l5D
KvOn4wTTNX663segbIYWTx32msuT+HLmGgKeALeOcIQTVB69RrLi+Goe2bnvlqWeFk6XoMMHv6qB
/KZmO+Iz+Sxo04d3W4kvoR1hY6eiYBCzRQK6ifxm9MaAZj/LCsdmfWPyEgtMlChnyWl5+eKKycSF
dmvJpyWcOXxYIH6Jwy2NRMg5N1oT1NCE4aJ9xpskfjO56L44Y+47jBN/XZvqc24SzxtZ3qVZ0Zd7
DBvNYJy8wYrwjVLBu+nlA+hdnhTD7JNFh8wPhTrC8P6/0+klMoVmGsjY8pzjnoPTjcfciPQcN5uQ
rVqh+iIU7tJDTpUU6NvosX14uRk2wHS/keGGKsjBxXJkmTmcc+52onzdSdOnMoFqwKNbrcQa4Qcp
PpG/OaGFFK5Ec/TPr0P3SYAGBNvYjOe1+OEu8t1JfRFMwvaS1x5UBDLXEfh8ZKM64IPeq/mG2KRc
mzKMr5YwAq2MEfzvJJN/N4uiGNKUNm+6dNGvYr7CoxMLNKiDIaWd/e6iHFvP2PC2prhaF4/jWfH9
XZYrRtrtxV9IFQ6DfAtmL/ZLX+6gqyfkncCl6lkS2m0eLrcQ+d/rPUBc9pxJ1aZD9fuCS/xlTif2
X58rWrkX9sn9M2XnDpgOjDo0WuyYJwKxWVa2RDkU6lJq3v2XctImACBebPj/vYY0jpWKJipUo2+T
C8pWzDotX0HAtmLzqfLMj5CRfDDku6ISb1tlsqZgBFq0kTmt3vCRnUxuPI0Uz6XTm382nktYVdJU
qcYIe1pYoo+pafG4TusBKQAM904HD/4tDrUH87JESkos5tbwtHGF4V5u4Zu5RPcKT1Wa1nuzGAD/
jpPEWNlz0UiKf0H7I+Te7JuEye2zVkoW2/tp49qLi/3WBlQ3cfLZPuG/tUtBXRf1yHZrttJSMxMN
0eK5YL6Itc30PsYPWdx/Jz2eO6b5Fa0Y4q6YU6o8wU1bAOgR10s1x2JjV8s2izKwNtU5OL5ArLwk
F6cqTBUeJBMD0d3U5vo8s6jddnJXYvQPdeXeZkSYi9EcVSi5tKjBr0l4fiflH4H6vwzeemvHOgpx
h5HjOyym5JH0VlHo7Bb8V8Go3QaLr4WqFtglP9FmWdCuMY07JKqr5mm/xhm1voBPIkU3WBbuaRmm
7i7oF3AlIONJiFmoGEZJHeTZQ1xX2tZaeq5HR+Zd5jfuiSwKSkpHKnI4GPkncOOcyAodd5EA9WTq
uEhFvvcQS45ycHMgnb0G65tAXBDlSaOZmUFsrtF5/POvqH2+6VnMGszLvq9akFOl7vMze4jYcXZp
9Hm5jGSkwKr3tVzMcHxF5b0mdA5RhnTSNaSqO9JQ4DLAJyMd4DDXwUW61Fz/+HnUxHgTi1D0KDZe
98NXVYWu27PDxuQKDzZJrScT8sk5f7kn74F3SCp/wS4bnf+/SlNr8fACYJ3UF1pDM2s60dXc9Q3h
vQHuDwR4PoJ7yvxRlO9O2WEasEsSu/wRoQUCkRYlTq1pmjSseOX8qwh21h56MAM7ZPRYXomf2mTv
sLlERDXv3QjlJZ5JbEk2Yj8iLfzXbZR4o0GlpHlP+pSgEsGHHWLBI8mmJggSqJxVhHHHt76flgqh
4tRecQJUEnolYl0TmITNJrSBrYYXLuKt5iXhwj4lOzzTu4/xiK2virFH8ilEtD8sOlLyJRhtFFgp
kkKw2nUtcZuhLxeXF3f6/GZVHno0PsPMtFTJuSWLvWGAaWwQoN8QVvkOd3+Tq4EzhkASWIoncXIH
leLKLGDrh5ZLOVknvfAs/CvrlSXXHf6I1e1794RogUz2pcSVB4/DHpPM3Ij37Oat+zd9PTI8LmP4
yKRUvLObbI4JfvS4CsJ5qjE0+mynvdDSTr194PIJJGxMQQ3WLwbePG4u2xwy+j+nG8oHB/ELbhHC
hxtyRfliJmHP3uQAnfwciaFxMA0HpiXovQDce2hSnb/cd0CN+M1j0V2F4VNI+mJOtfEFgSn6zX+j
7QYCQ1bAO24dUe4fxvHoJD+ewYjnvUy+HlZ37a0y7siHvOZtghKR3FcDidgohLibnRt0Hrvrwo4M
u5yMy0ZTYs0qnton0SJ22w7grhSvdOwHnLMBw8D1dD7wM6v9A2LeLEQKU7gxAQNFS8LNlrUWwsQy
OJ4NMsth/lNXztYO3zmFPCkyCBWS00YYOOV3TL40Ubad8p3jbjQm0jNPyEpaTaFBzXkIE+h9KoVl
KhB6tCOaIvlCSCyiRyYCPROkz0Utua3qAPC+BlfQMnAiaGVWSoJK5cbaIxsEUSJyG51m2kMpmEhT
Of2zC6cBnPtZc9GN7S47TuYeqls1ZdXqNOe7BkAC+1JgsWHEplq1T/BELdqvBAP1L9+XaFm/+gye
fJmShZ9uBxI0c9WH2vkI1MxSSqpF76JmG6WMg24ZR/bzvOUytDOkKj9ht6Uhq8e2VgO7xmiAOzxL
n3EmwG5hTY+uA0FW9ICvOiGxMGqA3xbUn7Kh804fwSROZfgz5+ByaSmoEkKIG537QKJXPDKtgwrH
R6ORoqlA8FBrv4/5gD9F2CCy8KvfUTAUznTUROIxFONv+B0rwNKdgtvnP/s2GGtWAzPo0LTe2U7j
heC7WtZRGEJRG45f/T9c7amcC1yVUI/Ja0PwjpGaY92/Of/nzDOokZ+YaQKkP0+p5NlK/81lLmGj
ccqJ0n/YI01rFrfRY909mKi0nhGd/LwCK375ZMs3RRABz5DNhIPHsh67dpvH3s5qwsGUsl8h+8w/
6xzAQfQ+iK8LJDICROiuZATXdhtOgy6uhPXPpvnNagf9UvET+i7MWKCpSRU5MbqkF7Dtl4lZDAFi
Thj8HjmG5/gs3Btvz/P5pBaeIApQRLBtJ9Wxm1BwjincpJ757FwGW16UwfeqPNxO6PwH77U+RyYs
3JjLs2eQEChb4+41F7IyhHFOEmqll57JVhowunTzMYiWV+8D+RAmmbtrHz0L7dNcEJB3MLn1Zyj1
82jIdJj9m0kQuLOaUyeAWD8ohzp1e3pkK23p7JTSLH7GLYznTpOeQqqtKG2DJrqjEr4Ui09B1ttV
0JuxVT9lUGFGCp90g8WdcA7xToWjt+bIDCHgluobIdyCukxx3s1nhZfV3oYfyunlSDKUNhK6oVfA
lCxIIjQg971BJasBnKfBOoVu6SV4fTDDfQdnRVC0dOikAMXgrBek6eaux88jXbFGcCwpHdyoBwCV
2FkiPKuErMjFLy5BJUpyBCWlvwJh3DFSGvGbBV53XcMgQjv4K819uahqDb2Gr4pkF6iSjlMeXgB0
7t4o/67GMQqdFBFelzYDweX1jhTUEstfrJ2bDJTquH08aOLRLzeSagZaOAQ792O+s32iiFms/uPy
yp0UE8zDRM8VJ9N+ElezMfxE37uSXftlX4hPphJ5TzZfyQW5ysiB6xI8QhZv4YxYgmB2W4y8X7Uw
Ud18zJRZB8j7J/1d17olf/3FPcArQI278aP95zyM3AIIpCpgPpTcAdsYZUIbPGB3OagmMQUKrpyO
r8ttq1JbKKBNxE9XPBc76z/16tpc02AiDXWmQRszSMppfhcNDNn8QHOmBfaEwrhIArzRqe/B8aHE
JHe18RxOmBdKqSyh/zMVgBjjFRq6wboGx+w0XS2FPjlPU52jtkp/oqsLQZL+f0Fk24SPNZvANTLX
OGFtigH/DNkgPVW94Wn86JcMaUJbOXjS9+p6+M9ctIUTy60ld0Sgt4ldmp3VioH0ljTChdpHrsyU
qmMeVLdzBq/9Pc0QeCcnlmSL6zE4p/UIDKAJHtNftG3yRXGngIl11XgF4B75ejsQjn97dE8F/86i
vdlEIliF4BKafKROBJSztHLYLcEppXRpCVV41gNokFHtDXX1HfsVldNyM+2Q5eDD7IJD+SDQqkJq
Q/nXBxZQrG8ZrRj7Bl2lbotbvUne3LiH6fxmttOlfjheVRD8xNPfp0LrJAzOhXUd30fXT4RbVluj
Lp8Syk5rZ8kX514s40kygtQPnIeGxyPbQnfQNZStkcxSiN4JqFkTQLYST1qglXvJo7npfU+BJFPG
Fbsn1mftMBdQSxVndC8nkXhiFLapWWGYxYu0VheX1Iyg/e5g0pEjbNWsGju0+LV3Fy7GzJvVParz
GH4wr60DL8JXDI+KbqeJGYRaaCFLnFYlOC4br9FANb6x+stbBu+ZiTmpLfA/OOfQ53tCdnqtMTDw
eQ9e/j+ayhzAdNfKgiXYdKu26wKo25sKKZoDYI0N1z8lHPMC7M7S63U9Q2V+9OKFzvU2I4Ih66OD
vyj6QgI/kXk88o9yMz6uAdFJfNGt3+Jl1bUL5Gu47EAA/ToTqT8vT4B54vAfyutsO9WA8MJON3/M
s9LR9DjTTEkhpwP0nQ9RzRv6sShxUy4rP2Q/fYHguRKX8Cc5N9KQKBoEgDezHX87bPnoJmc86mAr
rd9zLt2iis8sn/BMHfaAG3MN7pxQotmQSvjzU83a2pNzh5d9V2Da2BLv+BsBiNCpmmRA+nvyIGEs
3K25m1GZ9w4J482mi3C5EHtT26pGmYs7XzYXSHNauMBAka2gkND4q9HPzyK4eKO1yARWAGKirFc/
8vAu/SlkGhf7aPjGolU80B/zN9C3KE+7jdiMXt0nUzbr37LxsAjFhHxzInOEN2YUFIRwINGZPQ33
WcibFVV5iEN/MTP9geJzBvBiuvx1NJI24ReoE1e1guuaEV7c31v+NzT+uRhWbnGJH4PfhU64a6cn
VpS9PcUu7no9itlhi0sknA2K1UF4sP6s4IJOJazuuW8uHVdyKufdjDAdjNQ3a7t8oIBN5Z0nPws3
TjATnwWuW/QKIflvAnMqSNCR2ZFs8WRSjdBkXgduV6/VRjZRfBRCDCN4JcXkSJjuGsmNkp5GxH+v
V04XMWTn+d5z5PQrfqhker30FQAneh4rLZsbagl9xSdq1VQFNedUPDaRxiGC0at/iXy4ZUUSwcWy
sbB/R+ABvYdJK6bSKvFD5wYipUwvdzToNZOYAN1IOo3uVxTRZLvA2ibQTwiBdMvzBwaL0eJmf4cZ
AndbJ1TZJDlu62p87S7RSiqtAJMsNYCmstfarEstWQhq99Eh1rcZDw5Yf1ips8yI5p7XLyp/x1V2
9uIR4z2lDTLg17gWV7/sv0SGbL3tNerFNW8VtTJrdD28ecWpAcUqDv8C/Bn+mkJJjFVWGmtbCZLp
RKtQvNcNmNtjuLj9FmgUvQmCdlNsJK/OkX9G/Q8vcR84MpIbeutu2bcg/oq90VC4Si9HJXjO+98Y
dazSqx3vWDY7AyRCdHuwt/xscj7ANnxgfI+2aRpuRlh8uTvk3aWPynvowQ4Dmmdf1Pn8MOJF1IpF
VXRXMweeTtcKoCVts4kNlHGBzz81uacZw38t0UPazE2cXfsn7gg0kuW0po0Shrf2JMDZajb2a/Zn
fau4zdsFRNP1KduaGgbbTAJvZZLCl9Zome55fXJ3nim3mJaFT4X4WzmMbFFGwOlozfOfPICIDuAx
ESJjUyPKpCAoJwNEDs7I5YKkPzE8FiYSyvVQtfCnLEhfE+axNTenFCtmx8Fk1dIATAoGwzi1NTf7
XNtcyJ5dAE3lQGYT4j8HnWiCsXXK5f9PwWvGHIPCkTxdSZks2kmtPIAEtz/Weufnben4HugMshcX
b20bg6Dyim56k+eqXXmAsyNl8OOG832fdrAE31MHk1qaZ+OWfe1fOyBZPzygK+femMGBaHC+kVmC
sYqfrUTXmfDUemIqEgZ+hQxyxWA+vRyo+NjnwpqJY4ZfKNha9Mhe+6NmYAQZTuKd0ZugB6syWYYt
m5YWsCpelZ56J2PRblYFxn0Kd9v+XeMpQ+Gq2AXFvCy/UptcGNdJsGX1prjs78B2moJzU3JamHFd
V32p5KSV+Eh53uFCDFXJ16UiduR5TDDIQDkJBGo9EqVgbL40tTziTtmBViIJhwynrHmFIvsJ1cVe
Offl1OGy2GgTXMNILhFZwpZhPT5WemKgVObAsjiBjNIveenRSaCtbrve+1+FRkmFDqVGMEsDkzNC
ybKV4QUCrvVq4yzB9GqlNBuv9P7ClECekz1kxrX1LPx9spkzJ5JjQG99aZc/Rt6W81kWdZVSZvkn
Ttsj5UFxoiYOBwNS4qk1pmQUHApU18xk5dmQEwcuTDWxmqvkBr3yPXbR0oYDrcc6fmZsV73NYdrc
lMRiXeJczrsDdlaHKGKyUM46fSVTyovYQiFZR6EQdFcMykUfI+Ba68YRD4MzX3gqAZqtqHWXRUYl
p8Kv4bZ5xpLgeohyff2xmyGxZTgO1MRYedr0GSgEGSCUC+pRNwHoYVCZJt4xc2wSBHMtJ529fjW0
kXE/ghMNwsVNPaFdgDb/yP5VajEF0xMW2uEahNIg81jrwBZLy96h/BWC7crcd9jaD0D8eALDZqEb
BhsHw/9K25z5ftLpRv7HRDUuk6sRcDY7ik+n9eYWamy/5V+tebq5vFIY1xzRMxKbuu5rxE01hwo6
OBfuunQ4Er3RFUhW6SdbV24rXO7LGgC5YGu8AdTt9iomlp7ed9AnAiUa3fxxDsD+1dYgDXjzvSaN
3aekKHhWuvaXHBeT0OuS++XfKGCfmhMlSLyaceBzrjIgpkDFY0hJS+BWqPpRVwZoQqeju8BGJ1ch
8FYm/RFsF76P48t05GhEegGzBibsdtvXCaOvqvidENYaWMACx46lX+B3SuvAzlZs+ErLcYWZqZKd
/IRjwfiSnCN6YY7H/o8azVWMwVPJiq/uuBkugbgTuxNGsj/hnn3lyhP3wcSfTyInphfwyqvG8bGs
Rb810gxhd9773LrXpEyOlBBecMglVAQsoQv33l7Y/qLBU2SV3iBDII9bq+0ku0Xc3DHEWas+5/ST
8y31wYIT9ms47ATcltahIlZ36Zi9T0FdpPoRYfJXuhFwaFi2mvsa3jp5F6jrn7jBxxjHjCdKwqK3
t52pJcsYAm7Xr8BO0SfAEeXBfw/2O/vgKwIho8DJAZQ5CTtaiWIr62qRubuYnj7bVtcJdMcEmxO8
fz95ie3l2aPbtMzHLUmjRsdRVCQOwKrTltwGZItW4n3Zi7X2LTulXV4GoPx/f9ioijTV2a/XBFAn
IcIapk+W5CnDTQ2X0Vod+/LUTzkznHW/IO98s8n6lNRkV9Pbbygr8MZ8BsRcBFhoZB4WwFpQY9Gh
N/krpIq4CFr3rgy8Q+w8t8BG2AAy6keDecNuX/DNRourrGtCMwBP4Cqr9yyB3sIFFUf7uGXGj6K/
hBKuzm4XOl5ca+yOCkHgLhrcG0tMRNCG78Z65uOdXGti6EArVkvdLIJEtr+Gfnqh4poWzZs4EImu
nm8D2aJ8KZOfiwqRwlawew2OHRtBZTO2siQdIqoh9FzngIcrxGwjXihLRDcOLx/A4YCr3xPqwSUq
iNtzW1en3G9UHc7KdmH8e9B5UNqK5IqZav7oBgCVabBPsOFYN2Tpv6hSvGFUq561sW469dZ2umta
9HaC6F4+gKmfUki4kxv5S6/MT1CL10lppU9Yj+Wvudh8+js5hzQeCK+Rfo/f65N7PLd6ntiFLJsL
T/LddjsIaYfWx3m+LrcUcWj2xfIgeOpoOqwcHUGSiOt/L2uU6oFKFTQ5q6QxZSrkPVNPtMdlpQ3R
bYKiU6OETXVJI0Lp2uZvqMtrZea6ejQCDcxF7qZoQMYZph331kDD+4IFR4aUtdAd9J+TNIOP88LP
vu1MHHO21rGUrJ+MxhsUP89FnuLQSKRTJWzcjw/lm4+mMW2drvxyB23TpPunIIFZO0vlZktzT7df
oT7qVtoGF6aZmxbsI7GwyXewwPtOiB5MVv9yYgOGXPLZwpuW2txWkv1xnPUDut0xgDAGVWE3hmgH
gpAYKrszhWN+0TL7nUwfnfFhB6Ut41TcKzgesgRJ/saAghdoYi89+GhAmxAGW9EiDIPr3HmrAAkd
q876BsHXzVdEYtd5vmYabcBrj3AKm5DBZ0g+Zj9Kne7P+nrkNzFTl6gqUZ+Uv2T2EG8RAMBRPhiA
EiCQ4D/we7ebYS+nkj3HP+xXJnRhL2vrH4V7YzDMmHygpf6jzGf9E1xfPoHAcDy+QUngNmn6SAQc
J0l/0OMiIYYEKZS8m9ukhd7KIJ56/Od7K9Kubbrurvd7GkLz5dXsIfhN+BKakWsyhB+byDMz/SA1
a73ufoOI6hcSOgB2OeNeYBPSs4joLy2acekELf27vAN4pVJFJ6YhHZP4EWuytVc32XrRNfzxgPcw
7kWoxWAxkjyYohHi970vF6mPEbZZ5efSwO6oX7mfxpj1npiH8RttAhYxx3Gvd/CWtxd84u98jaoX
lWpa95YxjBB/hxsykiIZlGDzmvS6Zg1mXCqHOuVTpNQRTopS0w/dpBXbXW3C+3ej8K889/V2T/lJ
RIWVJreG1jpWHeJLTnFiM86IBttaFYBxdCBhMBAr+iUFqX0f1Rq/NRNC2trUM7QdRN8snwkLu4AR
nNQEqBqBE09+pThMmiNSDTB2qB8OnO3C1We7r+MEb0gQCdlJUu8a+91a4QMbe/xeR12prhJJTBA5
SWQYof0Uj2rUKRyBP1zapavWFvWjCRn1FrUv9V22xtzGkMfxrfxAR7uZw4OkympM1zFeduYzjB6N
cDwDeSEa+Z8IGSvsRiVhXmcYplBpaaGcLNZlecpkzbUKmia30mV4NUVfumTANG1sYOzy5nLt4cEI
bzUFKTwniQEpLISjM8yPmqkniA0XFgaban4EnawGohMNFKg4c+fL5WFR8hGREtRW0KxzitPlqFBy
/ZRQi5WPGvznP8Ke5STbpsLRBNMYvVTohLeKoqBF3CRFcDhHNzYkRHhdQnpby5/RoQKyLBDheCp2
PPS3gOY5z5w5HIqOxCFIi0K0u0AX4tnYU9kZljevDwLEKJXvH53klKVyfGL4qVw6n7LjiXjmD59V
PP/VwnbSzYbcgHIpeVQ34eGqDQv9Q3nsqbp6amzIJEvEhQA1YAqVyJcwo+X4YoD4jATm5/UGVFcX
TpH2tu0BYJJPF7vEQiVdtGg3H7j2ITmdZvYi4mOBoFR6hFgDfzZ6+gPdAyNMX4qWYWUKPVFeCYKL
JvGJ58ivXLAE/OzJNMwbriUYAJ/FqGbhZxvzoujZ5RDRoFrLjitKX/bJcYKdJaWl1HlzY1Ru3JNt
iiksQjkjYEjeNZ9s2TQd05ZMU1UYbdGcltasY4x0Sgwoy7P6QfT4XKEyQqNK6bqCdfUi7l8NH87B
cF87U9jkvNXgSXkESY68N0oqtS8/D68utTch7ttr3DFSeRdaGpBBXyOjDJ8esJfaFneYg4RpIVPH
KAML7Nj9/+iSitH0/WTEK4klLWr1s7mUMVAEV58HlRYQ32JwTY1ScEq5WvQKNGFDGAd1TaW4GoE6
jedKsw+gQcwP0G0r5LG4UhAM+RF/CcbqPbeTu+DLdHBcKYmixQk6Wfoh9N0ysEg0tkfoPsHIdMdQ
5SZ57hM+riwc7D2q7cO+IUyh2b0eRGX7JLI39dd7zxnN6WtR2gmtW4sN5OOVZU0wTbgC6S8TKrkj
exlPi0fId4qaWbx8zmx5rytdUrS1wddFMxWqEZyrchuJQdz+kV9INU24FRsu2qjQXPBjIE3IJJaJ
4tqDGo4JqTMIqhcxyslrFXYrepzGsCFj0NwL3iJ6tG8K4TfnspUDw0uhUGv2p25x/XpcmHnW/Bsq
/VqQTQJDRhApC4HfnoSvTLJzahrwjoEwpTNiTUaUYZeOF0bp5aYVq8RSd1viCJO2QCA8rIhHh3XB
87sKKFmxlML8NTVBuUhZKxZeBFHwbdKV8oimKWcADrOxENZK5gGNodq/HEIb0VHNT56AjMfJKS6R
IP2yOzw2ZROcHW4Rke67HXNsBoLYSLtEF8oTCyTty6b/7sArMMFIicLIfGc26Crz/S6qTmDsz8Ui
A8xz7f4l+1T2FCEgc9NonrupwoTSN8uB/N+2EMhOULSktUM/+oo6g1QTA0Thd6pKrhAJ2spX253l
D2TLZnaEz8mEc1lTxpnjldTYj66HIpc7M1d/wk00rp+9Sen/I87v53aQGGqMd/JD+UJdvfWw9VS4
Euj3kMcEqZFNfx0Z3neu1+ynV99nMo6i/8oGmtKApxdCKqgX0r0TShlFT127sNvyUrzk/GOiIcs6
WM8i7nYMCvClw3sBLLWXi5HwurhH0g0QKaO9evc0pT3KekKalIV1Xo8XgnrKWBoip8UGEjn9IQ5a
tXpmSjlTlZW+Ah+A84+yk1fx6HP6gpdZoQfbSLGXKD0jMa01YelJevP43Hm2EyqD3NnmOm2q3Of1
0Tw5SYXQ2bP1xDakXK667LO1/DKE3aEwlze4XncRlzcMYsZaZqliLppWKn/dwBE/ZptDQzKzdY1c
c7Zu+efEUUDxOg8Ys6HFjaQHHt92Eiu+2byLAlDHWAlZ9PAGbQWPv+MPIJ/wgI+cmrUBCKluctNp
x+UH865vFCOzTPiEhIEFiYgUcdySFCufrzSxsWo8N0f0sNlSvnFETKml+c9KDVUk3Kqu83aYsjdS
llk5e1xS7V0mOdd1mltA7MByfhBEC22Fze4g4U57SJpdmq5wpAhl2A1ADqmIW6zbW/kj3zZfTH5T
Jj0DCzYuwKNGWom3EuHzmpuMFR+AsMd4gwUQEzJaw9FMb6AgiMxwbH9teiaBOXdJ1fbQ8bQx1i2Y
YMtm6ZO7yTEJfel5f4bNTI7vy6FD4x7EQyhI5YdMIrM/n+DN2Nv9KO+LOzT4YuK+KK8FcPVOLlp5
ObO851nxzMZyBBFFBI3o3Wwo3A3Kj/3ytXNjf+vLYrg3bRxWpaqEfyRsBm29sgvz4fQpZAA9nl15
1laeWS2hUi7rsXWD9TgiqIJoEuZ+YQPkQ1np4noXGJ0dxTwgaT/MiB0mTDRkVES/g9JcpCTsTNRo
pPOcfnN6D9hDLYMRETtTYyxraGb+PWAyK9cfrCJmDT97p7OAWcdprx4xxWPfxhKGarHxGyTxsLg3
CQbmR2DOJp1WMJiBf7aHHKRGubdZ+1LF4ptxAO2YJNjx7XvqQJSBbSZKxohgK7No4RNqxNzzKcrh
2dMNha7eQIbGMZLy8t3k4+9E8mcazmNEl2WcHdV6Lt9sGmg0tZpR0sYHN2VbKOVK5wErzldkwZdh
ZWdP4jMxz3U4VZmo86V+JHyoFPHNbiChBpSIDA7pzmLmHaw6N9abGkvFKwan+9kwpzqju00W5yJ0
yn6ecVFi+HCyKY3xp3hlS80cy+Gdkq1qIY6BxNMu2YFyccUf2Xkk1/zOXl2DHrUYJO+QMnmTL6Ew
qQafFkxuIbLnEoxhys89pCDOywO0NOVf68DIC2Mcv3nOToQNMah3d4zOxcj3zUgzwUjNiCSdy95O
TFHwEsYl+iTgHOjaHqKhcH8qNb9Bd7JhZlkfCn/KeavZCWqmmFEDCoowm8gacjGLeUG2us62psfq
BQuROUEvsf9IbIlOKYZU99oX8MrxprFnF47m4nTqrvndVub15UAwi3A07lQoyYsrsHxJhoCPSEbY
oWvI9BqvEcqaqC3rIxlOP5JU9CwBwVWV8rKUkQ0fLWnsrSvSQhVrgPL4SzRMbtZU7eP3F7TAizle
/l7mGzavxuZHn+H3WP7SLWCKbJAVLwgkPLpt7p7wVpsgPWWuwiD/VwMgTzD/D+xhiH7FcfuHmZme
d9xGsSookHC5fZxqoM0ovc/7+eJ+ve1e6Z5CvSBFep6Wg3fjhGa8WPNY3y6u+YvfEQp3d1MHzMqK
yQsWC1lnISbUcTC/7v5B7SnJq/yuRa3LZQA7eZjPyWiihid9HHZtNxwR8s+X10xznBEBo7ByM+QV
1LggGi/mV9qgukyKXdkt8eqn5zVDteiY8XE/1lNkQoAlRyxA89qAyZotbkkJA6+8AlrBoJp6qkVc
cUz2mtaASOIqUpsulUKh+eAhbfTqTI1jurmXwr353DreoQVkm06WuHw2KTcLwLGDrQnr1F/oDDGW
NODBznhqrnt0i/BR271p65LMTaf748MvPvOtPRNyDNTIVYI9Oy9C+HWLhT2VfFpbVSYMDNwKnsEF
ThianvjAjK0vDgp/+SB3vwO+Sdpb+sel3wUCZf+E1UGciBzZ26+M3R3c/vtWSjHqBPmJzvzy+uzU
dVTLmBxkSNC4n2ICJPvDWT9qFYwji32yd9mghUis7Q4p598ym1fJN5hb4cGEzC5qRwcAYAaRjTl7
XrzTbweKi2vjgkWOHX8wQyq+XE4jJaK9TA9o1IP+RdDc7z0lZhhGAH+cqL3g5RsfmEC2iyB9VnZX
eyd519HNqew9sIz/zfuinpVd0wKVZCgUyTU+6mVAZMG6e98UDNRLSShd+MKuTrI8DF7oGQdnYea2
+YQZKB0lfgXD5B6ViR79hbSgPn14n+PE/Vu7NrxTlMfAUL5gEV/jA2c0niGZtwK7TSeqJol8IMPL
Ldgttt48YhjtCpFufFcCsIl69wHUpCX2xYQOZIFDoT3PDqmKA1RyQ0Jye6gzPu+xcPEZGtLC0oz9
JmqzyywmX8Jq+q/TlylGO/oR3visOqfISJf1UEfLb26VzTnNMUi8i5ArnCbYLaXoh/8jrLpQAOsE
dMNk7bFqn73RR7mMhewMnQRdpW5lVssgwN5IAozXCVoBl++5SgNC/KCrFqIhBgbpj+usIZb6TeQf
cidcwCp4hEKe6R6V54a0qYcSCEbjIjBB0vXcwaOz4s6PvNFNHS848CyUY9wlpbNEprrCAZs3N8WT
mhf+s4EElczyV63v+8mTyoOcgFec1ECyCV1CthGb8f2evQ1fYD0UEmU16KFESR5PJSloBoOtUrzL
BaQu2yD2W65RSsapvRZV+au/rNv8lgoIA3w2rUAvmXyaDdWj+1w2kaM9JyzXEfJGvcO6CsqRHew0
vY2vj/c2GS34YmMv2klzr49fZDwvO3ja1kIKcn/26EyexEZdD3egumjy9h3ugo7j78cdSRXkND6y
ClKlnYAQ/HB2rVDwJGUBcs7s3t/a5GuKm+DBK534crfXEL2UPSgtE5vi6ADRrZX2pgt1mS1Dox/8
Y6QnHwxyT2GLONQJezPOClDa5E+bfKJHej8QQFKgk5gY5TlIMD9Pgk6josgQ7FlVduyzES2hmumZ
WSoGwmf3g2lePAeF8EY+B8MLdGTrKU+gojQEF0ttvEJ69FjK4YArk2XMLcUFOLmPNvAMw7peoIhy
O8h8ugwwJNQEH8QOcpwi7TIE+56BvZ2lSMb88vWkPBhfIUkCfMyCTDMt533OsdVr6T6WIyB6Amyh
Qw00ORLsLRMvlTjy4FNZekbsoNikFOcBTEUv2Bxs4mk6GpZWEmxDTvL/6W5pZRRP32HEi31GgCKy
1dMaUGJOC6f/+m6WBcDcjz3Cv8IiutGMMe5qq834yvoqSm05SM4jS6YldM+SLIrzcEtusw5s3ked
UP8J4PizHGiumjTjTQiq/MTWu8ci2H/IK0V+V7dBKlpKcSFo48nDK4dcbSsgbUkyB9jhOgLQlGIL
uNmO62NRNExxKOH1M6Z1JKVObihZWrVpzNtPA2cO/xWJyqao8N0IlB29Z/OdmXLSAK7V4AZAuGLN
uLk9pntMkZCl97N/2epTOHBlLw4ZGqnMOQf/CphdJDOGEW1jQ3sI/xne8aYHWHDU355ElAL35o/O
tXCWj6Lmz3oBNr73msdvxMzsuHvzhfOF6HxVSoeepiR0jL5zt4e+lWeUuPDoLzeOZu/3aNXZ3DEb
AoNQWe5DADr3d2rvD+dZNkOQWCvu7+a2VZbHDpqSoBPr/xRVpnMhkhHm/Q9b58iemYdEBxI0lb45
MDyW/OTSQXlWmcPV6GMqc1aa9rV1SUUSvJur02r0VUVMjntfzv2qYx+kPyncYd0FgayzMaI0dKDA
TcrI27/lJIPaUuOaEX9TrEYdNBcD1s1D1zmStUfZyF1YK/svecIm+w33TUaSfQPda/PqCVqm1YL1
jbmFPWh3gX9Fco0F2PYdAn6P+oLfdLVzz/diW1EjWczcWoboz1hPVAqUm/Y3S64mWQ/6HRWS8JRc
PFQGjYpqJHavRGSR/4S0EoDEMg/Mz4qB3WbI3r2PedMDoyJnJ7j4HaVKUj2EElk7d7J9E6cCWpwM
Kkfuy10GzgeZPxoWbSfzyQqL8D0PnWQm+0RJNZ6qTCgispOB2W/hyNgt98Ea8O+5+tTPTwTvm16O
gHUhDULqCsTXVptK/Jto0Rq9B/um+mchTQ/afc+PS7KY3i+qcLaaYPzRVYqu8zl4hA8cmlykXoiB
B5UiUER3GneqXCcxmjq0q/PZ0OWJ6NaYOy/sIJLO4fJf+bzQXeqarltcxxzJxUo7rxPF3Rau3uJ9
k6Bh+z7p9QedFmRoGZal9r9Lu6nD0a4OmdqUgx+mMX4Uuf2Fk5s1marj8UMs1SCh73EYO0Rfoeaa
2ppoaV7Ljpujei+Fe41EPJ6D/DWcSASlbXvG04/XaokO2ginMCP9bMb4xhE3tSjj8cO+OR1n+7U7
+VDURV4X/aHtO847dULv9IGDuEFGzup3nd3/fZtZuHPAvtTAAVL9ZoayDD+kVdSgOsTJrbLeT27U
DB0VJICswZY7n+tI2KlQQsMCR8x6aoc74qpEiYOsZ8ARLpe1ujsOObC5AnT75XnQ0Y3beFbcQUoj
JtPolUmYgZ8Y4kowgwKffNmgPcWYbFgDGcs3LMeRdSyn3eIVNVqGQP2jhx6nNEUfGFR7xTLf3DdG
+sA8VGQDiLgaLmUGiexmg0I+pCIcc2QAJsHzJosI4v5S6P40Usfta1ACfpEkf0JoNwLEgYpuaIem
B64dTfVjZAV4Zm/g1P1hmq7s6ePoMK894AQviqM3s483uPyLLyjoRUX4JS34CplldiLByB+utzCx
mbUTY5iIWThyt9D1WNY6MFv4WWk5m12Xqq8/ICx96RiRKAXwELvcTCpA0iVqSVDArrALONNoTR2Z
DuVG1UnndaLB0j5YOnppxyVP4nLCpKHHbdrzHDsW/KEzfvkdgn/KQ6d2wrkly5IWdqS0CCW7gOdm
+7PHJ6PgIUXqWNnKAB4sLSf1wR2iZbhGb88JsvNVd20XrOvrQO2/6Tuh0vec0erTF6XmryPPY6FI
WrZ/wnaljKk8qP+51E4cx7thzSi7jOqTI13mZfIsqCF58aSSm15Kd118y0vahUmWkJ2wK3cmQeUZ
J9zvcHnFHz/S/URlgSHiZB/OSCZt2JLyu9Fg7VsM7pR2BK0/x8hXcAoiYCht/tG4fuAMLrTwkBBn
szqfoHPnOt5aj2JnB0RVPDSTrx/j4E+o/yNieYdnatRv4fd2vJgaWziwaHTnhkSygvEB15X+QSR2
sBz+cSjjIw2/tBC6ZXmTr4ut/IXDgR9W4k75uqthkmVUEAE6QyZACoIaa1Q61M8sZhmI8u2+bGXi
PwIOgorLb6XwF0DpmqyvBiRFyAU0ApzxootKgPa27tuBX95/W+/N9dm2u/UpBXTzK/BRC7Y3lNgD
EXviRkktNgNAK8yUGk06G0F174SwAYlxHE7UJUIb/9UKPVPCqv7nwOjylR1fVRzCamm0b1N4iQT0
G62+2h4xpEFt99PNLdykJPPBqFgOPqAuMI40wIHOz5YVnnVkRqJG9WXyyih//Kd5rNICn2hU0Y1l
6Qj3YvfcEQR631iyXJdtiNc98wLyLzyLJUq+RaxgSUHlAU/z4uqKXrZ8WKwR1gUTSPpuO0We+RKa
e8AUQdTy9s64inSlVnBf4qVT/5Fixd5rgAeocZpMENLEcmL1hVX0Gy/6kZFDsTs3AfpaoWJ2gZbn
+8pAjwTn3lCUC3jdJbNkrdvRE7b3qa7RnlKTl8GyxsM9PSStpzaiNEry2fbdv0VOwG1oWZxAoR1E
T/6TjRU5aZbNC3TI5XvuOuCvuLyZtC73A+Qz6La5aiT6SxTF9WhKwpNcowx9ov1hWqS1rzpia+Cl
NBqHmEVep6Cl9q1YbAiLj7ZId0ptGCKwXgT0Qcn/kivolRMzKidHXsIi6vrygLS81KdBXtXpEyfH
QNF8mYLpFu7ibslCThz7XfzgSlIjWOjDe0TTtoUf3q7VlmEqoHyLAJkkRSHQ/Vk/p+75e41fqddm
8aJQh2LAkZaGsyfcpnTOQf93GMNlbuArbMyS9MzVLqMKBmCgJPTC1UVp3fWR4EHJISi8vbckFbq5
NaKrKb5sqyACadSXnCgfMDq0NZBetUYYFciwx+qUrXOTuXeg4K4xU6GHV2J0WgTQkBTB56B33ont
+VQHXkOPy5iAaLRfVS+LPfMkm8rEevN7kbGdUVEQF16cXXk51x8GaXum5rUU5Pe8m36ScEgUeRKg
dqtn7uVpt9w/UkjKnoc5lnXwUVTmkeGnjrLvHrpfEXR8ljFihzGU3RuMRhaQ2cn8BHKwT2t9pcHI
qZ56Yp4hWNnRPKOjpIwqdUxMKoAZy+SKqjbZCXDi+z00+lwYPYWNW+YTAScUxv6ySiwUXZvM/vdY
zNAI1l3vNohrJGc7Ap1cx30jFsdqrDoHgv5iW8ImK/4URgJ2/h7sAJCPPtLLw3jRj3K7oplPrs2I
maE4+GnIYftjo2bbXuHi8iMVKPCS4sGiUC6wFT8RAZ/Hs7XO1T9F0t6t6DjBomus9+uzjRYgmXQ8
vpVF6vJ6YqNBX7c9Mx+E7jYiq6Lo6Cl7iJsniU13mKZzqBbgffdFHgOs6LV8xk1dPtp/kEzkEbCc
vdjggWRwxpO2+TbbWqBhLqhixECJh6tRYHz0tBzQMmkpuBShdm2QidqzqkYPfaiLD72yvrPj27af
5EoDW+HVLQKmdFmANzty0FCwt7LXmbYpku13aVEHXPzYRV4r5nVz6ol4o3sG/ZRkgerYd0Rhn9Ph
4iwRTtyF73lJ2Cb/D4TsgnhLA90RS4DttW09kixAOon5UF65ACA8LNdo84CtIGOxQ7zGMDsQvZJV
Ztr7IPsNykrAym+TVpd+LcBG+DbfzEpB4PRgoE9gVR+//FxLDFuPDTFLHO8az++BOdVb1ySL8aGL
sdAdLzYcergcRwBr27UCyiuQvmkIYvvRMSt7Opt6Y2bt46BnYd9CQ4k7+J4mfsegfVy2PFIPLQL2
likcd+/Iktb3X6iohEohP3iagCxg9Md9tKR/E2w5yXbJjDKASzXwg7IiKXYElm1hG5+MZNV/J4dh
JYPdlezBmPZTMc/3MZV/RbAEktRkMW/hHFy/3V1D4DnIiDw+QK1pnrVvowx0VwGQPVlOJhHiJFKg
z90XyL671eA32YCqpfW4foxrZ+9Mtll390tqZn3jH+B/dTMHoQ3Z9B46b7ExtSKxSZ/NHHwrJJ7v
/wcmGrEB+QuioR4bB152ld9SxKMb0hhDqABGvsq/dc8pi5snbVgNWRFsEtP9hsBYZwkuyYCuo21S
0Vz/ZYRMYhco1H8c1F1q4RfLEcQvNg+tbNFc7xD6UIFsby5CGwvc4js2SnQqK2KAmLY1lK4owYXY
+68QMUuwo5STsuBiAqVVDDo+IPFW3Wh1gxycF/ltIg/4wQHsVgfTnaZRWTfRVmFkXcVrIlivEDsf
wceiDhMDgremMFvELJBkS47fKj1/kQMAbP9yf91jeUJsZJrrmD1xKQP5ksMtb66LS+drNAuKzd3I
W0NKS16WNZqOYDp3tP5urfcyDY1ZQWXjzg7jz1N+WCOjs8kfb2pvs6cPoxns6moodY+0Eqvr2QrQ
+KZGZW2TSe0r6/spSotnt8Xdqwnc1ne5zvqLEFdVxLp04WAXdteTweJs8nL2+P5VAap8xZzD94cW
ogMI0sdJlkQulSPfHIS/E+88Bu2sUjV7Yk865E/9GzDUQBnNq59ukmcRdP0Fd0ZkuWiQjE9oRvRJ
y6EnsKn4Evhcx/3n15+N8PuaMvauqNPSoAtOllp8AGHbkhU2aeFY1QlDDiGegOvDenLRmgapR7Go
ES5athJTwgrQQuHjIxOwdbQCDY+WaLWgwyQWR6qCVY/cZL6ImrQdK3xMBX2lwiV42gWVAKp/AWjF
v7Gug1Z16T7pXoy/CxMK5SAvaIhr75NBpuWJ1c/2Lub7PNYNxs5HFB9Phd3ABSG/zPAjfSxeqwgP
WlcKJ8wGumru9E+h6DzdhjRsPoSwTtmApURDsvIjyxdjVtpHuDSbrwdHnk0lb/7ldrRmzlNS2+MI
v5kC+OdGXsmgjQRzhZg1+D4pTBokAFSZQ4dZst8kXAephf9yqfEA7JlqK3l7Jv0/pjFevNBQa9yl
KgsVJ6BkY5LEUdDqyh4pL7JdbuAdIAic3IDO9ERqtNaMWW30WKekIUTBfZdH5VXWH4LpJAZZcjto
Lm2uPVvkYwGuvKhAY81UvXZoau5vsXVMmSReSsgdzFhdc9EuUeuFqjtxf2/CmWiljsDnv95emj4A
vBA+s9ZiJIo5weizqDOi7QuL00SnPp6WJmcP1foFiP6R8lrd+lH4Hg2PCnyZ+dxU4crtgAUMc5tm
UdvKoq5RNR3KPcot8H6uQajm2VKU221wDWMjJ+07Gjxg4u/Nf3IoZwYvL1D4qBf/3ogV/Mrm6G/o
RufovdA9puyvBSPo7phwNdzQTvIEQodikAChRN9MKEhF0qK8D4n+cD1GT6eP/aWMvFMkW7yvPQxs
pUHUIfkx4svTpfqmPC21KoPd7PES8su5soSDwvVE7afokTI8X1JbYlBMaa666OTBMNvp+AWy1joz
DWFEuoa61PHSP34wxUHs4wLLxjIAmU60Zespa2JTGMzA5G9+5oPgU7pja2yvcAS5ISmCAtuSQFtT
KWoRH4YwpmV8tOvtiwbInJR6m3g1xMcBRUf7i7P+G7I8squN1wdFk/9VQqHxn7RUcLbz+s5tVT0h
efcPN1IM1STkU2fLCklvaQkzxIAlr54FpuqcLJLy5Zy8u8hb239wPW6Y/sRqJlYWYXj3llBYoXkE
fxbgR1sDdMGG7JbSK7gtGIIEEStKvLkrm0ClfrhKZqdHdq8/5utNYwskHKg7clnFWAsls0h/wjFt
0+ogFGSOuLHQ4y87zrSuhktXfMay7+8YeDEuIoBpXWnjYlFIpWO/MRsGfLuA3GSrJ2YUgv6JSdbi
HoIzKf7vT+npjm+TcdzBYwpcJIxbeCxDxNA1g6Tnk4F1+MD4oARM8QC7DbRU9AZsHwFsltmCwTHi
3Dmh26daCb3hX8RZqpAi9sIGllTRPBvhs6E8qsNsFPGkGg8S+ATiGV3m7mwW2HHBnMq02MU9tTk3
ETYVhPrTC6ZnN12HQ1KKVEBMjSxmt6Ar5d2MYG/A9jbWEy0RpHOl1AeRdAb1z9shz9uvVVZ0yBKT
rIQSiBkwfh+VVgkuNZ+wCBBjmd+JUx4e2qX/Q1pjxHqnUOULXhqWSUuseZNRUiy89TkHsyKN3L+9
SJsIBuSWZDQeRtjNk7h/xpvN5GNWsUnS3SJrkkWA947lbk0+1l3x9erixegfg37WT30SYb3pO/d+
ZdAy0kdewmfz7r+dRNsLtE9orl7r10G/URFVlpA9Ia/vOq0+p+t4SMVz3atxOfhrWUc14g/3uBNp
/JFVsre419vf0CXL/5tTeS8xM6CECkEc/0UWnX3I3CMGkjFBrH4ClKgwccyAifbEzSrS04RLt3YI
vQBJ6YF3jADWwUkQmFRpmBw85X/OaLEiao5wahhneTx6GnQeSooLum+OmCml0AT7yzgR4KIW53LZ
A/X5K30sAFYlTsfEts07fKJ4vH1tT0tI1SNO4/p7MIxbdHkBgYO2QuYWnOhcodYN79ZLWu1hPpb5
5FWo5e+gG5rcl6oSadk3V/02oR1ndAefrjTkq3eEJ0ZwavRmJwMi1YRzoYnJPB6vF1/gv6SVJuss
t+SeajiBfENaML4DZz1hcgnABkECStG62grceN+/Xo+52UsXTr6gDruILCfQm5dwNZypOmpme0cn
79iZvt/Yda8bnLUVIaesICICbe5U6LuDNrlDKWY0Ju72+kZJgG3ErJScHhdX9HmGYktZUrnXgVDK
g3IxyLYfOavK9W8zpr27vgaybrda2QQEhAY0UVuGBZRPXlZK8wOoMtyJwKrHlqVOuECm92d5fQxB
S2nI2ETGbqCwHLyACd3mE+OoRHID3qgJcQ83Fp2c9ozYNjI+9GA7RVzwpo9+aN8tr2SqBAQi2ia2
DAtzY4csBM669B3OT8VWZpHqTh/pURs17vO0B7PM5hcp8BYV7deQ3neSTFuJqJTIHn4Wo3Ty9NOd
3El1V69/K5VRBGTFZY6HRZucZN6sh9bOd8zab4TayCLAJ2Qc+R5lTqHknUnVkNj4vTjvSZBr78yi
hjjSkhR6iopkKzVWyMS15UTYDVg9NYvazRi/gcJ4wI7kjvlx6L9iMVf3MnAs+yd2xJOv5D8qi5Bj
C85RwiNJHtfL6va3Wxhl4R7l5noB6mVR/PBiAnUOzyRpOSFWYvMteI866So/dI3A7KBQcThUhUur
WBqmtMUROnBTuPzQ3wMT177lgYkYR6kyp+9xi2wu2BxBeqD6pTSDUvTZ32uTua7eK5CXHQBN0nUP
cV+WmvpBgKC7ykhTFH7YhYAPr0vKmPjQZ0hRUyS4Q5KBhwjXmHhc2WH3ztuxdPuG0COckm/q7ZUX
CDMnAGODvFqjt8XmLyEWNfBkhUTE4gOf8f5ybodpme4fYQRjK+Fr1eHTu0NFyknOuCz72qf7z+xf
2kLvrhoWqd2CQo+r9Et1eLpFfcMbY66bPuesLpxqPCLjTeuo3AMaTgw53cx08AxhhLDNgrbg+bnn
n5pzbfK9BVpA+uq0Fttc5RCc+gr0zkW9n+IkSCJow9LY4HfjbNh2j+mCO0qutrfdJGh7sh/PNClC
vO1xhWlLgYL0zBxTEcLNtg0LLAVmbBqMfqpqmo3K26Mv/TUFbUt5tIRTdsf0kAo4jNKz/elmVFZO
ZTC4vsx31Yzad66iA/SSm1HSbhTwhTRga351Ofgf+I7OAHrcf8MIaiM4H6/i9RuD9ZH7OBgNIjUU
S8OVNhJ9F/6Z7+nyeuUMgdPnHFKLHEMNz6d4ytHhRANOfFky/KagLX6lysTES3BuXgaT0q1f+0l1
XRln6dU44Xus5oRxLafN01P3ssRsOM19GctUq0FNcX71Mg/vLcsdTmGe2WNJbWlDuOHWqFvAtxEO
fqzf9Wa6h+Y3zvmCwTo7E3RycsSIdpvQyTjJE2ipXo9WPeegx2Q59s7uCAobpBTGgz/vK/FInoag
hJtTtwvYPOZTozOtdSRcVZo4YaTBVwFgqylGanZHDwFVhgzHXdgrTPe620FBb8r/p8PDJMTQGFYd
rK7h+/e8rUWQBM+oMjCnd/Bj9GZKPEZkYAMfz5xgymPlDJPfOU+6x79/Avu2KbaDXW3+odQsjLm4
ft8znOAkxWl3zHuRzHtDO6gjCOfpKUDxelqYZiIwxvAIY4jr7PBYASyc0jfbGQBP2Yjn4WwiE8QL
C80fUw05RwnxkfH+mRwlpDjhF5m+6M1I+3hfYfX6S/6U8PwVlb5FsItTTjTha4B7AmBwKuxFFfXe
f9A0azXD3hjJcQoZNBKVIQUEi+WQXltwBz9lZCHTuZjyEppez0AKK5e2c6AVCCTQfTwoBargDTQq
EkTiFLqaOiAjmWFVKjRfbLzwndWNNs9l4f9oJxiMfKeRxZvEN4LMiaBCiG4XX8okV1OK95Jg2sHX
+fOj0Pg8rlw8LbnVVbWIiP8GZDW93Yp0PQBzvpP4j6k5qk/5z/lhxf/DJwvjnV42IA/XRBO37GfZ
nrpsOxu67MIr762/uGMXvDaGagwj1lUjXpDNbQed1C92YmbfLPR5VuxGhoG9SJRZqPNN4w5UBe14
+RL+80P5CKzJaPxXZxlRX0XMSTWiSZLNM2eBXFQmQ4QyjCpaJC0dbsC4R35FdcgH7JV516AdjXss
1s8mITya1Ajaw7PMuDhUyhwp7cHeyn+jOYpFZhzE/vLazhjhAWsT3joTW3a5KpOGLLuRBno45WAS
qaLyz2VYFUe/AcgHdaiSM7HCIi66FKisODYNTzSWmVMVSu9jJUEDN2w57gnEZ8VB4OFUE5DFtFe3
OcTKiVzoWZ6fREl1INPpdSTgmy2zMITFI0cvENrZujTsZStmQlKBWxfQtMZ+TMKTddXYqmnknCIt
gMdpsmN/KySAOiSgEJwtEO8lWZIoybp79K8orcAXKJrQu7uEuHhhB/LXk+F9W9Rp4hRDrgtOLPSq
9NntScLsOT1PpH6ZBILklZzknZ62QzaGKKxStSEO7fVM179c2S2ozo6abye0bcKwc7cox++DoAF4
yH75bTU5NAW+KVOQmzDcOZLmevQkOcTmJbkGj5Ek2iwB7mFWbNggwITBq3fPHpiVODfbDlegGX53
wI5jRcN20zx2IlUMWNOMWRdLSZPwEvFgehRnEf9lX/hiL7O+cRnWz7SQwrLhNN3wGtMR8bBycOpY
9VtljqNhrpCFOpmWxeUBu5prQc/maRDRvG9fdgvsjjVHxA49uybGDWCA2XBKn57+h3LrC+84iWHC
Fl5Lxxt8nPX+vciBY7vnlHMkDP/sYNjfgMd+1TMcP4tHm16KZIRWKaGc0siRWaOhWLich6NaVMYL
8Pf24UtKruspKLUc8PUofBA6o3Wdd/4lDAOzDbL156pRvXcAGc+rYE4W6lqtr2/PXecag5J/NPdw
v8Verp+9SJQSVvkUI3nU96uW0m3VCribSIthDhsU2XbBFKpLVsdoZ9ho8rNdl6IgbU7J8OReTXxE
PE2x9e8uf28c55LiaEn1Hc6TdNbtnk53wh0b/MLz22QDeqyPO+Q37/brcwGWW5/ao7vFnrLQaQFx
WY98qMHUlhrY0nFuYgvJAILZfFyeYez9pgbMAXlbYh63lqunwyCrRUm/x/2WWtcCPalsHkCqOOgO
RidkkPWrWc85iCQD2J4Jw2mZTr2Hf7KHJgp/hTVvkt1mjAtut4+9+JVPpOCTJlrb2qKPURh7MTSc
io89XzLXwouCV8B73/cvrOPhNTbHyMzaz2pKhSG0gO2uqMwXu8LSHJM/z16YGND9CxmSqMQR6FbJ
rs0CrinfFIU+VDu5Rwz6BMPZUOthxTzB2J6KqhCAmNTmmXxOHx+rPLAhqIWWvKIGCP/1W7EUaPYI
lQGCIDBEQ7EaLbHovB1OMEfIJrdwifw2OYc2aqWV1G8c+3pILSp2FZpU1Mf8g5uQ2EBO2L2LGqus
y30gJaZpoaoA8fq2zKc5KSk3eNi3xbj2bICbDNm7EyUVjyRm6MZ4cCYYna6o6m+8QP0AJCnOJMpM
QPzWMLPbCVUwothSTNS906djOodwJ/YXY5gZO5UwAw9HHKZ33BzFBVnf2DRs0h3i/zgTACe+vIjQ
W2DIeFMqzJVbW657N1Tfy8FwXUBm4o0xAGwfMwlJgWcOxZwxuIvAep08KwQHrzz6x7qbFCIgPQN2
XOc2rqwjDsV7AUcjvRuvQNlK//4Wh0WAYCXW6GjiltGblSsjjNEgQr9XRtCyhJaaEpcYrcmQIfIl
N5XKXpZ4YM2J/MP07ZqFPQhNZvA1UwT5MmyZrxOMmUSBgKQJ5vgSSILLemmv6VR93JtuXEkOmZCn
Mo+D4hKyosHwh6s9L4L1IGjpb1K71ELR30sMwk2JMs7830y79ntQoPDdmcq+owfflxEURneripFb
ygBf0FXi+U7ieGtprGSNndIJ2uIHvMs9ywNMqeGmhBLWhTh1Ah8Is4HivyrRHjIbtcz+9BqFdy28
5fdENuye3mdBiN3wrYCDNHHcyIhfmxGcr9WPw4/XAbyHOZjApf16IRhrBI7X3KhFg+N6auZ6CB6c
sYItk+QGG3BORpAKf6czbI+3NS5jvurCVzgq8eZ6/Wmuas5qaLBn9VsF12QhoaIS2F0K5QjE+Zya
1qWsM0FUTBCgai7TeD8pfuL/YtSVf/1Is6dJuuaAmt7dXdqBpRgF5OoaSSOmaGJRizkt8Km8xAiR
eAW1AFGhxhGcZ8hdVXrnWc9KD05HF6Bl+BVRw5USacRxICTYaWDp6SqPtuDNBFsq7r93cXC1aM/s
6ZmZV09gM0vfrDTiXOLklrT4Ety3T4AKfVJfD/mCrfcB19C0qofy7N6GoBOFUIIKsETsKRt41m7u
HF5BqRybA+NqzWHbT4HhLCsK+Oc3GlKrh2YpC09Nm/AjyusT54WaeW8QRBmpSe0fhgNok8YKBhHY
KWBNiaP+qxQZLyvGSGs7on/vECyB/6pvDXjwvpXlZ3o3oFWQNaeTkFGNAqXd6HUdOiSo/G7ksCcM
RpVkHZ96XcH/nOc4j5DMVRCs9rb5ga97GZ4UyNX7Q+SeBTNbRxB4Qi/itce7LtDihpMRCDH26YRg
6cxntOXangRzLs4zZfR6BpXyjzwjXzg8gwvfX8GFXKkh+XyEfHPGn+7sgurhMRxIzorg8b9VdmO7
y3LSAdld9ZaAtYIpT7QeIQYgCLsnFaI3wwMMj0L2oChJSBF14txgutqYHbw1mBoQMVQIz2dHLLwk
On4sgAaOeTB/CS6qIoKyEeM5TxeJkAvxhKPEScFjxFUll7ZL9yNjPaHA42epmXXpFUI17W23N9ZT
LMLrGekuUj5q9+q8W1eK/1qAyNNl1V8V2yRoO4F/UB1zmyc8gxRQqPYXyVRfmIik90V0HD3I4ofo
RVsVJpkWxD8BzHAZoDYf4bzjEn5/822po8dhiYzczm2k0v5LK0RFHZtmQ+ZEpEDegE/BOANvFExE
SeQYGwydPsyHoOyno8DLTYH6wRlYalUrFDdN7JByRH1aWBcdleOUoGD2TivgQvSNK3raQybEGUhy
DjljgjJ13Ocr4mcowsLym/z4c1l9lbWhZSx7DdWAOVZ+Zjgk5uebmG4NfRwNPshg9wQHS4LdvWS5
ZPeJx3Ej7qa5rvHC0Nyw+Vq83CxiR0PK/kxqVNv10Z9kSeFEYDPIJvJN34w9a1x81/PCXbGpbg0t
DPY93XFqKl6sVBICL9x7d0SvcoeQYGnAHjwH+PZB+2dZ46/9fGtWL5O+ODEjM07EUxGvVtkKCost
jtY8N+UG0r1XhsdwFV+0L8aXDR9DAtg2YTsMJ0mwg6tgBkZ+HyXnRryMoxqZKoYuXxo2bdsvIfBK
ZJwNT5lDnlFZT+IMZHg/F7iWXJ6FXdsc1wnvl2Phv6YTcqzqHJnNY1U6DxloJ4tqlhG13NzMqyEd
QlMZm8sGpInjrwspwrUlqzURBTC97dL3PhWfl8vglHN6T+9pmL3ZgvCU20sKSNgpCf53qY7d9b/b
WOMxBRjl62QDDMXTa/aOn02Qfej+zSDH9Qr8nMMa77ncNxz7PLmpEDbVAmQxRlk1W5dtkOdJZ5j0
ZAjI+r3wJVxX73FTW0HguY5IhkIXJnd9epDkkPO62QMhz4pmBszY8q5A9GikX/eR8ilZ3ytoBcdD
STqYzqhrmQrpvJxNqwJ1tznwPKMaFSJjsqzqdq0LlRe2bwqJB7nlgIK9HHj2HpNxZikn3+HogpYs
aqoiA+EfikRXSqO8MtnUrp5jVFqlFUiJbK43vJiI6j4GDBKqUFoYP07Ns4L94DsLq2cDbDvbQLtL
wl09x+E/qUwBZmAkTXgR5wf9UCYpnTX4QyOdml+tqUKpZjMgKVML5cTxWlgfZD3MwC2aHRsWlKYC
a0LBNP2hRSAnCUA4jpHjQdRmiyYy8avEv3KOmsk3zgmZj4M6h6tpTsK5LgdFSid1K9GzOY49Y0oV
Y9S9ZpYakWOFC2Zq2ESo8B8iP2LjYZkDe6iFEaKlohX2Ob503ezed1DviFeAsvvUWzWFBRtgFDSs
Lj8LVe7YdOK4tX1p8EQOzHkHPeeHXZv3Wkz6YlyvRLEcQ70i5mq+DIlGfmL05sTK66wRc1n4lW1V
kfF0u632butijyjFo0JNW88OR6F7ufZJ4vhJEGFYmYxZ3y+HO0pQl+Im1IJSPNJ4kU2jCGmDyl8I
FcaK3oFUwrB/Ch2iOOvMualkB1TlKyBfagQGMcfaz3533zvH6pwAXVHr+T3EmNBNiyVbMUPfJc2g
4Dq7L8yqaYz2kKfDljx9xcsJzV5inPzuxMp6OhfhlyeKdfiBjNuxsmvbZJH5PfZkMYHRe9HPoC+b
itB1q3Nk6Gg6pStFB9JtVhCJviV9ZR6nPcROKvGmHD2KzhMahgVA+hCdAW+LcDx0EjcAcpzpScUj
mEaNBPVpbK0tgiS7M1k107+5AA/TC+/JBg6F5vafjDo/1Ek9YcszeuGRdCDqSAusxg19iFH2RVvn
RinQ+rGFEdnqu1I3bJLIn3rm2UGHvjdC4ZjTf2aLF9pz2WJOwUluCKjfj+JdomcyiSTsawVmIYvL
Ypd0cjlgrvLhLLrvqFLkU9iPzqDhPHeeE2m9GdAMBw8sH34K7VKUCh/rgwgBO8EEEkJJCMdwzn1Z
bBfbyn3lTXCPBeL7T4GarKLf2v8KhAkGoa82SSaYMIokUBw8G0fq1HTcd3nZSGhm+qWtAPsQzsjJ
JGIHUYOruAVGfXLaixJ01ntz8a53pKgYvNGIdnBceo/cJWGMskcw+APzJ4Y7McnqSKWnS/r3Bb7Q
OAcjIdRqBmPYG+a7MNrMAlGpJZn7xSN8pR7bRrKp4htJjiQKpdAqo8bYD7+E1QDSAfVJZXjj8kO7
C/ROvSh0uBtk7flwc7XoL5bIY7UFaKRNUHKdV0JFji2HZIIkn3T6jcsNX56Uc5glUlXpV8C9vMl1
pS4HdD+yFIVyaI8zbOmV6EMOD2JUolFjHhRm3pBYg7M7vpwcdDwzc6VxWe5M50BRspWRjDY7rMe8
RYWSjs0hzilOIApTaBJzUgIWEfvsH0iqaN7gX/+rrD38D5+EJGzY6oQR3UNZ8seXJSrQGXVQCE7E
IMBN/iETzU/m20HjsGGJ1OvwPgow5o4w2odTufrypNv9rouYX3hFoA4xPoUFrHZtUt5NtGhFQ2N8
dDK1AAE2HMMiDVL/zKU9pxjVZlQ7pQAU2lggQ8MZRwruMmL9VOkhs/9BOU4CJl6H2ahIcEM46X/1
CVo5+JbTeabRcyJ1A1+Uuu5mJYlPQ2BlNaIGnDBIkiIG/o50pKVxxzrakZvNXwBB/QTZIJh9q7/I
1ARauIyedB9qI+JAcna2lRE+p1IFleZIDo2CSJ/xKUAqUMFv/khtXkNVo2LfrJInQI2VrTiHsrbu
at8xp4n/YlvhkOq5iYM3T2Ct0CE19KU7dkW6X4Jpt+Po31Ix1evmNRZiZyNl0UAqIsq59S4MXjGx
FI7UuUTDf20o8aQNul4fxaxGC3apXtmSfnJUhOgGIg6y8dWmnzalRbHQ5YpYd5dQ+rGRd9ydTNG3
I+D1nx0rlIjxDZek8wGc22vMErXcvv83QOQCRwOWxnZnO0n0aSx5p4gLFL7x0C13hM+6dmJURI3n
dQz9jzCyrTsVCaKrmxE8Xf45NSh6HkXovOc349eg7aD2YhAEdlH7aleM2RwfgZeevydCIkJN2WHs
fYXkgR+SEyPzBq+hPOzrFLap1G/9ESRy8+38bNFcWW12CUJ1Z+iW9aQaRBfbDBni4QB36kilSBjI
nGWXM0SkEkHYF6Xbffi1XCqe0T0nNQC70pFhMecrhXaTUuvUfWmvQZXMqx3EuFZJo99VNRBqv0Zw
23u90qe92Xq7rX1DCGtsKAlBqumwQs7EORwBQbzHXMCvlA5X8zcuheO/x0VyvrCVU5R6TdUxxMo/
SfUnZG+6p6woGUjyd+vKGMU/MBh9WFMkyRhtPR/hkPo5zKg1wQQkVbZ+8G6UvFzRsPaPJdphcQ/G
YuPCD2gim7+iQ6gFq/4LLj5eLCuaIQyCUs1hgNJIddEqjdhDr1rfyfsGdB8Yfexi0t1HiN6V99aR
TM/ZIB7ztnQ14VhqX3DRztoeA4UcCLnifkwBs+EDRZREv0Eqd+vK1aSPmGc9f15ViZQkOrAUq5d7
RHdz34WGg7GhCKnkYLc8AMobEexrDtLAEb2gJRxPal1OAbZQ5HZFMg6NpX/5yu/9gRIUoKyRIEq1
zwbb97x57QQWzZzZIbfn4+Q9Sca9IfUGDJB3bVN9+JmyIrEEGS3yzr1JS9H16G3bqN5sO5K4HP/x
ay1CfCXqLwP7Juj7YSP2aSceniEhPGk9pxVf/JmZLZ5FbDEMqV5XjC+chCFETh/fGBuHrLJjQbsG
DX5J+qpzm60bY0CRmflH8RnV84X1WokoIUQ1Q9l6AzV8/ocHv1hTlzsGRSbQ9cbLBDRjFZ2eHGTK
a8pT2GofATSJNboosZwp8th89+QrxFuW6BsMlvhd14+Tjs7yQGrVEizjwFPyJO72M+6glOZeRJkg
LYDKVMHq2Ftm1orRHxtlpEhPRryeiuQpCiLkKXTxUOLUSWfMxe/GnNBXrO0AU4+JyG+PAjPgkdTf
z1Qn6oNrIw4DvWtAdLd4rQJJHXt3koRQTi3fQo85T3WCwfb831Risga0vNFGqF05RbeBbYRqSowI
OFKKJF9BtWblNqwQ7guHXJMSSfT860SA/VZaV2WGstuuUV7IJ8boitDPG2FUsHKc0fWSGSvN0J/G
wC12iHNyXwEMTVYMmzVSR0hBYwkZvcs9FYXedaDde78NH+nJ710s+JNK+VwEHD/PThzJPcJ58+RN
dGN9X1ALWNOQ5h87gftW3KQRjEmF8kwEzw/nB23wJPh/HpLcgnUdezjV30cgB9+MwDHnCqYf0nwg
Ol67NrSC7N4fsfKJlP/uA9qVMipwYg/ZCx5PX0up0OE7rwMZVmCutbZg4ptn6ej1WsFMzOtSA6/W
l2LAKDjMF4nmyAfCCacUv8+TRo3oJTWd9TKc9bACx3OBhOFk0pmLm6OJ/z69b6zI96Vz1oOtTdC2
g4lL6FjSY1h7g7HDMd95FvBW5cWBCwHcN+l9koj3BIOB0jP6UqY8RJSKUyCi8G2FZIIPhMV3MW7p
UjlceJa0SBvVYIgBgFhAnIdjivhzQ8SwUpjXgflj8Lhf0nmRVlX5+QXJy8SO/4gCanmdlffy5S+D
6WY1Qptx+lFJ088tsooHdL/BE2xdp9pksIRmqMXgjnNs0aiDCHbfAHaEco4t0FBPDtFH1V/pPe0i
Fj+m60TCOtmKghzQlFhXRChfMZt992pup/6l6sZrWYcz0uAZPrCgKMAKAvb7vrl/w4B2KJK5uqOs
uAJhXWanazp5O4hO+sn3UaLBrrgI2yaXUhvOQKVec33ShPiNAM7gervbcy+Oo9NFQ0DjEeRpKUT/
/59wbFJxpLSkQv3pSP8mKEfotBTHuPtnTR5iNMWxFzhVPMmjaeaEfSTZ8vvqW1dAWm+tlTmXthYK
Wo4Z0pKx9xQN2kGJl98/RpSWmQv+R6nh7jC81wEOutcEvNr+D5H/QGYOfXVcHMSVESikIQ2OP1Fb
cWqkjm+yEbvx+QXyCSmNKYQF0581x/dhduEUxohD/NuYm6IqisBI6CCkXNqxqrsXRg6nYuM2DWXL
maizy+3u5ZAOMKl1biCs64IE+h01RfcL8JHdWECQ+E8L7da0CoCWw3puw8pBNp4wWMv/wANKVPMF
GJPcsgFIqZcoHzkatMVqEWV9zP0UAVt8eHRtc1+w8wdRlJ00k3i2K8MqwpV+uUcgc6O8pIuddcME
evtjFE6EM8zJPrLaabf0us/wC/p4/RGqIV86WXCT/cTFT8Md6gBOPaaS3WKdFVs3WCs9l25An28L
maeIpZmhFIFD3dp99JRKd3D3JRIru1RS0LLKjkzZh3v06iq2YEHVYn6YhoHooauIv2UVRAZnSDOg
lH6R8O4kVegcn4b/XGJEPhNALN+a1u5anawuq7bqaQT0BUuA2D3yHECLCBqOx0gNDCNm4kdfHluu
/mPmET9rcuOYwJcWfHN6vv1U3uubCSK3AfwGis4y3CQ5PeFbwK5l76XFYdho/1QGYVhk7s+7a+cR
izCOEk/m6FGoFXkcHcCshBDNY+mgQA77waAyVhu/jFE0vX6bhnXNox958i94tuP+PNtvdrx1fgEN
xNSzylI94lEeOj7Rm4/cyEOX8InqEdiw7wASmZu7QhTaei58uvtnYdAX2QuVTwS3hmNUaeAOVqql
toN+YGdt01L+CIsyGs1bbH2tXfD3nUEoARSaJkqW3bLEB27DLsTMTDnzEDhcjYmjRiK5/gfmt+6t
k4/J2OtOO2CauLLdvGX8OVl8I3KpIdWaagl2XH5/0rjkzh8SOE62mu5AyXe1CHkQHVF1qkCjR9jj
+dHni97c1iTA5W0AsPKWXWsX/iVCkkzEuIdJqZQu3mwtPp+8wlFfS+KTsr46PzCQmsjzvkDLwzhv
duo6ZLsoS9kPsoc8+fGf+JBg2N1IF/Yt34utsv0NXeqG5RXLZ6KHUVc4Jtw3u449yqPCUnw2s5dL
gAYy3IlMhgRfXNfetvbGTgB6PTV1h06lHFHHbLerJAQV8aJTD/Mk/McxRnVT4DFDQo2AJ9SlsFTJ
GN4raNrUXSpctd21Jtox/YAbSlk+y5GnH3zCqn5dxCTUoYJncgkrpJzmNdgbllxvben/cxtOr6aE
36r/S5yzjbzlVhm2vFu9RfX6mmrXh2jYDpUnKMwXHFPwInY86ybXnSiJ40gvq6IukhDM1HXR6RkF
bvwrMHNKhgdxbJ+f0D2GeICvh6nO8FZWvepbQB8EFgLSYoDfj/Wch01G6nVVjvXXdJfXzHaE4ymd
JFcEOrU+wK4kxyFGAXPCRepQig3UgTtfwnBgKtRIcWw53rm8Vi47R/RIorhTMoexzLfCrt7VSRPF
o+ORH2AUZgdLq0MaTII06+FG1N8DFU9p0J3sbtVbNUJVGV87lKklyzEK9We1LrhlKBeo99KQGqIm
gO7Fj+zwqOdjXUlaJ1jnP6NMcelO3rzBnJcN6p9jbNj1he9Dnt/lNVkWnbUlseSZP7w+Cm+rYsWL
TwRMDquOJhgjqmoNL4Bk9qVLShJnORzmViPASNWpoZ6HB5W1SvqB2ueoqCUPP7pMIc5QqMz4pROQ
Ho+/Ve80n0Nqtbm4S6F6hzGNqXsF5Q1QwROVdme3ckb5R8eNE2anSiz8n2qLPZclSsOeCp43CXlm
BlEBGIUDD/6VP0X6ISIlQN7vZWCaW62RFOKMwtf0mgPywhgtMljokEO+yEKzG+cn+q/FO0sPCoFV
DaG129/hzlf8AdefbNqCpW8fE5mWw8e5fm6NF5E9VLEA5pnSTOAaB056k51gsvB4xtAptHU3JJjt
pA+MN6lgdIf2bTDRedZfNNoUFmbZQmf/JT0Lz0Sigwsi2tYhNhPOxhxPVcRQ/xXAizzBruPQEm4T
0M+AkCdioVLPS93AW1eX2AsEXJIxnqAedtC9W6VYDfbyZ+hNWnccZMpU3PbP19tQ3XnE+4Lgn7mx
TfsqfUYaFiCSqIJTa5kIqgtGBh16VQ4ACWlrKKUsu39KINreoTcIunn/o4rc9OIlcGjdUdFh+C9+
gVLQYPd3nXVjVhxnMORvZhtUNd3jomkqQ00JNiMaX4d7W5lbvnEh83HglIAnFOL0TMxupy5seZF1
EvIRijUV0Rh0HO5Z0E6us9N4uXaVtW4n12sVVj4Cv/+sRb0yVllK1kFcdxkYF3GcpVfmLsXxeIdC
5voxKVOM4WFpXyutGCvgA3Jy5UpCYpqBMIr8Z/GmGwIGg0o+CFiEaqywOcLZx0UmqAQ/JoJ3+B/r
+THtkZvQjCTX9uIZQAD7TitG60omr01uCq2GJfT3jFE4+/M3F+d1mg4OCj0u660LzRFGK5zesVv3
P/PZVrP30r9prMZMppI+qW0YseFAa6UsAVTaKcVJSdYojkibBc97d1Hv6eFX00SJfzR+uqW0RU9w
1MP7FXp4Glvc6uLMPuIwX7Y6rOPeaTspbdtw2eKKQYypiqJtFfGt2UoM/Ly96L5j5uSdQrJwAhBA
ZAGmjsJgDhtMLf4OExtN0/G9GgXmrDIiezjg3jKyTifzd+iEaLejVONfjKpcxbrgeJuyMvxidrQj
HW7vnNTuNUrZrjShrkJ9yjXHdnaKz+0VBVCHG6mk+9tlrtb40ODSXhd6f9TbH8k7x5PmU/1iWr5k
n6fHa7mwRk0XL0oimeRRP5/eqYab4qXI9RY7eLxiLwPNpvCQX6J67W2/Lo5MFXeOHiJVAgSofzAN
O7zmLdAqEfTPMo8JMPcWiQ+tyUYtxu28bIFu/ull2PiCpAWwKikgFgOkjJEPEIfxY01p+uO/0AY6
eRidMMEuhubiMn2KCmViZ0GkyaYP4NQt86oJhb4KnOBbhNXWI/QfIcCAY3BEulbhsoaF3dIwZf9D
KWuq2hPOfk3Q3P2ralGq5pnqf21cX3qMEQ9feTkM7yV/a7oe+T0imrypofdS2WA0BRGiGAxlE4Rr
56Fs3hA/U2PY1VWxJqr4FzP+ns3O5EFgfpXKqeeLhHAfK24sGAsEPZBJuamygO7ALTCynt+3oPT6
yb5CoTEkAfmmtzrsKdjteAFQQNzzlvzdTxn5OAM+e4E83jRsq2TOuxghcCuvN1ymVTQIhTpjb9EV
7ntbYSAlGpVxZsKkaIEvE/rA09W1IO7dHcfwyMHmJ7j/dY71vZoVT9Ql4bg1pM86DXoiJm8jsB1Z
oa1uj1PHLj7y1lxLfZl/zDNRtvehVDoq8m6y3sKthmYommxISx4fuPvhDBHs2Mfscc23CGRwFJdv
gaBX6iaBuM3WfBUInpX9h0ucohsOsC6BAFsi1NJapf3TOiID6EmMs2QjxmtGOmhzYJSEagSmNKN9
AKxC6VuFrXihgErW0Sfk5hwsZCZYMxl0EqeNeboYvHG9L1I0mymbxIww6Jk7rBYYdr6msxHXvvxs
fSh6N6chgC6YwctgMcik5DmM4+kRhq0Gye09+w/8gT7nnBnyvqBZ8RZ2JpNcTjXQ8Sd8HGdQmqSx
Nf/tyF4JXpGWj5tV2VF2N2omzLc6qyVbPAtPyJpK44Ob5JJHWJlBilBUyTO+DxXVVdAuf3mZSdKX
ioLkzOan2UwcvtsBZd1NP1a5JGqnx4lUJyKH9UD+aIRmckFM9cIIjXi1ki3jmWiQD2jH4okLt+Vz
YmQlPSen/51rl/bgXXqOiqEioqO9aZknvjskoGg+L+qW6SlUdgf4I4x13+Nz+3aMwxff/SAIr3IN
Pvfwd7zq+ASWKKoa4haMAS7PPOImP1KPTbQDTkLd/cQQDyiy3fLyvAbZMuJIilh1gSKT/fH40Q9m
nGlNN33sGSbCGC9gUjWhG4VJ3wTQleErqmc+CaJ7dxy8SVWvMN/RuPTuRD6Hht47zOCs9DzG7Z+a
5LMWhomU8vZDEjUAZ9+UmQfVXYK8aE1q3FG13MWVdELQvMqEmTf5uYYRT9Xc0yUpTFaU8yXqJvQf
h3g9KMJvPPKk7WSmvofNEfdb8Xq22kLNED2WyxKnLhk9Yhx81Qz1jSW1frea2n9j/7bnG4Iz0EIN
/G77kKgcUxkfflMduU3Or/hGRkI3af31zbVon1F6IwdovrbyViStYlfcLkhtPpxaexnzsBEsIKC7
b1mpq1fUY7rLqaOmWY8K1o9aSAiw+kRifOPF0eTY3JOdecUB2WNUjSfP/LjLjcU/aQ8xdmuP+E2+
WV4K0TFD2wStsrLP0OFhYqTZLknM9bD+lmNgGO0oSGbWsvOiY98RNuhEcS4nIC6A3pUsWpmdxKVW
mSWr0g3xwhSQeo4XQz5q2NdMg+xEVln35bBAECSvGMZ96AN+FlZsP0plNWduAHRtFu6rTh4wSM9v
B7PoSpgniKBExpTCzJ84cfdkCcqIDPdtlWmM0FDNU3rHCsv+0v5KkWBGfotkUpTFhx/4ktpR0nRx
Minq6BB8HDjZPP3PZNOzq6ZsTiEgbjxoDys72DtQ8+MBkhvW+/z0RCVe4183hIwT0Zkm1mnsYFf8
XnR7S3/dQs28833qmFFexK2qXPNvMi8nF66VVWmz3stVtY3RMVJ6z93rnhx58KFCmGobUd/bgPCK
Gqy01O8UaKx19cJ3silB5a5nJZanE/Wq9jSCsW1iydl1qv8DiCUShFZkTN0/nwC3xNENgRMVhjRC
xu+elDWaph/2VvLr9z5fA5z0J2DO9wUBTXoET+Wv9S4CDkd9h7W1qL0Tuy6gXgPofouwgjgosvmk
rtUQ/blcsVyLpHbNn6+ZKQpaO4+ouqG+8bcWpqnzg2BMdHExsscwa9mebRybxVMUhGiEMaQ0B8LT
3Zdp/6q47E8ObiDFfGoYn4A6aP29NyLgMvIMXFwnip1gpGUMml6x7n1m1fO4DMbBjh32uG7v+JF9
QxkKTPNaqjt0bIshmUNqKRFZYgioD+HNeNlzBMRsL/UYCn3EcM8JAlOOXA7zHMaTqrMZ3iAT885G
br8MffC8xU1+IaShlQGCP74Wfnju8wEoRfynMo0QpPQ0srq1TFyrw5I2PMCyhfGeou97s73m6Qio
45+TbBNJo0dPqK7V+GE/evfx2D25iZuqtoyFdJfkcyLQRpaG5lj9vrtcJA94iBo4gGNhEJh1b2vN
3vMn2MweboD8JeqGda+ORxx7R1zhk3Sdkajp981Jg+cFSKOJ7+wZlWkd4TvZtQjI6gD5+1Dj2UHE
mMzF+aL4eUWyvbfuD7y2Tt/nzh41Knt/TRkJ2r8u3qEa6lwbIgE4KAr8ngtNreJBbTUYwQUrRhhE
DomR2cnsmFvjD0dWIfzMuq6yXWYMl0lKgNli7wb9fxb5tUIoRzcK/iRdNcG5Dyn9Nzl19JosqUUW
hQZigdPXKbzlCgEwXFsAMl2A1PquvY1iddAKAsAhj+75GhuztYCOgRN4+5SvizjuWcQir+e3QIhb
Z5cgm0fuWwi90UvXflLtX0ZxgjdQzO0HOGLuuISKXZ7wRok7/Z3hgCE3x+EQ5mXi91ZYAGi18oWr
Es9a2+/AmT4e2NgeaX51RjhL9CbJ4TF25FRzIQkEMgSjCn5oApKUF66V2DAbSJWVOs9dDmnSFrle
LqGFZGDAQu4UN7TLSmuQOrKwubt4KcvKsBGgu/nsPyXTTJju3u8UTzoz65eo2EO5+NYI/JUdvIrz
TgW2uuio1f3+dfSwUojjXY7qHVK1QKkHu8chvx4ukw407WmIQwzfEJgiazu/9hYBxZDj5I+AT/HS
UNZ/VZVkaUPqmVkcc8fsOkeQrVD34SQVE0RVXXSvFKzHLG4RkcRm3Y3Z8Qt2cCB3TdWBTK0qb+A8
lD7v3bP/C1AorYYmNMQlpbuqBopSZFaARIDWO+b0MSvuFvDfj96TxCjXbY1Ta0EGTJVhipr5XL2o
N6tZvSj9G4/sG92WjoljqqBqqalnBx4ROFCZ4Bg+veefdRxVNB17GlLDN5Id7+zffHslI/CkI6gy
KcVgz2yGeRB9fb5C+bctJkTfyvL4tS4xPkeHrTIek6XIEfc/NTGM8xs/FM/2XZpiJkC3cxIzs1YZ
/QNTPn2HDYsk7DIXXd3SWVSXW1dw33CENtPP/H8D57cBjLUR9FZEQjo/5vwECkkG2Bufma7HLNeJ
2F4v9U4gW76u/+aK4gQmSewNm5fRp4jxZlnoeygpknBEtpGN2HIkE5vbkoJTOiyPUg8SIn4zT0qJ
5LboTIRbo62m9sjj0sE/LaVJ1xp6FkH1nC9zDMISwn1xIb1DpLYCSuYMy0qijtrY66tdRqgFdbXs
PnDGgEP+2GYa4KIrWLCPt4tT3PPlN70X8DMSa3sMeiHJkvpWb/ccPm1k/vRAaHHG5QP4qQORzO2L
wMcgBZdesxvxlbVaXqKsqYDZDNXa1yYmA9F4uZe7KzdNClRyuMRUeWu6uN83wQRNXtBjrUwbwJlD
mfDh/I0UuI4xfdUoE9NzT8mejPwP0ZZAdjFsxxRG5Srv4zI5KLa/v27NeAI4kJdhWOOT+eCi97ew
1shdUx4+4yNt+4a9KW9Zr2OEh77RUFkMZwsBadQ5GGFNuge+d3UCe2rSwICVRvbCYX8euUO8XOWI
Wlo9KKU008aqb/raebQwoRdclDe1B4yVEowx6pL58LiZO2IVszuZeQzhIWbsMWQ7ATBi/cdYEXDJ
2SjKFhQ7IhL9Zyp/knOSXCrJVaDvelhXwfX75V8FlMBVEOTXXsCA3xx2fYkPsu7E8oa8+Tc+lsvm
6STDiz7bRPg7Frfs8TnEJISaK0x2kRBvY1maT8HGbp1uHqQnNc7Crp+m88S33mS5LGR+l4kfPCBv
sEJH2b1kyCezAyWiRYQ+yluQ3Alku6jUOdGb3pPbtKzqceS4CKHcE2zLzsJxFXuv38hYHi+lQg/g
WqCXtfx58WxexiAcmLhd/9GWY2S09qoa9T5VxZmx0fBUsTi32JdvdmQeQZjqKOLUFMJd6IMoI9Vn
m0OAVo5KuEHYoWiNZb9UquIVT8MNTm9XR/v9wJXfmVM+E0PIMixQEuLgpfvycVAVfeuurNqRleUV
bYJgK3AftHRrnuYnlke6IEoBvZVrtfMZEVu5LWy1ppBuN6aYpGBOMjg4kdBRsyRJktSKvkX/3fTR
8ZS+GFR5mZNt7ctVbAxLoih57uPzhGpOYfe4Z25kByQBSxarPMcpY58/Wki9dQFQNDy8PXA3f8DK
GllPkvhR26O3Lykz3EF0ZO97wsdLbyKeRxXDDWww49ZfWLbUZxdhIkAWDr6IWyQVADuyoE2rRvVx
2mpT0trzn6jtu/KYzUOKeSqS7WIlzIU5Xr5s0Qw6Y9p3+/1is1B5LCCq4nbBskGvj56JcQi27AbE
sDShewNmKwX6tIR3/PFxprQ5CxyGHwpteUyv9GxAV474UjCaDYiJjUFL26gTWvmNEfhNXqfaSzRf
6yMbgmTAD6QCz1qhqpR+36m0WXUO+mTwy8uEHERaPADIcGRxZ+gVyr8xDo/M9FywUnxcfWA+X6KA
HklFD58CMQYcDofuw2mQVJHpOWAfS8nF7bF+vNkxddGfhyQ6vJwa6xT6D6OEtc7ZFEuQ0BxUCwcp
kKDybnoDhTf0mDfuiau+kwi52myxuHFDgZPLrt/7RBKMfrTqsfBXNtT8vfIcWgUJJ990lic3hqYY
XaCh+unFc0+qtStuDfAGw0xJvqPp0WnDkF9uL3TFAmKdDv8OGCxjcYQYhZZmEgy3HIAESlo6PzRq
ksLF/fljzmHe9xc8/V9haVMMh9oSqsoLAJVCHm2ldokSlcHmWJf/eqSoTqiEZgVNELnG6lF3gYkQ
GTBFSWBuzjs0T+nT/QccEnJXcISLeYTOg6gj9q5b+rh2tIxZSynyF6iywPbwlC9pz22Q1vUuMQGI
w7vDh5uvwsVm0khQQttId//Qhel89TX0F1HGRAUm7DxWz+qowgfO/DkEFH/A2qm4ayZ9DlqWM5A4
Dkw/zS21Z9CRjeTcH50Cb9vxkbTW1tlv2ylJd6W2UaKT5uK52d4YxgvxqJjFEyS6DzeMlVsN796w
ZP2f9i5H0/LKSFWKiqhtSFHlnHxI4vIWulBvx1q8Vdws4VVUMpBcuBEdVlizj8HdxKe53ml6BLZQ
FY58N9UuuaLsxn0EyL7OQINHSOdTrDJ159G/i6tJSooSeHHCiAg4NOkyF5NPraiF/uOJJGG2ubTj
yoSFXlhOB/cff8k7C2j04SM7uVOrMi8YVthShIFJl+wmT4gDqTd2zKLyx/crkQ68430K22aT36Vi
Ln5TOcdwsBbJOk6tAsaoIvMOwvnn6WDNiaec23qwPJeBcPuKzg7+Up8GnTvR7DP/hTL4ArjFdw+o
AVK8qes50p8xPgRV0hPnwBNZzyjfptwCVMbH7WfKc+kcEqcyRJVeUDJrnQke7gXsdFItWlPFcCOS
Ye0fQmCJUlc9/c4exO2s6XVCFJv3ONIecwp4qgJJ8eKN2Oe/h63X+XHeANsLp8FjSfFjLLiaM4Kk
02NORGTsxAbe6XXI/k8hu1XyrGEJdZ8oruy7lGVEH1DC2/Js2eAvOw9SNr8wmwqSCPdR6fk1Q58c
zeZ6pm69SFZyoH207LehwxMUhCkVfvXZoUu1lP96RB0kxjuiH0Hg8ZNX4Fz6LkaG/WFj7ljqcejC
o2ywo+U931mu8avg1HAQTXQcZf+wov90OsoM75bmI7Se9Z6gb5dkQ58OOlWFsg3pisWqU/D5VTn0
WUleZMX+PQC0TH4Ij2WkYgGPFFW9n3fov/6dqEejrmiTT8bDxqZqZcNllIIsJEiS5I9ztJKmF2vL
5EoB9nIHUJFyNKZItG4wGFIylyI7O6nUIyFiyNfvOcY5JIYAUPcXA+R91HfSHRZM5P0rHHojVo34
mjxK4Bl5mBbmIY/XKtGfjkii0PnGd00m+t0nSCNo0huclYe7JkkyIgIco5lJaZSpsh7F73flgGos
Bs4Vti7dv1FsS8v38P2ICnmIpzJqhCgUhguXq3m6GAVGMJJYShk/WGDInLlgvtxGZjheYgqnmTUL
dACPIpMTTjzOcjdDeYyL86JbT4wyKUm/rLiaptSdJL1gLIcl2J9I9/lALQP/AovnrLilA8aVKQLx
zdJGcc9QvcgMAOim0RypdZjUDSxL/MoieZrFps4exGhIYQpP9cjvMd5OlmY6BTelZKmABfPTwWly
qjKxmGDp5YxSyJ4x8h3j0cQQSdKFyOYGYgUEeIDKIxJHbFjuxrWYbM37NQTVq9n216MoebXwS8Vt
XeunHMOmnZ9tiQCb+ujkBE1StUD+vXx5FWfhqL7hMf/CQeW8a7hKOqUdRfVP58gx8dlw8w7O2Gle
ckdW7bigAQy6wn2pl5XIWURlyFWM4v9akZkG24BbNzRg2josQ5OrGjR10egJIW9wOrU+wJL4RhlT
ODOeeLCsKwASTeD7BribEr9ewqU0vZWLzTm2Nw6QNgHHFvbb4nC7NKxhB54e62vGEcrLGDSn/+Nq
Vgrij7Ht5cYY5YY+29SlGPuNijF++WdnHXDte+m3ViM6tGowJJ86l5EhZ53+VfLwju/gpSApQxna
P0E9Axn60unkpRKrm327n+BrbUj6/SVDnhpQpr6p+0XV6/LyQg0Vbs+Fl7A9wONxzDKeVjJaYe+u
pbZdRkCjy68OKkQxQF86EmMf8Pi0KvtLEUV5rWjy7U53MnVIkN67hcXiF/ceAXtWhdew+fk9C4dF
uMYTu4wbsBm7Xzf/BTscjw4kxMiRbvkMxFkVzYMUkOGboOW9U0OoTD/ZoqUOzKExsqL9yRBGsdrX
BY8HffTPK5fWIdKq3HJiVYic7QD8Z4V3nxzYhepfiK4XEMeEld3FtUGJy/sb5a2FbHXV3ClDhZVd
Bov3337EfeiGdkyQyMG2leNRc66eTkiURXXHHASuB9PDEpptoPoTZomtXXlmC6qYy4VSL6Romwu2
kwA2nZGuzoIUgeK5Nq1d38b5HoOdeM9FmZeEju+4XcMs0axzF3GfeFUx8zRNplAOhS6fZI2nEhFh
C7ShTwqTPDtJiR5trQFqAzFiu50yBWhq0ahnA1SMZRGAEv33WD7kyulpGmQd9H96BWEzUyFXvZfT
AkTpgNT1QNK6TlGE+Rtoq9JSSlenW/7/o0L7bmJzFKl4OMLuJv/uz/lteNHxw/j96NQL/iKjSQEW
+0zSiDZoR23jExpwq749P93EyMLDsEjLbxZM/4vSWo291WZ54OdMWIeWh/q1Y9ym5R8ZXi23sNyT
DOfL1Rw/6kQB1WOdQu3yRD48xcTuTRT9tLLl2C7SaIYkq+/d7vUTLWrP2ZhQuQIVlQUQXQr4Kh8X
O74PRCTFijoIDpQhbxLI9hbovIz8ur7QvjoKqhai9t4y8L2xJnRC+AuElWSC7iAgnw5PAGvqqY/H
2KpY1T5iOKjtSAtqPHZQ3qyJRStb8sCeNDGLEKteKca9JWgLQniH9kn7fDaJKafyDqVJhhggITdA
kVhIU01g2XRIa3TlO81uRqn7PoKW6nSoZekpQxypHE+xEVs6p3ham740RMFXOeqk73BybuIOL0nF
bNTswFdMejdbxYN0w5WMp2/hL8KGgHagkneMIJo27PDprT8IydVPR7LQRP93EM2QJY8W5WG+T5N3
+zJ8GN2vaLo6vIeJda7YTw3xz+hYbMaT88pGR0S7oBHdtWDZ2wQuGSgUNPlWgnXtO1f46A9JVRk2
tvsqdThsvZygKu/mHQ+iSAcdbPRQLF86ZQEBFD9+dRrpccwLhPnSYtYZQKPIYkRLRuJ9UMLIoTJf
Wu4hF+EWumc5v8icYu6fzftjeMqQiXVtzFn7ek5FsCGyAwGb2+36jf4WuL+aKkaHjRygcg1QlXOg
rx1Qwsa5hhG61CJwmCfal+VqZz32/UMqc6zYJFqqGdB5aNhXkZDAjLn5RUn46s5iP9xkT6z4rh+1
8g5N1FCbO6wo1e+vaRPriD4rX0W21HaEo9jK5Q+BfGLwV7Q1ijxKGncn6LWPHChCHgWkxkFDZw+4
fcP25L8aSh++uGIHao8htw+c6wRJS6YcZEdn3Gmy85vRnCpxAt7PhhWwKSG0ASIU60upGY058zC+
EPXsiqGWEKBinE0YTJgxyB0Bg2fQYf53jr0SyC1EQShyuR08NIuyc1et53uRodIOZ1t3YwMaUa3p
eaWxg0D6gnCsGlPsg4hkAINpFA1/OyCx+17LluTXJLLhWDWhFiwCr0z7UfFQClc53NkRlDpFdYnx
ZG/CZrLHdxdWH6FPbxiFccApsQGt2J+sfJRE13/Wq3ctNTDaO8mmV4ZesSYdiIJ0p18/hwhI47AA
uKcYtQuER1Z9+tOTSV7ZMNXun6Djxit7QF7zKnu1NUsUDxNw2daOP++PYiwEmEowesExBru0l5sU
NJ7/5dKpeqMze9bKxutrdQepE7+sFbxIkDy55MypGFp25oqoNVGiA2pF3tBIrtsT0cXVPSSVKZGh
kOXluX9SiJWO+IHaA9ECPxbHofoVW8JrcNPzosWsB42wFPbppvWxhcAD76vEZGGF5hbokWtmLbjT
QvYBGxj74b4eKySicx4rIYL9CKLZglwSzVgqZNjc2pCnzsmwrXaMS3n7Jm3kwxTzrizTCz6NmsS0
9cC7LcntER/FkmDXDAZ/2A6stF71RgNrrc1NcpEBPyqGtU9zcKbvRlhZMEIjm+MHas9zKU9A1TmJ
gagwEhTbQ0uPCAqzzsdYSPvC+4BoxDMU8ytOgkaA2WtX6QB1YD5nc2VilAnzsQZYJ44xHmNFkQZO
2onj+imDLF1+iS6E2sOSM7aqriVEN2TcjTCfu1xQGXyrm3DafgVL7ZL14RWZWdA2im+lsgTr4RAP
KE7So49StQOtSHlxNynvauewxWO7PCDirIG2jS6z61IkkIfPmUuNzAQqj+e/96CnhIquJ9gc/tq0
Zo8rT56At43H5ivqRHnkUj0dApLrnsq5vp2p0GgDLeaUY1lrwpLRq5oUEb4oLXwbbK45J5fPpPbw
72Ak+hsfZ2Jy5UIBxSYEDOBxNxEe69E7z/G/cP931jNWuhGvL5sw2bgHhfInqJIi0nmwVeCEXIko
WjrVS9TGI+UOa8cIiFvmX4rDc/7vZiMuoqdgZYzMHoJBIZ+XnXVtn08YA2G/nvcyszhqLvJB3Ogz
zLcyy0B1DsUTFIM3zangMscN8rxb97BAlX9HjLEI8c58MorgmnR4Vfku//KJdbpFT8+8wociMTCI
z2CVJ140v8Obf39UDBp2x3qpcRjSE2maIj7T1RvI3U2FfionQ+ehM2kZUnF/q74KWfGqiYnbqTVd
3uuOAVhrP0StLpzeFNzm0O3lBo26uS6GHaCYrzbEwLdqL7JBjol+Dc7JAk3XQw22nRydvMuaJj5z
eUD2sm+m8sJ2mP/icf+H5LEApf/S98t7C7pVNk3lX7bScTmQvKGqp1Ekeo4SV29IpF6nAS/6HRSs
SHwmy8rZ5uv2Oauk5Xy91yHC+KqCRaScXpegGkfoHOD5GkJKqzggSPE79Qp0oLCQ7rdNWpmNN599
jhKA8LTTQg4gSoImtgJlJRIjmA+ysHU/NAv9j7Ewwx7FfR5xpVS/Zl4Jk+EvVajwOEOBZZPYtRvq
SB9KQ+WlXFEJQRqhSlG/iUFLoCKC53F4WtCAaCE7EbA5W8OOc9QVb8bEomL/xNJagtaGuGqPRz/a
+bIBk+Fu0i+/cGy65OhViN1aWQkw+khMqzWniK2f+d5y2a79AK+8AvBIDCG62rYMfYI6vUQ2bcSx
MwUirNlAHmIIJvlZhWpZCpCTT9g3xY0IaGsEosQMt8Od84F1R51SpXWaKuiLnB2jBBlBLK8U0QVe
7R5L1BOIDdY9p7YHR8PhpmWSgJhx0roPLY+iBHJJiXAnMzu8utTEnPKY4OQUtAw+qF/YwXMhGW4Q
tHV4+Ym/6f6teOWFpseXEaMEW2Lcs+EmnIeF+Feihbcr9yu/bSXbkr6Oox59dHbBlILtUP49JhTn
N5DKfvHFVMZIpw3Y6ymHko7gf/ReUOrK6zL7zEuvxlKlRVUr+TUlXarAasTWuOA8mPLVfxaiweKD
VdPMR80qHqiyVNuh+Yt7Zq42SUNE7EqAEcuUYNnZ/RclB2rEM89VvxZXCX9HTdaDB20RB3VClWEt
zOviYRZFBh1egVWdK5aS5+CYCxkBJCnmy8TgNTmix6Yx770jDgzNN0i9rNtjRHzku1Gx6xWZ5rKj
Qk/6YmSStNk0fVTGVtwmjIkzhWeCjzmdsuD8bfpzB2HkDG/byjW2nR0curIjyw5gP8LU6zkotKX4
dktcyN9OqfCd1Q3HjBYN0tOlR22WxVkzy/MswDTsxK3gMohg2YbNyjC60missN+oXMbz9ZQs8P77
LzEfnvgzn18xXwOBamT1yeeRXr/AiGdpSygk5kTswSYN6q/Y7eeG47ZAGkZ7pDO+6XjbuMDYBCRD
OHrr4BzmA/CzEy7JPiElKL5LJrOxGg8WlKxiwy00lJWt4VEgbugp1fRrw7tEflarbFx+T6MDxgYp
fK4CnBvp8bkxfkRLC+j2F3xZly4hoB+ollnlt/ota3NLPpJ+JfQv4Lie1PkrR84E9ZQPLB1t8x2f
BmNNrnEwRSJv/0PmfAgVbMuNwbibjLe9pIKlbN4gD6FR9TkFzIpOCT6P4+IAwjJ8wwXex3quLCmn
GXsfaHYvScKvTuj1J4SuJyQZjJd8QZhHgcn/fvBZAVz3f/CdDExBU0CNIftHzHk9A/036OiQfZEg
QHrO6NG959jvIP+mBN1MAii0aEH/LvEhTuG9LQ6bcevBIhDvYl5LhZMivn7djk73HP8USwHK2CqE
qwxI4Xx1guCHf69+HDaYBWDyWTve3u3jYfVrQ2EJLm8X7mU9ikIjH4A1M3oQILWJWzrRK3rl2VT8
hTai0QsxtkbSTG1TxQf4wtjWsFgjmstD24Suqo/y5lqhiOTV570XgrIVz3hSqcALwM5BH5kjivrx
lwq2K2Yqvzf0eoIJ8YAuywv8upyclZBbU2oPx2jXPzF2RET/mHcRqxq1AX3SnmNcLbSIasb911WW
ew1xu4lVkkFQWAHl1O6RAgAVVwrfPDt0KQdF8gnD2XzWqlAloXcgUh2M2RlQFtaFneeQARJJrg/Y
xChWq5aSJVKUdTwY554aHES6cptnqM88rRGS0Tiu3zitlj0RRWdakMHDAn+pDwAjxbPEo90sTMqo
NzAOA+B8yr+XJNo+C49yKBg1E7GttdjK7q3RoiuHhf+TvzJoBJculjS5MYn7FESlgv+M9pAcYe5l
5Urq8+elg2x6aEM1drG95GY7kKe3dBqqjF1q7Zna+9dgBVQjG4hNYLlecddjA7OVohiTTVY8SvYF
oxlwBj72+ypppEQ0ouVCiNo6V4D/IPh7ulFW1pZk5NxZMNRU10Nxhyr0udYMCmsCE0Wrks5AqmDg
mqtbmHlhTFLCc4F2xJ4yMm2CLmzFOBZv/2Y0vMcIe3CncZDxRd3LQyMcz+4YGODafcyfT+oBr0ZA
fJrS7lhG+ib1F9ELY8SlNlcDAI++K31kmRJPYBD50I1kTaNLeCIi774XJYe22hUVHtwt656hb14K
xErEI3JXtRM+s5U6t+ZoJ5e0t4wmcJXz63+V6HAVLw/PGNCcD8NUQKGs82ZuNTRoV6MzKPg6Qzab
69uliKZeWZ84Tez/ECP3MROvKZvkWgWksOSa8RFZIK/7EWyZSryAr4txXncmPjqepXvTrVChJlcc
RsMrc/HELoHodnXv8hCeo0UvcaR3AMZRr/tWdl/X39i5HefijSDMM8S48f+IFB5g5JW3qdXpUB+S
h0QNQLbUACExHgZL7zAFlC+KnxVWk7QEIZMMRqRuiiqvrYbu/nOwbccXkNFh620w5fzV1pTjLo+n
4OT5LVdd7OWsLcnQ/MkawBsAxnfMUv4FfS1Il95mFpl1YcEwlx6myutkQcy1P0ZMvfzPmBkNd/KZ
C5fmBzBvWINdXWekPxHIYcUpJvPxm4eqmOth43gV7flW55LztqC7pMjt0kvXwjBq5Pk+5JO4O/Iz
J20EWslKSul/j8BiZ1bL1mTkxKAJB4KflIbap4YGbRbiWG8PQF/r68+lHEQPPD2hKkMPGxwF26rT
jyWOAwnHuCk6+fzy8vLz5lxIgBF/l2OfbEuj1zV7VI2+JfCY6ebFnz+p12G6LRX5lsfPH7+D+qfL
AUItZ6+QVR8UqLgSS2jSJsDw85gz5I8jmj3Jv/RykFUmjHmr3TyuMmVuRmksIQbd7v3KmCTTc2l1
062U3XRchKz/tdt0XJMeSzwQbhIr9+HjVqZyWwKQR4w8xJPEH9KKLojor8WCVrNPwmBpzJ2+ayxN
mjKet+VvDdCGxJ6uAOSFkqJEJD5kH1jRKMU8g4jbfODMj/0UJccuW1k2kujzMgVMg/mmIE60NYJm
KO9v6kwUvor6bc+ANCMYwrmRLMlenT7mOPQiszmDKY0mzVugUeN5lSv08wnOS/0JkS1R+uLOfN3o
GOl/MfS3ArkGqmB0iYW9ShzvHB7jxHMJKPx9uxUKRO81cZXqcBjsTfD+lm1UD9qs/0KPu3tbCIUO
tcM1hpRG+sYUdNWSkOxl0xIYNL+9JUBT1O03Lq0XrZfVI5cUbMZ91ZD04vHq9FvR9LmKSGL77UTo
zaP97wLf4n4u/zz8/D9JQy2j3j8qNXvzaLI8h9q5Ow8c3lOx8/qjGIZEr87LdTzH1Fq4HQ5QNElP
CnDDyPA+gasMCs0CTxeUcISkl/V/uw9UF+i8uSVdP4t12BWsjs0BYG7K7nywgxrmIdBaA1OlwraY
QQKpBLcmQJYPkJXe2CVtLWbRKOlYO6Xq01x73qNQ0SxonDk6X1oMxsnvr3DZ8nX8eIcNREzE16vl
tX47v60P6pIbow9dpy3H+lHGSf5T2EsGgmUdKERyV816C3KzALSKPBQa0tGWplNpgwCRjhV23IOF
jGiaxNjxU5tPzdbdpiOQeM/NE2RQsGpMwBKGGYXjkHmoJyR9lbc8SDymbGG+fMNwFJF30DYFiIMb
dxL5QtCmxxHvT3lhH17HAAP4dtSsprDqurDwSGpBAEsJ/yd5R4X7r221cpCGyMRv20CYzeKDEbpE
ve+tw8sImNFbUklYD4vxEnXnb6k988Jt+DRVIgCUFOVUxNy+eY7IeQqk3jUjiUp9BC4PbmAR14Xd
inBXYxPRhtOdC+3jf9JgQbKdJSuGRE7wzwuclihz1zHA6fK3Tragtg6xzlMCs6QZ+PJzhwkzYIRQ
cfjUzhNCVYyZK5IHIczya8ATcwF/WKnYS1p0Yi8qImzJNQ2xprJPeJI8OjhzL6blowLFhOpB06wC
oK7s8sQog/cTlJBUSVM8R6n06ZQRl+Ai/TAgFonvPK2lIsvFgZ7OeTXrWt9fuhf9DOWsGu+yuprK
YRn1BoP62nlgitXx0ZoRyIIK4+xRp9gS1gUJ4nJngLBFUsAq7Rtl981xIZmt+lXpepZUuQC6lLvt
fPkWV/d7Lu6kV26OW3GARD74a6RcGYU5sNNH/exqfUheMxIaJPKhD2+kQX0Uw+9iakmK+meKFuS7
ItheMiEM0IZdakbHP7h/T7pauSVtBeor+p/eJCJFRVfP2rx1FJSSZUugLK6itEQYV+9Fgkg2Dxcr
6SqHdIu/MfuPlvA5D7wLb9TujJSWXTDyr1qAmqdGewbWAM8R7i0X9avWy5L4MCNGUAJOX1KlbMXR
FidOwKyph1wGUK8+87VhC9U5cBeQA4wd6owcHaOEVv+d73Uk9m66VBQ8Ci/kPZDxVF3Rkm12rY2d
LS5Y9WwkNWsuIrbQ7UHB8UU7QiFOVm7vAIJKMpYzVw8Hs+OM0t9SdNkIxeXX0A/QLzyOoGBV9J4p
ZCPIhKMDYbPtQXspKTMPTUWRPmcl2GC4aeAhxRB3pcLRDbtO8xIINKNm/a0XXB6jFCgFbhIf2Eum
jNqEqRXHBScI9o2TSi8bf743TjsZTnclWA0p/zd71zGUPg8PYjEt9Uv/o2uSqDCn7B2oSxYoNAUA
++L52qrsnAmEFSo+5tCW+Zi2HcIFH8P+TEBMQNVMjB8OuPNgmgbmnJ+JEl95iSNLBEISImpXcv7c
vptttTjZOXNQUAf8YATk+xMACAq43vkCCjwqvKnpKm/v+vlvrUYWExtlHkcw/qb7TQDfsTCYHa1W
0CX4/0SieT1dzHWF8DNYIsU0WSSKyQnmCwDcMk/g+qlq2NNBLIG8DGynQp9JP1sMfbcTfJ5oQg5P
/B2iU7MhfKgzY2RBfwJF895BE9zF6t0HtRENCcrukxUKMcq5CR0QlMvIPZ2dNwTwpkwF7BdsjA8E
LtGtWhAvEZqG5NKaMpdvdGm0kJyIlK7v2GfhpEGGCNNcwnF8WrN0kOKxm9Th3GKf9Ou+ktpbmUdJ
GH/GIEvsEfZES5GVS2rkRASH9LYtuJSTrF6oF36G8lzn352wm3uwhuXDHQVqfNX8tpm7rRn2nsdC
BXvzt5InYNFy/kLN58ZeS/9YjU+nBvZVl4/vDoi6SQGbTTAu7vJXMZXd9z3pAfLPgr6Tth+KUKgV
KBBWp/y7L060vn/u0LJvd+bAtzyhSXXv0QitjAMthtrVmpAktttpeuAS9TdeCZm/giCfxpKxf5YG
mvR2/7Q+fiekhVaevHfXjyWp+tnf2aqg9r8F8F7Bb2lcuSroHF3w/wKBccXeNk+ZBnZ/1rujLgGj
E1BDw+Ews+83Bi89JyenxrvL3deNgdpto6ZzICnldStFyy6OF1LBkdR1IV3DxaHY83pJ8uTasQ6N
DnehXMH14QmAuT7qM/nlvDIcZuKTXAdfTNRUE3fhyP7WDBTvHC7p7MAtoDr/nuBxBqb5vQuob0oJ
1JMWBAQzvqe7Kd1H2NazlgD/p24XdWsTVJP+Tg5HTrgX7IgNGJ9xRCBBHWrWOvPRZjw+fPfvdh2I
rDscM7BOg52k6zieKly9XCFIcn5gYjbZRUXwfUFfAYsCDOUzJXY8tSlFJw/eo3GAe8qxNgk9c9OW
RtF4EUAMj1cEEk9bExcZjxGiywbQukY0v3EQcTWVnL6tbXo291EW1iEnhGEBW08mpKe60kgxyoyX
7lf4GEoZV/l1nJeWW5D67TBH48YmGIEdIjVzBJR1KapOZqIRiOw+N9p5mcaSVBni0mRjgzIfQ4Wc
fKtT7l+jNv+6OrcRP4KHKekPKdn+0W6mgyrjkQFf3GcL3TQCr2D/nFuYL6kU0KHINQZscGyqBLlk
AaMVdizvqcGAy5AwxFA8E8TDheUfp2Wvs7yYkDapob4KxK7g5MB5cLnvSrm+USCDSDSeaVobOrnl
3A7XTzKKSyuCBPf7ZqiamN748UYAEoncg1wzr52G1xW+PA8lQ9FUUd+GZqB286KOLBIx/GeqOLUl
aRuSxXhnz0hDa+iZ3kqjmLj+o/EJ9M8tCQJ2qOaWAlyRROkqo/BVvYiYYUMRPkaznIsABBZBIYVY
1PzdPO4TkYIKH8IvQxZeX4ISWKuiXplT/xK529poKNEFxVnGB+cp3I099efswpVE1P0VYeS2NFB4
vr1V6a2DWvuPOnSqVt43TafurU0lWLERhQESYaB2RT162Q2w+AO1NTPPc9cIk+OwM+OM52V9vOjq
cGNUVsA0BiNkKIPMDttwXknoUHzc0hGiJbLgzdUBZ2flLjSDjCoPC78lKlleUIuxFOWCT/Kb8CFi
020mTcHbuVb6kSn3umSTSQg5VFfdPCtgsUn7tG6il4hDCgmcbjO0YppgmAHP1vY4a/NsSEobGF79
ZtdtkEgR+hFK7AulPlm+KMjmr7ZnjmR+RDaAaGTivkWKGMw9bz6RvnH3E+Xup6UPn5vi2S01dDtf
IIM0tstebiu/S/UnJD1aHDD7O1b443Z0X4/RjF1XbtDenx7yKLWElT9B7zA0w2ccXbuJlX+llJEh
WqfbfouaAMoMm3/fjmlS5Fq1ivm4Lv0C+v/qGQW6HWH8228D4U0VOF0oFEXGteY5TRyDLME6SSw+
Nv8uVXQVW8/wkqhujc0IKMdhRcjZ0DeC3kmYugV5zwW5AmKfwbySuTiCEy+1hyZVos81VEyfvJmP
hkd6LFF/jMM3c+qzH9csxpFzkl3mZmIsoAUbuvHHK0Ggb2rGcoAI9aVyRqT21kPXwJy2nf7bV4V9
5yuSFXqbm2rZ70OA2BebYRhjd1wBN45pIDM1PA6QbwjzDYSDk4zObqzPGyGb5djWzMqI4hZNWOgC
810ary4aNzAm1gLtttw6mueDIbdvUEsuTB8uP07kYDOCQ+IpuGWiYiuu/vcCheVIEAcgpWGhxPPR
AsRD+r/RFRUBUxIhgqzxDEgidADZfE4i5AoGy6xUZtWxBSek7GPHqgKNLiUSKFAzBqU3EMSny04K
FYpOsQXy0PZ3NjC2S4WstrhHcg32FzGkbtKU/T7HBVZmiGcjpMtbDkj60MSVePo7lLNzweAhRRSg
b7RRP/fq3KBnPk9/UqD1wKkm6vTX4k6CgP+WkwQfys0vmKrS0pk/K5poqxpm6HK8yNV9+UTo9PBu
rHReKL+CKsS94ryRuq8HovkRH0yuYSyBQwzFenc+OTMqpFJqiYrAbwbySNbFhgI9CyRZZvR3kOAT
1xi1VTC6j6ILzAtB3Exv0zWAj74jCrfHawfs9fLW88WxspR7RHRMXVAG15SgUFC8jw3oOmJl3+29
abQhQuY0KXt/JqRyjzDwGfkxNuFcMdKu4daDhqbSwdC3Zea0EP9cfk/TZ6nkUSF//LbIH4nql0vR
bRKIvrcb643itrmxGVytzdyrd1PXDyfmFKzwdL3EBzH6ZmjiyorJ1i+feuEbe2vXGSvJ2OD3574e
Jh1RTREAByjSR+BRbdyb+p6aBI0MDffU+ZORrku+IpTY9Nn1mDs2C0KfT6fIuL9/aNAQHIUdmkZh
XYpRcCM9BlBfDQw6Zu55oyUTcP/Mlp1LUIYl9gWWhIa+yXtoEj8cMYrkCO5hEXxVh8iv8+mYKA1r
LCO0HGuVH6lU2ChTRLinYRXP5pAci9ggFlUE4zv1aI01CDj35NNsNNXEjxnp7vRykoYzNAunAfqU
RMt3aAdf6pKRflNE16tj+vKWNSthV8ruBrs9gADGwv967alihBEG9K9O2cGRsYuIMkbN4cZfuwRA
iuCTHujqvUmZSvZRLW6MLCQE8Am24Cjv6zkWAumysc0QH40yBfMqe3Ilob2PFGSw457QMDEZVPNl
2IR3Mx+y2NKhdcMXfpJu6jPADe82ZWt2j01bGhhIvvwqWzBd49BEJsQvKad9MVgZDNFEdyrkSxCx
4bIF+84tjnjeT4I+HChATYTNC0Bv/8Knh8+B3QHDmfSu5Eyno5YcZSbwvKY7m3AzwzZDXC/wBmTE
I5SnOstnI8PhK80Jix4BQ8UhSVUhe3iQf5YLrPmSH1B4cEsyLK36e4Rl/C2ci6PRqGrKJiF6FQId
iiOfQ4j9B7lybcM5aZKGIg9k21a9V3qOAU8+pMzxqmmgQZDUicgsU6f9KXtZyGC0yZICIeWhrd8Z
Ai8uXFGtCEQKcRT2fJAHf6FACY8OYkk2Ct+BofEFQe41GrcPPpeAzR7U7SSbWdT5hSXPrqKgqL76
U9AwhwYbv9T/rUmb1811fmUloUUVqTGHAr3rqBQHjzjyCAru91VKGxEhqDyDMu8FUBCoNKTDRIuN
YmXi3scuSke7+tXN4Ek3Jis8VPM426ZuE1gQka4hN3sp15rUsmD41XZopxKLu0Hzc970whBHmorT
WGDOm1smbb/ew4iN/A+t2qYxBxo8iYMNNz+/yxQWCdRzspTtOaZ3hcPgpVPb7GZzCGaHGB57UH+P
4uS/fqo2E4ScXPYM3X3Jmz5fsBz473f6K3A/HJITprsun93rNEmpFn1HWnvlJO/P2stVS8alrK6G
6NdE7JVJpx520pRIwBeF2j5XAp/pdZqgfgbUlS+zBwf+mhddnCvtBnqDCvzF6eQjuWHSGbN3Ks1z
k4iEMp29PllNFqDb476uuS0gv19j+T3WwItaCePmIL/6CNdn2rHdKZgsNp0AdetWTRxek1+n37hK
KTPaxUYk1OYv3WXr1q9v9iPtHBgij5nMxrxcI+cIRtUrAwGwRC6PO7yMB5evCoCumUAv5O0/RLTU
VBbFBUIJGItIgdUXL36RPK989AePn2wVWMO4DfX/p8TWp3eTfo1h4GZZJgfVkrRSeLPRvXwI4oPU
7nl/av04vpjlvxpydo6227m4fCyecSRGrSgxN2X//l8/PuleGlTTNz7XgoHvrBgcHg2LeJ3QCFWK
cA0XReJZnn+W0rOt4Uy7b1dr2C6wOTNTpEaTOVALNkFsNx0yhKT6O/FAdO6mULHL6ArGJDEBdF9W
KU9BEVghsmCoJHjV2Plx0eoS7ZJKiy20LBRaNtdfM6k3zwdv2bhDHVKVwz45L7uitarEe3SDNUxo
ZeSfardEW623gUl9m+Cp7T7VT55R+15abF3fErTHVumYrmMPyJPXg8Ojllfp2iv5SnQ68OwY2mFK
IOh9uyFjRSLMb5PlrmuwCi2dr00CZQDJI/hBYW58S7owZUC7GcHqkJcQmKfqpqRt4PD3EvmPOYXF
2cNl/cUZQ48LE+vmGcFMgn4ogGPnuRmr5vRbRVVr7Fuh2Uxpkp8/yn/jr+0gX9ceCZWagu3ozAiW
byGrVzlB2Oc4D8Oor8eP/ldoAEvEOfZMJIzlFCdnN33ztZsT2MKOFICreX86Qdo8q3oP1bW13bU3
gcHo9DvADRZtqe62afBZDEfZarXuXCGTk4l39vhZe1oD7n/xM0gDrzMDe7sXwPiZeXYNgeK+qC/c
FJaBq1xNjjdtnJ73XJX6cmLGUB/42w3NAGVDqLsWwivAiWTA/UI6Ol1yvqkfAw/bLz5RKUo4mhB7
/BMxsw9H5sXF37tFJyn3Ox5HUtbAjzFBHuSjSqgTGRVus6imQKIF3i2jBOP4IByQhQfdifWOjZhl
r5vq9N64K74R9CaUBCCrpULm2XIOaNux0Eus6+U+5YuOkPjymVQH4WayXnqMnrnPqsxNVhdW54Wc
4Kl62nERfUG1U5MY3tnBiOjQCRIuf1sKh0wJ/U1C65t5o8FByGVX5R/45VT49g016yswEHiwqWIG
pMuR1/Fszuddp9XeSPgIsm2IaUClMif1w64aQE8l5XpHxeWaq1HsDKJiMoJb6SWOrUV2R8IGL8g+
ex+bGP/1uEbvaO9qbQ3l5Acb8IQQekFDXQjrPmfWdkDVp7NkoeGyU5tCqckeR50CLMemZA1ztWKe
LRdgfaG5fD9o9D4pdrBbR9/eNYnKRjABQzq7g5wdwux9+8HkSdaZHtUA3VajHnIFeCBGsA2Dy2Aq
0qNAreNz0E4Lg0dHGwuig+MX/DWimmFlt6l4mU/ZLzurM3jL67AL/eoCDxDolpCoSlVffGsZMTVg
ZyWed7KbO1EEmVdtwzmS9xIl2AZBjwtVdUC6nYDt4WdvIoKXalDD59vdmSkrgPVvMZO42TNChtMv
lKa0cZawrEKhUE98gOIxt1xBvaUzRGlDWChQPKmT1cSxC6TbcqKyTVEZyUqJMA3SUGR/lUmn8zll
JTusk8WCYQkcpCONWZJh7m8G9bSOvPhJQ0KOwTbTLXV5o+KoT4qryqSnJj2/ej7bWJTIl3Ylt/fG
bmRfLx/d3InDkQCNE5amfSL1m1MEmMK28j/WDpmDFSa69iFihWPER+0lurt0+G+GYpquFSXBYDV8
q295MBn34KebtuMx/850lQEl4CWmkTcN9g0Sf4Igh3DKS4saziNMTsF4F2tj9r54q9p7oz3fZeKu
7OJx47d/RJECvOt6FoEA+t10ykI5E9Jqa1deeV1VI0zEfCQ8GINZRQUWB3El6uSPsLWRnr6W0gfr
WGy42IA3SmsKUt4GADIaT8+dk8aTu4HTyC0kqE4R0vFyPhvonYKH5sLLXpbqN7WuyXtVB0KYyf7o
cXVnG4SS8G7XGzvlZZkhyR9P/R2H33C3s06LdiSBY8DRYn+InVX8zThT1r7K6HlJ+D9MSr3+bVax
ZTgpMcLP4XGOLyZBIpVsZW1INph3qcCJ3g1oQWfkVixg6egYJ7XwBFF5MRjRF9dBDnyjosRugrvW
kRS7EZ7+tjKL5iUlW3YGX1xCPWvS2C8nNbP2LmniWaG8knk2eLf3Kr4IDPyNBWZupybwgYgrcf3r
vhrtDvFn/7+AI27aDl/HIJg7gVb4r81rFKwsYitO7T83+lxnJdWd1IzmTwDegsXElVcKq7wfS9gK
8llsgPUazHgPvzEE2PcPPZOaJExrtsG6YLhdlRDB1RP0mXtOY3kRI4IlBi6J/aDjZz0PKP8f5UnV
VDBHHArKLlu3OtIozT8miM5Rk77K6qOq+EEfGkly4/yPtjFPtYlc83fonvWBhgj5E2m1aRwSerGM
ycr1kst4k4XNkFRfNVOjQT5ND0iYJlX7YDVN9x3qhprS+5QjIMArg0i592RE2tD6+VEgqUJhaiiP
oeWibwdbWCc1YNRq852U9VwdIou7Yg9u5rV1pxay9RA8cKBYEu27jMG06hbER1TjHc7FcUiId99r
Vfqp9xioLLuHaSXNlVeZcY2kLS3rYh//pT6wOchIqXWtOOHFcqxBFPjtrKPy1qxKkM/jaX1ZKN+G
rEaBPU5rx8mNOalY3Y+/bcH7LkDfemPm/0mWIrb1GBz8s4kNydYlkgAwt0/XPmEBvB7oiuLmm3ih
AhpH61YeZZ8XqpCfud19itSiBHegh77Dm1Yg6XIHjBtPdCmx+SRqjBpJ3aHEXkyBff3U0+ejxV53
lmB6N9Y9ZnbvdFWfnznSc1gCmZiXPBWC7Z64u37l7yntV9DWN7oGHXYw4D8ZB0vDp3aAgb75SmcC
AbKMJhd+qYVm+3a/qDM60CWcCfXafA0ewIN+XLg6PdrrwbwG6Bm/F3RkVcp0JlonUbBd0I/y95Oi
b8YaleVMg6u6fLwID7lJGTrftWowSt0FKP7Lekc8OBOoKHI4T93lmkqvBsu8JOA/99Dm/O+Vfs1d
QDyEYztcBn4JCPHO7pYqR/xs9Ie16ZUCgiWjnvL+9OUNhWgmJ/aKvcmX21+mCYYhZZ2XtXzsrj2e
Xev/Irzrw4BrVHqfvftFQzaPxn/SX8cQUyhko4nWNZ0baZlP7pIm8PHzBb5xlD0MdZkeoVqnJs2q
E/sC0ccjnM1yDeuwR1cG/TETFgYVO2N7NXupl9/VYLkv6dSZ7/ZXr/2wKqmj0epKE3V8KPRk74P/
kkByevE77yZScLo21nArwicqUPylUxbtFyX6jFpYlnPSKvlsN7tP0eutKJT0TrnqXvyKWgfsHmod
OpDm2zB/kbIaz+qCSI44EquSyJuduNv3ip+WvEmZo1LbpbC76ZlwpWO9eu+8WE/ACghi6ESK5inH
XK3H0lnX5r8CMS1BFnzwSvrzcR8hE3b17DfL2pDfeKR8PD3OFs52u6Y8Mu0yUz7yX0i5bUlb2Gmb
sTL4etFnwzjQlh0hXvB9elCBxzrKVOOuCMR23H2d5mSbUZrqrncljcEAACuLC0XopVeKGim85QUM
TThcsWjLyrU0n9+cl4+rALL1iejc7JN6h104p6RSEinunCMqtQ48VyGmjMy8BReupuGptmRLuVX6
+6CkDtqrj7qhPir6kIXt1TB8YD34xiLYQqQYOzIo+BAeGyFADUU8mifl+XC78FEQBfuizduRwhgd
lP9L6MyuJpkUZDW2sJkttv/rZf/Flq5ENe9Hi8r/5DE/pguFJ9n1MfEY5165NNOJmZjI6oY/KhJM
SWp9rOIK+DEFet937lnIiRKmmT3OBz67s35tmAk5AGv7G9QIc9XRozDo2/gldN/Ch/xH5mXm1Qxp
KMqFIuyV7xwFSl7/am0b1RGq4nF7g5MmXAS6NJK2up6zU4sNVwo/EMZiYB2XGpgik7vIj0R7vcsr
G6K1IiM7J864P1aJj+SfuDUgC13vMMHh2R6yCPA/m9DFkxoYthygexpnoSpvUjdmXxWmA3TQTbxr
aFcwTUQ7ONQIXyadIk+whYku2DZbTkHNJQ1rX4kTVBWRcmfwzUZLeF2SO5KpZyHZqyOQ20lA2ygs
L85gd+t756daL7Se9yPegll2UcX6CeeE8nG5r9Ezis/CgLeFWlKeT3ziT2GcUxkdosJfjZKJQAgy
ICIlA4M6ytG2OBcYH5g5Mwsp18MA2o7phekaOYfqJU9C33q7uub7nSpXzsdEz12FqXteiDvQeLsR
/RSDrpA5DRJkfyL5rZciJTNFEh5gnrFCI2UEkQpgTJDSXKTj7Cyeb8Uu/a4o9xNWUclDGo64NByy
dqHgR27E6fyImhFGeCWAxZimzsqRV8U0eiOoQkwTrimIyCTAgAjvi4jag0CbzdRsua7/ewC2FsKo
PdBfSdZvxFJ1xZO4CnegOgLEc4jabbDrwlMPq0cgwGGN1qpqeFA9piBVsRMHNoqeGZ6EqZV15e1e
+xKp053ZFAGxSdCfLcwRP6Dkwv7NF7NqIfYH0VAwM4ByIdzX9O+CfDvzMU3cdzDEDyOthlg9vkOZ
mPwbXhe7/j1VI0sdokqI/fceMw1kWe+9oqQHaedLops6wXsbhKpItlxCgd/BJMcjzENzU0M1XKD9
HO1nL5NA/0ywJjtXvverHZCenx+zfEGKB6xcl5QVnmEY40Bu6tcSCfGnZXW33NJBGoLbhngOMAcf
uyiB0sMtca8UuVYPODLm5ENSUo1el+mfJlhdSt8wzJxT1xbD9Bo00/Z5sOpSN6jsRguaneHSLUZu
+eHydLmRyKL1p8jmSpkP08Yd9sppzBbWEdOePpZbaD1AnLNi+zQK5Gh7g9KSN5Loq5i44j8xD1/j
xVJvE/HMfD0QBlNMBh261O96honB3vXQ57vAyicxtHQJ+9Gy0ntM006WWAfpFyEAGqsaQRHtRCgA
Tf0Y3IoBPW8xUyc5JAaTlew0Yga2L9bTVWkGtaJt8D3YR6YL8xFLiJoWEVPko8ZGvnADMoui9iQc
SaTEcI9Ya1wvhnw70ZZ1z597wDNFoWqg7sHRPiHANuO/15mVSCCXeVEpvABzbB7XTzY/ghAif0rL
sBC47VEePi6dPHJKlSKtsTT6lskhb1eWsVrS4CsV/CxKpcLjvqN0Rt21U3jDOK+gBXEWlYYndGJg
qeaqorYjpL/wAOiYxmq8DZIvEgZNMqK0RbZnMcWcHrc0UjMPZZ6hHWNIgtXanpjS4pCMt9YNCAEN
8F47BUz7D47zPAq8zZ7xDj+pHpxAlMcHsuC0f5vl4SgP+cSz3KPeL0PHgm+z9jFwRRe1SyRed3KV
BUk1YtxdRSGLgcatKW87R4v2kvEW7j7JaFv6amKV7J8oDr2EoWrhDr9FFzCEVsbn33oTkos7GuZF
//9JLLHEW7O+o1548ZbNPBJ2cWkGpnw0HxRgBhKer0y2AybOwLdAQD+CQh9ng6wFg3xV8Pa9uHDO
I5Kf6uPfOkX4vLPLLA20zypVSJooDtbgvAzSinFWWI3UxCTgVPmNbKyQ/Jtw9g7Ei0iC9ikuirhn
m46BgIBlv0FkOn7U5ROSaQEP+hSCyh41Rb7dqa2Hu4k78LLPr0bTAS6m5B3/aCnkhn5BCqbBr0Vm
AQpplhKjzev/izH3546Q7IGjL8VNxAQ19H4rVvUSOcjkLjfBsK9wwAXMbQFVNA4ZNtYJRlDrshLt
IBfEVNXrL+/8hVtMy4+XqiQAFd5yZ3oXWUiqOOUF67FjhLBo9il0fsr02/FcuuSYepEkjLcsNBJf
QVCKC7i0BacDRxhzUH232NOvEfe1oiCQvIxxMAaaoA8cBNvxLJ0tGm8SbdIcSJBMEvB/wXu5bXsP
g/An9V+19YwSmuQoegdA1vUQIUxuRvh50EqmmsX0UBap7/x9EF/b1/tG+iAsfkXEXVnmzgI8xrhI
YBxyixvlFK9AImQ5+pv0vpBP99/ZwjdCjcGi2/ddp3CqOSllDpl0BS2L0SI3+VAgJUQiJrHd9uec
aSWAwtNccsJNIAyOzhov9O/JcK/WOsu35oxRO+KLt8SVbgg5LiTearmPvhKSvDdzhs+iF92mlGeT
7826P93qFbAtGy7UqmImbXf2OTB8zHXYbmzQ/sFVtgdsgSqFWvr0l4OwM1AfTffnZJ4+iBioTZMf
vV4PxfxBqK4neTJFLkzQQhspWghXQicTa4omPr1wDU1vZ6wqVq3v4Jul5fn+ze2GMa/K1DHhxcnr
N3Ts1wgBP7R1qS456zfmw+I0iGwWFB9R8x4FdjWounTweWiPTial4vpkvFjMivIYlthCVF2GxtAD
E6Uvv9geUtk4Fxc8CET3h2ssh8VkutcZyJrwmzzoT7BilbegiaysAm/sLbpkb7WXGibg+pgi7d6p
UIxtbiMJY90BMppJ0oGfcQQNR0YBktsoTlxStptq51i/5TRaI1+idBcyrhWajJFaXrnvmeMfKyKi
NpHjbutk7MnmcBt5329IdwFXXNn03uphshrNkuthtI8trFDkg9kDdxeHyhRZSp39Frvkdo7Tmnxu
kfbs2YaBaqgmApdOZtsIG6KhuxHT+usZwqBxygfy9yYPjtB/p1Ides0EZIJEB7viD7lEQTvW37tt
rpKthZkbFgX+fdQtn+D5P4Qi/NrBVHKd500AR15zGAVcbIXQViIS99u50gpP8tktYOU7ykomSV77
BmcLgEAoy/viQdQPR5/+UXuMBE7hNYFqOuS79qEuZvrRh+pkRPKhD2ovuUX09QEf1gALXssjVNH9
XELhqSyOS0t0AHfyX06f1PHojerdmw4yhYcp1x4BZFZs6xhDa5I0uS0qh7UaLrhKazoXidc3OrJP
oOORaVVOJDQBjKmLX3KKHEfnWKhrb4zwKxzCROllaKdHx0ME95+vPDVkqsTBUhmv4/t1LeXvjYQg
vrbMkfbZmgpPpJhxj7V4qO9KHmqs/0K6ehOkLPW2IGKFdiHGqQt1/P+NgSbdO+13ghTMtXME86ka
R/bAncz6L4b0RcIOuqrGUNbhCaKAbTpi3COXwC1p064TgADdifM2hjiGS9SVEbX3yCPjFAGsIJhG
RAoDds+uHF5+DFECbJ4VHyBrsY9V4ihfbAGPnIuu6qTKIz52zEuO1KwFpCtvuqEhkGoNHMgZ7yz3
NRf3dsxMSW2BhoC+0xvhcxhzDrL9j0DtNAa0uDzjXqjfKDYVORoriSiiUcAsh/lm3hI2+Fu3Kw5L
ylKTCPlyz90ULLq/WaOoiESZwFTAMUpguaGejvAyaqzBS9H00dif2afZJmk226299sEsG/oq7bIc
Sc25wv3/D5VU1IuVLYJCJ0zkgThrvXEFcchiGTzs9mU5w7fCrSByt+c2072LMZUozkhsrru7mibU
+fx/wdobRtyvIzloQf3qb1R806o4Vh5j5cBA17P7GDUcMAtqJnVHDVQKcLBBiDfeeCyH44qeQJSZ
41IcGm/wtEwBI2iJHErU98VnFJyL2XRlxlpimXHZV13Nh6Sg4of978Q1whXLyaRr0ds8u9UjWQV0
eyvXD+4ENadD8s/bOMA7FVvHvphVV8xmZYpDGXfc8Rnl4FNTWhOpRqxBbnbEya1oC0Hkf8/4MFN+
ugmhaM0Az+UyMUwwPxH3EJIQZ8IW2w1EFwO9gpqeXMJruxTMwlvpng4ObZBkIk14Ah1JjcKAHxhH
UQk1e5iiVMg3IcscwkLi3v4P98S5+QOaw9wghLWDmOL7CB8N6siJ6WSGWW3Ri/o/4oZbt7GAM0ZN
COTXXzYb1N11VEc5cPelzNM+oGWKFcFH8jAQlCnwDPQ+vJCvh/k/P5wju04PH8jyo3FMU63CZLpZ
nHu50yPr6bDUNelaefNZjKdPmnr5th4a3HW80TqmCjtaP26QsZ2vHhoC4lafyLvTl49797rPPvSG
caf+2iZmwOFzbTdaBifV7mJbTRdfBZ84thpUcsHc6Y01dkwIn0gJiuYHVD0LgBsTE0LIytyxAeqk
5L67t8w1s9u6KE5wBY4J0N9DMZxxQ4c5ubTLTtBdqrTK4bW77fe6TmLG5NqwGnLDxpL+OH7rV7hw
NMMlQt7nz0vYyHXtdw8+h1UMlMokBVZ/72v/VkRZp2IndAUMKevF7b2rwUd7hEwy2PgrIO6MBnK+
O7bYIV4Tp8ZON2LcA3Rw1qmpM+P3J1euQUYV914p+9ng7iSkbl6hz74IDIULvXbuvTs6CVbPUxxh
3tYZnjiYNqgBLdrBaJxCcA0u1x2eMwN4EzpISbE2MjwMMxPpA2zhyYMzbn+FEWM/xISN9uoOWgWq
UQMjE4dVjcx/z64TjUrZ1hRc9rucQAY0SfhcFATXOMTZ2ftgfzcutdEbr2mSL+wEM8IBivrPvrzr
cHKEC3LnvnlJiewuujZdXvXhLhu4vo/n4V+OlU0h3XP64zGJfS/uXf+wzBiKDiN9UEVanGMaQQM5
tNnLxvUeLXRVUb6JqCl2/jsQWLpz1648YGBEnbx0hoWHte5K094dPxNsNJj3ro+jwJ71WhRvuDYG
ccROnSYTz9EZDnBon7Zr9R1qEAeR5qtN8DxAu9bdvtlHCaFUITvkj+8DIAPnTswGE+7s3aAXjnpk
V6+baL7bPserEwgCj23JEQeK67kDDG5pAY/ZHaPG1rWhc+42WGEPvbi2wi/n+oCY2z2ph+qdCN5p
F1ymZQsoaKJVYGNMjT4SiQjXHZUXFJJCEWb6/zfS1y9azfeNs6UA1Vx16iVXOyRN3Ywb74rvBEIw
3AHEXbq2pe2/8E2xD6V2pZEMNPiPtxWw3PAwN4gFT/8sXbnxLuCi10hdvieOxoRJ4i1N/1RS+sJF
2FbHk2W4t7kMt7e+HK0BDz+bkK0zycs1REdAsNTt7tTOA4Ad82d5vlcL6oeP2pVDaizILEyeOzdu
vWMKwwdikLCEkzbqpr+zX7yn/wOZXKgzh76NM1N4btxBCS/VK2F5qf19KzSgBDblR7CBXhcnQCRv
3Z07tkidz5dwCvhNDPY3CCMYe7D0Nx2vskIL5NM+7IXqvbdRym2R48N1745X+t5oR167UI9TVc/i
+YmUBRL29leD0pKc5j5ym6Tl1aAjYFA9z5429DP6INzd/1i3NhMXeB8A2phOjuyc1iQH3V60dZdv
P2qcRi1oILD1QbS8vvTMtTk7pGThXHEIicd3pk+yz71PzhYY4dLFss2DqGS2IqAsiVWbh7nqj0E5
OBGWDm2S1a/elreG8Id2lgnFkgmpm7VEq0X0g5/HsFWGnSCtgZmg7ZOZrzoK5jejsNox8egVvdUN
3XBFEkIMzvCl89YO0Im1bTI2MqCS3Lh93MQTHXt+nORIFlR5E9jBkUeNYpXMwiTW8X8gFxvPxSGS
5R6JTxh9MxQzwwQrlvTvs768JwQ5JlMoESq8zO1MIBqXXl/6DQrK7TS7ww9WkEeiQhmHnWoEHuFd
FoeXFbBxmEy7jDLxq09Y5+1OG+IAmz0mJYFiG1SX6BjEzx2WsiYUIPZq9N//OzDLy27zbRFVhyTD
0UBjU1QnOdIGHYdAW4BWQGQmbBCURQt34iwhC20evBDJmvgOmlcjEbxsVJ9uhTgyi6+gWLLbQIbi
OICgKm6nRGbHIzvCCgQks6xZu5OAG7lTQaxSRCEjo4cC4boELCYUgqbyCDrkmc7du5h5EpH5TGv9
Z+qrV/mZjf5bUkvalia/8hDpSmwu7U3cPXnVsTr5e0pOJC3KIn//yxapb4YdmIlxCcWTc/tCMi6D
KprI9n9mNnuKjG4b7juA2ELGhM9TJcDE7autxVIrrukXTc/cTwFdrfom5VhtUFfaSXqgUi+h8hQi
BPfWcdBmT3qjElvIWZE6EtPSqBrgIxdVgr0cvk3KcJmcXfPMUkb9fOmnglohmvybPhA3vs40LYiA
HC6iE+ZaKUjg/0AxM5a+amvROEMXAmmFVri91Ss3CV01Pod1lFLjVwaOJYzsyKdwAp5n2EkXqsbP
ao2Kh9tiPVv6gbEfXYzq3jLk5v04tY0qE3fPAtsSo/u0y3rTfw0KrjBlufuU3XVItxrt1RcOVx/f
BSBdfudKK+2CInDC8SjT2GBmt7WMYLAppPSzm85K6ZTchW/YgRRweUt5jm5G+K3l+c9WB2Ltcso/
dgb4qBJp9o9127mr3TnuHH0f5djSu5tc+7xqy02jvVlWKdCnhCkRs5tCG5j94u3zrduZ4PTjtwMA
QlVTa2viC6Z/mWd8vdZwhw+zIPCVvFPtynoEMXqRYSzW323L/rdwqHLyG4dc4hjc/J9rD725Jakd
MwIuBMAv//CnKekSS/VXsAsubdb+3/gbHxGD5ydVaoIZ1JbQsae9vBY+nTwiWQJh8mjDX1EYNKIa
5BdkqYU4xal6RiUf8HFZ5JDarnB8C3RsDPkVsEFbLdukEMndPS0Tu9Ttz5Ghn4nmxas1EJxp0gxt
m13ytTvjskvLYHXPWAhjEUtxfV+RNZbxpBI6G3PBl98dnU2IuAVQK+2z99MkdCEpuvZ9nHtmirGu
QbY56+rMsq5K6MJeSU3Z781g7Z1eJ6iHLKKkfJOa3pfgLdK4tAN8geXe8RA5G3NglYUsIOJhGSct
CeTC9AJsExL5BrlG8Lkfddy+cei7/23RZK899U/lyShWgKEEadXgos3WGCyfgrhYqWUfhMQrYQl2
413HFn2wslrZwwjizSLNSGC4Qbvlqj6bCIree8YdxyOiLoADA6iqOVaW0V60eVyAQ3jrxeT7x36k
V7lB79GjNnSPHyVZjD8E3vQHQ9PeZ02X4Xu+mXSBpOKG2Oi0FsEDzbqiYo3Y+tSZ2vfeNpN+8b+0
CIxMfvMLMrB6+5+Ix4amt1C9Rvj8zgFEmZXeoGk7Y3LtN3AlLfDGxk8EzMkB7SmQ8DUMoBo/v99p
LA+qvroCKeWxtb6PYn5K/uQcQf+gRAjg8TfYV3A1ZDzx415HXcvvHenEhC/0xQmfHvLFGGBgiVDd
RkBUKYLZBcdeI0iLj15rwXbaZm0P1+9jvnZQkn+qteA9M+NuZFmKGjmx9zuFUTEOS5nx5r8vUDJX
9iO5K4w2h0tZ7H742jKQ3wIyQRQIKPqWDrbFC7BfumVUXD/LATpd/TowZF11SOU+HLvqR7+rWSC3
jiAzCB6lWO621/CECO+4mb+vT1i0/OUxVYEfzPFoO/Hh5TaMBLMDuuwKZ43A4uM/syIDy60iUYIf
98JKdEsdY6DfylcrIrsYsAUlj6qzNbHQp7jOVZwigZZCOZdILqnpvXs8wzejKW5ynGSuQ93XUqPm
E+KiC46r1jeu2Al7+UKaJlEJrw1iwKxZ2EwGsoslGWMLK/6WJ4JFFtVW2hbZgj5D969vRQyaYxp/
r2zrjg3nJvBLwfmsFccmUJj9OnvSE6OQATfO2hzAhI9qwlFffDZb6QMEGkJ4krvQDaT3mz25cSKj
cG2laILLYUrkZWci3t/vKZ0QbBU+K/YvMkd44Lg4vIW1vZZsE+VosbYqVe/Pg8BD3qvprKHSdYLp
Hruhqwo7Q7m4FMr2jKdO8NQZogBGXvO29F8kRL0fD3G9woZ3tRDUmnRRYPmCsKGkxKkYNeQdbbU+
QDWB7/2LWSRZPiz/HZG3qNlanbbhWosO2e8oo8oUdEUJ2DCNDh/LVvbMbht95dI4kDruTN+ZoHnS
dmzWtMIutWcMf2ujW3sWiIs1zvhz2BYPbD8dXk1i5DGVS/mAwd2KZrQH9Xmq96XK3hgQdne4t1t1
Z/DnfVcrpqdvHV7QWQ0K6gaXmXtyUs2CjFeguysO+m51qxrC/IqVDAboI6KdF+Ds3vmLVXgsPyGi
ZHi/Wr+fiqOv+IcltPCotdOWg9NuJ+hecc7dKWsJmf3KFD2O+aLPIuz2Kv2UQmeyXhmLNCiDCZZ9
yOyT4YdtN8HOX7vocdrlCQhqlZaI+dDe+KsK1RORxqh0obJplnCEAxeMyDbrQQJjz1WW0roE0e7k
BNoQsOGJl2c1duPrS1COL3v3Rj8aMLwx5U0dgOdF0Q/FFrmGxH0YogVttaeZZcUrEbtzmP/PbK8f
tnaXSfiaCoNygTEdu9HoqMuOjDFvNOBZVpc0mX8TLNiMfnuqX0Oow2bHqNW5mPk3owvPs5YXqgol
PdtFsw4Ji0y9B+pBTwl+dw26GshIVRMtiqoQbmutZFp8xhj33EAMWeJ6Wl8/xTSd+/e4VBooGJPk
K9GNs2nQ+xl24k7ewxQsXQJH4mrZpFOb5ncZtW25aGqTZmaJ30BPcyYZLi0HAU5Vhtg6z1YNx/oj
qhXyM4duruXo/xML9f2D2Kk6i5+9WuO7C0aMEEXC9ipCt1VkIBbGqBIpubXLeJyQUZ/r10blfyZz
MZgCeL/xrBUOhKn7QkiLSugmq5CJdjTCsNoOqAMYDZoE64ApQZFYFQ5WykMIehJOqRQCaVX3xsPX
Dz2DtqeNF/vlh4OAE2DmqVALesZXQJpq1udbP3piMwqMoiGQTdhbMd9AaO4QtoYCiSYbIMgF2qW2
rTjBp/Qqz4zm/2z4Y2OSTehmMG6WRbin0GvkHTTMuU5iSEcl+cwHPyhxXmsGBZlcsXLmJr1QzHUi
wvPWVqQeq1j/r7lBvrI97k59Vb1DGqg09wTt+OkvvgEVjWN+AylPhnZq0ud7S/lv5eaTyV94NkEx
SUnF9VHogZA1rHtfPASd9h2jECrWI8LNVHpsMkHJZ+HpFK9Y3MZCxtqNI1/di12JD6HbQM1sDhAp
z18ZqNAlUII8Pgd4rVi8eXwZRhxc8cE9ibnjjQjTMqICCdpt0o7ETfXb+hAo47u3AlOIcqiVLl6S
mzvot4/VUiZdHI+upE5tkeVwGEJhvJ6Q1F7jdNq3oZ5xFDJaUZCrdmWL9mlnITqH7Nnc8+bMNK6V
vs9cRzq9I7o5JYwxV/zWspFwLnLY73YhcQbgqnoVwA6I3CBjBcoId7UxXW8nfbCxAMPyT7FN63Pw
rJffEOm8jL39b70zrBTrQs/NlrQrRHwsvx8OQU6EThPG1rUzc8IaTo0rsjD99iW5YQtJgUsXL37f
iXvlOcswHmiFa3ymj53XEv1oKz83DM5A2sVZ6gb6hcuRvwNYv9LtDabMxBzeqlYmjQI5UI6qcrkQ
/2+DtEgLSO0gp8Cm6yNKPUB0Lx/21fvKX02OIGizL69PzmAuGq2pw4dEwvm4zCHjLuwg/g6YI7QL
UdFHu5twFjyu99AQjrcg8R5aK2rjLAQHYuKLlFnl5I8+udu2P1RPIZVOIfdxR9OJBIBlPIB6yP1n
d2MrxejOWIfzuA3mo42BgdQeFMz9HRfRp9jBcWSSX79ppcKe0xbfPpr9P/FptttE/8F11s92/Hhq
0gYzwy/+rU4r9bPv/HYp4U9pzXPlZPSODFBvGt7Qzd1WELeRF+Ul79e64S6LBevZqumey81lkE0a
PlVdcgkRLJ0ETz6Y17QQXZgId7SSWGx0uMVrIbYyoluN54yd5PuEnSXaOFWzKuQlGv+9dxLV5MIp
qMRzEgHlJmH1R32XodbRfdNz4Ny19wcNpF03vkUpZOxYKQyrPvyKBcDgPXMv8rX/qiGZyw6BjBFP
R3415zh3Oi2MCB4WI5lwA/KPLbB/EdohTBAtazjcGWzDvClpkZ2PeKCtkaLwatbnEF83+8DQcUKx
kmtW7aMrDSgCeKQmCmEEyPWv//NzvXuhSbw6qEJaMcE2cGwxnU5jobnp91V/MTtNM+IhxTW9xCVh
/f80g50rbGtAJ/g58rvKf8M60X3GCxxEmrv6GYJXgpK5/e0bXI1XsfHRmM0mK7O//ixt0LyU4MIa
YOTni/6Jz4z2Uggkn+TSeyRGB5Qx3ewY3NJIh9Kk89ItfTAHBo3kD4pvEsE1LQsyuHHdXVb5rSPG
x9UZdsdpHlwUVIdtqhTxQWHu+oWDJDs1E6J3HjbqbT03HPRgS0o0jzj+3ourgGyrUmAveI55hXgb
YkGczCNY34lyXm5KIQPppD7yx+SlN2t8UxudCK1uIcEnIOPPgDVsVfOzYlNlJun2q4HiuPO0OZZK
+qdrDspNnrP+WHSLw1Wbzfhr8BLiBL7Djda4b2jHuTEQsXkAk8ojFeKOG5WPxXZvCo1SOaFB1FTj
2cSwN1ec437O0Lb6E7Yxlg0mGDobfy3kXQ0BuLvHDcUetkCMHrNZrgzHnaWY2NziFmIqJSGkn+d2
0pt0IJB68sfH6S9iOqB8tnhjmv8zcg77R4axdICnkVcvE/ZVDCWUqM0eqxLu7Zf10voTplo92iFZ
oWlHK4y5nnAFkTEWZARlmHQ8wYkzoNouXwA2scUmBfr7w+eSAPPZ2HnBn7/dnvLXEk+53W011UXD
aI6brkXGCj61taEBvFNRYVDaXEmSgNYZFsxpmdLQ7SEZOfqYZp2NH9qtlfnn6W8HOuYjyoT037w2
PSogMHqJC6FNv942UQHtvRofA+KaG3V2kCEu5eS72TqbJZRboeo0quDHxoZXrFvYjJfGSXkDs1RX
Q5P6ROyOESGvFBUSeWyzZ8UllBKhG9xG8rX4RImbd6g+v0PSQTrB8X1mDvThnixE+Uv50o5FPD5z
ke4fiz5l/MJJO9Z6/I79teCEddoSjndF0CLRK+wsIhLS8pdo+JAhORjsFXQGGO+fRTrXf1fArlup
eh4LjeKcTzYlTyFa5+DEW7GEinsJFBtZ9Qlt6sZVdFZImHpliNmQQWdisXgbc2dWbOF5XVlkc4El
9oFqDZxfLD/BpTvhEVvQHniucJS3y8ZkZ4Pl+nVliipQt3+HPyu9lWvElBQKb2FMbC65OzrqL6bn
XYKaUfKkfZ39SQ7SfoJcSAOYP0p5F00DKcMjwzeBnydxXWjmEbhba3QYLKzGbsM5Upkn85D20d+e
XY79Eu/lWKgacEPB1OF89Bdh2wmhZGWjraLzdmHjBqotDxS2Poa7blSuBGYg/xHghaOCjcufhvLY
d1fRhnLhBChMQ6tn09hZ9isqNoOBnkMpEQzg3Multhzck2SkMZ71oHQbUwECJZ6JTdzn5CnmTuUO
HDo3vc+pEMs1cIi4xzp3LIuxE6Km16KyZjaUjhD8c/vw1mkQNWUQAcQxdnQsBQr5j7+/aAXRdVTc
EhBWDzje9YDeowfk35Y6fSFIvcYyb6DT9IORwPF5kWHXCSNoT8obQ4LhWCqqVKU0h1w+hechS/Xr
dBFA7uyr26JmiJLEH88acoT673Gijg5JrUyPWsT5fE2WS8F+CJTLqL09eLPMmvLph6OiU1TfjlHJ
hshAYOT2ZzPQnCaM2yHd52mv7EspdtcukNu0oSZaejR5NxHNr91AiIWGeWK0QlSRftMu3b51NTzr
RZ7UqgsPlZ7bSqW/Qb1xI0oWSMSPFR8yn6+WULQcJDRjeEFTnQK43xl3opkgkf557NI4ES1ICbYY
4iqZP41u0qG4XnIN8Miug1w1RMPuYBs7E/wjneFISmpwqObajzo/V5qFdn5VR75BEdC+crgTe5O3
cpaym47u1Chef7EIo6S8sCuygsbigf4wd8OQwt0RWoQYrdymPxhHjgVdEP84s1+YsHmcxIvhf2Ga
5/oBg735KhKHSIvNK+LUIfTdPdj8S3JRIdkvTgK7woqiu//vRulxBHLPLXLqIYSK8orpEI+te0+1
qNA3p0JvvnHTKg1RndkCjFqPy51Qsr62rXvaE2TFZ2OycPjQXJJ71Ot9bLB8KYUpY5HqrlE8tLTK
Szl23TQ+5Jn0JyWcY5jHJkFGehyU5eulmTkrIQJpGEAIzDnwCnpvLWcj4WMKStk9BK4xvftPtK9A
EtjUDFzC3XAlfiCL8LWKj54/Ib4rEPWoZCvqGvCfyk6LPq9HieJITCZsnanl+lk16mT0/oscm2nj
MtDeIjQHjg+7XdMTvu0AAkJLpNzK70BRg/4aRSmTQ0E4hgKXjbXZo6EkaIgPAUaM6bVOK81C5GlB
G0wM+bTuXxAX2Oz0PTteEaAXUZANXnLFoFzmavfbtiicaO84/sGT6ptnGkZsoOh+znr1HGht1kCx
FQn21BYLh+GRrUVmwCico6AeV5VjduMKrFxdtoWY0jQWJz90W5O3xueA2DflVU5zIAEgqbH2iDjB
pvtSEtRzUWhUKdnlZ0Ve75bKxVwzk0OeharKcUp9dYpIy3dxvfK31fDLQHajj/veKRqtBO7+Rb/i
cK3pXXJFaUD+E1iULhVlRwEBG0phEgt4POj7walxDlSJIjtWF/sUKxLHJoZCYeaPaCo73AuYsyal
+CO3zC9T2mC0CkGAsGy9r1lYmaXcuqcclhKbwK7VnrHqLakaTEXtAEMyaauskTjxf71BSH48azfr
YWEh22i82B888if0lf94jeTa+NeTR+sbOOIULnybyHvgXALhRQ27T7Rh3EliaULBQ7EZdBK7N1m8
lyS9xlwGe33y45QBvWbSMf8L+nt/BWfANdyvwgRZNt73k8EMtYNDqVeIRu+yg2fuoDmnA6riISAG
wwgQyETSlfe6LktgPF881+RivOinMLLhgKQDaVFU8sNsssYWwnKzYjWNDkERnaCnZbI4ygvx8hHf
qB27iasteueqS726R3H5HbsWbkiw8ScBY998RX9MBrO+zd8dyq4ZJ1GhtPWC2wZkZLL+0JQK3MtV
wqilrzq0Ug7dDQ28NEeRuzl+vp3A4UprYVTa5kHgyxKXmW7eFy+6Wqs0rGOnD9OFR+i3MnzJ+PO6
CJ5RQYJ0lX4CHtzdpqLAlyQ1LBMYXwmBDg+lFZ6A58Aiibm5gd0hznE0pY5oVrtHxdXMvFSYvO5l
qi9jrJGKDQKQ8PZ7sbhDbJcwxkMruE+8kqnVqRLsg7+EzJi7bB/2JdO7XgYQ02woIpri2L5Jcu4Y
5F/RVybNMhBO4QSaXOGhVAK51vhcSeaQjYc5lfY+8nulimU8QCFghJTjc77/nvj/dHKkAbGbJBoU
nvVSCQQC5vyaamg15MYtjcJXsXL1MOsBVOwOjUUWIy4DPY9iZwFUgYyGj/oH6N61J7XTUh1yvFks
Mck8pgA3LpoGS4ztYS4ciuarXXPvnCv42zOGVHyL0TglSXm0FYgK83xA0f1ztwy3AlOU+PlUp+IR
nJ360JZGpAf7W4bjELUvNFVHtPtwBReXvZutrjVzQmT4skfKh08U9lL6MnUPqhsniUug92Uet6Tv
Vme+LNP6yg4wSURddZrhl/vIMRS4r3EWJy8rAbxh7SbKDCCDwIJM7H2GPMkDaBbSMl0GmTTWyplo
eAu9juumowdTce54909sjRxSbcvXLFrtjZo/lAsn5wTujJtjXRyw1ImV26IdJbIrqYivNYPDhiBQ
IIcXky1fMnV0sj9JiD9xzagOAHqb/tjb8y4i973oDYyG7wbVzlzas6gYtms+Vz6nQ0klN4UMFO8T
9MSRKk+MowxktE005zEAa2nIEX5Gvg8DOPrLeROWW7jAV58DEGG6h4d3PrUuMtlNtVbEpb66jhfJ
Wl59jh7bz87djuW8kCrzo0unDpEEjNay2joSqrg2nxLcMVoVZEXXJdZ8hBSdmGtqtiFel+kCzMdC
7FMPSReh4waM94PH7zwTDGqPTa9/Sw5Kzj+5/072hQFHYIudkV+H3EmyIGWRMixFMcolPOHxTsrJ
4Mz2tX6m9s+8T8lVEkw4MD8T/IC4HmfIWHnysRwmTp5ZCbR6c1bi73lJIHTVCk0/ZqJTVomg9OnK
kMaUwFs59db2GkOf5CuIXtSQ7W2fcdwsoRlQ4Ewl/iMI1EUhPDK6kWBGAZ6DqnqXLSb+BxHz1OL9
UIGniyrDgx4UAZSPR8KmBI5qAopf2XlUx80OQw36SNNsW+G8Do8rSBJHVRYLYBF5I+M7bgdIpfML
n4zjmnhctQK0P7su+4WCzqOCyvzNuM6QoNuIRkiv5HFE4IGOaG+Yh/nFFnGZMpf9yVfsJFwpJp5O
3WxNiE3SZjFqADsEwWzND8J/67p6WIYVbUMmRRIkgcypa+p3tDesm/j/MIwDM+RGF0D83izu91L0
QURkKaLnETcH7PcJrGUrZsFfUI2CBBboHtpKA0a5XXNbvuv0cvwAxluQUqKbp3pie3UN8uHf5UZ0
Hv0nKIcqP/V18VqyosJm/l4L/ho0lclioTa4sYIN7DK4eeqMD0CivKmsixVQZJQ/A1Rm3JNg8rWY
xLrEJ7GJgTkb09m/y8iZh4xLNHd/V8BbFy894Pzxg4Uu3b7vr8mo2ROpCp4cwinuQ42nuWgOuXWb
Ur+DGtVZ8tF1ou2bnI4MvE1JvYTdWqBxVtCU3GUZzRGduWczDxlauQpQ0ODNuCo3ha+eSBZxHDgV
y/g3HKxNr+nUrbjnyQGWWlRsawBUn/qjyBAg0p86GpQFywybVRnPa/VNUiB71OsvezuBZLZdNXWs
ilUsbDHMzL53gGy7N0hKs0k0OWOxYodo/rUHyvIr5DQt7DeNfLCHzYhMePz8Y6lcgz74Cn4Oy9kx
gLUmvaujcn/wJJi2//F9PqN5C8esqEejp4hbqk6EnoE9ynT443JsKSJdGoHtl8xYncvWuJiy1h8m
88zKzZSV7gLf3zK6t/N+/7p7F2WuodMieLMdX3v20QklpvTOPQEHwVc/BoFubSE15wH2YTERItVV
X3jPoLzkH9/0qvneozIC0p63xdULibx+/ZfKc46QvJzrlMw6GEx2nmkRdqhiAZMZxTW1fXhu9Eo6
SIF+j4sJvvWCbYaVzRYGlQJsif0OlqFWsNtp5tFMcK9ahBSc6zA355J2fkOQcYefmymDcyxyvHqi
hK62n0efudMMjnyyuDxR0o45ASBojrkGPSvoDSsH3LFdh//v9BOX+UXo9A7xdKrZ4vENk6zf6VNM
pYwz53tV25iP3YVXyDotSgVoAYf3gj+JOoLzb7hzrhOkByt/AbDrsI75sKKONrv+Pczl3B/xgzZh
iSfMFhbRdyn18vPPs/f179xxRU0ipPq3egWFRlYOOuohAgAYdOMA8KNDp4WgFtdloe+7qBVT5PX1
x6wuOJLHTaAn01uVRUSH8n8nNk71Tj1EP7n7uiuE0cyyVkYQ+xHJNHxqpDJR/0a8QqwMRYJdmiYI
GvYf2B4Tat0fzmTSQlJQAG/Ts3BpxH5H0ZdgHiGtB+JD77nhCEuvXEGPeX84V2vAI1ow3QLbM/tV
QK0gro0DXe9+zN+lvP4xN4d61i1+YfsE6Eh92dQaEg4fdpEA7zcf2ymZJEHwQcvSXaZ/Qqx4TYPp
P+OwZlqzJXqWDXxnyqdjopq+xcV2AdDc/QiFEfBwbNpleG9lq2mKd4rRwA6xYcQw4Ay1O7ciNQzY
+Ft6j/yq9VdA/uolXHQCoSxfTCqKM/chJRKfl2NizoqulK1zxQ26rNkGnzgNIppz8D0UVIvftR1N
jTaAsypgqlg2WQi+fXXeGsN+VHyJ85ez75mFchnNeiRFSMDcv5Y88G/jpfBqhmRQls5xwMbTxIS4
0/qwNciykPlwF5dkvR1b9U1ovkrx9Y7XGyM4CB8LoT2HDBvCwSkl/tHsq6pz7B3/LE+l2rnVL6Nl
6y2VpeHPqs5bpyqTJ7c2+mTzgCFZp7GdgKK384n3axNxl810OrAlZj8IgEMMhFyDGHgNUu8lTqe6
Fp05ZLO6dQsi5f4Sz8uuXGharzR1dqrjwPJ3wBo5m4YcHzJPo4WnKFaYTp6GWJVVPGo8jFaZ2TxQ
e9aDPihe6XLVxpmIR1y2m7w+KDMo4O2Wo+sbebB1j/XML8h7vra3GhnWkJh1+chwsMGEMx4gdCFT
Q1pbgEQPWwoHAIq9atjFaILQVvuHWjpA6C/wIZqrqb8ZYdo7fdlHYChXpPh+3qKzc3uEQV2p5O2S
Q/JB7Fz4goLSZhAOiypjZDiGbViT4wCKlMKKNo7ItrS1Gdu63mvycw9LfL3l5wZs4rgJzGDNZVxZ
x89HogvUrqMrJzT6fGAiq/wNnLkYlIfSxJ/Hc/VbHpti5S88c+R45h+bQS9b7blFAcFL3EN1NA4a
CfTeEPSugo5kiwAsZe8vTNJC5rEhmw7ktGKnHd2xh6vZy3Li9RNCzCID1Bqe8VDQOvaUcHneffzg
i/e4bvQv+nK4X2FvpJz2GVZEUKsLdrXGmnYioLkof0haMdxe7vV/G4nyJrNOM2amnRYC0RdaybxS
ELwkYLgYzdukXwaOjVzJ/LQ7Ru6fIZ9KGBqlX09GN7pJPPWCc+zP51aKrtXkDgQ/oElNqe3we5Vw
vts1Q++kjZZl5sya5z49apKc3cxuywhcqx2KDesvihbMSCNUMXlhC5uwi5ZkOL1LKJpiDEKtm1Ob
2VhFYvbUam/1qLOcjbeeIXkDKSr5JquDftDeV2dTC6JMIXaVmKkA2kvtAvVDhPz47bqqNee0KTah
Jcb2DjQCyid8+gntxU+BYvcetvZqn/rUYJ1Jkx16y+SfXpr2Zf8petsw9rKRwi+85WTFUavxx4p2
f/H2QPG2MusiVmf7IZkDMEQkn503Ckga2qbj9M7e3CWR1zpX+8oaFKpMwpmCRO1orfT8dbrz/Gji
wPp507XSHuFRBTTfl7Qy7KqXY/7OYkWO0/aTnOk7wHIjk2c3A0BnDLwO46lbGOVSt+3nJNntJjLX
0U8PwhX3gQxB03ABOdk0Jccc+rhfJHZsFWx6KA2sFTLNDsB+AnlO0P01F1ZB+F5Blcbg/gLeVygq
++cio0qi3F/V8QPW5TsjpJTmeVDtPg6wBcHtJlEYDkp4RJLRhWanDHS3NsT2wTQ4+1QyxwyQXo63
6ypuoCKa2vGDomaZeeX3teayWsY18r1Gz5k3ECHTAiUzXIkg09F4ZqYZqOyDSsuJO1HszAAIObiB
FFGFVtg9OajIMoQPcNFYxxpPQHaqkFR7N0dhcrJ6Ekg9rZyeVEai/JvS1FycYuYN7Cbihdor/vmY
aXuTgblLuualbWXbu7Ykvkse/Wztpugn8IGuURgaU9qfgwBKaLxGX5F5ccv2oyxwmd6fIpLH8LPb
tHSReQUAILtxM3Vu4RYPBsLlSoEMh1udY9o/2DnaLd1meXa92EwWsO3Y2lECm7T4QUKUQqaWnuTD
LfqlYk4UNc+SU7DtsTn76c5HVDUWfHJq02dOLwdYXqtOh9GV2B1XJEkdjW7Ok3MzlT/bX6k4Z1yZ
zmDzgGutOCPvZlL0ZbzIV8Sz47jKM8Npiai5FCVD+xrrZi65B31QH9uj1BWuhy4WB7KS+OP4C10w
kos0GXI1i1zc/usS5uuxb9QxNOb9W95G/BWTmjw/mxvUBdunkFU7wFvlVb6hFCq2gZaf7XpCQSZw
ItHUxdKTbNnos7ZujF1iRuK7cUy62Zzm4Q/gdGTcXf329sa8kecLn+u/ih4EIP4hxOMB3Tc5N7k7
flRgsWU+uRCQ6RMz4cei1iVMsO3SiH8kL2r3p3D0uM8hw4rEd/omTKJvRWwMDchEnSSgtlzaQC2h
9K5wd5yscNBizRdWHF4FEbZjaWG5ZcH7QJlCcqyyx89BfTk6NGqc7GuhCuyv5orpa4H6Whr13abM
k3bZulDtEkqXypu48DiBjhbpqokcGc3PfImLFPFV+EPPFFK644bq75/HnzZ+qCQxo/iIVOnK+XXn
DJ9NXsU4QB8aDh6PZmz8pwzXpGBU7sXwFF/A6Bg0YMTOMTQ2W0DOpluFq6o/eLWdwhcsWeX5C5CJ
2A4apQZgEsCRU6gIMuLQNYhTiv0jzE5lmaoEw2xO9J3n0vHkVMMIkIGVn/jwLj9oYlqgXqnHQoSO
NTwmeYbe7wEBiwrdkTgEJYjeV7wka16WqKRFj9smc1MojUXJ+UExVo7wGB4oMhS7YNaeuV+/OICo
gExwnr1e7c7kETL+I2YWod/Z6VoI4Ak1Sovdp1reQbfHCtLk6Cn5oNisjV1LNr7rQ7Zyhq0UW55W
2S1+lFKB0Xdv5w4IiO4gODqkNt2zIcQRW1QzztWrF9Z3km6wBRw0ylC5kkohFq09S3EitGuGFgb6
UKx6IZFQ2KJUVW11dNyo6mf4BHllsA7RLJSawj6Io2zGn1HjODRfNTN7hC3g4D0KP9hTJ2SxvshL
WPrhH1c7mwl+SlPrPC5VRSaaDMvUpY7zi/zSTPmgTq1vX5C+315mmbWeoixM5si8wTfw77fEGKBQ
zIs3tjwM2wYO+24vQsBcN8l5KYqbIvwljGaE7RiGqHxTbnFB4Y7fL9tsyZNAmfHOmm4hVxBMEYII
pLdY9KnCWAiCxOG8Noo7bnYTELLx91oB+9D/y/IHsPdRwSQ7T/M5H1Ih+FhsDstrlhjzfMkoqzcr
HJpBbjiTxdsozp3dj+3FzDF23mqGU+eeBj1agd1mCxX9tZ8YEs2mNISkh+kmcs+7mHsC4gArCQjK
mAu+M2/6j9vHVczQKhOYlmtz/tu4lGdXrFW14uNN/uaY+j/+dYZfoLRO5M3jWl9uuEcAlKmKzMAP
+YELpIH2w97J2jZs5stfqZTS9J06utwx0RP64Y3gIiaip5BUOIwHOYkriWo6ExQHC+I8t6QPtsvN
empnllva6CGLrFjmn87YefoqjOlb2aSo/D/JUEF98jfj928rboHDoV5LiPuXJiv3R8yoM+HqFffc
pPyAH+6apKmbQA6AyoJJeJkByW01RgEX4JPrxTL0lndsbPPcNX0UCwojjiphRqeF5XENMuXXM7R4
zOpp5zL7RzbdNHAg6PCsy+wV+2fIxVN55ImMMb6nIL1D+WtZmLqD4hceD4c87w9Wbr4Gw0vJBOaV
9HkIsj13KZRA0EIT8QfFzWkbKNy5eiObQNUSiuLL4cMeyFxQ5qimeVzKoVq+e/eGh3Ps0FlQ8fIK
iZsUbX9G9f4j9XYOjLxmCof9eYDYtqgmd6jnoYXGBPT9pKieUX7+yyf/EDhSxJdL2Qs2ELYwXj9f
lHGnMUuunSUL1e3D4PG7DKyfBuPiutnJBZ7jIFkW1jart0eoRjHHTxteCGmf2fUDj+XcuQq/uSNp
uJqaDH/r9XWZ93zeFq0umRwD4JbYyncKG+5FzuuzepkgOGGLcDGR23WV01tA8hv5L9LNqB4ykrHX
MvYuPO7Lp0Of1DJphcpPgm86tFyWE3YIGTz0hd2qeXaWl66AjkJFqAlxkTi7ANFLnnRlHbp9d+x2
ymkWh2uuSxf4z8kvjuiYY/xlnqIORz4Suz1mUX0rlE12oyqr9hZ/gqZ+72JRK5RaAXog0DKR3x8B
21X2GchGtdsfRDyMgmth3AaimNBfd07D3pDd0eK3ObodgCMC7JXNNcgHfUqirWvwTUoLoEbsNV5T
uKa/6ruXqbTKcWx8PYVa2KtsK2TxOgGfRTRpBmraqOurj8gyWsWFL+832YsA/iA+CUU69N2aydYr
w4FYr9FmrnIv9YzrwG904bdjb3o3KGdjOvqYQHgAs8Y/hTuRASLLDEiRunhOM2Hoam8WwET0NLev
lVfVdusVDjf06mBx4j3cr3QcnikzlOiA5r9CpLT8BR+AKKV2Tb+++oVae+4x0+B1AUI0YA9tjMo/
T4CZfByec9AV7DybMdevoRqueW20mGfSb0pkohl/QSBn7y2to6zFtgAftn+K5ccNJHKr/mJzb9qk
D6oVNHP3g/g3w5jjyZgnFwzKLaNG31EVc8UnLespxcGv8e2usRjSwTrMdJUC64Zmy7gfmna6sJql
FjSRV8VR6Zo+UPnrVwIpnVOT5GPXjUmkoGQy7eSFUQlVS5uFk4+C/PRcQKxLgoKAp2m0NPAw4A8U
Wx/Qv20a5aA6dvptptV9S/ZBhvT54tkvcLeQTuOg8ZCQN+bV44wMVJLuIDdYkvRPEW8iKI1X3OO4
TKNvP/jXZyNza21Z66BHcw62lvN2YDDnkUq4P5QKPWSMbr3U93Py2NAD7WAakTa1CzbDfRexq/MU
BeTqKHM9YwXzRAxGAiw19cz/LEvlOgqAfKmMI0+iE7vkRZTKw4HueinX233Na3hpvoNZeM+nzA8I
Ei5+GlmzJKWDNdPkekrhY9rtGmTFgfmZpZQ/8I9u9mkcNDt9qYcFxyIT0n7ZQ/VFdMvd/1WRgNHp
V+KGHWmrfLuKeBJkjdG/mPYW83lbsQBA0vO6LyaJVY6nl30i52/X6ijuhoxrJfZY3Gia7eVB86K+
fJU3F6+u0cxZrc4t4Oyj9X058m1ltrTE3o7BBpsQ55n6ckWwgiyrafYKtCWljkVwnO3MeGVGBO56
xR7Hdyl5urSIWk0ZKoez4+BDhmRNheAQjSORXpBpwNGMZ2EP3X6quNDqlLsbOEJHXZHKU5mRKuIa
EpbAtvTgopYMfiYjyWE0ySGi7AuN8np8DxrbKj3ytPh42ngVIImVg4Y8tcm+9/ydAFNYgdAHeJxj
7J6qIXdrHuR+u9K4WtTbKMRADrZzvRO1Xl9jIBj7Cv+IbCOEA8hySurZvrH0KIUzb9YlibuPf3qS
d5CNvUaSJ4KasWJ/pG4hvkF6fabZec6uISzEtKIhCul/MoCfr/+lQi/PEgOgCpRYb5k+lM0eMYHn
nBDsXjdwe4t+7XDPZAA9QnrtNwia1DlQifxbtCbWRoEr07zP6mMDjdF/V099tBDEFs9VHDj8z/U5
4mGjTWYJSv1GEIQUzkO+n7Ww6MddXnisiwTdSLTd8/7wjzGAk2maXCQwT6A57kO+q0R5Phtpk8Qx
Trj1Ybbw/i7NEjlj3ivXFrfPckICgb+ny86Stz/wS6cClF65AoveySPekle4PYzlWyowPlscZTFh
HN+kl7pZTxJQ+7YEETaLeYBGg1pqe/36nG6BCpjjLk+owe/bnqV1fzxStyzNj6FmR57yBQCCg9f5
n3FuFAh+vcg4pmx/MQrtspLQwKTqMIdxfnFnwAhXTWhEMH1JSrgh7fjUh2mHWejzw/0W/az/GEa7
89XWm1Y4b/9EmIg2HMYck6xZTvU/ckuQ3ADe7l4UtcBPv0wELs4+pQ1p81wD/+/TsVXBNgC2Yoj1
4lqR2jhNlW4muax/iqRDG9UM54xX2pXcdNMepA6o8uvWKJXgGC3bdLzO2H2ckoEF4oNddodsODdU
bYu9eUddkMVEBJUfngICU4xlDOQRX9Ck2Ya9KxqJ0tWY4Xdr7eYLHtkp7byvJaP9FoHLeOZikU4N
C+fNmo/CQB+UagSXiWezKUt3dT7wBsRUlNucPXRqVFlHY0iwlPGu5/X8vv2UNMXhp+dVnP44Xbpd
Idt1EOJAhwgufZ8HcefPIJ/9K/Olv8N675ezr6W5De/uTEF4P/pdVOWPhhWspYSiZh8iNMeDjXwA
3TALosLe2aYwwIpLN8JyrqU6BwHyC2z6uT5Q7SfMgfu7DYDqWsFVnXyNhfBwdtoJbJiIoP1Aj/Ay
qX30czB3Lk5K2VQnQ++WHFiO8GnkZcCgtzxWMVKpuJi8G96gJAV2MKf3i+alxTxJUpFhikEBTzQ3
bWz5d+i8L21vin00i8D+kLTfUJPou+i3W1M4OGnQQXWGsNUwC1rMNTQQ8n+ugXf4y/x8dKL0D5S1
tIul0V9VGnfRgIXHPIYtnT3i3r4DLt5tsmwemhjw0H7fTeNPOjDagEevNH2TBeKPR4PKg3iTI6kB
1HZlQxnYAQNc5vBB9w5mw64jht+bmbFRMwfbF0MV7dogOM0EQoAYTIx0iZuxHJqv7/Dg74a1MK3m
q2jSaaT7QGiQAuG9ODxUEcRFlyjUNAJcZHhBMm7M5xKv9USlIhRJ+eTOGbtSHWYsmU1L5Q8h+cA7
QbIfi6HA6Zv7RtAoj6UV4Ik4AB0DIFILqSNj9B7lVP7sd2hAN4/0vaTa8mQcW6bMhxxNYA47JEBE
pJCwK0nVdYaolpiCwF9y1yvVR4ooxWh6OONRHLKIour0732xwU/ovY2dDMbK4VBq0RjGvFGb08+e
8fbJxPB2rFU4Mccl7uRl3SWFRL0z0c1InXhQtScVIJ0Bj0BFYhf+/b36iEd9DcKl68Pd2RXD9zzW
7N2a91jVMK7aHzxglyji4SCkmiIr+FHpNs6dzo1CfxusQ+HMuQAgywkFWvrUiQzMKx/yfvB81daG
jz2SGtHfvCvnJY7Xpj/4PX22npJtgm5fPE2T0Ac3YE6pSWMsNmU0JdUtIDW61+8zD8Jl0ttjEY6X
pLRJnprTCEss7viBgCmUIltnjZs0vacRx45P3nSfgiHltQ7/BvuygxuzJJ6wly05E4jxhwimjBeH
uVB1XVOPpVQV85Q9De5RupBII93fIfjlOrRzQwRiQ3LXBdR0VLDkKbGBmNqgyoVigtgbaw1cUN1o
qzBMmXWTZG7h5/Z9QVfDzvR1wlponbIgYnKEEq7n67uQ35mTkG7lC8wExkVaHG/MU9HfbRl174ZF
uAJUbkc5tDGGjLBKvxH/cjHcLZUIQOY3cl5uEaPPVOWjmJWu/IOTxWTDul53DqslUo4RV8CcyQ90
W821jrI/j6uSd4HgVZx/Hv82IiXwedXneCPacFPghi+BSiO3yzBRY2gSydNju34vF3JDMaKKbson
kANYOwSdfnVyHRdh7yxuOV0M9G+GK+3cCGtUb1u+/JNwD6/OgQaILLtsudFvDiwC2Wy5eTQkjaJq
PEA3RtrquM8By42YtolnLe+qir/4GVSYz96CnRK6Lxh5xA8rkZrcBhA71sQIGJxQ3qfZFnmovPuu
DoXHoPoVQAyzJl4U1FwoOV/8ZXyO2IlvHauwNvc16ACAI8O+zSEHpXi3X58+51UoHWHf3tAxQWDB
0OityvNI8gBwq5BaWk5vN0QiODnJ/Ur5G/+T1H5oPIxZTLLLCol/NzueJAGqSVk1vSZye4a44aek
Rg1hKdMWL1zlxOfczjTjeIrUJwb0Wg2OGdNi0tVFWK61qyMTfOtYV6aqz4uBlqQcjs/Ys9Yu6J7U
31EaTMgkHRaLwTs9V4LqvqAlT+vACnshaz+ihcbe6/dDMn5CQBegISfhNd52B76z/QXZ/P5H5nFG
GMiGpyYDlH77Zi+Quqr/X/yTbzURnzj1gJLaObrMXoSu188Nq7FaEaS4TZ/T3Wza0GI+K9hr7Miz
HtqA4Z6ERkZnbRn4T0kjZ+ijsuDp4ZulqgSGf0IKgb4ow3Yw15Ga0uk3M0oz2GV8cJdNF/Xn2/QV
fEaUn0NCL/VwmZiBTnoqjW28bJI4SS0efQBoRiyBsBv612QmKVYpPunQ1DV4JS9jwmBGm9nzlwOT
3SmlQRR6BWCvguEHRTksznHnHQ0hkcfutzybOggwLhNhcXuCDFCFCEa8E/UcCv4H7D5jFyhCrUV3
Snq/tcMO1rr44+qCEIl1H1moY1mhav2ecubfiZaYv1CfdHOGnT7Am5lk1B1eHkgBJ0o4vGdsZw8h
89+TAVaJFcpDwZ/2YxOgp7+T3+eO6WOcUPrLblzYcJwq9N2sSggJIOVBQMTWVtB3BapU7wEzlTkE
lPuONNafyZWHPWupRbKt8bsmhWThvaruwXtFCn7HnCNBMrzm9t7ikMF2r01tlwrEuXBJk0qPUXFO
sp0FO2Tjdalv29zKNiU1eE9dH95wUyo8EeL4EBuc2bfeUsP1nfkGY7x2VuazWIJmd+RjDn4E2EAn
lKcH6qtJOLxo++qxbzXvMjCh49f4b/GDqOz9hCJzlZbEVeH1WKmIYIVvcX0WBkYeTeTBMBFu5omU
9lqLPl/1ahaXBNjZhZwbpNQfniHw7yMYc+Ga/zYN5/lGfZESsX1ZagVg1JEdIgsVqzwpI1VrpmqT
d+ipN10awJcfKGotRu8Bn7Y3nWjZNIKLW2xU0KzThhPaM6QQSZx9LhgfsDbvIYGxVZowlQU+hfMV
5lGwU5Z/6xSIdT0zgts9bCfZqG4VhkaijECLxFy0sVOpwHWEXPPIs44tYFA9/ULSpWongioNglPX
dh/B3ZQvHf31traBVPcpGLlebsgx8Fe7bQYeouZFO+D30tpYg7ITB68tFvH09AlA2KMWVsLxDXiX
+gkjJnspzido2x4NQsnhNpHQtrpQvbBs+/pEtROMGEmbmHoDkUia/fRe5DnBT21Q5FT1S6H63wlh
VX0v5RHcrcE+wZVyamYpVZekal3S5h/+/HbT150muIpylOjgsRppNIqTsIvfaPeea3rHMfh4C+5H
nkxwG4Os578H0NJMUU5AvFHVAklzvmXTxBW6e7Jlo0ryywlBqYazmtnzAs6MSUDwPhC/HEVZU5hd
1QuxQ6h+IRwMU8DGqjfMbBaNkbKqbVXkNUeq0mP4q82JAaZTCmnqNk4qGITGdyw02VSeB8Gq6URF
b7RCqiKSMzczdUnoI2neJOdGCE5fOK5qfDt3FFwD7RuKPKA5Xd6k0W9emMtmNQU5mmEenJfXfStq
HNnYKrSa3bGYqbYVOV89V+HfSkWgVC4filwN7bxb+mrIFyQ9Un1WNQG4j3HWIQD9WW88o8M8g2yw
N9vNdnbVI+hC7d6zs7RAkawHNTDO5qC5v+TJABJa3VOcN5nA7wFI3jXpwdg9mfPjK4cFx7OO81Bn
gLJ1JtNedLSUMJP4UircBGMJ4VPM2mIyfy7tx58DNvQHOYGM6rj/4yx22jK8ERR9Xt0yRmTY9dnb
duc5Mj3UrXVHYafELnNprdaxozYoyv9z2UgWeqBZq0ngJ41NnBXw2158J4PQicTaIaqIaeIOR3yK
VNp/2h2yN59PwsmojcbKdPccq+BuAe6oyQ1E7vLxAaGE4+vl3lDr7nhxceRXUSEvnJZR8g0PO0hy
1PLwUdKwv1v1l7Q1pXl/W/jTgVv0/MZSGqNoTKle/0sVxOFf0n0HK1NFkSp7D7NpryuqaPHo5G/A
b0HlAgayIfCbpcGaMNGfJDDSuhNk79U8q2kmxD+SycpfeUhh86b32xxpLyziDdfh43aU8PrrOhR9
OKhjo8QsBg5cRXAwTQ4m4LdAVPH6GndA8qtVEeL4bgdsHIzjFVFe7VYDquJd/mdqF4UCHbPUefQi
+ISqyJEEBsZsZ4n5OBO2hTLCMnTW/cikN2Bg+dvbk85k+BPAMY9kzZjT1JvJIWM/wyNJSttJ9Zvh
FbHK/vimjcWRvVj3P3D3b2JapGqSDb1/qXpHMWRA5G1FzFLfoO38OGowo8tKgyRwOJem6dUsvQCv
l0X0Zg9EnVPNTzINMPic310e01AgXdqA5Wk7GbTiwlu0o9gvIz6MBmv0RC2XkDfff/qAMPeaCe3r
4vpw5Lcf0o4iZovrZPD1XSrINvv3cC591uazyOWL5tC2VHRtTeySjEUkzJ0+vfvgIE48mimPZnsR
t+pudRnnctBMizGQvR1vnnlXyl4ByAvd8Pq6IQkucyMbTu5Y3ZU3JFtERXsVGxs3vDQzbl1+yNPm
g5X+MX1OhMNUihQ+5EVqZP1wd/J/eMUvfQGBnxXy7LRopqaXWbYrLioyc6a3AMqr7Gcnt5LLy963
uSEX7jA2oGXTfS0BdImC2GDxB7ANPLPkTcqamdXm/+SXpVAPLss2kW0zIl/NEJsJxX/lUeys7f5R
qGu9i4PXwxuqVfWv1Qotu2JvKYCAxFIVInWcWwO61/Y66Xx/fooPryNa8qzOouGiQXbwsaHSIpKQ
2LOY6K4EQhnAK2FzYvDqQ9Fq3raxqhNfiahUgI5IO/FWOqAwndglw6BGmcNRTc76k2UFqIxcWO0O
dyeE6D9LpXYtWVUDz97CWETtb16rzhh8FQxHvVftFnUXP5C89Zl+CjJf4ceZbpRcK3VJuX71pDIF
io+9+jlf6ajka8rD8dH48+abC8RkO1mO6snaN0JMrxB3SFY8Gk4QCzIb3J03S7VKeM0NBCg3oId/
eaqIqxMBwTZK2cmGm0vW6HLfa8zgkefTwrvkfxVb+mLpFRFT2KdVaWGctA0Jfa0OeiZ5KR8IYzxD
bhvXihtUJZDBbV+dMRSNM92BE2JGp34u+gUeGRMUjtFLBwsyglgHQQSGLQJdiQbBbXTXlF4ZK5Rl
Jt7eRdkJb2jQrefhp2f3YayAHOPXb0NtTYr97bReS0Rr7igABYzRHaOsmOgZmYTsIgUxk3Bpzywq
YgSAj+PNpeagen1uvrH21UKIYTtOf/k70Dyqey0giZMz2PfpZmpxk/mXGjnmAZmIEigyVF4Eff+A
px8q2zDcmxsMb3cM8kgKI5maNvombKGdL48lrZASpXnvfWQeW8+Ca6QX2GDgt3J73O3ytmb1YUbf
LV3YFPbfMdJK5kDykz8EdDoMUtCn75i8t3ShFCSK3kWLDRvw6PxCZVxBMK95oSfcRJtl5056XKsH
+NvrYt7bYyV4kTxpsNVcHpYtPOUWONYHZIv2iPkR/9DwMw5djHhI6DLW28xlVa8bt8e69KYQ3OSM
iMy4V74QcOBRsvNN1bZrMFoKOsFFsLVV+4P4enLof8DPAGV4SNaLo5UAL4j/Z1yQl34MC0wI8ORE
Mbwvu6nWTmbODDro6ujRGb1ZgG6+1SiebF6oYR5QcAWaZXx4UQXspiwBptwHiXD0Obmkbi8RWZ2V
zbKApVvfNeVJ+Ax23r9Hg66kUW2IJ85jyWGfATp0y+29wGJVjLVsCq8qCT9LTps3+LHdv28Wt7zH
0AtvWIs8htiaBCJEHgwrytUy2HJYDXILLdTJRsNo9xIQSGC4F67g9h9e3PWTzVwATX9h5unb4HOF
n1kXN2Zys7IvBSO3hgVUwADGIqMkTVtzsMFO43Taebz8UIfnxnjFap37srUIs7cGd9uviZR6xw6G
BQxs1spm/1sczePJ/jOEyk4X1Yt846lQJ3W0h+0xdroseOejXPd7Vx/pR21LpJ9NKdl+omGBvxro
cL+KIhVAAIIL3CiYFshIRfN5RSCewEao6Zg8/B4tA75I8XBrxXwn6NQ6EwZ+ZMUx/uZLKfyEfIqZ
wcu7J9Rgim6JxMSVmF/gZggfeXBlMkbNHft6LvbNaFzYgqm7Cl0H9kDVeFJikxszfgYLsG+9jnnf
sP/aD7IsdxMIIAM9Ou3uDwlQppMoNleP26ccJc4bFdwd/ikgRS2j3cpS4dTrqWfjYWEIvK/jqxgI
pE91VDG9a5fyNnv+Jbt6qgPnJ5onXdlRqr0joivOkgzAYa0B9KAwFMzTSG05yTGH67AnqDB585T/
wapuZH2Hs/p07Sy0Smh/mpSkv4oHtqGAZtTMEJKLS2uzQjMVdneh2Qx7lA67F/T2q+FEpr6JZi69
j57DBYFOGSB1uBwxtLlpQ57LkV/q1KWzO9wXvIWwK32u7KtSWMjnNiwbQcuV1zivg+/sn00A9QBz
j5McVNK+pePmYxLk6ms+5cs9rTwKdOJbqHhDbBENET4fkeqHiqz5USAYWBCsnr0/e6ycmjlrMW8u
jzYHQE8pe/IZ9+vD22J4Gh5auhCe3yS2OPnwcsOIsEL/0WczomiHMgUCHu0HT70vgJlwM2oGzrgG
sNn/gyCWPcUZhXGy9ljGQsBxF/+YxmyDUp7rNdI1bX50crwNy2pbJOW4QSgqvQwHagL4JNyhAOQA
zRnvz2mE4HpVEar5+hffOA4Du25O1H09nsj0fou45GJcYYtgawClaHwDMQmHLWl3+09Vw89Y7GmN
lemat6LDGCGWTNdGJ87mCxXpD5GDUvfZuvvRu1Ojg5y1I2Du6xWIxXvYrNnyTBr9NwUbFctjF9CE
TbRcfym6p4M5nRSOa5FFfzG8TKgrcFqzqupcxfED3tHJ4pzqlprTLWhOcVTbrg9Fqf9pempC0SIc
00cBnvYvgjCiFi7e9UKeNNRM6mNCUTiPGOTDLF3iqHYwEVuAgoAKP76NDJMZ7ThyRDxXbyKt5LMR
Qf4H/zUwAwYtGa60K18SCxumIcZ4DQIP9ojvEV5IHdSJkO/DCZfbOmeYxH6hJwtJGHMBatGfoJ8F
sT2Yh3tcmJa7DC1sY5STWf6FVMn/FStuyVM5y8qAPs2osHn5VFFOuBMfxWu4lGyx4kj4pprwTqdS
7NzB8uVNEMDMVmnzgBMGT1tLuocVZGYAFoi9qszFz1wHQQ5UgGcygQjkQ/qVPvm262uQsJUQ3efM
57lcsDaHRvn5B4lMbXqZS5AyanF9P2O0YxWOM6tuM9Fh766MYBQaJTbRsxxtDX3BvbT5dp2TL8qj
12hVFeN1jGANgJwgWw0++GCRdlFUTPSo5uOYXnnec34xrO7l+ewXavvZZZzK5vBVNUkRO4ywD1Z1
IVn2n1jh6BfmqYDMsMJ3QY6PQMHg7g6MhaMMZLyVNXJLnXxH89cKvQyT8N1Sww+7e/fHgiDJuOGT
QIGUHmd2iY+SOpXDyNn012aMCwfTIJ+cHQZDlFwI+eUeRaensB+fUWvTauWWpe3jqaPDyNwhcl3d
qT1Q5+NI9cUge+n/0h3fCfsrTaQ8po7U100tORHzwyjQd6JtXaMgrMXTHpWorA/1yWKDVGvFCak8
ZXbN5zJo75kq5wQWDBB1IZrXi53irw13E0ulYGrHPRLVQPGV2H9v0hc/RxWeQpWHso5Asj7wtxUD
9IDw5QaIbMlR4VC0wesfVgzaNeYP+SYKZdUy8wgTtI+pUmQkn8D+pfSuC0fm2sY3PIYFMU8+GQ+O
6RRYS1lhmXwHQEi7nqnleJuGTs5CScND92lsmD8XaTqEQWt9vLrYHPHNSgN0CiplRttchdk4LOZk
s8rqxWd7iSxfqiJo+MzQDdKGbii6DSLsY0z4lBpqEYQYuy/wSEnNt8kR8VWaGtQZt+tmaiLKYjeS
PBhDCtWMg/yafdevgZqgQgN1V2g5DjiMDwJbs2wa/HijBA/RsNoxYQjVlmVIGcjw6RadiiEeyWpX
GGie/uSiZWWhGCEQIZYpQvsNtoX6b0xNRXMk/fj0Mf+Izce/9O+Xqy2pN7OlDxJwOBwkxu1wlDTx
4f1KzDqK78f1Lk7ME2hQlv9lksBIENzwdJtMXEV7PAykKU9O0gJzvQKGkvZFJlQHNmp770UWEWm9
8r5SISYUP8yK3DDFQ9CcKWeVs27Ml7SXTAiYCmAtjOsCnXoQ4h+Opf33CVTe0nUgw0wUSPL/wcsf
Col9lRc7GpZsk8SJffsNwkv3k1dU6lWcNus17TkH1TbE1XOWPg3guq7+mEulsUOmlbgjzyCUW1gK
8NrdymfsnKCG4w1wYj7VhN+IIfDbZOuel7x3LPno7AmrJGV/buCqxUzacE4T1ufZXrArkZT9qS3L
pPwARHmhu4e5FEcOD5uj5Re7YBCiFIo8e1YR5EHO6xGxAzpGapudQfzqVnuI0R/bsheQMLWmkczQ
DO5NdKnIHjVUXeI5fOK3kDH1Ph+Uahwlyvz3fj0llQLZFobKlHAk3nAh9eVAw+58nye7nWajBPB5
kjhfZUqy7pH9PS7SHDkOXG5crvlPeS8yvTtHbXXqIARobIitn2+KMhKIJ25bObWBYFri3kF/CuTO
PP5U5opiaGm/Nv6jJU6HCihGJFLUYX0rb6IT9+Q3eY98gtzhcNA+Uga/tajdHNgxOGulDNga8CYp
fW/ZWP/wccoSfCVJ0oFqLCRtnxZrgD+RKR1zvOabUkwO7bMZK0QMwGLfMny0h/PsoKzMvrqzZ9oE
D6YKcQPVYDrlKUXgQJCijaZeR6tEIZ0r+j7i814xxnhvSeol/eoMkzvt4Nzju2kgNxzzGn/+dTBF
9N0RngtGPzt5coKADdxhmN08QpIEJpcH1TsztcNZjnihN/l7dryOpo/LO3xubNE3LvbQdXuaDcxv
oWCixSTNgU8WbeptPQb70ipP8TMT/xHlo3eEKR5fpHnKKEuRRCLWoyl1dkRkXabLmyA/6i0LErpf
pGto2Z5IDYFmOmluL5t1+rLIq8A/XjVKvysX+zi/sfVBeNzamt2HNT0zHh/+2bRGmZBT5kviqXrg
9/h3psuLZC0c+TfLxqN1OTrAa6EB32n52ZX5FNcyUal/RDzLW0AlPSqluH88s92PNJZrTbVC2IcT
eijdktUY9LLdGpOy7KNDiv9q+2yDuHIJlY3/+vw2yHBP9/bd7vLUVmG9oVa8k0+quv/6e201txGq
knL2+Cl9L/TFg08Kw59HRsMzTsZsTGQLVZJcR/JgqwF35rk+dDGtXmjKbAem/oqKoOgSboToURq6
GKEE8PImfh/70TSa9Xg9zKODRDHVmIKgR2SKvUJv5UK5Ys+yA4WzfGcFBIyaWqBWVunG0Ur0TmCq
xye9ZOgDgMb641bqO9dID1VVqqeUjaz/YbJ7ZteLb1pKsZ/+eDMkV6N7ppbZHo2Fmple73I+YEel
4X69rlvgnqzW+EaCII2/Z8x0uvnV3NJa5k38fVdiQVbUtFTgdZEbATgZ5+jA+hMO9TrC+8XJjxlu
VZk6UVEzfI6YOVOZJeRz9/vDedvLCrWcuodSNR5a+DQTmo2PNPGBT8bF8YNm3u5YVi3EteV2gWs7
FQ1aZoI7zMA6V1vO5ivS03cpt19T+aCV7SVh8aQIURidIYrTCJZOMfB6+OBIt95zBT3DVYcto6Qe
U3DHqbF4nUusapnpXQS0Gv6K88CEYakvGV4tfVlD49iwiMa6SahsLY2FvdcuPQ37hUywQWJsFaVK
5sc5aOIOTNayySzWLdbXY40tpjbdORfRul56piaYFo/Rt5R3duMFW/Jm8zZpRzs1tG+FViwqO+fv
wtTSX1aY8kxA8I1PrPVRW5q4aU04n5uD1TJLOBAx/KkXlUIOJP6UKmVaWfPDDk/PZlvDK2xq8tq8
8sAyhWVYALlup6wzZJa0A6NX4aTssROQhYJxOF1QXQLa/7EJTjjOF84WbZcQxe8e6cA12qyuu5+L
S5KCQwNPXc8CVYzntBVVgdkuPh5PL0Ri/DJPRPdZ+npW1MdoEFMB+NSGVHll2TSjSscp2kvVCvRL
DZmLrNn5Q1JLX3t0qcDO9vQCQclUrG6QhkLlpZhvGIubkagKYRfrLFocoa5PQ2lGsGyt+LU4hAEn
/LQYIkQw6mY0pZoMPz5MSjOO5deq7hAsk1D+9yPjLcTACt8e0FyC4nIa/ecbZRT+7/4i/s5tRA4z
E55c+CJYC05VMCZJZTVahivq9dSnWiGRvzL1lywBb8TCajvvf83NXzrrj5H4aDJyfX1VM+L0NyIF
Y+MnbckpYCOsj/G3G/1W9VQ2mkoaGH+XTOeaL42ruyLC8Z5HnfYYVIcGV+ebe5g7M807xMm0g6vy
fxlJwvq5vdWUSfYzCwBbxJNFz5DEB/HuEHNRKn4fit/0kxTM2E461oSarn+nacu1jvxgnS5FbcTA
HXGr6d7ROhZpahH/sdgE96AKU9GzZKXZGCJVOH13zGBiEgMXNRCskQpGNfiVaLy/zpS0KsLtQByt
z7i2kjw9Gy77+Tx71RaWfluxyDiIMBm3qCsz2CgF7mS8GbUsc4OLV2eyQVBgLCtI3PNg2BkZeHDB
UHjJegB6p+Cu+Oi3Ysm1bJEREt4CQr5qn2iv9efBl36ZRAR/7xcZa7K7LU+r94yQfG5MKF7lypPl
TinR+cTb1zdsHN0k1Ypz7CrZG5uGFEf6D/uHsvKWJC5wY3q+x/uzRQt9Qv6NOqeIzVSD1jd0uka7
aDv7lp9E+jFiGod2qBqFwM5GqrbaIQ5yvKXKMWFGwuZg3zeHk47B6N5aFrLMWSGLfHKeTT2qK4vu
rtlTJozdo3wiuDjGRDD5hY04xE2jhYgDBwfi4NvNNbt2pgad8WJAX3JFho4lLQ7eYnph0VVaxx88
FrNxra4UjdMhXuheu9+BnUAGt7uRzI+rJbD8ysOH7RI8Bjn3YOcrhQsGYICCsMdThHBUa04igBkn
k/Iw2Rj9um4sPer36u9aln4YNEgJHB9f5qrkCc7RV7U5TFmDiXMitp6g2Pi0CQIRbiV3t4TCOa8I
bzhCRe4NKYBG0JFFk9kG7B1iVW6SN24+rtD0k1l6O+qlfxFE6Z3Ks53h0MYPGcwikONvpfm4hNyh
E06NAELZiDkgqweuZKmhCXe1mozmenMeRR73L/kGvFUabP7ZOGAUGWw+wSJS4QvYOEzqJl31Pa3y
lE8kDv6cuu8WBgh2Ng/O20QlFogGWlcgUwt+FcLXNNdfWn49zCASjjJTlo4UGsXI6hGxaEqEKDix
EgayNRrfL9nmWmRCg+wSWhOMZgylojrBLJBngMWvIPCrkTjwQKhN5eib1sbYRaGWL2l9uzCiHwgD
cldN8A/J+oLlKZSTIRj/hEKAMLVcPhh7EwUdypXCvzoWQ9Si+jzmvV6RW11Uc/w3NgGXSHCzazzb
1vKJ9Av/bR/WRhfjt/I/skRbUi80zTcORSois5WNyOXNT76h9H5aEyqwQMTHUx+WNZzNxSkyDlTw
r3X0GGjT6r9HB3GXDn+RitCC6VFs2Ho32+YWf72jJsKoe9wevLUhzXJ9I6z/QuX90CqRq8wRbv8N
FBv9FFjtP2KbEdTnwya3kiWVix1JZVTy1kwLxlam9Z6rt9eMODF0gCzYJU/a7O7gMtFVLgoBGIFS
vo+RjeNCFiFGIuxU8x34qYX7eNSu6/UsLpF99/K4n8JLhftMCqLyAv2vbiYUL0hj3De58t51fhcK
7EKsHFRneGeBtVSsxZFnZEu5dsrLYVOzFgwTOeTgScSlUnZ8pohqJXSOGKB0sRbko9DpzimJpDoc
RfGePoP+3gF8DL5iIEv+W9YGPl4MLxAxsEMs6FEaAD+mEfwAMg6aY3PWhJ0upPLdxRJqvzjOnMmH
verYlOz8bbgBov9S/9eFKkBwTAXstZmpNs79WXaKdwShhtZCXor9Pvs5g90j+NL3dvSDrbKEVB59
oEw5bqgvDwyzWwS1SvuGqZ+NsrLtVu+tsV/SboWVZlz3Mm1Dn4MyCiksQmmdKr/p0Z3gm132snCm
UYSScYjEC21Gy8OJdXAxtTT/EbFMa1xoSh6AdxqJPAprSXGEstHE7or7Hh3P1COKOtIiHeDATRe/
k7mRKU7T7dZleT8uz9bT6hMa+zRZmQ9HbVcaFNAXiKzk3eiGv3e5yC0znJFtdmGM/jhtm9fUn1+k
Tm6ALMPrDEVTL6q0P4ueYnVH/W4flH9zfOy6zEmPNV+UjXcU4irBnmhXm0YmZl0BJuIPtGqP7Tna
W2ll2sUw0n2mV87wY0NNvvPn406lmqpm7Ft3pWe87Ctx6A29LCtIG89TUMBqAy2GO7BIFwzfxL1p
zXpTczTgtiWyqTiSZYuyv+6M8o/UHF2Qti4nTsk+sKUFTAtl0UYJ2qJPJUJClAx2OSTgNc3LecXL
208xjS+xIDqUsuPgyB1RAlcPZet26OrWkWRcNjqLRHBUWZkMDhy/PP6moJHafb5CSIlUrDTPlydp
Va1y3ADXtJyjzTOUGtPYLPqF432GOI1Oj5a7bzkv1m0vodMT4XUduZNEeW1eQ2CSzb3TD//U3CjX
lHPqoXMjRqQ9eAYZFwJaaM18isqihGuv5/tKrJy8rVVI8dt6G0imgDBM5s5wXPKz+GTyOwROVyRf
zcyTLSmTFzzrT1zE40jYaiQcfVNgnHoYlbMppnEJVeunNlO9rBeUVmrsKmS7RbvQeUqXEGbHxgtr
Z524dFtYRo1QIN4+UZUoUuLDHKZ4r4/hzCEkpIncPss2EtT49Zi04RRmX/VxjQhBjSzGhUMeuwej
jfb7OYazK8DOtQCoEHuoygHY6HWJR8HFW1tuMxPBLch9D7773xGjCngQQuDcQgLRYkHsjMoLjEHe
NflWyqRzvovdFW/bxeRTOiXuFVvCNrR1iheAhKC1210oyrzT8FRtccVVtoPMFf6w1wugkkoJ2dYm
hVhD+rPkNEy9dyUcUq8JfqOmXGJ7NM6Z//KWKA+FTHfLECULA2XprFo8I+MnyNcnLTFM3f/cZI3Y
BxdZnpAxzPXGFjlJHPsyKKTnUK3mr3Y/RcrXvQQJoyemMz3x8t2W8jWyNPMhq8X2CU4p2/vFhbdA
uod7AGWRWwRd7ccxDQ4w+sipSZGtd7IcdEzmh/d6N/CaIui18pTEzMf1eQvV4lQrxL0lUi0vM8/V
q2zs3nr99BD9DPpH2HVWpLtv/BK8nNTGw4jCK1bELYekQMS1UyKYWfSWVnQE57XGio7dtBH7sXXH
8vGzOJbBlHwwnTLIlnQh/SPibr9aCvhECguw9PP4HUH9guUpp+AJErnrJqae2iLXBHGT4WEdCxIa
9VL5mtRfMqwDX8f0nI+TeKg3XIvc/ZCC0UA4TwefKIVww6xC1+mL9M9sGuUuqRX1te9IDzrMfyVM
8Xx+A3DbBgSE8ClIUyGpgPmibaQx4Kjkj3eF3J/547aWlUTo5IL2vfXD3nSX6Ge1lRZsF2KSkiUb
8dSQGBmgbleX5L46r50B2OA+w2ZojwJMXW50dTPtfCeUGOULCjZz3wxJn/RvxLpmsYhDfD5qFvnz
k8XU38lJ5K42fbiyBnweLdB4Db0mkG6aPcumYGhtheTu8pLNVZwx0C/OmXMVXXF8mZzCzqzISudR
CBWA7k44XyUTvVeAKNyMjdkX05wVHf0BJK80F2a+WWC6eYV3tXZOAop5sVI+nCIsFXC0X7Zk+s7j
jdwGsHP3b83LX4E9hlCYCaJBmPlVqwZqBCjmJMqsNHNrGYHf0HzQz0yR9rIeeX2zI2BzrO8fthiK
XhGa08IYVKennIDSAhsJNbLGqrtCnOdpEr0P93R2CQ/hHqzXimtJefBfY4TSPc5de28Z7tgjcpR3
JgIna1tHhxG3/++6yLKloVK05YtV9oEO2qaHhFOSbmrEN21uUuPrsGjs03lf7bajbboq3Gtvd7Zo
DW/Jtge05ORYqYzMO5PgDck1Tzif5rSte4xcykBxHSFHo8K4E47ZeioHkscXboEpLgy26V7bzJqL
/QEgivTIGuQvNvnQfjUEfICZ8EsVM6RICeK2ztTk1UdFhepqG2vREZGh96fvB+6+dONyEz4glrN0
4n6NyIxHKjtVg0IvKq+C/LGWBORD5XBM5aAkWQGayu2x/YWSz0s2b++hJQAGvf/j+66R5+gQTewx
ix4/yQxfbFkZUbds4uPDg3VmC8VQhmlKZ7N5QqKGEKRnwjvoPc3SSv+ZsJ/YWsE6hG1dLU/btwVu
itN1WGEeEUxniTpps27BSUPbIqUrX+olpcAy971vrRCw1vymS6VZ4Wxac8yCcd6u+11EO3e8NITz
jD4Ab36tzRtUhqoK2hoU5DaAg9NLpAp0dOOTZqWfh0+zj5drJjaDqf6UBiqvlJdLmVeR7l3AVIbZ
MGXp4eKh3RqG+A5DsHvq2P9POsF3UilLTuBxulty6+C/LTnXa4dfNbNZ70ggRfcevjTKSKHHz+Fm
4+SQzRGH8W3uxRboLBCl7xJmwEwIFd50b1NtDMs5Qop3161oVJ1yWw208pfkUmwSZPuuywxolq/X
wSohk9L4IN/cZzbnsL4n9FiydGn9qS3w1QRFWpjJhvcnqakzLpquyMTVfvqmSbD1x+NxtAewy4vd
oNq57yZw/nS/z/SiWx4o0t06pCwO/k6lNDSsKHfsOBbu/k9QJBwfcsVV9nJ/RJfCgE4kFJt0Pufb
HrL9NmyI3QtKTCLzNHBtW1yUFzTa1cNpczTEy9nWH6ImQngzGUo+xZ6UM6HaU+sw9NgHD6k+ywHZ
8m3YAth6/ClZn1nw5KeAMAEwVSG6OTQIeTiBEk2n52i4jlxizFw9wOjciJKaSu4wJES5Xmtane4I
sw8l0whh3SV4Rb7casEL0Nm5/T39OC9m6CG0Ce265Vj4cYPypBW7a9o8DhfZYw6eKE9weSalThvA
axaMmkzIGFl6817DHRey5DWAM5/5s6jPRiJp9aEuc8El7GpyP3MOuMfEpJQouAgsxpUoAOac5AN5
+f95tDzcM2vNDte5tMfwWIjbYh3K24bqzsDiSZIkXcmkBmeFNbp7cPNFveQf4Mm+ipFx93EiwdFF
5lK3o2BWCepGuXi747RDigZGAq6tcPBDmHrbL3p0rfwZgtAFZjo3P+AkUw/yYkHMAoY5bEGBmU+c
bt24YoVTrnBIKfgo2UWHO4zl+XzDPUVZU1WyVYUGGBScwCqNCLx1V+zvWjQr4fW42oemeEKxmyFO
FXAnTSMHsMeTPfBroMYu95FI64We5d6X6OViX+F1w9UEj+xZT9tpkakh1d+i1MKQhKnTdHTGgz9N
fz5V4QVuWBWOksGkPkzvoXSTxDqPLRSZxYcLBAQgZf6yWbIDfmJafBiWG6YgWKRuN4ug+cW5TFrZ
VllvbcPKi0ZZ+vU84FW9O3y+SujIn1mTUQzEpu1X62pfwpNR42mAUwqnVY1vnRoMb9YmR/E/Nvmr
v15au2j0DzDb/qEdQwGaq7ViKU/QiZ6nGpYuq+Ptwp834oKDwQrYRmetUGEvb4MAMYNZHxdQWF5n
OOsWsOOEiHC2SIRFzW0P4AapMUsMIDDqHGwsIk1wLou3eQJZX7ZxmwLT0PUko6TFN/RRGHAJ31K9
k9ZbRfpBbktTyCx9pAWUbAyDxxzyFSNiJK4Z+Zei4h36PIexd2MnulgApJUEtgy5mpcT4zVSA/I9
l5tR5Rxp7mvOOzh4HpOvtvHDsHEcJfV4U+yVbNmZGk15Bblicvs/WCwLbUee4V+QUFAhlmoxaTVv
s6XCqad38CURQExteo2uJ1tszPHbt4bsj3FvOmiA15sHGqD51EPF9R9Lvu29IUeTzRZFK/LPv9ZS
cAJ+1y1yjzp+Cr2cbC9ek4UhRM06QLZvzyGlc8FVm1zh6gJZsQgWE7aeqUBVDtzoh8DaGOp2N/xW
lascccEe3vTebHfKkw46rT/9T3M2PANTu8LK9/nKrqq7YTWFsZHBriMSoFicpsSu23bEdg+glqyy
xE9ktHb9qfsbOU4JNCJwa/X9y9/VdJDNIsAM8zxVgnnzydIhe4GyEDxD5qiuhCVeNcsUeYBL1p+9
ka0Cuk/A1xYUfbuax0vlniIezeBbhOkMvzQ/ebaBjFiOG+ts9pEYpY08zpBkWQj7k6ToIqKCPsK+
gzFk7/E5B9qGvcy3Sjp2eKOZmgWvPglzqfU9RVjpcAkmdBKZ9qIl/aSS6aHf3CelrbVdOLEoFpkk
Gm/CVyq/SfmUET9pSeyHPZazegMUdEeUdsF1vCiM4prMmB/us/q6s/OPeioqUu2nbJYQypuhTkoF
L2TLSy6iD55KeTVbiPVjLyt2HfGQdrTcANpSrsODXQegSp0xg0T4ru6ysNAIvFeV4IKmR3scT0Ox
r8T1kQh0RnSJI5sRbTypx5gJSytCLI/y6TXYizauClGg62g98zg0sVKioo5Jskn28U9p8Y0BrrEF
aVN7s3Vfi82HsDMizT+5Jv8+6x7DevgIupyOuwveC9nRx/E0ZfNMMHw7Kar4vVpsL558Byo3qmGV
9tzVjHd4SDS09vi2+KWJr4t4IqHpD/mEujN/sgIiPBQf8ycWkUZzU/h8jr0QpRfoG2s5qS3v/4G0
ifpyGYLn6nxt0NraC0nh961dYRw+EgPBRQiZukd5EL5IgVQvqcbgguAFAXscxkGKp8HKVabiWMs7
JbAXspuiNXbib6FSAczIWcMPNy1+dec6HuKN4t8jUtJ4g+z7JzpzBPW/2VjztBhe4LntRnp4JDWe
E0wqhHBoBqOyLZFDqplKfaQiMgeCOpkBH+sb2TtB+LhBy3Y7CoZV9wjjddITR2ZZ56xVHjwBuD47
eDXBJ0TWRARGwOC+/mK2R2gmBRfwx1i6MMzxozPVjR0wYS6TYcyDQWBmeH+pVGbBLUFsqtfANKlP
dwONW/tNDPnuB/C8j+7ytfqsOYvCsITrOdj9seZJJnD/gIkvRvDm43CfQShjuG1Wkz4zKMPrMUdJ
BEPsYRVfQKT9ICxOymi4f2PJLKTEGAUmf9Z9K/FZdN/Kar/gXKFdP9tz2vyHDzHKnwr6a5PZo3bh
V+vZllQA4ouabQ+VdBCxKoCwC2W5Z3i2snfqO61BSbbKQgWbvb3m71P0h7uC9YA8XnhUande2Otf
7s2ZquoLlLd2j/MGHoq8J5AobX0KnBLkJNdH8oqJL3kExJnS0EvmdO4EVRu9o3rFus/4dFHBcHdc
vf5frPY8PgGCswms2UcsDirkCqPclVTtGwTmYDHt9Fwdqi4BWk1uUAntz57e9B36kdT0FiPoJxhk
dvsh7k+o/Eau+TOxufoXlO+z+E+3TtDFJLkH50Fv0i7+D29U8Bwbl4f2xMFPEni3gnWtuyhnzaHK
omR/fhtvqVvLj4p8h13Ef3wIj4FxOURYeVzk2zI8WskTzB26CCET9G+5x8yuJN7RNWj+AMVz6j8P
i1Pdlc6TJWpBXCjXWu/VjHGOd4VdinM5IbNHvsEx8uEBY2LFCvCDSRzhK6JP6tIOP1keyD0WWIIH
0GTGT5vTzEi7mUwQAHwWgO0Xh1D52C4WO0rkN+p6MrKEfLbRV3k/EEKL9z8T8SfS+tIU58OecxWU
v6dUMnc+dOitdBYqQJfkTU7otW25j9XviLXEdFgzcK3aamBPQmUxiP3yg0qOQJ6k0HwQ0mXOKMle
O7bV//pILN11eJ17/O9m8I9gnhq2yakxG9zqUxBbzd9yWDqrafZclXs5jSf8hVn+wOINKeYXxdn9
IhFucB4rz3Dkod6KNtmBUCD//n+mf4lRR7hxWZpDpUaOXmkWUzwlMnAcjuQtvNdvioAZ5GTW+NVy
GEshb2CwXi1jrCTUQiCWMn0WU3E4kvich6MBNOICSGzsVnp+cXUNDVXbhdXmoXqEL6fzCRBnNtWU
3lo06xVVpF9jrxAyBOgxEkbL1Z6Fltr9xD7cmBtnunAGPB/C9rxwOx9AMZBPFR/sY/dQSjnQqLNl
6Fkx0qWHHblsnHCEJYdNirnbN8TANkqwzuliHwsrv+YPBb2q5O10BAyxaS052EfndaVRRHZizXVI
dFOq0KB+zKVu2au7oHpAuWYJBQ8Y4YUQVeTahzqtAlK4RAkL+KbTVROvkxficX3z14vb0pbZiF6r
HqMF73LTFPdEhN1Wm2J8s6pMt/HIQVsx2y8QHXGNOKPXJAAl+dJ5ViwM8Ztz/1nckfG2/oEVUujL
hiLOJDzu7ileESmzOagDqQDLQlLCB1QmyoZxZK9E6tnurXvQW4wFf+TI79TNMU9J4TsK7ktM/blP
RBAczAbjOCExLeTa95Mb3RPjDCqX0DFjwwiHSv/s9ptsWQTrW27SNbEh/k7UWjvlMohDiecahR41
lwmhuMVF4ExotBtPmgTTOUDYEu598pZs3iNNzKAsQzcmJ0ljFHj4gIrMbfaFHQ6MZrQ6UrQy4gmj
fuSVzAfI63rBDOiV7xOR1+nVwa1lkwvw/R2pEtxd4wzTjqzlfOESHDLetLlsDGywURkOXO3bcrO2
c8U6F88ENPJxjHepH2g2C0BjsFkct70yl+9ThvhkZc0/34SLqG0vwLKmCqesCbEjBly5pNgw8i0q
JqhjVtjbnM8W7SN5v6OSl/3MAGWHPSEizqkeA94KuwmgqvpudRVYmJ8XW5MG/ftjJEb6+ryg5QL8
nUkjkoP8W9ndYuqkwdE/vnhoSlS+xGbX2FcDQZm3PS9fcGNNJcfAqBacFpL0HL+C7Y07YoAcvFL2
kf89X4Pl6eqKrDA9IKyv6sabuPzEjwg9SJzsNE/h1vLsfKHQ37d/fnCWGlkAGhp+IoFM0GnwSLDG
PO96zzbQQDhMOYJQtTQ1fpGBb28R3F8peHOTxu6+ihZoqnrZ8YnfjlRid6FR8PUQqfijEisR5VYz
eNDyZkez0vNST4yuPIX5Un2avu9ajCOAnQAYwjiTgjPqGzR0816i0pp9QbRYsxQpHK7kimOQ1qkS
3JTTRBHp+N4zBFzJkjXIMlrNuL8Ar4o1++qdOSSyE8Vpjr0qZ/KwARVlOplQXCPBQaJ4BNg+gOPj
fHeQ+lNSS3BCUDvFyqqvUzy0YvyEKTDeJspY9XYBdpLjPnauRCdkef6SXhmyFWNsg7lXkbfUAOr9
EpdJlMLskNRR6Vjz0vSFPiPEXt0sswxDJE1fux5IUbKqUJSItr+//NvGYqZhrS8yhQbJtpdi6Q1I
JUbAOUSpeVhSwnLZZobD+c/ncD7D6sMK/ondpVNTSb3oxYqFafD4v1bsvv130SYYGVjHsgRyD7wg
pHm/jgh7LgZg85nvl6p83ivxJ/0fbnGilakqq0VN4cp3qXBj3eW3EUZJ5DAY/3XcM9fpSD3QIdAb
Kzaiowu/BfMhrieHqo38t1Al+yPXJLP40A0/rLebFnA3hJ9LN0eYQmYGGR/F92r02He/WDPxxydT
uMbyCI/gs9Po7VpZYEZsqGKHuqGo9n84epFhI2367X+0jreTKJO2LUr03FAsW/rolTDarV5P9bps
PfFsD151rnNXPF3issNDXRwkHpEvfZHNc+8AIye/eEg5/ShS8BQBJ9E/LDRTtEyCLUY2xQX0e0bq
cJYdFRxkvbdjlbby274TjdGHLNBTRc5swv3LH8Rcq3KuDA+JX/Sz6I3PgKcYm0zfr0n+k5/hcM7w
6PPGPje7N3Th/ZUYc0CVeKhP+W4S5abgHx5T2Sw9gi2JKJsIvLMfgqbIJn1g2fCkw0sgnV+u+wIM
z8LBhLO1hjVnGoidmzqHFOIlclBBEfTrAMwcUriX9zzy+jd7jmrNdeQ7NWH48bU5qRlDOx5Ro8e+
q+kPsvzYZ9tHa79nUpa2BOwbKLbzhr6d5h3gD9yLRh/gdBL8j3DUgJxii9QUTuQLTw5N4Dn65iKZ
M3woywX0KBmgCAd7l3qaDc52eU5x57eZJCV/wG8OCWJxMhgTPKde9v2bRaMnTpHSWIyDH7jxZLNF
uxwDfDHBQsDnysrKUlOOTrED3HUFGKG+ysgbQqyeydW1WzKWhWkxWwcWuEt2XS07mLfzbSEqZesD
/baVQi+cuYQ/5IoAjgBi/y/UVxTFvjw5G3SDiH4tuKQ6QEaQas/3Ezq14RR+kwvSXE6bA34CKFPv
vmfaEyVbpB97VM3o53RvWp+fb0S5aWKFXH6wfgWqA4kubQ46M3BxmE6R622xblTtmS8/2r27JvGY
zMjiZMyBPAWt93tZZ597DvWQHvdaXRej/kWRNv9q3SY6WqNmXWKUqeEeNdnk1oqv1axJoaMxuHk5
tktWPQatNJgsWbmbn6lzNslknQJhvbixU2aicwwZTp7JCigR16uU99WpKVzBAuL0U1gFu9Wnu4vh
RNxRN+E9gDXTmBLkxFewTZzoeGko6J/Iv+Ee5/4m7vbLVmhms2z9G2lcsY20oYYy7AlWgOyNbLat
cNAPEHqroFIikPG/Z81fc+veOfYdMoIQhGMrBJi1jZZKSuaxMyrSh42mihKsaFsoUscm3wGHMlkB
MdXWYHFLgOc7GFY8LssaKc61QDVdU+vf0ryS+OjdPSUR0vu87+vcTgeF9ICt038TJtuR3MMcd1d8
lDGjb+ZowTME0AbTiF+DUlmWZ5Nh5Pqn+IDuiQTgvOXy7iJxOMmUjKyr8/Tv4y1PYjsSVjjh0SAe
BuNixnB0nBpUtNZ+i9L9plP0jNBfnISUeu+XL/2jxGEDFyxD48Cp/BowMLrDK1lceKoLAX4sWrKv
EdQfEmMZG8I95+jjt7qvtuQNGOlTN/mVq1XGmxJam2Ok80SyKAtlxkkBiLsY6jFnXIJhw4kjlJpG
xJKl6MHVlnIWmICFIcj4dPxUZbARzu2i5cIlWyADmoC9bqRKbCwmHBnP/rxYYkNif/MP9BP+lYB+
RafXIK8JA0N5ufcxNmyaeruAhpFsyDSAtOSjPqAcIXNpjF/yyXAleip+jlSWIbdiGdTe7ZKN59rV
H2DyKryzbzZz3Obx6XYwQ1hniZ1EVB9Bukl39MtSU84oUztB3V01NeJ3+9c6+dSn2dmLsoKXSmrI
gB4QhBLGbJvPO/p30+IZHYHBMzScgiLkieJZ2OiH6Ddz//eY6BHgfkXhYKKNMwN7KKo7H5D1sP0N
4TsAUztonLUK/Z0a8QPIzs4eBywjtnw9niM0jog8W42oCGDXZnDHPCRavpK7rc0EVv1iyXc427w3
JeqxGDZ5ryWQNnVnjAuZbvC96HJeMfe4FzdvS/xD/nwL7e64jdE3yi9YW6L9nRiD3IZS0as2+39q
CEgZ57zZnNtpCH6IGK83e8rkeXEws2LhLHEpvHp+xHoVpwHMNE5TvHOiyVLjgs+jBziglaLE4LjA
lZ7xduzGwMDXev/Hu846zTx6r75jDz6dioQvWxaBzNaK1zbrJVeOBDmMARbkNX2luLu/VS8tQoeO
RmNzSfPWmjdDqE65vFRZzX31KIIIBCjdauSNeQgJ3IYwFmO3pybERVMhAEJrtAYvyJk65rhvf5Iu
dbk1J/biWTMWLm9veWnUCxcb3Ae9U8oiZ7u1JISK45N7RLy8WcafgmkdqFHoOMsE1TFuW/vmimUr
NDqIBoZhHlBmW1D4yWeiDTZOyBmCW6ffkEEG3Fo2drD42IvzzQn+sU+ef6rfRPFSXhEBKKMLaepd
WXhFld9Faq5sPlu0uYjy4g09keFg276uCw0ymgA35mzcZ6ouFDsJJstcbZVR5sl72jxrZ0qe+FCN
gH0PN3v2wmkSAFZ76bf91MKccMYQ/JGy9H5wS/BkWXzG7yS0/8L5+n0ka2AaUM3Pqv0hiKt/V00h
OBsHsyndSEhbNmW7TETvyfGXeyrUyuB+yNH1GAslc7dGe26ARJ7u6zY11GG3AuwMb+HoTHn/6beW
UlR5ElD9cTefbj73fNY3uUh0QNsFmIxSdrz3MmTMT1FjjTy4Gis76VjrCilDfYMPOw+khhSKYe2j
eHGB3lrqekcn7Ha2HE6Ml/Ndv0c+2THezh9FRoEEPD7vJPf70NBYy5gpqedYyUfoNSQ0VqE0Hm5q
eiPHb+sTwba3bZpviOon3g2wmlb9x+HFy1i1pCJIBGgGhZ3qVJd9WcAY9QSACJMvJnGOZbD9NDkz
hPeuXjwLqBmeROvsQQHVScI3AEdMhk1UKFhA/tIJ1XGWbQ8NSyf5GgWHDK6epEKz+Sxx0XIoCloL
ZCOb+dM3v6ViqDfN/PRH/dy7ok/NE3fuIht7emAczDdkKM4DbKnRn+lSzNrOB9PdC+dVxuXF4aMg
80xy8og6+84/5LTDpkxHhos7PSErLqxxolzAP3wSFbwKur+FbPvUucCApWmnxFOTvbpXYWBHUJfP
yjKvvuIQIBbe/l7bb6Mdegu8hBWBtEOW8FixP6j88dmWB3B4GPfutSsIvhFFmgxj2pXMRp5SBdfj
xsyogOE1MWuQYYEEjwGqX1d2R8bqHgtz8cIq1P9KWBwSxIIgLKWMF6kGejFVhjOlvcfMOo8PyXgX
nMYW1H8lyP5u6mO1GYvoYsA3nwLn6EIIxP0sw0QwtARWBXRwFyyknFeof2My1F2aUtHat6SUylw4
JeUf5z4+rN1I5alH8car5G8X8tNkj3Rpe2dndsjFmVuOQ1Av2krortNqi2Z0W3xxs1wUKJw+atzL
WMiyG6zOYeaY98ekPc30022eo65SmKHF6ReoMlx4ry2EnIgH5cougxcCazfes6DgjVkl5FnTR4bk
Cqea+zIn2CvYCqL9ibQsRHKUEjiq8fTLhrVmYM/QC0OlTveBDve5ABU0Nzx0FYCxrr7bB6juLfcv
lwNU5Z0aTc+tq0G4Roibb2r1PjOIgPVpL9Dm+HbrzuKL7TO9lwrilF2JsExVadtee4w7UbCz20bl
iQtZD+Ae8aELXxoB3212hDXrvwamE3TT/gAspESJyP/NDNHFMzgpuTHnVBkhp3F5aD7pDe5tpP+d
VGO4yc0+9Gt3Ohz5ZJVPLa5/uXZb1giEekBu9iuMkEXw/lvKnVFg5QYYCNiZLHYGLJkpSVvpTbYI
jn7WKa7dXXPYyTyJ348F1+cdFs/2kWlm99lBOlonPnhPlilTT0f9m5ZAljus6L72HUuonvld2ZPO
V9bRx+l6Ohljbg2mHlpwW+UUPrLBGMIkPHRPM3AXxNNYdjxPSP/bcXi9EL0WqNITW6a+JAVrQGPz
WL4mc5Xb0tAywwYWKCUg9CvHbbNMhb6hk9BdY0X9+XAIE7YoU5JxCmJri4Xhd3/HUvFtaiabISFa
p1XXMN+0R1pupQdhpHsSeR2PtemVN8Iss93neJHhery5CWdiXKrYq5gFEL2RCnncHEd4Bw9ZIH+/
woeHOD4ZVGQCO9pX6K79e199cmqnbYRXUqN+aVu7Nny4WyLccajGk7vAE+CxrxsKdJUkM9OVtT9n
E6AnqT0HTgtXHgXKs/d0py+JO6RH8anX7RbHeXdolBir00Oq9aMwA0TMy+vW9PQbJ3XYOG4OOhsn
aEAs39PdOXUYy51isDlwsIwQDiRV+XdaQHAVGRNvVeZTib93bz/+OeDMX5HcN8Vupp7N21eiKrco
QvJSL0WEK0jz5lePGParlf7ceDlEq8rIewrZ/IJacffqWxe1+Ai4tAyNkyPwCndgd9xXfa0Qq3aV
YiJnVSV6hMOuB/7WVV2/vIv1oGJq2+rx+u9q8adE08FfExP6rWa1ormAYDbw5SVBY74sel9/56ib
oytJoWc4RJ6Cnv3gq/npWCBNhWly+/lMjdX77HF1M+onUSL7sSFNI7TRU/vcQkUtwspmzeXPTKJ7
MKhV6SU5L3iy5i8ue4Y86J3zwufs+4vqdrtkolYfJDejj4TOsbv7qARwFTv59aEJftMYnJkV4XAI
VSdOGEwES//lBe3wiQJdw1CIR7ncL8w/ylIR9ZyzgkDSB2t5NX3uRu4wFJTwnOS4oGSLK+jOU8dp
WskMMkipVQA+hxMpYQALNQZ5XX4DMYbiWZr2g18XHx4ihHj+ocW5BC+XelBoPdS7SLOy7eGsUBve
26b3V6qr4fVOmeL8E58vLjSCo9zpfMEeI/7w5RhNFXEkPEyULueJFKQzStdNHzV1ysS77BT4TK+E
BSdd0KglMN5U+5KbdAdlsXqWjVwBq+RZDnvZE7nWv9mMwUCnp+Re181vNnforvC+zhPCNqNftmi6
5vyqF/HEwuUZBa5SRJLfs01GVkILQQ5UysedQE+FiDfxK9QJWZ8Bn3Yvs1ZY1+oFRHcb/xf5XEGL
p65de/ToP5lBShuAta33MHr1s4YZpdkfz3vadPyqnjR7ShRQFlaCwGUNj3Y3BVx59F44ezwoXFaL
VUxjetwmjmS7CfHFwXpGwG3I9woSJawlyUj7cI9gyzEjEOiPN1SWOyjVwMZYHZS1dJw9q0YCSq17
nBonumZQOi8mB+mDHhoFc6t5PWPJylSCZWL1N67j6AXnEG+rN8/o58D6GeUoxRO4WI+Brv2WBgEU
CJMphmA+fOBAf2zMjN+gchj8/YR2Iq4JBKbBPqxlgm1QfankwvVuMqP0BuI7Vk6l6jrfj9q9Jtkw
U5oPaLEe0syVj2HCtK5P2jZ4RwK/FpFlL+NGGe3ScM1evbPSBNgBg9H9/waJj5ePIOaWqd3wi4+N
RoRv7N4DXHqaZhFPFlgcudEn5S/YNCTWVex/qJenfQ+4l/SaoIa2sBIHWbZkFgZSHQ6oY6NXN6h5
7dlpc4so4VLadsSnkvnbVcxplizsBNE1i816pTy3muepcFzaaBJrM4o3hhbjQjX9cw32X+21CcPW
5wSNR+NeyhhZdZHSoAwhBh5jjCF00Avn/FcJMjd0rCYDtbB3EAy4PXHHQ7kpPKis5L+C+6XFEsQV
6l+aXARfMmtg6JzMBBnSGCX2dFL5RIz/vC3WXvvBvZu+VM0dctF7OEm3vLqGhyvKzRxGZ75ON3Dt
4ckiiw2jukw0YLu6ATmvneEGkWuBjhjAUMe1eBZ37Qvx1u8nCGu2E4Aanz/NizxuJb0rok3DdkoF
P+B1CDiVt84cIet8eFuNk0b4tlqkEa6vxpEaCWXPbz9HfAijoiTuXTc5M6VI08hPYdYULNQSWEPM
e9A9OqJ37n0vfQ74f1svi0OyqBR/5EawbYqIR0hNcCYIFQdc33iv3gsLBs3NA0Vsu+QGeTx1FpCi
XuUQBqBndP6f/PEMCXdGE5PvlJUX78j14zahub/fKfsE9ysrSzkaCZ8aXlY2Hm9b8aX088GrSdWt
VB8NaqY5kEQrrp0S8WbGQApOK9aefKRZwTRQ6mTIC2UtYDZFSC4mU+V3U8lYUTDYdgBBcX64J8DW
9ZPpdPxrxjvT8uAL5dqC8f/tfkJ5yXMpKfFStudeDtE/znWuqIhRuIgoIooy6XHuOMBGUVXWR6oh
LCz7R6gke8sfxo5ugVfGnb1hwFsCb/aooPsaqwQPbHhE0YfJHDtBvpZ4/IpwPYHYdyodSzTmM5dw
RJ7M2HHKevr4t5naozil0vRWOxQFMSGikl0yg7PhwPhHoOs96k8TmAEJaBdTq/K72BiCXm9dKLVM
ke+j9NmD5JqK0EzGhZW0V70O5rRTSqKVuQbBATUEufwdiApm0P/wupAYhsnJ9qFImyV5L9UU/Ra2
vhQYbZdQRoybvocyDspLJl2K17wX7VxcuWoR+6Od31dprjvPfuZuXdRhDVXIKsfixzuLStgreFNL
tBP4Nm1G5dbz1uj3pqRIUihsnRgQE6qzbAB4iRVbIURBZ25qahvff/qgG0zKOAutaeb4OOewEyAd
ygJUJr2j3LO1TXQwyni9RySTOIBXK2ikvo5/jo9knHFGNflmsQuypT4y/Gt4W8qO/BYDWO5AAqUS
xbX5C/q64Ci1n4Dfl1p1CuE7LjUOR/Bw9PCCyC3lH2KafbYvyGlXymUbGTkulBBSSoWHfj1WMih+
iJBj6HtH3bTo9f1f7PTdyMykQjXIyQi0hNuretvrGEmOYrE0phXmmYj5EfeoFPvWjK5+eq689qUy
jbJd0J05EL8rZwN6Hw/WDiNw75E9HS/DNInH5W10OofAMgPv+aTVqloKWhlbjpE4JlDQAg+oZeZu
p0pxUSHaMnmjDUhJg1MhloQcWUBeKHFiz140r/aqXhEcf7GeSQ10hk5u8iHzSSxaBFe51mI0Sor7
q2SV2xnIC4qIPCU4+LdT5dHo61/hlpeyBOz0HGbKlPZqnpXw7ITeDC4/VaHUdd8WVeunsrKqdcdQ
GxlnxQQZn/kzDWTARbLS49z3qUlUVFuxkRaVQQPSEwnyw/bu2ame/zmhfjUBs2FVczvEkT5WE9y/
HJ+ADvTCEE6C5gw88xhgn1aVCpZqBbdh6pio3DPBKMPlUHNfR5+sQFJCw/goi2X1DiyJiskTMzNS
B8NbyFYWKQjef8QCMjnsl3iWZ09gFlWRgbWtS9DHFtWX0XvEPrGp2yjxfujMwGS43vRgTZXO0MFO
bEcNZw2zcZ7zkicCnOepF7k1GQqivrXG6YwqQ6Rt3zDsQ7qFe7N4GCMoau76An4kp9LN/wjcNX7X
tBkp7k5wBG66zglYokVIaPs4XSm0kXkkgQ9FEClmE2F8KCaqrIVv6COXy3u2phPYTGG+EhYytNoj
OvTSLW1T9LfuwLhkspirYmTqsWWhfoQ24KuSULO1quns0d5wa2k/FbZw4Tl37oPk1sgCV9ZzOvW3
21xfMw3+CLz5DuGCRKe1D1udgXR189vZo9eXOCtetQiKYCYBd9y8GBnHlmow5MbaxF7jO4hVDS6t
9DLjekDSNjIivq7xtPJO4ur0DLkUDiurslh1JHSzqpGuqDqRfF+9VVow73d+9NBI7DGezY6o2G7X
OLaJk5+lWceeYm0JPKXmwJjf+gQmsrq9m0AbU3y47w1wRGvduZz1j+EFBqjOZrhp91rBlOyqmeDj
vfxkeblPEFZu9iBKbexIrCHib92cf2322WAlHbg4Ba24PN9X867YsmhgOBagC90IiP+lMt5nESDa
jQvSzVbbPPGqripOylXZmsvEN/VqZMt0pOqGihL4U6X51sZo2RrFdLXQMTnOrDNi0c8GAJKt1/l0
wKOcYhLGMQKjBKvF4RZ3BHK83URPx+UrjfNZs8G/LbfToD44ixRvHdQJWvPm4JBCQhjbS6B78W00
KHis+KLCyrhdOVpJe+/FynmggqF9zSt7o9DhEsOarkTtjBtYVF3yJ9dF08XC4dX/+DjwofJws5+8
AibzyffeYHMCejVsGTdlNhUVsFTHnEwD6FAcIEXb+7k4LAceCIbFN3BYK39uaHTkNu+8j23Kes96
moCRkBQOMBTOM3liXmQM56n0/wdzNj9bepl+CtgBWrApXA6/PxQcZE8l0OHIC4JLGVN88DAh4ham
PAbLnrn3JUZmxicHhrwp2Zzpp4Z/wG5z1Bh3DSp7kQdhJP4Zng/kzHPS8Yvbcuga4FJGVMnuAhRJ
XgaZVdoV2hjTNthikvhtJ5ht4RBMLS7t7dua5swpAU0oP8SsX4gyjXVjKOGfKxv0QJetRMyBNPzS
zP9ckufTZ3We/jSFiUVdjm6tVtVoirroyY+78/AfZMz2zUQMnqveSSo7T1TJy4ggtgsZCeEagbkF
k7qQXJBC/bdNDMlFrqbJjpw9gEYwtqlLl9ySdtRkVuSpRI/o21Y9maxUlQC191CpcmK0JCb6qTqY
B0ThVC8T+GMAme62lJIamZDmxzrx07+Riw9p4GQf9gOtpSo9pZAoU5kp2xdn6FDynFxSekzvN86B
s1MWvVR29bIwOSgPF0IkOE6IxveORTo4qhR3CG/b5NJIOq1cfN9x6PQ1VICT1nqZ1HiXIXn9sBq7
BWaQgGz7/ERgP4VROq5jwgQJnB6xF9NUpzr7e/vXRdQ5PI714d5en1QBhNXsBvWwsCC+f/tAMSzy
EfdTpUkaSn9IvKlExULZmt2Pyo8XQxKcXavFXNhsNXJQgX3+A3wRvk4YqJazrb/T1OHvVsrx1yhq
+OdHrILi5yyxchIn5JtdGMVysMERo4AER5yzFVmWElnEvyZJ8RqiFyLX6In8/G47sExBo4J5u17q
ePsxRZOAxksVWaBA/pwD/x1sHLCEdW8OzZynaUf+Ml7FdH3Pej5j6S+OQf1/arbhVxUqtT4dpUhO
DX5dszh4/0fivyBHqVvpTIf/smqNobR4aI619srBH7sJJf1hdJ2j/5YmMlk9lefMMeO3k4jig+6x
+/B+ih+cNwnqp95y9aP/Qlj7Fbt1Qi1yn7c982N7vNTHUI8KwkwCwB2k7Pb2YAvJCgVH4tqnSn0J
ljnZYpLfrNQCY4I1iz/8y/XIE6AGbjA5dfv0lBrtGopPKisY6TfxX1o15qycp0QHnqNwJjuHRV2J
m2G24srZGUCRyBsANpvp+s91wtt3UR/1DGB15fyqKY0RDHqWUq2m4gIj9yNwyxlfchCpcBcM1W0d
Io3oLD5A6c3sHekjJmRri7eB2VI6SihFSKyeTF8e0+CuJOfWjrZZPvE06uE2sf39lTd4Eahl6cP0
hVjj7EBISxQUcbOuT784b//pJBxnh5Olff8Dv1IdhCObvJffOM4DBcNWnh7itFie+Iw7mXKQG7js
RVkLBhAFo81l6hjww+anNybfI9cRjsIiKdsBeFRDhmieSQ+843JPOvDS7dxv4jRNjCtrewwIsdDh
RC7mRSKtCHPH1nsBuXZJ/J25zfrXemmbeGzPf82H4qkyjD5vOkj0+u/gXbqzTgV/xQzB5eKNy1UM
LDPRpmPVGDLu0Zv6B9lWyxSshDVhKcH56qBjJ89pCUsqCrUbhkdE1t9BC7dqHxRgqSQBXUK2lvhJ
i5CtjqJoW7kruJLs8bl/RXROCggeR/toZrhrTaCiKiythIOmW4nuGNr8VmVLOgFtfVjcvQXuX++6
brsL6U5smXpIm7cqsBUiUVYfx7slHTu7DRT6yq2489Q/L0fSDbBEs6f8AkZVw65PhXUGu5czOdMt
o66t+IxEXIx6DIZhd5JQuAGV9inPzofu8YCWlLgVbak1XbZIWZMWuy1yaZnGEyrYbkAa071XW+Cs
1tWQnA62XWXt6SWTzEg7CLw6C6iaMcTmJvRZrBfujKzdgWBBYWJsExoctHwVrBpzODHxJjmTQECy
wt1anIGjNJlXQlCt0/3vuDJa7H2eRmAvzPLEteTog/xg2zz+dB8Iq31tRZ9kWrk0ryCiYZltyWUD
rOix1nSx90bZFeNFUyt6zFZvC4afwcZd7xZl9igjwa6AOG2qezu8UG8FHaLRAkRV9e1V5JR0oTdI
ZotheZ1C4hJfG5nHDK7l8PQgO+0juRgUm9bfYLnn78cWBj6d8hxTqxrDkBZXkMuWFD9noDJRPSOY
wGhQIoDzfNkyDVA9qkbkTTTB181GyVUlxjT7/VmqYTS79ZSujwOfGTyDErBWMTCKf9ZMq0GRAR1c
a9NXsZisic6JujVfISKWXgVymqRyW4aMoYHg6hN5qCHOAE7Cd4d72divRk3ODXpkhT2O6d0gCRNf
zrzNyE4wnn58ikmuOe36+CR5s1SNPmdiEeue0acR0xM4+Fai2TrPp5cwnlEsFtSQ0RSPQzRTm3OV
aCjvBslttmQ6jmUxCW3if6MUEEsBa4NTiPUruVRGKIzXFMPKCPbxtYJQ0r8/NX8+deg5EevXMA7m
fCFnLKdDWk6zgR2AIUTdiP86IgPIwPgq6QPvfbEJnuZjMiC9hzlMQ3mZn0/41ne9CmGJvewqvEeB
7NLQMTYqBW0IazrAej5D/gPpIS8HsWp9eq1LbEPO5MKyyRnogGEW9g+nRI/OOCoerG5Zpu1LF3E2
SEQilg35PZAzIJz0A9CuI2owZ/ijaZJypqZMoc0gKTWg589M6Z7LtcKkTovvvkVylCBvpJwZXVjD
DNFQkGxjuExBW8K7S9UFmCIG+0I8pfCw0KzFxqOjcAUoXKI4rAyJt+U2MfkT5hqpxBEe2toO4U06
blBJiovwrcJft8XyCOuG5InYWbF4EtR1gN7ET99xKqEsd4eBaeI8Px0b4LLSxDl2sJqJtF6wn7lp
HT0iu879GS1gQShPTBOZOddd6h4S+6UpYpiQNws7xkB+t67NVIucRJsOMwsQ9TGFdpbUUpHjGUUv
7x94JR4r9h7x2PuD/Q/zDh00x5Z5bO8g61RC7ulBRwds7IFvdepYd/UYkwuYCpUJZPbMjZjjl8mS
c1tpcF+WIprvMscPNrorZ65vvRshZzFF0oEwcuKFPlhyXYkVmSU30BQozRozMer7Q8UbP9ymez7E
ZPWBVcrlkjWEzpSmkpf4i4YFfZsu4fIFU4VBbimpXd+9XLtK7ESEKh1P19Rw19URLTJsTiCEHrFp
zYd9J185jw9/4KOd02pEeTISYiqffN8JzX+dBsD+mE9vEDyoSnpoObqursU8qhCJW/1ZunhqzVqH
N2fDcHhVWXzc+Wq9w1ueLM+O3AoCTxvj5ffcs/MyHdpTg03tqT8buAPzpRg+eJJ8OFQRO3eaA33F
Q55EYz/s49rSQPNIPcaPXMBQTMf+dVfNUNBRMB0nH2OKIazJf+YOoh1Z3hHyWrfXk3q7ykbipMen
LtSARW5bBl9q63WhHcWvmfF6urXMK93cQufy7a76J4+po3sR+fkB7ISWpK2QFyCAU+z2dYXPipDE
IFiO5Lb5dRdHnxrQgnbsLZiUwPu6+K17+XUL5lrbx+rfzOrcD/bR9t2/Y+lGs7jfzuz/JgsGWl5L
JlgLrGpt6YoIyOHEnVccemxGwQK9wQtr51xA4jaofma9jWsKbMtE5sINweNwIhYVpmE8WrTcTL5d
OvSulmSPpXoY9aLDw06Bu7wcqKTRrAMuRVFEGIrzKjFJxwYiDd/A+DYXZbAGa8Ykw41YAukLTO4j
jALGYRcW7CoKIJc1c22XXEnIIewB0NYPDPe17GedSmwXkdHeJZmX20PLThIt9dUB+5mX0vcNb+AG
M/myyAD1/eVK7VZHPzkw1fnfwmLP6ALXwOXMWT/7osycE0oixByCVA1LVES/wzvHUmWmgwwoaznq
tUZT3GPmJuXO9Koheo6Gxn5FiTQHTwR1+KGN0IIi0Cmuh0vr7IIKk9hHrYhyDeht8yjkAFk/3GO4
Xv5kOecTZJ3FeS2fqXP0Gs6qL+p2Cars6VlK9nxO4kezb7WSHuFACjetDlYc7ojgByHYAMRREXZd
bQ/dTYfYjj3h7Z8bxF1peUyrqoi6BOkIsAuMT4iYBUfTPKYsGEb3YlcI5yb0wXpb4DlW+KQEK2d4
FcEZlJu0sXDIxcRL+yevVzSUO1et71ahSqYCMkyScHbb8vaKC8N4zB94Hv+rZaEplArsrX7/LPgu
4Nv/uNripJaqPV0IJvfcO2FFhO1CeCqamruxX24OinxEEbhhBFD+KGlVOUcA+QmbXaiZUdQHyAmT
AK/SL8ffkpDHlCLj9KN7ek8iQoCKPv8wQ+ipcztSUNQ/n2jNnMnnmkCvVPXFdbRj6qQlJI/hgJp8
4Tl2Wd8pmToUG17niKPeQ83jfksiCP75oyWYanfzrqdv0jQVS0ADa4QgAwp42kCnaocjzybJr4Ge
pJgDGafkYjfLJ6ZExfVmd4oAKX5V6mk9d3tamIY8w+rASMeKt1mjJqBTTC/N0cI8xdIsai2tA313
lRUmbl6MP2Jv4yrPcVzLvgbimlYPBkuvS3uKcprnY7XFlO6ikWV7CAfYMBZ7H05evF4xxRPPlvjY
arj+5Oqjg8kjsTDwzyYFO8Yw+NOj50ZEeaM+n3ioMSb6x14ZlOjrKS/fRPe3Q3TyLbhOOv9vX+Lp
6gAsGU3pbEGfFOke+D0wZxuGSKWTCCyXWvzkGqdQUMRrmuVLhm8+u5vcCxJT4TmloLb1uh4ckE7f
iuXbKLjre2gmwDooUle3XPep2K8jQmHnjLXXVKo4AeeN7pXWVEsqoiOsFqcQgGyhXbdzlgGiZ+2l
ycFBzTB3OG37APG+9blJKSCRl+7D9j+wuJgKNRWyKgjf9QhfgQeRXJGvqwvN3xUS1ztPxQr1HFOA
BSIH4Cl/EB+Wz/pfw32u10adPzxve/oHwQWOmgBtSS/4S93Nmm64/cm2V1aUleEJP95SiuOkQHWm
mhl6KbANtfUcMSDUBhwiAD81S4Hpj3yh0925QPTcIjaP8aZ1EnhJdaBMRxN9uA9NF9La29p9t4xM
fmaslJtUGI/Pe45KTc2Cfr0e1HuaMli8QFY8FsbzUJdxQRjdhr0e2GMSe3/AUs9HRoGX8BD4uhmM
bo7hkAQZcKX8JiXojR3JgQjfRN2OFC0yUQuVqrjtS3z7NuICufFfHRyqO7w5a7K/8HoGvH0tEDpW
qRlXBlIRE6e7EIJeW469JK7aY/aApGOxK1PFVWXecJUzprh1G82nTwwMbGTl08JPmG/LVIgslv16
3izuKXbAhT3cQKoaI4/NgkZpiNHXPxPYXfYF7ExTwX7KMgDcIz2o1ZJNKMbDArdemZ4IyDAHaPwq
fBPu9N8a2EJzS1TNYpwYMNGkPqcLh96Q1fhnIOSrbiO1fHzaYyxp4qu4+M6n9BDZ069UyFBUULmb
fDk8o2b9CeUrhtQ8H32DG1pcvDByf+QHJHr/TB8bFqbbmiQ4TC0yzG3IsWuq5u3Np+O+n6j9RIpE
oIBel+Q15O37MFTr6sf1zBRqgYBPfNEL1hF/oTFcmn8KTQzr6GK+ZaIeujdL3OXQSxD/0jsMrcl9
TgxaiY1UsGlfboiZOhmY2s3CBwYMJWWb7rJeg2dD/srJNooWfwTBJYpn+aOlRV86WvijkmhDaXK1
/TYikcLqk4XG7BRc20pbf5N+YEw9HDehEx3+TIJdTtQfitWNJR1AN+2vSgCkFqY42FTKfsByY5E/
7cbSxkeKYFgFQnIevq7QGKzoeDzekw9/t3rLt9/AvjI37Dg7ZcoFNpk7dHMRihB1TeBgo4RcGGBE
5IwmpJ6ao5nsgezcXyrLNvpwJ1XtTItR8a4W3ePkx/BspZb0LXc3IzvQObiiLk4OTk8uzUUjtFTa
Iw+a89hI1zLcLX6q1uTfjgnd6s/iUvtXrcIqoSar650KNi6n8vN08GPXcWIKSsKvcKhc5xxbf6nB
OlNh/laqMckgRshGXsbaZWzZp1MgKJE7Wq2knT8UlPJrqwEGXxwDVORRYoSEZgvmmD6vRdYN2y0d
DVjYLx4YlLIfaOjdcnDZTNYxbB5R/dhOfF1V4adqFvDdhfGPhgRar4/zHg5Vv/FYcqiW0NiVqbiQ
5f0jZ2vFSchyHtIpzIr+9sKzCS0Jovieprw0I0jHhMzzUvVYPhgXs+olGrHzB8kgutwoXODyFoIq
N+oHiz5SbyXqrg0Se6M1GcquonnRpyOKDXPj29iKT7ov2XdGhRlRnX9z1DpGoJRrVSOL0MMdMSeZ
hujTDUl26oa/7RcAcseLU8iCc4vp2Rre6Il1gLv8EA0nptxBwGQRcnWs9clUZKhA2XnhT/tYcwKp
19MMy1mfK7BxfuwTgFS89IAjSOMhxK3flg72fj5Nib3XBK9JrLhK+ctE+8uUsMqqlV/JPiaUul5p
mKdKB0dHHUFASMDDoymMxvW8oPfCEnCibEQeuo3Iz3GrRgKz0oSpg1CwQS/gY++Segy89baFPdIU
4VE00reGdEJGaxoDWz+bWeRYPD8c4ebJpG11gh963VaF+MksU9J2d265tUDVP9PXCVb3o+p5VQ1H
ZsR3KD8oHuxaSGc+zrsqcbVypq0ji+svRn4DKEz1wRFKQlf/h3tkLuR/DPB1Bn3HgCINIug7jty5
a8GNcLzcITUtmldYpC5GrGD73erluM93KASJ6xTmifR36Ngjxq+P+IwaAuyNJF8JsPEjTRPoFOHb
/CZ3fcho1SGb/i6S6vrdCrcNmX4sGboe6kPyDSRmPxSFIVtlEoGra04TDfpmX/T5gNE7D7l2cT+J
U6TshCwgGb4Ztz2rVWXGdHLJnZvI/XtZxTmdKBwXoU8m97zviAsizTojY8jaKvl3JJOreDW4vyJu
hvPPuEDvUitkuwu8UQzoz3373Qf1lnxmTWbSIcs/3GsbLYh/6PPz073uzOK/TdWL7eYpreTEDThK
0NzomBsLMg1i6JKr2NspnRsJHyrag/In6mNc4D5ru5FgejJmeAW1ha/cxN1SSHY5BaxQNMCdkHvG
vCp7SS01qk5gYK11aMG8tIkfb9eL3WcrxVAqiw5FyH4I5bqTbeQ9kMYTKKVhDV7VReFU70cV9/Sd
vdE3J7t5obaeb0Q2NhFKjYv5AtjiaqtX78DlD9eEc3ScmsJ2UGapbTHyJgR9lqblwCT2yhgrAyAJ
ME9TMH/8pExDRBZIY5rnOp/mx2qs5AiquXvytGJkNJYsfeU+/nkaUkqBd9QkpEYrOt3InxyqJnVh
1I4y1klbnIxEARnZz4UFqurvnCWfQ0PGvuh1hodUJGPK4oVLzhYDsDjtxMUwc2SSI4DkbgXp+8og
aFMMfVVJHmE4cVL2wxdeMEgqqAM1swoUa6sEyph0+w2QLqUs0u4aXFRSdYp+bXaLidjFhZD/YNLv
/ixLaNOye87hzq2a3BqnS7yFNBLfXFWftpLOos3idOQfmf17WQo3mVwUerzI2OfB+VdSy9T8+G+1
glmqj3ZkoNVuYWLW/+2ozVXOzzIaD4Bm00kQnz2NyXjLTS2mIVqNsS/PxSchh8jDX9UUu5CuLxwQ
Z6FbfOVZMuKtsP5bCXS/xVe78ye27g9v6vnQ/KAAXhhC9Ph7pyHeqZhXxDcwmmOK7A+q07qKz9y9
A5+aec+YT4J3iTfRV8oE2/no7DPjmQ9DgwCkyNlrthnfOoWY/IP9XwIkBfX/cs5LcXz2ZLtJHyP1
El6ehSAOL1Qv3Pp/Ipv/+qsuuAfBnMEEXkzEEtAyhGZXPAnyao+FvvEu3bDzJOzZLMz4BlnKr5Z3
VGWMd+U0Mch/vmuBpcLvlq2lvet0Y7+MaO9WlwlgZ6GFmfqQ6bbpfqKUh+XSI1GRLJs3oeopAnzA
8k1BvLCiHbJr2UPxaF9CwcqX+L/Y40yawtrFKQkKLHuF4Q6LdGqh+TPRmbRc0394jGWCAJ/Bribv
NFEKvSoAtrnj2S3VTPbY7HMJCQYXqJTwtNQIfgrO0XEFPcuGfyMnwQi4VxsSfj/rONxLG6atD8iJ
HjtcHPCgZpuJI5LIC8WoaUeVZxoEwaV1pqvmdJwjH3faeG+KtSUFk0kdmk8squ7lXAGSC1qbLn/U
tPXxG/XWYbRUo/ouCNPdqUZjvtlckYRGO2v7HRxkhgIR97mrLgrR3jd3cns6GaEmJTcHgeg8wYSb
ULozMC81DqPzyAxYvNvtmNhYwDs69nl3LcZSSYq6yxlxVxlkfebTMIozcItu6d0f0sqPeU0NmyvR
Zms+7wT80YrKYqXAp/Aj5tTsjzjNsfEQdKhWinpSeA8r34bxl+kw9gkvaRLVNzxe1OW4M/gwfdUx
2KxP3ivULTd8wfFISFVIMxUbPTh66MUpbDMTCGfdvFAy0UAVT7Ucalj24uzSM8Zoeag1N4aBemC8
ybNxTDWxmAMJGO6AtiMmoRboY9k3kba8idxlEsFVQGgoaTkxkTf2SHcCOJHG0l/IDQ9Q4UoR8YF9
mMKaMJr6OW0hZYbGm08SyoejRdZ0oup1sOep/s7H8WA4Emfz4P+KvGpBrUV0+gvfS/MBPjs5KYLg
rQkABadFYO/tde6cyXA21CsqYMqdoF0FTP5mdO/4kStYu6hhTLCVXxcheVZLezNadmL1DGOKc3ca
IdggacHnr+FNcaavKf8dLEihE7MC9Jf2MosS/rf2sNEDLaNL9I+UUUZv3cjmcC33lsQVW07j0nPa
wX3ErvkF/qYvnFmpSsjq7KAbqmFp9OpGZqADMlkDLPbwZXLkdPpu+nMmr29N+oJs8VmF4FmeYEWS
lsz05Y3QjcNGBQ8aEfbz8NPQ0NtHZevc8bw/nDUIg2yzluLsFCiyYkiuEgX3aulYarx1/Nvff6BC
sa81tHJZrT9Iv79JIeZqzpcT3E9B3xD6fSVyorPJQ51EcdME4dGoY59Q9Bi9OYT7We6RMrq6C/Xl
/MjvNnyR20rdH+NQLpsyMDdGnMArJHiHB3xFdb8+RJ6lptOkAG47HYBbNPpGrpZ+h/fEElV3FnGS
KIMQ929OL9s7sKKs7o+piFKm1EfrxpX4nRIIBFc1K4A9PoBu/d7YO0r7UhLu0RV2FTETIeNjdu5p
pqMtstKdXNNfDjljE4R1+shd1L3EellS7JBHRFM/Mzstiqi4N/uNSUA/mUw94qx/88FNxrx8jSXv
utgjOUAJucaWt4Hi48TaIFhHE0v7GHaQO8Eeou0jxyjJff2saMXmTXP59MX07MsSepJUkjaqCEhx
qvpwXlCljO/Rabm8F6XEWf3ngaDgoH83MG9czOMF8pjL2Kv/9goR2/SzBsR/JDsxjo5dHRlOIikq
mwZITNnQQFcVgsKnoBNsaRitY/fI1WFTyDp4hfW5brdL7lZhfwbe0bZswByKSmR1uNvw3bwOMwKo
Lf58+4LMrNUc+Ot1xLGHoV7jC5VI2F6dSWf3F1kmBXdj6dhDkkOpqbuH12WAJR+s+2aFXzIuW9uG
gDS0wf51G96eNnO8l1wSoW+IRcrl2DY1srYrY4i7pIuRyWTRxV+o+xrao1kmijmGHusnoVhwLm9p
yCNzvm8iK4N2d8UJpBNAVJauAVztbF7n3OB3zTI2Dk/gEIllpKDEojDbq4sGVqz4li6WFBJFqoCO
lA84VD/dMv3sXM+DT9Ve9Zwy0CUrWzPQSlILN4FLZcrzzl+gOX4v7i01ntSu96DsoPF3UfzdY0vP
l1WUw1Xl1dQEE6avMD8rN9l6kmPSdwNejQ+cOMwMrq6hq+wO3tJHt12vove3md7ONe1dyu5fLeKf
qh1LSfiXveH6IzY/1fU7SMJY7ZawZU5jH8LNnYwKrVMpNTFsnfPo2CDVkJ8v148YcBHhWqhb5UrC
5U4sJfwuf0IHinc6Z1gvpOuFK4MZfX1nG6FOdJBVZQc/N1qWVDNlGcDrw+bgn/85Hi6t3kTYsvL6
R4MK8ddNznyTc0/8gFyYa5HFnFksOf8TCsuVMDW91yggwazVFX2uVccR1G5EbAmukAX3k+irw3C5
B2wWTwWnCTTJ+dp5otH3w6bGXKYE0M9ImNmlzxgi5XX2y+5wuReD2IsPX/cwlQS9rXr8vL5j+GXE
CR8Zd/yxNLaHrKmRzs+jjH0K02wpdzdhiV7tL9v9UCBzV/WSUZ/mMI6EmWacnsQ9ILt4YUTjDPTJ
TsFDKxZxrt9GatQOC7JlmOtau6ttHxHItoTxk3U/DKVvhjJRbNQD/CYHFIT9aRYL8dg8iqr3cWbL
UzWBaL16WaMAvkdbQ3gQMfGnPScLuTxKE3QnTw6gwCuViwEvGxk21h1uLI8hBOwnv5cX6HZqkfQj
EFBLTLm5ivUqWafVnMwZnwlsQogjWZYlmUCBHGcddgdYe0ZMyAr46RFVeXSXrN9UQ19Cmfm9zKHv
pUHXvuzMqVTVRve1dCl/W04VEA2hQjp1OIR1IxC8hXIDavEsQHSp0ps1Mw0+wridire6r3NMNVvj
USlhGddOmJWHOS1QxumyEcHvnuxBGW7QZ4IfLcohbWvIoIr/S700n+/rjFqvUnIXxYH0Wo1yGCWc
Cmhq86A20kiIaFixLyacjQ85BpFqxy17qOrGRYdTZh42noMcOtxhgTii//c0w0mbSVuGTaAGjnej
Q9NwCqllJAkg/H/tLacSzQdtR8enquErH7q8Wtn/osn9frwR+OzHcq0j2lST2rLY8HYNeagqWndn
ngGfsztYiDjdwXrminD4DH0fGqUYRlM/19uMActi1TlLT2RVBojVwUtWUkuKbk9rVT5MN0l1xdUf
iUrfv299pJF+P013r9L2VSTxtsL6sk6fV0wPsvWlkpNLMDBmO+zi9VK/5tp5fi1KqLyYdNBnG+gt
zfkC8qdAbNwoCM7t123iPd0V3/iX95p+Vu8ER8zWuwEN2rV6Cl0CtUMVCW+wEYpe3OdK24WwKMB/
HpKsy7TBzhniNf9qbWdMp9l9l16hED7iVs0V0pHW29XjOiIjutw4pg+ZeRljbLsY42AUWm0yOreW
aDX1dB5fSa40NOAIMVqEp0f9udAmZncpdao7hnLRKEW8HMK682NoHFIVBDianETxpyN18fLIhpW+
rC4qZVNsh86PSCJxVd4Wyw+8yqIjimnrdfQTEVPTstrGbwLmiwNrPGseTxHz4CLg7gFJc8xs6Rku
KT3JbmgLWQRbouAn1gnMwd8rTDzHNjRk6BRH4IS3cGxEIm/A+SvpY4zgTpSvuKf/TcBeb8z1T4zL
4qmUT2xvxz7OZhZL5UNgPKBviBVGnM4IsYUrWSwChMv5Rpr99uGhIB//7P+zX0iWlAmnxunDwSZZ
p3I8ogVk2P3lNN/lwkYh9+X6Q7BAXyhY42CUV0s9c1Vfv5LzuD3/v/uuibFq2f1U/jSTa9GzksTb
Xnapj9JPGqso2K8OqOts34cFNdHHOzU3i673LKi+8H4vZ81fhgFyL64h0iDPqJV4udfOrFm82VA/
dFqOdMQx0SRzxmH62FgVlS90uVooEApgaFTknuV9ho/2KUxxDp3MQEXE4IZ7Bq+Ftw13PPqbGWd/
+Svc70X1s034ooYZdq8FSASL8S21NUzdAGwOY5QHvGecLNqvyzrwEwkFrLiJY6v4p+mukniaKE2D
PrLDpzTMW56v/ealYQpZDC+FWMjxVt+LfGubaTezHe85ENi7Ly9J5nVQ05gpnQ7AKBsL6Dyn7HUC
7CVjQkilhLMP9/c6kG+M9Z/PNGOi5gghu2DSkro9Gn7UfOfzF6cSk87muAgx/PSczgDH48eAtj81
bECfUyAhhilpesNysurvzNDDSWwbnXp0fCa5bYYBvqijh7wk74wbhSFosGB5q1bddlFMdV9fn5Sj
MVgkxqM2ObVqFC3mjAgBy4TzxCJm8Atos9fXESgZa65VNfnB8gVanrk1K3T5t8d5EbhtfSO5KT5/
dSzjIKTX/kNQCxEbVBr+/Ridhs/BnY4IDlU+g4wy56i8+kPVPLCejCQg/nexmNxSgJT4Y7OB1pZa
XLvD2wRv/tvuov/SLXxLX7Dw5sDWoIqAsQHLnNzis4/gxJYAtyvDc4MsFzkeNwSvUZE6Cg2s52Mr
PQx9ZIKnFQpOAD2WyZm3Wv30stEWRC7b2T0kfX9znoAoAK/HhLCNyFRkxlEN4dP+MYrLnwtdkdKn
DHGaIgVJFxCOowAkIqTSxYIQdeXbEB8l9zdHIEFjCiY0JKXg//t1XevFpUusAP1p+GZq3HUSsNUJ
Elggle8q9lQsIPouQ2BjR/nSTAFBrFTk0MjfrgIlPOxqh4XjzvoAi4fJhtJOMdpLWVDtQ/wRRiHF
v44u5p2sV4Fu4RuoFCSiIgTb+ZHTv7EfdbiSSkuPPwNP7j+gUN1CAb/qHembuBOgdO34b05IjUsm
UN1ioWPWvGExMioxWI3QNw4gzZDbxYpc60oy3wbDg8sq0sMlt1YVsdmyNwD/NPNuTxOWho8eXKzh
nJaxpMUm4t5GxlbEkhCYYNdFdmposF6Wb+UYNVEiqbrBwtW/0UDqVyKtKo0889E9uvFv5x4fzbOL
9M1bXhwf35Fxysw9TBxYnxvD4HbMc59J9Vt+wjgun936fnWrfa9zsdvO2ho7v513MyjxvkWJwTAd
nFhNF6Y7hop6HTKMYvGikRxreWJJYCrWeGGlxaZrZOzFRvR1JJfWaDIL7iy17x/XnDFOGecfs3oa
AMoOGF2FL7QsGGBW696FUAbS3VlJfVI1/IWZ21m+7uCPJsJ5dYK+QfrlGFKk/KwVxEnIP8yXsLur
vB1oXOMnkHjiDjZY1XhkXEyd51oikMGGxyqKxYDv1LRg8egiGqkHwHm94CzCnhofRFNkBK50BiyN
3YtBT8LjtISga/Nz5d7aKp7bK7kuCW8ynkfcRhISQzGi9d1c2Hx7clT3hteWVEWscNsjY92l+RZZ
2qqaIEMUWYWeHV4324XwY1+Mh9MB6IlRH+e3c733dEYQynxrcVQakol394IK9U/sMZCZsxDOsRfY
rQ0vjDdoODJnVVrIzokIm+PysIrcFRx95ewG0sBwsD0LbA5nfi53mJi1zMjFH8r2trejvak7jVz9
oalIaFWvgcwT+7J02h/E0C9pznKA2fc1cUutfL4FP4W+LvGa0XWsyE101z520A4sxzLjo1ioZSmg
OObB+t9FoWAw8ZAVD6yPv5Ahbrw4/ORWgfPmRr2KuC83BzOYn0MU1tOmOs3GqgBFmNgxRUODtacS
0RvffN8rH4mtVmYE1wcr/o1+zdlWopnrgCUqOiv5urC6V/LT1fUDGHPhCDTRnTMrI6QOFMbMHFIc
YwEL2gQ9qeyeFoGFG1ZXWWMBHmF3lrPGU4rtbPDClur9OztqpSpGlwtv9/bs+AjRqsRP4fWqt8gB
KVsEwbfMngx1giPWcIsJSJO5PFXCZsWNk/i3jVL1b6CXwKFyH5g9YkBJgZU+D0kqEMYwfEb/4Xeo
NmYioSuLFpgCB8nKPgktpFGUlscPU+jpvelJt/KF82k1AJYDL3fcbAhbVAZu3a88ltInlkH2kXCC
74FaEKokiH0zpVXH1NGdHWsJQJW4cv7lpJ/3dxyJoJG8FDuwHpPNMPNGKwqvNDahnGO0x5+uxP2k
76xMZcXAVx5w5xSqZYhcCsz3ft4mcsAls2zfYpUrC+nkPf8zsSoM18vN67/CwB6IXp6iZNODmBtK
yLC4USgcck65MtlHXUHlzsVP1GuQ15IHBDHp8hGdDKYjgw2hD2G8A5F2y3YgovcJ88wBOmWCFoH9
QcBXyIpoC7WWujOPJaQLdb9Va23UYEFQfvEj5j0k9V3jm45hp+eQSzcMxCVqpb7QdNWoTLdocsgP
PqX0oWqbpR8rR8nwoHNf0HPdg3jFz2tSJFhDvfAGrpd6v5WrhT8xzPWKOQ7lufT9vBApiTpsksbu
CH/VR1IZ9pWkocJpenbRBUkwWmgR8Kpf9FE2QEakGNcb0S6UpKLyh32+cq3i50od7pLwZLDt33G1
Z+SQD+3Hqa7651gNhNUXlEgpf/NB0lpjxMY8+ISCCEPiDGOmDaeQi0iO7IdkssUKF+QrkmF1ts4k
fjzGB4EPZlwoA9xlAl45Xy6dj/cLq2Sa0vDAeGdW9sNyulhfBjvPVzQ6n45fVzcqD/Az4TX3Mlfb
avjBo/4k4EHZwyiwD8wfdxD4YuRRFGEUl4M6EOa3LifIfhnmGJYj/mNJqoN5Rnm37Qs9GSBdXyUN
F9p6VVr50V2Vjkr+ZGH468xkb2A6NmBsve5NaOy/+fpfTNJTgCosMYQLnJ13G6OjPSflMrKLMiGZ
mLgKce8VgG1KnVgwqkkPMGq+N7+6iN1jZgPOOPL/ZuEGsEsoF9F/UeSCbCj3ZFfWQ454fC9/4ktB
Qd8A0H1Z7KmwKf9pS/r5ZyHNrAd+SEADFUYge7kvvcJkB35Dzr7c7zud1/L9tqqMYEzPk83jZ66y
cAiOZtzPLzDa1IFJSJnzvPm8wMt3NZkmx9IlPdm2aZUHtJ+TfYGdAJt1HrdyoJbhADE8mWsnDAlT
By7TOg+e6F92zpwmR5wNbYE1uIOu6+g0zmCkjKyiUnhbO7/3SyrvJNDBphYfR/n0IOtLRoe7ERRh
xv9KwooXdc30qVr2KTZkBTAR/Zb6ns1ToczzRqsJbMDra1laBU4PDXpKvDK5j06CSQv7HmT9h1t7
5LJAgF5G8qm4mcEipkVsLWKGakazMgYUZChPmp1jaiYX/CTyXNWesH7skkvF02FgjO50/zCOpc4s
zYJfkQaIK1Y01Q+/VTcJifU/V1K8vUGCUCA6IvYkxU8EGwnat0zQoQl0oMLhu7tZxqz8zj5bHxLW
Abj1obMUUk8aSGJmuYxLW1qR1N121bh4JfTCWVNzB9TyZzsD7RndT6+k1qP5UVjrY4xDZNQHnQxH
ygRkHZPVoQu2Eyz7i+Slc69xYrUZIU8YEfutblbRmipwelsht3mAwa4370XaxE8LGvzezi7oo3Wx
w/3HogJZZ1MP8QYT6x3yD7rJ9d3aCweJToCC+ipjsHtKrdP1NSDGaLoto9Pl0kURCUTm58XIZR7X
5K5oI+WvuAVeTK139Gl6wsQVYIdpYSUGP5SVY5GsxkRMvqJBbh/7FhjObhJ+3OSb0blN2P9q10aQ
+dtXPiD2RUI4aIqDj1kq7xvYB4NW45WGOvfVm8nN9hAioC8PXHoW4MhqtgmhXon7elko1aTO5TMm
3E7nJU5MIS7XjIQMDmBDAAayRlbZW9hs0YY+cnSJf/oicBL7IM6D8nceTfH5gR3ZUUGzi8Uzys2a
lJhTZANhQB1X9Yvy3JIxrs/fDdby1UPRdjv8MdTreljJ9+HyG9nlJoaQE7Qqu3836GC5di+UtWrL
i7w/Bn94gr1gv8+0k8mvEkQ0dLZCw7B184ZqYQ2Igkz/6A1+jFBW+ubCEpJbRWDv4gfBuYfl9bK8
ARHL81d5SCfHB3ZpFw6u8ngPwzmK9jCnbqnmmlrkc8kxdM0dDKmyUJGOd+vViWjh9j2eWSxZgm/8
tYoYVnFlK8fU+UFHOh5zszsHHYIhqOewHIqXsCe9UgXw6KvuNFj+ELnyIBB6zutf0h6Ngo8DhXgt
hFlStAo/2PWb9KSgVNsw/AYqGJ9gj63bjqh/56jqa6GWUAFRFVNNq/44zr/EVS37TA+/iiKS91I6
eBqW72BNOR+dX+MR3BZ6UWB4eJaHngbimuhAX/xnxT/BJljL/C+1NWe+4Iew1Jp0+m7rLREL1yhe
0kkC0QfSd0K3FMv7VcUJe4V9EgrYlWV7eJBtZAlrVQ7hiq+0MMwygc3TrPokvgwUCc/wquLyCwB6
9ATviXXgYaNOo+uXnuIdAYrlrpJXJ7SoTcufa1coMiccpOfw0fGCQMaswrRpHF5C+bbvhyyWf7Av
qlnnA3OCXxn6hX2ixXW5Pse6AMPf4JsweVZNgmY+3ag5mmDYznenTaDqPWrrG3GlyhmUYKPdUq5W
P5SPaZMLN2ggD3nhICoyVq/RNaJRmfCtbvqkpFMsE6vZJACLcWU/+yJzkKoL08bMl+QBn8cmHTxI
Z659qcY2ynNtcoYFRbs2Xuwo688aD4qT0HIfjf2vVFpnE/GzIYU9B3KjHX/rUrcghyxO3QUDMYp/
QFZMwuzGTl29fSP6gR3wEzXfaKyJwRwCodtiWGbMeClafXP0ztZ+6XJB9LsQmiLf8TR+d4T/9S+D
DPRIOJoHvG9qoOtHF6R7SJ4Uw3eeDvlsXW0r2PKb/5berWV9OZPrWrYQTCfeXmBXkRZdQic06gj1
xB+7KQ1h0A/b/rblwj/XNsLr1ef8iOu/gK6tdPUznvfqrIQaC+3cwnQONvZM2Gue1oT2zmtYJIzj
ZFaEBQbzbCoa5ODVgVJBRd/SuGx6sxUfbBA2Yidr7jocmu7ELRa+4RguuSe5NlSD3NyAkntGguVR
lGfxCWgP2PqKFhlVg0xqo8Ro/dyIV0Vv76ZFdj2CxA+fdIZrs4Su3qCpgE4nxrgNbnUnsK5LoNBQ
rrzy1zs8XWTAwemqsSDHM/aLeqNp1MMzA6o+3DpGGs2UhnreLuigu3ggWUBaz+15xVdLzfw3Ux7b
08DLudkntv/Ty+MBcoj5nhERXUbpQUzTq3nXrDQNnI4iBiNONxkD2jxAWAIaym2/J3GibljijJSr
JyWIoKb+rr8o7JLPYpTIDn1MlJxSquYGSyeY6o0ZZ89rs+/NGbWK9qGXdm39S84xT3N3vT4TXFCh
llJU4sl2PyCQJfC/Rs4zzAzNaietfkvQ0VHCaBpaLGbu9xhpPlpi+UwX4vRj8bgvtRzKsYHwtZ0c
F5nBWOxLh8O5Wi3FUl3dJ7gg29sEXnsMgXF1gQPEcGxQpLW9WUP7qBucq3sAXHNPEZiN/3C7lbRp
aetoJwN9gCGcHLq26anHw95LcdvV12MuhUhcLpbu8XIiC186eivrOFU39aC/a98dJgHtpGTMyWOk
G0rAOCgaUNiArrOz+ZYHN98lRKYi9lT03ye/RffRveWKUQIb1tqVJ9cJqzmBIh5RDYza7f9lL2Qt
Z44X5GhqymIbyj8PD736P406QpkAmZLctgNs4ZDpfRWJcEaTtnCeMRWuYAO8g11WWDQ+LAehz+TC
5LBQz/bHzHh+8ZFg3j0uX21v1s3upUsya9MHWaU2UybUnNpsJYyO1ZGravb5c4pNuoZTsip5iUqR
eUkP0iqiRY5mOZUT2SZQg2PoCZ7VwZ49LahQg5C2hf61Ui15184CrkuW0AM9ZLloyQ3OAjE7b+q4
aTaSAwuYcUSCRC7r7Ti9dzuWK+aoj1uvxPJ8tyLNkGx2z4CtpaHf5j+0qZJ10E7n6dFxWYJzYpol
W46otvVYBT8Ccxs3WteRqbR8It3eba7UANbqi35Zqdh0mPydo3a1+jgBjGxqwGZyf9dMPXMeQdyZ
PyhQHFK1EOabcGCJZ42n/ioWZgch04sfQ7BW8G/TbevTZz/WVEyTLKLTywkrhHvgHzl/6q38bFz7
ZA6KvGbVoOXScwx1Pl9jyAHyPmsNRvXoZUN2k8pxJfwHrWYWdU8FuhjBUipbuNtf0oCGz/mCJ5c1
6HPfXDpzCdQD36c7KfKsh+qXtEUU1O5ozu5flw8026J4jVMQuHhNnljOJkwuGdfXTRC/4JzHN0Kg
0VtMGdoXD/QYh9wuL2OeFcSu7tbW72L3UMqc7WZDFCV9IT8PagNSFNKZM8ORrZelhyAMl172hdRP
SA1Bf/FuYBaiGcN4SwVaAx2Pb5h68gewzx3k8/6T0bzznmh2vLX8aXYfSVZzTTX1iSlpjIg5dz6Q
v9JYZjspfnM7thRtWL/XqUQlPh7vdRJz6HkDM6MTynzoTGvpewmt1nROQhEKzu5OhyK1xS8YTLn8
XR4H1yWCQIO2QgXYsoGcGRO5J1WAwMw9pBAPHV7720dYSCc1mwFf7GOfoPUV/QJtmJUnw4EBciEi
6XdnoAWDYHQVSg74YzqRk0PcCdn289O8os2hk4eSsX43RSbR5JX2vNFTEPG3cZKas0T+kwtT3fex
VrnAU8N4D/soxRWF5mZcxS40xI3fpadeD4f3F3yfxFG/mcEfZDwQT/o4v7EsG562kSuveQ5IHw+9
tSs63a7QWx/ohJoS5T40yDCQ//EDCKJyqU+i+V+3dW1f2ZrqL8QVmF7uNTDjt73nFwhcuobFaqRP
ah2jrmZ/kKJIkGks0USK2h1ZI3aBVA4oSzio9dEKXH05fPXU7hKSQET2TCBfdncwYMEYtpbEmQXk
l90N6TB6B6/0CqO6tVgZ0SX5I0jvgdGEWv8UvVfz5eWoWTf5rsJpu2AC1soCSttrwoUTBlEDUOUp
fvWkcD7xeQvPKFaL2QUOm3VUFC7kIoYREHt9j9xAaIH563Q689SKYQONa+JY4SguEeLudDTvYvgu
fpuM7Ja5HI3TSqnz4U+pHlMyz56wOTuxb2FeNJt3Bxz7bj/YHziJvnfuUO6zHPKbuqR/5EuFASHo
nSsgtVV4C/RuIKPXEKPO6H51vn6uYHHcBn4xau81uRQZQepZMZsd7FHY3EVjLsThHaUvci0boMUL
UgbLhLKrcdChSyupDcUzU3KyNy+95dnt3KC/LjzVH6U93sIzk7bVpngAU1pttzFqVXY9Sk6eE6v/
txwQEhe3+YoV1ez/OdFvC2HMCORUcUgK4G5exNeaZF3f+7E7nZDZ82C34MN0771BLRqRZ5vdBCWu
M7Nr+2IKZqOO8/mlkyrHYx+1Pw6LcFWdM5oBo+gYd+zOlRmqro7U7irAj93sNcExWLDbxelqyjVv
fviMlVYU//W2DYXJuVMB3AyQ9ccADdPxkwP6ChHNGhV+Gd6/k4ZaG6KwVoNGPruzwf40S8UxKgrS
/+ICv2VAGHnubC4TShZsf9KQ7dzJSw8YE1A2PfeAgwd5EnDfq3o1jx3usyIfCoL3rDu1ZKDS4xga
894Ugr7jUT3xKCapWJSoRRta+rLR7FgK/NaHTwuTZYG0kL+3XIt3Xm2tFWET8WqBIU88fm9YGm2q
JUDlauDSl/TCfgawH4TzD2pbqvd4KOS25lEOxP1c9iIZf5XiTCbTxP2Sh8JBDL7o9NpPWovM3/Wz
tfBnCifYqKVfFOKwQ37sWjj8SoQhfwCo5YvogEvdiOP5NpFV2TmEukgxq7fCEv5Va4vix/IfJzwh
lQfj3mTq5KKd+75QJMIiPG8kE38v3ydw9jTLmgmix2Woydztim4P1MIgXMpWIqX9JE6UjYIUb1GM
0dSoX1z0khSotFVVc9949F89qKJlkdmUMvTc75bs5xGVvkL4rRJ3a4PP8gBxDx4hWTfpRuh8cJFB
DfGKL58EqgN0utSsJ0bp+naQlFYSA5+Ex5lysE9eA08jOvGnfKYoMk/7uRj/Rdy9L1ZfKHH8Pq3M
+9e/1Rv/2wEyt4aEGF1Xjj4YMAJlJC1+Fuy7VCyLrk+NsMX1FdtteEsYuCbA+uef/k1nxpkV55yH
Wo+0pm+5CWk0QParR/1796u+jtl0adN2ZngcpYYo+6Aqzken69PKmEkXlGZZKBwHzup8lfJI1LaM
9GcaBCtwYFfAUD5334l7ttzyiXpQzWcB6vydEzTHEiVyQQjsKGPNhN59ISRlTqiHVs37hjRdjpjP
JQPdu1UzmXoLRBZ6V+ZBNQ6jX+F1fKzh/AkV0NdEmEU3geosgdgHuEmp7iVKF6UZZbNRJS1Zvhy/
9ct5lcvvzzATfLIeyasHNTbRCSP1WoOR6DfRLa6Org4IzivEi6Xq8Lz5bT3RjueGlE0fRvDX7Ymr
tK4ecn9Lsfas2XvgxP2wHtswvNXyuZMUGAfzl3rT5BJmo7wfLRGXS3+jDICf+s9xnqSy+fh51FYW
ZXBH0ww84yFLnXLjCevE+yKMHlSanS9rV4QNw2Fg6zWrvlyyDMgOaidvmhDofXr4AR2pxR62M+xY
R4H2/8tmrgTszkkAuuy8o12Bex85SCo6ksHiTWtkEsFVpqX4q1rJypZQ6uB95TCPyxNMK0A3xcts
rzUxyUMLfuFbTG4gYJRG0/UZCaVlWeqrENeTCbVT02dTeSr3LlbnNZj4mc5uKCCMy0rtl3bez3gP
Pzmf1I+Qvu2vUOASusSAsxDWAlL0ppFS1DdpS0SxzWHOOwivi8zZKNr0y7x8d4K+A1qn8RheugSJ
4gBEjiYB3WQ/Yo/bZhTJIlyYO8MxfpKz+bgIkwke4rmsmhqq7W0JpHfivh15vnAlmsdX1P/f/cLx
bsbpCOwnpZe7wQmiCt7wbYdh91M5q1ckwKrtzko/IxRc6QDpszm0boPO54CN/sY+Oc+DJJ06VxJV
Te91MGE8TcDYlC16lk2ZZIoeM2j468oeYdWTvSezYOwlQ8DREe/WGD3796f3rNm/mBcd0NJhX8tS
ycvJZ6Hyqvj1/Q0SzMskmU1LlenW9PKaE2WgM3B4mYCTSqGeeWJKTyc+zwMW+oW70aQMJjLrT7dH
TzV4oqUxoli0J65t/6AVYLGLeGdyITplfhVKmHfEmQIEPcqGFkgiWpD3Ehlzw/lP/MJ0uaqbJAPX
z8QNJs1k8bSVVne+Q8nwzHtD45Qm3Y/FMYL9HIL1MINZNvsyXzcmmt/VFsVXc8Yco90cXvWyUmmz
uK+6P0JpYoXWT8pCqlX4ACejmV76oZwHYB4qWbSrBacUObh/2rl4mN5YhQj1VUNqMERp6ztmX73F
sngIPb8JVEh5eF4aMrAjrk8tv9JqTEbCeI7DoiIs7LEhUZTC8RTWWY2KvbiFvcGZ8//JCLr2ZQtn
Z4mPP4FRKKUeIBgnKz9IZBdlfUsaf0s4LsVXi7T4F3czLhQ1fwxoNRUwpXn+/Mwze1dkpMqdzEx/
YrZPZJZ9oDzpP+vKVah9Fa9CTCNC3uEtxXdXA+Jnb5b1rsTO988A8Ut8AOH0swNCDi2LmoNfhd4+
qzQbbCO5UedsTN5pN5RKJK03zZKLLiIL6DRwjRrSrk5XlhqYUjGU8w23FPDCTp0GhHbxM7zbF97z
sAZqjVBUCkriQii2S2ZOWKWhFiePfiwleAuZMMPGpbhqpzb8ay8i2qkVtUlsjfioD3XNlY3flQ3p
6xtjq1ls1+vgqJOa2v8DR+3LFm6a5SEuRYga4IK/eiC/Na4f7jrGctGztVwGYWXzV8lUfmzi21gh
w2/ZktxoQ7C2X3F9WVOdVYwkd5OhQEbi5dpUEWKrnKg3cbynGCPsiPyl5ht/8D7sypnY4GA8X2hr
3vrElK+RAApUx9T8dmpWEzmIFMyomAKwDCf4s7lSh585D9lWjQRHuNLtBvEaP2Mm3vNIvJBOjbkw
RkI7dlFFQ+WFeE3j+gwO3AuWTmWF67G+8yhyeMwKNZT7kIYwZP58uSzE5l6z3drqVeC3OyLC6ZKt
elscyrZzkyuBTyh8jb6iHuDArshUW3fRATQp4Uyueiq6uYRj90LaBtvh/O5bbhH5HCayVHHwFpjz
LbRju5+kKlmiGSEZD5fU2icqug8kr+EfDk5UMTX9UAbGy7jA5FLDu8YkTac3g1cPuYFlajEqg3rh
3/PIMYnwN8Mj4kFxOKk2bTeD5hH0Fmzqq/eLsXojyjO9KjCqxGjKb/sPjeXPQUVK7TnHZEgHdimW
kJFpaGc/oy+fABYH9RPqobh5Tm6nDVxPUVq/GX+5sjfB/eakq6JHD8Yxf+fuaaXeqsIZBiGcT7QE
Af3kmATcCtGD26hgaV5YRJUmaNlYkyp066dPGPdrfaQ3emhUdwWK9Bf+HO+S8JTZJMd6la5yjN1L
yP5IiQdQGfpdOn+QoV4vBaOb8uUXc5c568QIMXbHb9doYmJOj01FJzObDxIAAT6i9QFJlp6jH8b0
porV623RYhcJgufGon6vxZ2s20MEAXFBsNPZ9GtrTWcQbBd+V8tEgReMjDPu5PbKdGHwQ/09EIM4
TEw13Dl4Go4YjM3R+7GpPNBNMiPPNl9OJgN1P1IO13895K1SnLgm59otoN1+gfb5I080yogQ2WAJ
AoKTb3Gz2iacQMIAlGIP/kIeZkB2SDn1uX9nVrIrJ1hsLfggQSMKiONf+H9SmSoqfZesxhkXXqFe
FYClumwtiGU1i4RRYWNDF/n94JC92S9Hes3dnq/x+iyC1TYrrm9V8hZJRNyvytvAuJ9sd5FMT1e0
4+2lbM5KWsCdv7+zuYG6mc8KoJ7qDmq3AZb/4T1CLbHtf4M0RdDcEcG1/yVIBVoOuNKbt4UScqVY
4xwbM8ANA0Z+Vp6afCZbL1k2eXpzTU8Z7eBFrx4dhqjS1iyhUv1MKbCQwTBvlAk8aVk48T/53KSO
ypQgx6ND31w4mL7Ahroobbsd5azBKzcDqlrRUTnVeO9a6M3d/FcnuXI9Fgt3mOd0PU99Qh7bM4LC
wJSlOUbP3TVC69uisNGl9IeZhFKM+6i31zGwfcdbiX07m9+mzG2R8WeGnHtw9QbznJSi7JTj2czS
S4pqSwo82n5IqWyENbrHJv5iO7A5jz9pbKVSs5zt05VdewSR9yRYBWaDs9v5oPClPDZtf+6M6l70
tB6rSYdg08YWUNxH0xsdaEpE+FFY1hPUrWazwmZitPZUjYJ7fxVKE4GYB01c2siIS732U+fvgW1w
ymg2xGIjxJo9uOP5hG8U0ryn1YS07MKE+ljbKhaI/u7j8O5Pwfd+mTptFI+hYKiWUp8dVzq5yfhQ
UcOypW8S0cw/xTvmISefkDOO55b8l7gVsUno61v3dVslKbNgrHqZ+tUON8hUbmx2vFv7GZmt7Zky
bkM2yV5x5R0LgQMpj+bZFNeBuQ/TAaixYkjaFYxWPKCUcc4kYxfXqmQm6H8PkmOaE7B9ybhghnr0
sQwfuY/3gdywaTWgF68wPrLEhq5cw4SzZlYqRps8xDT9/TU4vhmCgJTuzwKVQsv2RIPPeLIcujNl
WKvnuz2U2bz1uz8udeMeFQ7VTz5Ec/tZbo/td6uTXyvPrN9wChxLYhoPb7tjJoVXYrHiioLOCyWo
RM6GFwJR+ZZ5H0d4DUhE1u67iuHNDziuz+MV8cLI7PButhwNT0BR3G2zls626aoEEpwMsDz6mB/w
tKlusfDjZ5FBJGnnSN6+VjKqrBmtaKwmeha6P3u4LPwYVwhq4VTBwiF46E9ENmhAvtlJtVh+EWqz
g20pJRMRpZxQJyKscwZ7UO21BrywGuuTQvDPUcP2Q6lJeTk780yh9Q9z969+LRoi8i3bdUyMXbBV
+fP1q0DsLRu04ApLE4cjrP9fIo1Q4qSDuyqYYXc1+dM+TczOTcbFcpItAUvKvLR1xZuakDNE8sxX
5Y9oJP2nTtYn/RDtRljqky5ySLu+xeSHV/uS98daPZTjddo5zl6LKY5vKTOocRtF8ibZwlNFGYcm
SV8rNC61FV6C5KeVs+acYT2jCnS3eYIgLfCop5FXHmne/Wukxr/dnjCH2d3C0Dr1pxeSP9iBSxVO
QlDln8fBWRynpPvFkGCXLtiWcY+qo0dBYsEQqRDhzwHZY67WuOeLpcRzpklh/5PYbzRU258x83/F
WqMl7KzgJ+ZHbnEznKCr7bUDeLKgzFYWjva0BCRCIOzuEIPD2EjoVYtjE5+vh1tgjIh7mPUPbtq7
Iw1M3efsHCU1U8fFmQ75sQYVuRtvstWUS4V+viseb/BFfpUmbB0YlZGsWWPlsFwknQaGIwIAJiv9
Eq2V/rGohMmRizMDyHGWBPLSZgF8uKWzADa07fUjY/kmZvNqS2u6UDTUP2gvTaIZD2oDOR6MKvUn
iXVMITzILar9/3R9HcBPZqwBkB/alfYuGkYhMG+9N1kQEYOj+izWsnZgeNp5zginVqnodHKcGat0
wRFoNo3Z0ek/LM8tgw+NppJUH7aiMQaJFrMZx1WprHHCO5I0mfsY9OdXCoLe2G1mQGPmGlVElk4T
dEznTTDal1wJdnEWTC4ZS7TLTxuAIRbLkX6cB97N/0y7Arg1W4vFvW45WBwyyOWKy79EEvoV+nUf
p231DWfWmx0pZkl0MAPUje/obk4fH7LnewRyzNINYb7qxqBnf7oPUUDrz0MSE/I5nUw4mfJpZhCk
zNxJerPwOOxAeEpsR13pqwVAlpE2Xq8Ys5AALPTDdYRSFAJP6S8xoUlZE7W5ghg3Yb0XLrMLIoHB
naJHxQHzwZus1syOgjGax1lKicXXV10wx1hHTX5q9hE9fxFXtfnkuQ/tLjkuxcfv4eBpRcz6xeHo
tjtcl4cd56EjirQ7VpOuKAEzp8dTY+c9SoMLE8hrWMtQN2DfQUdC+OqvtFnqhRHDhCr/5bnEHSW7
5exKE+Kj6wBsoSEdrSha36E584i2ScZlIAodweqLpnrHxDN7okX8z23yAzfAWFYDQ80FGVhpbmJ2
BenosfyGtIm/eggoPZ80kEe+BvVMJlD0Y/xFe9w9RlPEo5pNYgQeZFIkFnE5l6b/01wPx1PfoSEO
UmYWJfpEYMf9ScEgo61xeJgGKZw+lK6yG/8RMDbwIQNPlbwv6rdvsJZMksfX64bnj/r4QpzNNYz/
0YMFF1YBBtU+pPKwTG1Qbjold0GPrBuuMW5gWvTd6CMiwz99v//pBDI0eBZ05+J2wRftsBi3HISW
tsaxyedgSOFpADcHnQwLJbdVlgfAal+/w556Qz5UTvwG4yp6+q+17ZDCBOebzyVtaA+or0usNuej
QZ0Ns6z3Rl/NvJKIWHLJGvg4zdxOGb0hPChHw6fB2ji3zrQujJUXmHoPFHsViCT/4JlhvANngftH
U2p7qURhkCIBU+TEuYiR2yQG2mr8DSEvjnUC0rNfdjWyijkDmg6KzHTS6l4vFNsGhPShzuZdruTi
9Ngyve2DEkfPkd9dojPP3Qk7+gcJup/SqCRYq5BswvMhieII83n3kn7FpG65OhW/Bl8JOdcLmQRs
g9lyeY8rQe5dis1WncRUbsqpf4BQisx4yE8sQ1aBRa/nRlReG+y2wXky/4/Dnl82Uam3OUe+V5Vv
vcEslI5FwooZiNwBmqH+/23bmuBjUKlSwsjeYyrGnyZTiVvT6oRLCW5UUZwJN5ycwHPqV6/AlUJe
SOsBMLdJb5rNUshXt+WnQOLKXPnUPf41X8P44/iqCYCLQVwO2SjCUoo/DU0WUl47OlDL+DveR1Rd
oKqdVRzv7piJFcWM4c9DnQUQlPyiFn3F6ZPc2m96H1y8OtsLNJ7qq0cYoy5DcRp+zLUgULxrF6sh
Xek060ZraziOY2dhjvUC+QbFw5GE84DGLjm2RoPapjJDmAIVF/WpmjiScbTZVWNPLSi/3xvZmfrq
8R3BKQ0Kjzoq2GhDwv+jJ3vX0pkqzSBE7zAobuVncM53S+7Touzu/78SsIcN9tdaF9KysIVvmwqb
H9NZIwON5t4T2ebKBAYLPthbpaDg6lKx/Dqv7vBVlvcEdm0b9KPx5mPK5+vevyXN4i5Nu0oAddTP
x6Zs474X9qkH6XW9aKjK09IedgGwYJUVFOddqbc7JatOa7EEU1iFgcecMFUEND+aU6gl9GQGD0X5
nDyDTo5KpnE3o+W6r35vnxjimZXMI/WAvOvUGV1tNMqVk7JDdWwCS48KeJeR3eXGJRpFQjUGG/UD
mXnb0udq3/aGrCh5cxIVHAv0n8+AnKOtKYdrZ3bkkzYcbIpaBHe49C2c0v0tkKpvNdiKGc9grDm7
4p8ZzPUNKLiEKEOsKmAJ4Fb7A5MYL2Y1d+FA6ooFveH42JUapf5MKBZUnRFbF47hUTGGQUqpHxX7
2LATcoq9+ZyrlnqQlkP/cQsOb6ME0c3nfcWr/B0AvdTG/pN1eGvKJPt4H5hoqlDt1C5AP0/rDOnw
RWJeX32n+qKy9+Ing5LagMxFHYyrf5IwycsLjoNb/k6mVi/oOoo+zmlGBhnqia7ZtKitHwISzUNg
U2lbzWVjmx5g+VRVUrgj5ty2rniw4tQ1f4dVjzezfHq3/+OMxAZOxIyrVLxVCqZAwB/CSkkx8KqY
j8C8dAFOHBlh/XMVoYMCPZq508m92x+StSacc/NTLDrZ/kYi+vLJ174VYMjVu4WZUbJWUQ0oSHca
++1lim01c+P1T/IfVVVoxBLIc0ztdvgRjOD8u3D8GmT9A1ATpe/FlRWLbfzNHe8ZVXlJxs/jJTkl
SiVRXFvFUJeGDq/BEbvY1qO0nFLPKc3Je283NLXZQjogg4M337O5Yv+4dTShd5KSIMaPipxDNRs8
s8FrkPVzU85tNIba52z+LtmInFxQwb86cAQ2DFAg1fcKDDi4TBNZX7S5A1z3udlUf7yHhNYPCbnM
s9cZBYpn26s4WPitF7par9FEGDyG9DZFOph6YHEkY8sF/vultr8+mKwCVIKCpv6f+FwBMoR7+GIY
AP90vfmx24JG0/mIsckbgt0ReO+wre/mjnkaA8ke7GJjCXvGJWlRUvmjaoSzLWKkIjYyTLFkRQjh
VM0hfAkyep3PhnRnxvusQoCJq4k7IyzpwTuJoyTE/EMzzBCXM2aTDmaeBxw9t5moN9uE6Cz5Asdd
aKnk0BLZ2TJUnnANeIVvILmYaxX4VhXde2zt/8YCKJsaUxhzQlW6WsAnT8G1o6atwQAvrcSgzr/W
z+sf3XjI1ik0Jn8yMN+WLhlJ0OoDgHLkIcHEfHJQ7sm8YxsyWLxZa+Tf0USNW6J51Zxxuu2vr2Gk
WYs4ygKBcDfX4GUdX4uztZnFROK0SI/FLha5hH8xCtNn18n8khKl/VOIfA+Zy0eBD5CSQVK6sotp
OB/eE5LDKWuzNWkpJgoIE2G4pCNKAC+GznI7FtVb99xjqH6sbGGVnYtGS0usRif2qJPWHISg7Iud
M2qGUAmaqXmgj1OmpLg5IdWpNC3Y+zl92wakMubwX8wGgGl+iuyMA3RHKarqdRUNvvsdwjBR1yil
0sLgSlH5PMgtCH3Fp/JqI0f2Egj37jw8GCHy89eKhiH+VNkVo6cyitAuhN0J6PyIcoWd/GQ72o/8
WHrR5ml5Qs4uv/PZShEqfl9pjxlTEMwUIe+r3HjYZm3R2IltJYspf4MdJ40bHoExOjA+9zVZ6weK
AH6pMkK4cbX3e2zQs+WadBEhFmOx9gZMU1PoKAtECdz9bF3kB3qWiQ5VhjQXCBlDB0EiqF2MIPaI
CkKk5RnrUywS5WFjD8tYbkl7eXajVTkUeIfIRbPaxuMMpj0zfFg/Cx/gjnD8rWerCk7wD1CcP4nv
te3ElhCXu28hUkk0/wXglNGPqZvfsTSkgfuTJj7BMihqgLNuxmUnbrrVEZpOR0gVtCMICvLMp7Dh
94nPQgCqr1WCvlQSBdKurYNtI8+G46W61GTHmINGA9KU4fS4WJtCgHFEYIkgTiwogLMwen5G6rNr
zRSd3u+xrtgM4G1mNWQqY8ionvRcnvNYVdqIvJ/f6tNq9YEOIXFM4Yk8J3du88W9AegVPVAXI6Ng
KciQmjKseaRLZ8KCXkSYeIK2Vug0ZdKZTX82hXMXi3FK7s0IHMXrupW8hRSiUZcFAri8pv1ZEUWO
AfZKmh4gyNdITC/SBUotZgi4QQ9kwkIEg9AjF2qYzn3r2GkySUThVELfrn5S4PSJst0xVhbiaaqp
PdJaVzH+lGDojjhvOXIcvUJ3Iln6O8sohDs4kX1MwZgvbiuXE56jRiFaLEAiQ3rRVgpJSmqH76s4
9nQN3svh5MR5Pho7zwk8SUyZa2kKrXOgdOAQ+Tk1dpubApmVEtRcl0bPxbltVAdW1JDKoiiduIif
jmurpF6fkl+APHlHSzJyg9JtgWPvoL0H1GuU+Y3s8mh8wE9v6dM1YoKeQFvoj5q2i0YwW3MzGacH
xQzf1VCA/PnTvrT3jH6bKsiplKS38ysR29AId8mStH6MOlbDIA2etI3Fm8ErFf4309TUq7q8XSeM
lwWEobghd+b/dVs+o7KUYLc/53rwZZ2szRa96JvvjqdjjY7i/we9BjOA8lHhrwNweNSu9ljmA1DZ
1trRJjdHzMP1W1uNqU/YINcGBepFUxUby91nzF9TqoaX2kdvow8HsrrOjCYQq7ukcwe+CB4+giJ2
BMaWT0lGMrldX8hYfxiKFtjZow4BoK/6Rn/qlW+uLKkq0THWmI0HfmXadGef/qpDjC9UV9+PKIVx
aZpEYwgArDWzWclQi+20JL0hwX+Xhi/UGi1H9GCDMwi30LkgqQNetGmiRKetDFcGfF+4AH1UaUSo
2JSEwmkvu0U1mwUjT3cx7LZDgySWC6OTCbqG21Cvbrve2uWkTD6cOqo5gjbeeDHDMhuhKMJ4VNwF
UCzBf+81VhR1oZyimmaG5RNxLiX1ExnQUu0VC5QsIEErFHoGuyVpYZnFhce2QB5bqaD5u+ayOELS
2Cm0107eRDGeqwWzUzZ4FwnUgyBYwmBnln45fF34kfoqfaclG+fDXGbEH1jNzFOzyLShFHQy1Omk
shhLbWI0ZQI5Y4wKhx+/VnslhLOlBFUZcppZPmzRzBoIswZbuTEguYjaNW7VtlrJvR6o5/epyQzH
8xWqEexJjZalL5jtcDiADPxDszrroppG6q40qzlctSXS1iPHmNNTvms/1U9VTUAhCZw/V1S3OCW5
eEV0VCnvxpKLin3FrCLaa+OLHrBrq+Cx1+E94qU6YgMYhmEkC1k+2At6QAs6FhJFjXiA7cAXQ7er
7STONPAzbH/frFQ84lN4NkrQOlFB7XKogGHxpdRYIcW+B9u1QA3mGsfo4q5rTYAj5WqiOeYH435S
QQHbnMeDHZx+LTW9katHkeAXxB0M7juROC1qrMQY5855pt1x7vbmo13QXHRoxjTAhwh2UdwXWgfD
3zusRkeJk/JdDIziNDKKPp52F5uNYGDnGSmCE9fV4AYQNG5bcw+2ceE8XByuqVlbBz6Wisv12ZSg
FGW9CETTuOjlIaiGSeRVvmIdF988me5XWOMmiFrW8ep/FbS2AeQRbbZb567d+gcgMwPYFtsmfaZT
tW9yhPPyQVbPrxw0t8hrBy7tHmFrOf61hWjYQ027wGtEujU3I21gWGP6rjpKqst3luHlcqwuXUca
2jghBwRE3rsnoDtYwUZMyPTaIv3ikCuurO4eSShPWYQToiWGqjwaqPfJLu0Jhf+/Y97GO6yXak+S
F4ORKq6HUHpAHxPUxH5lK3NbrqbLej/Rg0L9Almf+rZW7w17Q/QiuI1MHMH9r/GwOiGQ77daVUMA
sm40fSsk1J/b4WFeA/jeK/3GXjd7XbRzYO5CqrnAdjRbVA0+96d1tT1OX+Ra+gjiuf4KzihXV7hB
sK/i3fpRubNFdU9sPSutXhEZh6bZYaF6vjCaqaJoQMCA+lxMQzUAmkguaZ7dd/iHBBoP7Vihxnqr
nkfU8iR8+Dt80EjmOgC5bYP0sSj5nC3x6fjbkqhJMMIh9iJWLBCT+6iqv6bJFpMFMkY7TjQaSccp
LlNxT9W2nqI/3YwY6ncWmDaB49sy9XrQEBorp0dbrvoLN6xoa6bZGWvQjKsxVEH5XjVRe/PjK7s5
JP8zqkGSlUEIap3PjY8x/zMLf92v/jNgfF4ZdLyeNhInySZjvc3GilbOW22+CcH0viYH9S02mluR
Bbz1QmO1chZoYaNUpU4iwy3wa2ZCBPzFBGNnK1fCK8t4IbMEus8sraBMvovx2LECUTWJq2caY7zm
T01R0T/Kuhvk8CSZiRZyn3zk6twK8Lrsh2IJfB1ATwzP4XHwdNYEulf0mmyRo0JOIykuaZuDlxoq
05h9hhMEaIroM4jAcdoBFgUW/gX08o2kQK4IfI4fksIDgEwOy0m3yahn/76sI3FfzgeYudQknTQ3
d3cBms3NGc9wm5bwIRSeTztMD/h82Ia44CucX4NyJr1kZGyR7eumFc8cma8yjZ+C1JyRMJtjbCtx
VuiJRGVtszKSzv8Y7de3AAkCl24hg48uYRVWIrWke86CtX9LCnD+5tF1ktOq+deNODQgbxxV9I+q
xjpccCC6MPcgd1+TxS7pItDyCpkAUe/mOQWSPCyf1cgiv1hkBxH4vNiQaXztxNOOfQWZsdYlo/cD
Jw4Vf+kiuxSrD9xTdApt7VITdlaXAxB4npC70q8FkEcr0siAPrnretIbtDCBnnOjwCusB+FvsPwD
xHNKCrcu/IL7zWumL/woIN4T7GQnFwGKy5vt3zSIZ79WUHijaozhK7nCZ2xnnX8EF+e80EdX3V7M
zyJ3jOeihpcbcLkAzNB8LWdhrnhZmg9n7it1r3eSfcIGcJILFW91pX/k+3+ysCSGqH5z0Eq+ThDe
AoRyGTeS8SSxeV+BdhhumERSv+FFUxvosCcZtwsPQtKJCAzcdDkBiNPXhs8ZrnvG0Ve6xLiQ6hQ6
522/SJYQcFCMEPyR2VfcIXdHM8Tuf2UXrTzt2wnFo+MIcs1fa0yrk5v4KuzFo34vnTiXNCMAkVlF
mI/iCEj8M2hxawqbVG86H3OpqXMo6XbYkKPQM0Dl2TU2fjjVS1Hcp3Ja/YyZ2C8+KEmiOehnV2jR
M1501ykYyIfnZqsRFZewzGRGTu+s/c0xwt3LxQ0AugMHeVhzp2EBiR2+TUl4Ht9/vB6OBL4FKaBY
+xT1AqnJRx2pYUU6LSh8dDLiqt/ay/ZTDiuYxzsBalNes8ex1e0cq8mFxfFkaOjNukqlfEFCKUNP
hS7COLDbYxbWPvaO00BbSKPuaciDPXpieekaql4AeitUH9v3T3V2MO+XEbkHaAMpXgnrn7ODU65o
tNgBSXfLTTLNWeFcI2ALvlTQ4IsaISYgg2iFqdqAwbgs9lfqSXhOXIoZDfLbocfZXwt7UHA+xm11
Xz9f4xH3ODsuvTE9ZLGn8gUNYGyi++MWtrpGOO1RLYAuh5DudiNwZ0hzci8900uyfA7cyxSJ2+iU
W+snfbI/KzKiHnJQp5wYAvXCdJlYqQiOKvH366PFhbdDDr2xg8vaVwDdzRbaQcVoudDBXm1GwGm4
PJLqTBtdPgR0ZXLItoWKEquH9cJgDyz++tbMCKkXOu5YkP4kgVCvUadrBgn3lpG2pR1ozmKIoX7t
QQMHQiuKNL7GvZmavhgDvMgM/nw3MxcsJ+WbPYS/ATw9KTVvOUx6KeAWdv8DtvwoNmzorhJCgMEN
IFi6lY3/YrjGV3zggujOAh6SF69oKyrFEXvpf9msBDvRR+J6G8Ha7G2mh8m2b24Tru1AOtATsLmR
ZaE/xGh7gTduQ3ecHNxnj06FMlVEnbHNjeRwf+fUi1TjVd0MvK1n6u3jzNwrPpCM3bVSMAP5N7m8
lABOwIcobJAZjgWK5/6CIMQLB9Yye55Oq3zxPfRGv0Kf1PlX7sOllW+oCt2r06PVVKZNMb5Vw6hT
WZAt13lIO06e4Qdoy06lHk8mQJFnvrnh2TzIheC0ziu/iWASpvlPkIofZYmEH2UvCvsawipPQYC7
nQvgUxNTczwFmjsN3SgSbGCANM1KjvPGzD2D2bCjr0FuPLJyN46QN31GbuAl84uXjruTS374uSkW
rmPa0kcP/upzkW6A9P1+jP5s3VeWz3nLHmjml/QLEeh4ieAcdLdMiFccdideZAWBP+YwgGWE5N26
PY71RDWEaKRzeIVfNEg6MSoAJU1T/Xb+0hP5FzRpvyUUUij6jj2W74pixNhLAyXfvscfg+NdfCYd
zzpi4DIxN99uWKvS3URF1mjJKIP9yCeysoj0iiaj5r5CC8G2qkyorRIzP1B+kMqPB72c9b0vQFpw
7Qq4xOCKb6qsgs0LTprj/K6xhVkNBX+dflO6gD5th9s8HCxDt411OvsP9e8qUZs79Ij5tcRXFneK
dcXfra5upyUC1V2lzHA5Dt388l/sHcKklhnCEVpaybp78d2xdufOH2wnPOqWB3X+4qW19ZSYNMyj
C9qTjzcm6OA7Dz2JApCjnkqfGtvLPaWif3BtL6OqRUHb0nbvtISjuvKTwqro3JKpiFZo9Hvn/uuO
4JiQ1kHGVfVfv7IAzLoVGRhKAZE8A/ElLk2CgyhiiePEjOotL031NQYz7/R8Tu+TiyhmajiqdR/0
jEO56D0ohjgd4p3vFnPF2qjG2IsO+XJH7K2L2Ixo5vJMSzngsVGjTs3QQF7jfGCMPLBs8TB13GL4
ur/qfMc/BhGhCgIPyVNN59pJCLLxwbQUMKZ/l8spvc74+DUjXP2UnoQLOD7BfFt2jkARUj6G8s/n
JcJzBuiUAJzvYtiwrCI0CAV2S9Aj+IBrqfL0s0GsIULWe9aFe/JL8hBf3bbLgvdoW0eJC7AiA0tV
Y9XcOXtjSz5yQtU7Nhhmo/YU6KRv1uF6XH6NCQHambq7csSVzWrKvRHifhg5R3BTTh7ZmIsJs1+8
kw1k32sTd8Lbt5WONC3Ds76hipfwB+U1Qo/qd65p0cvPuFTd7quOWs1dzCZsKkuHSheHFdHVn5SL
hFkRoJCdlWGaJ/Llq0FKhZ0lIdBgJVguIYl63PY299jne8o3ugFTOHQJJbxSstyG4zbqRu1KS60z
GBQ1jxrAGkSFX65OdBG+a0cJWgPvY13xQ5hyq/mPncSDhDpYH5bZjX6pUOL/cLXSlrQU5FnOlzfT
7WO9v+82uDmrEr1z7lsMgJo3aBiVs8zCLvqHhB5ZpbcbOYfVRkb5WiF7gYbmbopJGszTsHJDC39E
PKzwgIQT+IpS9npK/OsUGLHTKZtprBi28wmDgiDiHkd7tBPpbC5lermciSizqGM6yNRspMxJVhDN
6N0oWWWoWJjjr5ryipPV4shgj3OH/KAAnF/EHM33OBmdvEKA2zAntXttSVio+sKtcNLBHCFMd6Iz
hl4TWQZRg4XitceFWcB6y3pPI9I4jg0TPWeiuGgEhzG+LiRv31qKL9rEHjYj2YrtzenujWQWDEsc
Q2GOVKelN/t7JIXz4+L9ol1cqHzflm+f84eXe+ryhlUxR7VdwTunxwoQTl4enVRJetVy6oIMGKcg
buIMXfkQBwErdNv+KHcEsYTWCIwZ/j8tdOqgTapzRNDJ0p3vLOQlR028/K8tDsEmadEBSbsMa/4/
K98bsTFgmfvV0LeY690QuT75qPrnQnlLiYwsqFVSqdc1galvHrxu08l9KWNA9bc11XqWgFWy5KkU
fYn4/PvwcMCtVv0eAKSRzXXVy2SoG8OIgLyIuYi4CjzgRQ2NB6tsukHEYPfDj+op/keGy83Igzhq
EuFoE2351Lg0PARJYDsNsOV3lePaqnHvQZaaepfVxU4ycLyjJUFuQaY9QbmwMKd8oUmX3JxBmimd
Onc/HXKM5gDVGG82bWMfwxBr5+3nWNApn/gaYWXdRpti2qcvK2CfdRMP5wpkznfFH1MIcw30wSnL
U81aWOIfonO43MmXqPRbWSDc15F/XPYq47kW7jhgH5ENaBSwfDkupBSzcZhGm1MC0Ytk8Yj3zT1V
mmZ/R3qVIYan9Nk8Hs5z38HfuD648u9eohqOuyB3e7dayEyXQz/HrvSs0sj6X1/IggLa0cTz7AqP
fMQ+vmKtrp1jyUNXgg2nTuYllptbp8UYhlerVn1PZ/ng3LwdIijUJ0udWduK/ciUeDbqsvUHynSJ
MyreuUdh5cdxfWc0Yp6o/zU/ymxTs9wqmhmOrxSYa4yygYBUC836AfAMg/nlebUi9l+mS/8a37/F
zgom0pBoxsnH73jLun+UebKYyS/F20VjCosdHhM8oZBCDtcIOdjIzo+TuYvAL2Wy58m0d1p1Gd8j
w8D8ROtLSmxjyRaLvkdAUgjIBHBz36dry8ZBEsnu9bvHaG9Satt49b/f8lmN85fjoNHLRb1/TUQx
LFKMZM9XCK4ADxB5dUz7Z9mNd6ks34Flvx55PMnHbnbA2n9we2U28HA9K1pUf6Dq4pFs7SdmpgKz
1hgZW8RkpWFeMi5ohnn34qRDncsdY5J6O3lL1NSw1EzLcCA/+6VriNvcjUEqlE/JpLLSlPMWCTQE
NQoPtB2kSAWT0M0bXwwe7to5dgjSc+xlV1dHzWwoJyzhDfDpzrA2xQ9NlJKRyOH7t+dvzwe8JKqc
SqbtOlJpIomPyAonBvbgnO55KE3B1JFKRPgw5Jki5EGRu6QVMo0IQSjhetwBnYJUgl6yWrfiC4ag
dLQM6X/hSdjolqPs6mhxhK6cbcoiGEAvJJ5O/pLVjaaeI2O64I9T/ybSQkZCs8kPMto3yIykIkG/
fBn6XKu00r30ZLDNxXwDmHGDVo98/Q8st9mUT1rXJxJ7z934s+QU4+i5utnMQCrZn2NbOxeXRupN
p14fzx8CY978+e4dbJYJuID7hzJuo2gwS/GUOGmaRFOlIPaG7NOTMpkBBJxbJsCFW9FLgwh1IWSB
beQwQnxQ8inexhkWSUqH0rtN2/2W9r2K8ksK18Lqd9VpaTh+/YhvfJ+rPFJA3pNstQLOaZS0LLBr
vLSjPHP9ygqrNDtLZs28e9ETK++1XtpigBUgSFgf7a3KTYEhogPEAa3r0VEX8gJs3Y/0BAnSpE1i
zeoS81U0aTehxe2dEr39jHItnHo3g/oEw6mQ0q0QX3IlDtze+E0m0qaNYNndxz76cyovYUvoXzNz
yv3vh2TZy9VShFyI+6cDhm2OtHVT2Pp5Z9ooTJITs4ODgjsWUK2R2ypDVNDsWTIKvorgkERWCghU
fvA6xJpt3+pTz8qRM49ANYB5rek/Gjn9V2OAu7odBI8BXguCE9RPUQ2fy7TnwvnGIRrdWhO8jtNU
ex1ihPLs6wFQV2ouUQ4lhXCY4hxgcqs1UTn9gyuZ5gEW8kxCNePTxLDhIFnHLxYEm5Rsd/9A/3ZA
S0gDYhZo9bzzJs98hNTNQ4JdFiq9+mOCoLPYEpEUiwCLc2IRsFFPT7YbpuTN36YRDkjW63DvC+9u
G5KOkjrCGu+PgZ35REEsTE8MIhXdCmY3t6aRFUMGNDK1atiX5MToIwmIAvJb2WL4Wb5yPWC4QrH1
mpu2I9mhY6uQ6qZV33ugLjkMdzP3GMMKPE5VG2PhGQfoWScr2hWabQjJ9ZrknP6k7/Q9v/6qdlOk
QHZmFY01sJ8+MQF8589u0umecALU2GxwgKzf/WVPPBGh2Jz8bHJ4TJYTuGYD8vsVfRQxnagJrPmE
FopX8Z6d6YqBOp8NGg7+eKjigNDZUX8bZY96tMSigtMs57u/PAnMA1iPiOgs3Nlx4zirp8cJxWdP
LitPHkkhLumtselozTUv/9TpwjwNCWEaoXd1t876SAi5RB69+gH+CQjLqbDTIDKKK0OnzpPs2a15
88UM2BrMy4M5cD64fWvhKtfOE5vxkv9nrJdTBsfuCsFDMhqAtS5ma011mPi3BD85b8FZZpxv6EG3
TmmdEGjMH1JA+l8Yhy9rGdznJqx+zQ5Ob1aQWEn4U6vIVv+3LQ9w3elZKNxrnM0kvSdJOmrETdyX
6zJ0m5Ux+2k2fg+0kbJIpcnnHiJN30mcp0YLmO/AIZrZJOF8KHVoXgQyd814Oh4JZoQ9gjrBzR0L
Klt9a/C7pYgOD+uaT+FzZIlB40wDHdHG/LN//EaNt8JPxfptICbmqehuDfuVOt78tbizRTqyGlVM
A+3jHrUz7TKRiHFuqnxVssRr7luQKiIBGBEdaH0NByQnigqv3MExzgPQlN8cD7SxrtOhB6tclza8
zv8XuuoEX6P7BqCrO/Yt7VNgIDwHH1wOmnm0EdH1YkNpmCy7U2SKGsNLq6Ps+oyTq0Lj5cWi3wiK
R7aGad2mVs3NFV1t31aR2/r+ZnaB0lrWv6mjPXS5KO4gn6qPweNfhoZ8wpWBi4L3UchAAEcU5H1b
82Az4P0zPJSbyv7ZYyvAVAtt2vKxkbXPBgHYWblVVhgAIn63CwXTQC6qFByCFzWte9bBM6HuOC1X
0oQhZA7r6r7qqmpRFkWrlLLm3ciW/Ng8hXbwEN2PpHwYpb40M86TdOf7xRnCil5LMgxejqi7BzZV
dX6EUaDZGtzgsbmvyd2Af1fOLVnXtLmpS4ZyL+o0iqjRctbrjaClVmdM7gn1UKc4vLqUpy0I/ode
sbXkDmJY79UoAm0B+59s5W2xqN5vFYV47/3rNrIGX2mwMtk/OG2DQ4yEfXPS4jy09m3h1N28Y0W2
mDNRMFTfU1xKWFH/hZxxPn+T1JMKLls1yOzpJ6It4uqe7+2RKWSim/mA4HF7ZSk3N1zhfb7ZSlF/
okC0smeO94WpN0Qv3bGUd7VMwpDL+m5QBnVa5U4lqxYT2EaoKl2uI4CS/tuLNSninBHnRbzLRyZA
oxxXYBOuz3qZznUIGjcBJQoYpi52+pExfceX301fi3+Fsv0UzaVlo7BJP0akbJnRP8P5rPAmUVc/
Lxj6HOmPg008KZDpMPuwL5+vNd4V83/JVng+/VS3Hwj1jb4e0y1VnB+nAgpt4dZPq0tGT7FW109W
B1GU4ghOrnk1VxgppoaNLPbD6FEYUUK8VpxWTV5xe4wUwpre+/SDu3QG4Ya+l3AP/GbjJlwxooj/
4JOOz6WRElFLJ7tT1sfBJzWj11MlYandl10h7d3FosnG6VjWkNpc4rvzNg58jgoRaVWgxxVf0teG
sahf0zS+vYAwCqkw9sANFxlr18A1nM8W43r8qSx0g4KZ+h7342GErGFkLckiDmKbLCo30e/JP0kU
JMWq9RueiWR+XLmG8525/36zQE0uLiQarglXOURsZDqZuqO+cwF9BgEPpDHRVzh7pYZSBKD9VK0R
VNAkL4KWZoMfnUCp01CaUVAdlfmZR/Ldg1zqwX6GcDtGUX0AlgcSpqhnJJAy8famesoqJ9VOSSbt
uBH3YuOPp8ut6cl5rNVumlt0sWzVSIxvauC1Xr8EWijasO7rt6pGbymvLhGIJrLV3+92Ml0vTwMF
JsluJUUjhjy3cT7eq/ZVz1/8WVnFlmJXzQYdoE/jwFi7vzQ+G85oE+NSYwmBzCOTkRKWIOw5iOPA
z3h6rbq0rfgwHbbSXC5XkyoxP7ODjLOPg0o205pQ6tZr40nSoAxVR7MoMPvklDXd0orEqNlGYrVT
isY8SOA5Y4y9GRrIm3m1KJE0dP+fJnGFvAeKagCx/C8gpDhgsLO8ra22iivX/yd5lTuER6RIJBtq
+Zx4R9IGRBRFBzlU/AJsffXMJ3I16vT9UlUwsORECGmTB3RtcDQRfr5GaCs39sCVUfLA2QXOItaD
pc0WIEEkfCC5tmN2IPIQQkh6Uwwdd6pQMexkNz1ba8nejjT/rVcDzXV7MYa5Vik80sNPSmbKvku1
AgAd89NQW+0+tF9YfkpA7Fwii79rGPRL4aftfnfAlm7VP+nHHf6cWndzBNRP+djp+v4WFFHg3lF8
DC9UzFl0rkrKeocYtuUYyaJ9xPJUmFkXvrrunVTwribjHLOndfVBGTzrWwnB6salv3i3umqKj611
TCaMA14rhFwYdF3xsGwnvM/1tXu9xxrWOUrOzBJ7PxTWG68j7WKHMgCVHyamTzes2LBO0YuEKYOT
MZ2XicDlmnlKQjjKbCgG3EoID7Sf9BTp5HqwpT3Ysvb0fXQxpSq3rxDgKlmXRX91Z6VEfs7oIxC6
cR+GPsUlilo8F6RH9QD8cdLdWVTGEwEY7CInMbfvtHU21qKAkV6zyo8xa/sPCc5opf/oQpE1Poj5
1uIEfTHBxr+CMa0ue1AwcnwrbxHhRa+uf7wHceAxif9J+orkW7tWzPT/Z9AOxSLnYOb1nWwLHsvl
vejO0oGQD92+zFn5Ob560sM46au1CqtEx/1rtogE+wy/IKM/IIYEIaaMZEQ6nJ2XqeM/2lfcUoib
l5RTOQRmSQjLoCe0m8VGgDZ/9Lc/4rXdJpQzMHxzqYlpLnxot3cJVa1L25PaD/T59Nq4F+g97Cjh
TJPa58XIXBTRlhwbHai+3szL2qm5Zvxt/r+pMrl745ecK/Bn3mVBSNk0umWjZmTX3w3y0lcr7dV9
zwpG0sJ+IsDrJNSNgL5090nz3SsN+GeUWy71VlusbfYo1/uCYcvwuS0RJ++02UmqZIXqFAupKdEo
AxcZVttjhYDMfE21xp6lcAqK4uUPVJgMFjlDhnMZPLr7lFI3Gn2bLg640V2yCT5w1XC9PIIFJ4Zb
m26fug7x7w2AVfSHgjNKKAU2ZF2zH3wI37Afde2ZQOiVIf6UpE/eCXrZPFb8p6r1T93l2NAwP0q7
LDXkFlu25UYVujLTGXP/NhJ8yu5xFcRrqIgnDpjzyYqzw6T4mAvlG6Ok9dXgDypbVcCOL3sR+MhP
IqgUD4G3Me+8C7xdYZ84x6OZ54jisdiLXOrwitdP1Vi1W4/bIvJLh6ZgzfY+4XZ6hcYuXOf0RfqX
5FDn8FlyQjZXXX/CKyhqiDwkhV9ZHAiSF0OzYpZw+M3ln8DdIc71uYYy9pfKCdJtwVePpkm7Ib/C
mePN/5Wlx+sfV3PcMqPxVdZcFqc52LhlxdPQ7SndrM3M+h/83KO0cMcaLHASC9Dl9U7A5KD5w8QD
+Ycg8ddillbW/7P90HYu0WT+f4XpL7+TPOC9oLJNXDD1thbjT2t5mfyM1MWDCpmE3BxRPZ9BQSRT
nxvSkpEU71P7aSoAAGv3Zom7G0+buwvvYCpulPgkLlBY5hEBRra0zVun1Uzb/y3u3IUNJK96J2xK
0f+0kg8Q147dW/ZGrmLfrrqmZBVq2WokPf4zs7UcC1VTivENo3vaTWHigqFlC9KjXLH3xBySbjeU
ECYA4oaH9TC0f9NfIGDDNBxd2Z/xbWIzNYXDvzidXjORs84kzb9LIHehXweozIwwD0gsAXt7q8Q1
Xzd7V/a2VRFOqJzqcKG8JcX5zxccZq2hLuLghpVS7gV2FokpvGXa3viL64aStxRtut4dmiWpGpfz
gmZ5mzBMHohOJHB+d0Xr74B5TOyeCFS1dfHyg1th+jV9xFrf4WrQ1XUOZisQqlpZLJpZJtvZJIRC
NQV+bJCU4BZL2tRU2VYf4T20XYmf3++60UhortI58Ho5mFHmTyyLt01R5SmzvEq5Upz8sNAz6cJl
DqCQQR1dPRe/8DoYZxoQGr3Gb+GQDPcUZdCd8gVSiInhhHNmcEo8T3v+KB9t6uJDPJoKZC9IWf/T
bCeB1qZlTgRTRjm1z6Du12PR0w/vogZ3bQtRcKD5Gh62zrIvlddVGSHXubXHNLxIxePpN0yYfRpH
roc3mtPuGzRf28f4/rdnUe11XpVNSJ6IfzmCcqbeQauzNgS0/876c8Ys1vyUM0GMrd/FNiJPgqt/
wUKYBaKfMtKaMW6kkEw/uY8oziW8OrrX0cJDhWs4Pcu6OKY8SYnkv3bjAFP2Qssr4p6IZQDHy71p
HfgE8s79q08nurzHxUxNkfzIwhkQ2IbqA93pEyySx2noo4AlBe81X0kMc3cZ59W8ArjVi5VbwVTN
ecUnxSAFpEYTxyJqbyTd6gfSguGguq0Ao1QlmOyuJTJf/4821mti4nVMxmKfSC+pcggaVqBkjGQX
iFrl23i1jo/FxBTZeEhLzKzX28bnywf63c8sy09emZEAZsHX42Qk800ktrihq6ed8aFgbNnmSHRt
X1uT3TsUZG4tmRnefkJVrkbECebbRAlCiB0ixxGLtGMs+i2Way3z41vyHQaoQMD0+tqpsQ4FCnwN
4doSmPTR/znhyeZrN50sTEVAsOL0PqkB83a357ET/DdYAM+BMw3d5b2x3HYfS2D9Uk3dp51IyzQj
o6cYnCbcyn9HGiVOrdQYXuKzSRhf+DJzV5lJaPjjO+c4+kmx8aUE86+w72i+bxNpuJeE8kPtWF1i
z0JCKhE//Iq+oBAk1k3WhseKQOrtu5cTEc7DdxVUXkWZpUjx7AlBUJ1fWF7e29eKAUHIVrPF8DMz
mSd+nDrtkHBIR69ZWH2KSxFawVZdvLdlSgdw9o91ZeUZeWOTsgNzxumcStd58CiyMD5DDYtHYD2Z
zarl279Vzs637jAKvhgcHnj38PelcyKYuF40PBQXxwvqcvd4XU903NO3N41/IYzL+LmTflH5Yu65
lYfJ7i6VpBiiBWZEudhqan6oiANbjcMVN8jsMpGAmK0QmMKfir2965WZJDCnuVeR/XtEpcvMaMun
01QhlqItJW65poJwGpZ10JfeJ3JQVYYFP1CNGPpc6Fw7PWAexTzzl/BoSl2cATbee/BMBrH2VLhE
EzJYT2L7oB9gmJKaoOOcMkBzuTzewyLO3tVnrccDJZHY13eLknmj2Sb6jN2aSjBXjRpVrNi1dhXD
qNMpD15DJ5+YIXYqOosEX55vh9tenqVYnqt9sBbvkzS3g/cG9+QlRuQwWbF2CwkKL0SF1KIuHoqJ
KPVassFgd+Rz9TbBKiq7HoaxE/OtNUwy89dux51LyJdY4XR+jxVtAOjdRNhRi+jB2fDaChRet7rx
0CxCncrJSbJ22kPRWBCHDLll/2fWEbQ1GO/XWxL4N0oFLTfADG0KtAXWqAnSBsDlkIuaVf+vX2eu
1V33PjM4a8x2w+r6F62qihAdtabinpG7bv7quP5wdk06eVjijmrYfIHk0xS1spXJd0OHx/pkxbBt
t0a1gUSunD4UAK/JHlcsCPgLIceDQCjCN9w9BSeRMMSpZ2P9ISDBo3sx/4rYjKctnoWLT0whJAIH
JytV84XxTXJ1Yw+lVSd00L7SeBZfS9zECVTolXYV7mdwPh+Zqff03sVrVD4X52hD94+Q1Y9fgi1/
zOCjm3QkwStHyIgaBnUteFNbacGhQdEhq+mNZafvoVVDnoWvbNhmXYqFu3q2X5SBIz1gR4dIyl+s
567SI+YWtOux6zcDBvDE5adCx1xE8V+f6C/Gv/qA3wX1qxY7c2NauPKTTA/CSXOK0wzheUFfv280
0GZb5ZRJ54plMFP5GkbDy62EbLHLBbNpoOmk9q9y/AxpZntnL0WX9uwzblkvf6eS/Vt2CxvTiRhc
jvsVTI4PIUS6tbsIHNHcZnP2fc/QYQB3yC56Ic38FMq8eBhrzy9EMk+LwJ0gt9PnSDwWJmWl2l7W
VNww8BU/x8peSLVqMZ0sN/O3iwxTfDQUaFiNFZeobZuxUWQlS7fXm2vzH7GcucNWbxpos/7P5nE+
EkDF/ujOUmG49W5yFxtvkmLCBpQne9k/YXMIiRQibcMqUTzJ+eavZEWntfixVgJxt9y4miPk8/sV
evT8OaAjn3CDWA5bpFENjHrDwqi/A1jmFhQv0/pdmD8KycTWQbZ0WdXsoCgutTd06WVVyRkWpAn5
GcoR7c/Uj5e83N+qhmFt9aBiF3uz0fUvOd9VeJRrWOq3jjhZHz/3EQRnZGDN1RGanZ24BzGZVMgH
kkkjayWFvmXTeViXCbI+1s2S1PJUJW1e9Hs1W4e36Rl7mCs2Rwd4PBSP5YY92QIlnmiaJUHzkeY8
WzCfy/0frRSCdqsVXHLdwJ/4BNLoBJFJsc6Ps2KQyCKB9J4VJAYiVcdE3GLjIo0c4Qm8JbOonUkr
ue0vBSD0j1yduV6cFSNU0WV2eVMtkN6kSiEQeeHQoO3luwBCSccQPZ1xstzBG8f/Wo3OYocosEbz
HvHJc3IWyo5Ak3BiJcerAWawzV9r3BMudH/t1vxQS4vmZO/0Ehb8U0zJRe4QYTPROIxjRLP9UarB
oa+o9dFmhT6yvRh2SDcJDv5XXqSR4o4WkODVWCFRDRYobQ1QjAPxuSF06f6gZ7+9NryjZ3PEcJLx
tL9NOAZLyMVfQbD3eYq502fxlojQ5VgsP7Eb9Oxt7UbAASB4MUr5Y/MiEGXnj88qA0qL4Ff1tCj4
xJr96gFwk+VjfxIKGBf2pCv+cOz9Zp1ikM+gMBurzD+dTgzt1mSeKwAL0U8Cu0VIZGlFdqpcqXIe
Shv+Bo8y+MJxTnqqvDYwKxzt+jybdEB1i5jE0R8460FXJYvi0GOq+7ZcOq75xoLXxBVn6iEF47Um
tpMNOejQDS7SF9d5CuF2CLOnWXbVFWwo9hArSm6a+GY7pY8KE6oRn/PE5iutMwfZYZ8xq4N/+HGN
4OBedV3caz/ARW51GopLopecE/zEYN29ohHmNGA6+eM4cOgzgQSXwTJy5b8G4+9RUZO+jerfpDrS
ItD0U7g/JiEg3mac5cYq7cD6TTQ2TLyg1jOxn+5ALVVAgNhQJIIU3JWI/Sk44qGGvRLs4KolXHfE
2QXH3fadUaKMvD7Ktgsa6NEeFS8u6hwQcE4pxVHP21QJcHTZimVPE5GRelAuc7sNBo+j46hMDAN9
gVTFqG9fI422cqX5AUCmL3L9PgRJh4rFZbp6Dvk2ntOoCsNcsIwF4Kestf7dCUitIGs6Puht0PT9
EJbLEbo2UuIXVqVmO4bk4i41G2O1plqjeuVgqCyLR3mgAmnYFQq2BTHm00ThaF7FxR0uCZSLoKCa
tOoVOcdqXLZlfFhrSmVQSiV4sXxK41YaBSESlKQ7yvvtuTExtzDhWBsV9MSWrP9XA8b7rUydnSEx
9worGiri/RpwK85GGZy2uOf0Puez2623Uxr3pmPgk5qLGQE0i+AqUnxrQfnIesFROAMZDByawClu
srBqj5xUP7Hy1IKYeNDWV2BnlyUVI4ESUR8pZAB6WQ1bhfQKFYreSekXWThcQbFW76hGGpTBORZI
oXNDPxxuLJpMpRSTe/22d5E7urjXEAEuCM7iO6Ctum/Gf2J4lU9YV6uiDralDR+izUVh/AqB07jw
pXibBPsLq7qjmi9AsmAhzS34EHN8x/pGSTtvJGoxX4dov6TgUq9M8BiYILnl/W9crJuHHmmD6PfJ
dUSJNS+dNVNYigJYkON/NLcfQ8y7KEnBX5/wIk+CencOPwODeSyCMNxQdxYjMZr1Of1wjtwsxWlz
HFeukVej0zJSPWDwSt3gTzUtqxe2/SBPdN1wZLkbLleDtMZIHA+ZbBNZE22FKtcPZcDz8U8xWzzJ
Tktv6LuvMRbfUYEu4tmIL39NwWSyFI7168HJS0NUtM8p3f7SrfWrMzxFSggNwwfWxMX91KQr/sii
SovQzIZ5qjoJ3eyXjue+LBxI5f6JAwzK4pMNqMHb9fEGpy9YtfUAlDDv6jRAe1s/YuqeJM8jFRfG
RD24Fb586viQaPGwaTBXKN7ZJ95CnbRlJ3Xiv7hVdNt6GweLXOiQBrYzD1dWJEBirCfRGWtQrVhp
JfK7vj6inEFySE6BHSbW+0Q6yas9ON6SJaSpBQlJdxB+GvB9mRIScYKjocBxTgBoX9P2wbLTaFjU
63Vt48PlnJZLXs1bEq2JNvv+GTYd8ivUJNKns6M4P21ycp2lk+OXiOyrTRzT34BD5cdSo4ULeir8
75RgPjx209z4dHGCsbkVC09j+3bkFvoc1T2T9WqD2vhtTNZkJf36W1EDyog7WoyKlt/oHS8rD1Lo
HlVf1+Q8X2DebQ9zPwERvPX4qFpngPtj73DUz9XcW9H4jXTpfkNFlxyFEmDNz1BlsZmUwvgxIuxi
Nlp6wqg2Y0Hv2IHOe2SUjpahhUtjG9oxxiC4xQiPvQZ5kOTZEbMEkdXSMvBjeZ6UHh0iNJl/Dfsa
uouzra48ossLt9IQtk2UC2ZlC+tnBeSrM07B/xnx30dmVS2owM4Jqz1jzclyeFCt/5wTERZABBO7
CLMxI2BCuPPoxEDpP3LO2B+v9QgbMUr0Iv0RO0IQdP92FmITvvgWsTf2HvHBAp19L4CoJEzDEr7U
EXElK+PzKkP5JfpUINeUiIPkh6Pc4h4P2lLojJgL4icwOSUQOnnlz69YluYoOBRoKb6uJ6cX/2GA
nkUE05uJHe+1iR/pDYMuUE7VF5QyW3FCkYsss8gXU+vVppms+k46SjCWgCN8jA2SA0hX8TG2RVa7
FrKDxtf+1U0mI7zzVMqyO9SNf0xfFKAlHgtbyCur8Df7L5H3Pfv/PTg+zE4Gnje5R10Zp27gNtOj
Ls63M/fripQLFPI+25+FrauvcLXmyGwFGIYBWAl2ijRmjBcehw3++nNdXH5Lj//1OAdD9dWNtK81
lJxCZgz/IzccYg+HdIsseRxpZHI9s8lM5Gvjbm6QvwHC47n4feksllzj0w0z6XPws57fjg+Geqw3
iLnVF+0zhRxQBeDi8V9uVPxBlq/6OJptkdv5Umos7ZIF015hBO7IYEiGdOMuN7bjeLj2jLt5QdOm
cJbCBqy5DBkeUXJVtFzC2h5QtM12Yf+ZR8f1dYV3XjzFDGIcfvwibSmJMX5dEwKpfZh6tV6SS9lp
QGateiaAgaIv+rZqG+gFus2i0vTu2c3O1hlY5OEgWMy+qXmVuqJDbfv+dYyaWwJMnKIOUMpr+Ykm
F9QSbWxpIB4XOboyS9py4nFdIzbYRBfGeP3+dMUFkdIYVfMaGSAk0NX8LHI0dTXoy2l7S2+2Bb4D
KMCxMCPxylK3otcEyC1+o5rZOAyj2+xsb4HUhJYQjR7vvZbDeit957zyVUtbTM+Xan2sa66Hz9qv
TLlS26KGPGMCytOG49vbx6+r/TuPe/Bttai7PUCNVQsl52eJSvLe2Kohim6T9pBBTF9/H1k6wD03
L1pogcsMo/1tWn+chInxSvd60RI6YdQKJy9hsnltKkl9skyXlaA4QQ/iiKADvxrX14AkQsK5jq5M
LtLf3Doxr/GwQb+hOIIbCKyGSrx/b/IWMkPVZF2R3+fCkQcd0NhiGG3y1oaiGqaXaahtIJSd5WJY
67bbW0LLLqc6vppW9IELN35ij0buN1EU1D55Bw8yfoYxBcN1xbc1L/nPVrwVlfl+GjIXSW1REUmp
c/LaeJdSxtEDGU7qVFAMR830Ip8IqUhJOVCjO+rVZtrCUeMbRR0mGAPR7+hmJjgowaECYRNdXz+z
hEPvmbzxkwvbXKJWGX8WzmRxRoT5rH/fjbLYtMqb3T7xrwLipwfaW+X+eFQDMijmuEmcqpJwWnCQ
ZXCTgTbLLwyLPLHxmZjyhvfC0NlqeeAtGYRjhhAymY78BOUbe3s79O+leMf1FLhvP4JY6h5h4GSE
u09Aoly1FHslf5fCe5HMI/EBmHfkBzuDEBTFYjllHHNXoQLVuQUNURbxlNssdnQebR1F+0e+7VPA
qTJIoPngVeNwIsEgxNR6h42rGzqeJp0BafbZvJQmDPDpRlzzk2hvEvjOH6pw40Pm5mS6CRHZxDgM
vG20FH2UBGXhw6dQKt5ZpoiJoxoyKiBIrGBqgoNcSIlL7xRsxPR8PCcKqOlMql969zPsrmSSu9wc
pXa6egTt1luyX4p/qepf6ezBqnqP90jZVZ2JOoinsfjq59VsOXVD4CADBCOEf4s4VX5/LNTL7pBZ
9L51v+E0ih1mG+N1xTlKs6qdasMRHd6f4L8bzRTBV7M/44KyJpLOfqzmgXg8W5kyRMgbGmBoSNff
Y78GG75bZ0PcstVzVUYdT3jG1Xp1Gswi67Z1PzBJ+vMYVkojJZ3Sc6c0mitUUABcFmDRKgFg55+M
iSgJCvJ4uhd4vJvM9xHt6cSVUiBQXRd5vPOvPtb/yrBOzsTIdQ2Lm0QopEAhkFpBpuLGf7+SYWQn
yE0budjotJhhP/Z+Bob6tSsNgY4P8M8HiZULPoraryoe9A3J6HCCROVqdtSfybjzmfPb2DqRK/qk
YAZnNLywCr2W9IqGtFSPk8K3Ri8x6nuu3feAsfaV2KhW+hGl+TyVLpYSp2rSQ74jkNqpOAN3GLNv
og9yUOCA1MZEQjs70Q/iJICNQl9/JHTWnNQKHhoC9YqeNbNoNgW9xG32tBR/vsxJ3hAVHElf7uSP
7N+BbvoHAzgPAzV6puMeCRGblfH+O9p9v/t2E8eTLfs4HrKK7PYDgBGPRzJZUKfm9IhlAHB1TWVe
D91afHUXbH2+P8wVgEWdbDXcT1sDs/u6RZLi9tkBwXoIZqvrRVIXekkQfERpSpGsA4OVWRvubshZ
jnFU5rLCBYCmbTAlxbJ2ibPArPNjiip48GtCXngYYe+z+J/hNNKHwNNUnaL3pomFzk1dFuxrZpBV
WrjTqnfJr5wdAy8VEVmENDK4m0DSHkA6oqYRnZGmTjEPsLVrSxjMJexVAKLO6ggFs5I6Bcd6GbPn
vEb++vu2nZGvcXSe8r6QXPIyke9XwyygOPTu+IhgaZG8U0xTcbTW/FdG3kYODe3+V5I8yYqxVagD
BE5D9AW1LM6tgsLUvj8Po+q5OqjAPQkcVKvPiqnJ3hqt8W37ajzPf2G1OgHmMImWiwMRI8feIz7y
XWfNlsi37ptQIqjKi2Brz44T8lEtE33vaRYhbvf7Yk8A+gdxi2gffgeScWf8JjjBirQ+xeEt9RjP
5qaNNnHm2U9oEnw2F/7AWF212PxS/TcMmB3XOqDJCZ6TnMrOhE7YDmTUPps4LLqp0GXrabnPJxpi
pOce1k+hb14A9BtZqzpLxgbFpQZkc47lMtuMW6N9KKp5aHSP6ctdZ1sBjiTQstctqZ2bf6x1eoCy
7LSKAHSGeq+E58Wx8QGnF0iqy2QeM7XRxK8b+4kcQ4Mb/B/gxrDjd3xaOaYSVt1XdCDaLs7gZstF
aowCJ1hKRcqwt0aBLsqHVGM/nzKgYjKEdjfU0Yv2X+nQVEn3Q95AFJYULT3CY7cltgBD/Bk6PJTg
UvH7hTXU7QKVNyMfMZG39udNqwVKLJ+iXn+MCDtSGDlFRXeHUUQIEx407iUNqYQL4rI5fzJ3bI0E
lNRFqBWkauR9FWDfIXiKIjjPjsRmuirCCD0ghpQpjnK7tmBS5FWSfXkXMocEJPvRTt0rS4I32d8X
QKCTmfYtkQE26zbiWa5OO99DGn8iWg6C5JGdAEm4aDd2wq1NbzEuETzdjY/ar8qcTUZGnQDIrGh8
xjsuI+0PcikQlrCDoqZw/rsBGYK/HSW0iZzRTVGXYIoTRYkmOs4wCAWg/fPSyGJTw51NYua+J7g+
qIwAjikf8RI4NEyxOItEVmUN4GT6Clw8ofqK4QARc9g3wiIXpPUfgCo1bL1daDPRCksIDvV6VQal
93PxkG7Xp7akFmYq/ybHrLEhCkxaz1cZy6SeHueINt/ohDBl3q1AtA0YeaGQGIrDvAJvx+vPgYe7
TWMRzCT+Py5Xj/Yn1NPGj5cqJKn/BYn+jdogPECGuC5gk+IyIKmEtKtN3UcOtI+PkgsuYaa9OdJ1
FASU7xRlKASoZh9Wi60JlLLRSoQsbDSdOpf2auKf5O3gmr5XlyegFr9+Nmysz1bqRy2ziG9UgEmt
Xyg2tvDQmrtD38M9Oa1R8DkVox+5eehZXEhnaF/n4BN+7jOsjw4eTIhsFyFLj2tTuaLusB9mPxDR
NYsZgBKcndpnRQ1jWQFHg1ris7I2EBLa99Vd9jxQ5YH2dc6o9OiucwVlMHJTAYz80g7QHCm9d7lR
TbT0GSV6Z8KEVwotyZw8aClOptYJTBm2WqKNgIp9LngkOBXwTRC4yScSU6JJv1DSF0kEG4NUNwqI
At/6g+jKE3oEWsimb1lz6Fvez/Bf3wcobqlf3BEW74OZfdsmzVn2UpgP6RH6pbhdJb4D981mdx+v
W+EKZY/m7320Iy6JPG4KZRHeMS6czV9H368tTonm+SUEgtcHCgqZ0bffpkA1SeDb3+IrOBkOw/DC
rxDrgXhrlFUrMEFliEbujvNKRnBYTGwhfJLXNBi/trSaGRiR2VkHFPfKfAJ7bGymrxxV1vrOz+S5
5zPK5R17+10zgarUG1ymStSRGjaTaoolIgXKVzNAJ0Oa178neXpfhu9zG688RUwXum+Jp8AG2Zmf
sZzZY2zMKjOQAJnF1sRiuxskcutyrn5fV0p1l2U/A05EqAIymRACpzxrud27FurW157bSws3bKk9
5s3RqJ6bnE2qY96Fhm0QOTR+uQLwFudKLUeWUMzQ59C8a/4jFdvsYTCusr8zjWrasSJsKC2LiXH4
GU1MVbLNe8liBnsCrP6ry9ZZNuFN/DiHqEu08iaoGePH/b/Gov4m3JOZ6PHez1ci743e8tUsx9AS
YCone+Qhy81R9+CXWNVmkjtKyP/J1spJ19jDOrMQmW8lTKmpw9Xbef7d+6lejGUSZJpzzP/h/uE0
09aK5WR4/5O75GcIHlb0OBualYKh+0l5ET0pqjBNnN1GOrKPQJ+zF4cdozkPYPqKv3uDp1TlkjKM
R9+4MBqlsFZPAtQMdeUZg0fAwDhcEzanY0+tDvWWHAIhw7tvuD/lZhbbVEFnwGwv34uN1U2Uutd0
gJHrn8E06AFZEMfmYOnUD7J499Uq3mQ4ZBb4p+xpimxc3ORfr+YgUkd6lN6jgsSNqwHRtFBc/Le2
EPff4AfTJndPlPh/PVQI5j80xNN938wBTTbRnvbnSBYXDQcEXGkRMN7hTfxGJTYrOQmrcQWzLnwN
1chfY7jCF9avCsi686Jd97YIQv4nJgDN3Mr3JZmN6RNrCFoMbeIK6Sh143k8rZ0nu83vFxNeQ7yx
+wyIOmZDW/+N3VHdzKVDr7oEMjlsVLgTF6RJDVlzTEOjAKYq373mQfpVdH8rE1krNRkkaFGB2WNZ
H7djqiemEkRxlE3BMauMrXuFSf0jLt5CZrnOtcZOzoiNA41C5y8xU/j5Q9SnUF+Wq4LWDjsH0sJy
22Fu7abPvVMxpmsQBKqowUaAkNPSVNfcl5mDpZrbpZ01RrExmxG9cT0AKw//tKCDrGeuFtU4bs3d
A66iwfeEZY530WP0V43k6h1SQHT83krTG1Yk4caQv9wnrASZDFcMiSDJnC9ACKn1HSgD1+JVx2ut
eRdqxGAeTL46f7AqKcP/Jopztm89hCt4GPqCkkJboW/TMS1ADuhL3y3v6Gb2lWSoy/V0twJgAFqG
3SRn6FesViMcCPQUIJ15e6J0zRCKHavXy2ytTJWxZuONqbxGuKJkY1WKIK0FRdGc8ccwKJaXUCDf
oIkaNN31ixmRM9XADQkAUDds0rBmx+Wg7hAyh8WHF7CEv8hT3RQt8kILytG5XW/9MmaD1kGbNu3E
ehHrEdxLhkdQrSsw/fplArwAQPGK86FT8oXb7Mv6EE0Tpilatg4bm1qmDHJnSDGznts9YBt9V/LE
yauTFox+CgCdGqVWPdPMQqpCquzfgz1i3pDpfW27Yazx1iWP1gfs8/kPyFsKKrSsKLcWsqsLikcj
G0GeTXVDC//daN7vkzERPaGiM9YcTVsogFu7TyFclfmwddbjemnJ68HYoT4aiPAIe46jT7hbbP76
Z0GsifWDGCslFW/mAhKFpwnpHXe10MQ31IJOmEuUIA3IA1lFdLrq36CHBaUVTarFjIcg6UeBqC88
ex/afjQrCJjHaxnI0OiRsdYd2OeSXcFQwc39/AnQzV4ZAHjlUVpgE9xb+jssK0cpOG+D2zKAwSan
cHP4CkiN9PJsEg42eztyadhXXqIaHgQZmaSyMQZZo/EagrBUwBEiuRdzM9iXa9Nrn3O0qPbVmUQW
4p/wLmrTIGpuzcpUfN+R8Kz874NcJStAPQpjwAauVYWpedYjjMuiqQ1/oQQea19hXWNM/XFgKe4J
u6dZBaIxzG2qvhOdL6c9shDPfdIGJklRW8MnW2dCd5iYs/6Bod/S0lUXYpvtP7pXz/iQk9t/adSB
xPq9kRkFykq+K7ojkmuXnQ3QSpH975KuitRJ9oPl2QTvrq8F2lzfIurftJO78QF/yZweK08b5fNV
emStLjhDPlTBkUsahPh9mpEwmMv+yq4oS3JAEc+kT0EqeOgF+bl2V4wr96UT7OMqGHIvEthRuzFE
VP95WSS7fC5xDdRE6rQBqkJnf3KIrlF6wdQnCWulIjbljmf9jrVRD7g/Xm342EJlW8zkT8yoBfyh
HE3bAkCXg6wBFqxvVI1N9+5GpNi1F/0qHk/HW/DlqsDEEdIsw6MDfH4bnYtA0hgt4mAHoYK0VkQd
19AqpZeB/bdF/uGTQwH7upGbsPEk7EEvgyDk42bWyXHFSoY75sck1ceXNQBrOTFRh1pT9iLu42GV
khE0Mh/BVZJw4pm4v2JxFzZiyPDSPkwoAOAjgMiFDQxI4018S8UGRJWL/0+dGH677e+wMG98X8+R
IZySmgTFIq2G+l1L2MPMiilU4B/byJsYfffBZxER6K2lofgvZYo4PFxGlnwJFWzWgVohwjLb71e+
PlLSDDLyZdpxWgCmK9XMqRB9X/TNTNQxv1/oDN8TwSBtWgCfGKNzln15dCok0vJnX78Pt9kGFj5P
kf/CH0vQSmO0vMSxRPgs9XGeef9Gd/WwJvXCPG+/ZVXsjJNY+dvUmYkEIIQqXxTAAVDlOXOaArP9
B5fYR3FkRrSiRGEN9ImpvZRp7EujJP1115gJ7Em8M191G9jmlT+Doh1+pgs3UsqUMQbfxc+Ghh26
nC9wOuBXnfkLFC/4ywzTwxarOA1Xt7LVa6xQG3BLBLa+9B8wMfabg3pXSCBXsI/KWL1lXD/1zXNr
mjh/yppE4qEcBeSqfZVYnGe7YGF1wJAiWM/FdqOQHKprXrUgphhbSMkB+HVRBrWe+6/N4cQ5F7G8
JCEQ+JQDE1VN48JLkCDMCrtsW20pzMHH+Nu8iSPt4ppkqUBMBfuCpp6mTP+8qR9AP1dhw5/wfzfd
WtZw53qO994C9d4lpXcXn4xPh765XqWgb8Xip3IlA95j3gYBLD8NmeOChb9bnUAHEfYIt0mKdttD
CIKtgb8jF6MBs6RkWOrLKCo8QvLueNSXW7UNrJw8+27ntRstw/DX+f4CFBAmJDC3Ov0K729htgp6
qfnxow9o3Cj69Ik6XJQf0SvkELc0AFfLJ9S1JrfjWIaC8trbr4NnTs40b458rYtpwSw2VfDciFwh
yvYCkP6lU+X7uL0RLy+zjAM2nk9Ibksggcz2Hej+H5QWHgoEo/LnEXBJyDCIEk0oU+768uhBqQBB
7M52K8Os6oCR99RyGv3md+M5eOuucJcHx3QqxgSqyXy5NXh/8EsI7j+Hx9QqH2jdiv6HqvqXPU2Q
C9OjZAY1C9OSN4Bvk3WuX46OMwO15FO8yYEr0W5eo1tWJP4Vx6TAjbJd5OVjCMSJJqt1XuNBkVAV
U0ceKmeYpfqx1weLxeWjhXggenAyrBG/4KuYeECavedTCz7C7Zk8gHdqfxP6D0q2InhSmTvTd5Qj
lxMgYa+AFh/ymtW8sPDT1b0IDJ+HepOyVfyzDzAbftgSZT/89hphln4ndFa+DZmYX0lrS+hkzGXZ
ebH/yDqTpIwaxscW+Y4riPUAF4g99Zo0A/wyzDSrRFkeyEHwILgBEs9ICp3+FMT+4yaLjE/h48Zo
BxSC+vPStofCoIosAX+0xQxRFeuptOAFhTfFiqVKkYOXCaJlLV462RpuN8WpP3vh1PVbqxxESjKX
t9Xisk2EAl8f8LR6Aj6jgR2FAlXq3QoyeV+YZchue5ezt6gyzyHbYMGELK6Ns8z2KcHV0RDwCAym
aNy2gbb+9P8DKW4/Whyi53bGmpPE8qm9BSeHm9yQdh8BHXufAdasfXdffo1h1LqxTjAXWZDIohTu
DiTNdHep/kGZfR0d0ncAyj1xW8VHmSd/IfzrTmhSTh0QwWfcS0A01g3VY/sVUCj3BDQl4i0LeR1x
D+2RjyAC9kftdEFvCUADcMG9Ns9IcM676YF3OZiMl1h5ntA6lvFGmJVltys49htT34Ogetsi0DV/
EQ+uKX9BWHpfxiv2nncAA7YOs31EbZN4eq8HTkNf1FxXp/25EaEPiUQL6hBI1eHNfstRBpbFJy4y
FX+x3Zqm786zMgWJ9UBrhRTBiCuWxwZzgNJ1uEwByG1hMDEhp5quDgwFwy4iI33WxY5Z9LTtC+fT
WYeFHLVfDP5+MnhZE/L9ZhVvcR8MTVVGiohVFWdHtk7MADOs6Hg0hNNMR3ku5L/TfwzcTjGoCvxY
2KMgOqGwX1imcartl/3kBaV9hc71NwDk5kA2zIwWZQJot2CvdlSkizIKAJRuOHo2cTv14r95bjnJ
v+ot+OobpAMVDGCKM9u445WFHVaU32QA03rgyqKlbw31g4H8lrTsd2BDPctDexH52G3gUa5UJRIq
0BNqtBdvjOmgyN29zpHDtblZda8aoNZTZjYLRwe5Uv/lYqjXGEjobCjgBmNzga61iGRXNANY+214
7FjBUr0xRM+G02IWIKsKg6y2T8GxUKL7cpCAx0b38Bj3vBgvS9oxFCOCAXTxMOQf5/RnqexPVyZn
N+Zk1I4xrSLLFa4wZPi6NacHcdpHzB69UOjYX/xSBE65mylBKmrz1khisFyBjJUqR3QptmR2J4nC
Dt1ItXryLh2ppIEfPpWrNnPjjezsrTYM3uDE8+Uzx1lOFBunO3nPeUcP69XL0iZh7d2e29iS18cK
f/EwUdysmpG+kZGSklSkjfkfuh1tA+zfzGZPE88rKGrBVygkIusyeT9SLd8RyP5EXP782ZvoaX+s
T9IqlCNj5ybmXNshkMKwFELYG4i8BbZb0Q2NYw4eh1iXADgospu89S+hkebG1jwzwXE2X4c7/t/R
f2uhU0a5GVKKpblUMLN4mtHKT4Gs5i5Qh4hTRb0WX1tfDy+nQUmFdEue8KrGE4gmFUWS3lV2XaaZ
k2cgQvjqGHyk3CQKgofY8ZXwg5alszhbqHwX9ihtgCV3kECDVHPihwAdzfwLxgOnBUK/LAy9NUDj
w4tLJbEZIRUnFpahM70fLhEaQe2tIJkiYUz2oX9dztabmg5j+nfxH0g6qs66nJbHhtu69N2IHV05
e6lyAaunkknoC0fsyLrbwnH9vsgXwoisQTYLyoYIWgvDuaY9Bia/yUICDj1+Xd63CrqhOmgyG5/a
+1nOFPFW/NSD33JGiYlhgHcv80+1xP9QTi9DTW25nSDsG12ZhHhxzbGSJlAvzCwMkv5gQxr5LK4N
qMamLcV1dHR/ivF+LAk+czjavxrmVGq5fr6c9JvU5Q3cStt3xupRd+oJmOEaIM7vfqqCBb0toAEc
qBvEQoBeyfYZltyZLgzUn4hC3lyMpqpLoXwWzIgppB3yk6Vnv6XQYM4rytzEMUqwYEmR2rn+Dxfx
mpjcqY15buhPLscLPd7MRimVzN7ur9V1t4c7XhEFpAPHafjXm0EiasOP3TB0f4W4+BkiJFBIwkv7
0BnUgTB5RwFPFE5WwEWD0jXaU47f31rmSH5EnOeQ8IW3mEwbmIVE/Zf/ByPv01Aj5dYhr3qehS1O
HenSjItAKQfKMMu01IGOIKPrXDM6wnNQFGgnVZnsazeuxdXCye6oAoB0j3BXTiCETquf0Hn88keh
CHHPycS0bmswUmZ8lo8yfnvBD1/MwA/oixdUaOljNB001SRIKZqffghM31m8gAZ1S5N8abMT4iBR
JbIP33Et5A8aXf54wxVn8fVu5CFs2H6GkPFgHNHkZdlYm5OFnS67lU7yxBk4RDqEcSDBS/Ph0k4f
VWNsqw7r++Lavvqu7oAb8Nf2OPMg/vctkKF5cvK+zyRkDosOrx3nzjbcUtfxcAtovIE+b7ckc8bB
IHCkMjmJlgyqHCxxWm3TceA3EuLqyfU3dldr/VDjYowuzFPFxZhECWEUBIoVNVFAsqauMQtNQKFz
EkQfAEIPWDRcNvd8xcRlI6R5FymWikSnsFaueSpBSeQtJxOiyOssfKTWhPpxS0Fs137fCv0dWHjH
lQoKjGpPIEH/yTroyqVOaywd/JmBSR9OTLQ7zKPOO09raddeG51VAWZSPMd/OdKfBRq2NeVzOV4A
AFn4WmPQdT2x32AKhD4nCdg5/PFfwA+onS5opaRSgsCII3hq+uz42zkoKatW6MGsiVEBb8pV3dEA
ZMSFMeFkQ0cBYI4INGXxxxAwFXAWa981Zu03RdSlwl/2CJDrmO/ecIfuDncl/LBP2UFHyAOC6aud
FlcpglJpc6RWkd9seU05V1N79/SR8RGc088lDZuBWAjQRJBhUh4qvNTfdfynXfMGBj/etk7zgHTw
0OYF3GJDzrvu00ofc1ZZiK+LeUcCETvUO2PYbI6X4J0eFNdtGGuq8/mWZIPH/yY/u6m2LXTuuZiZ
a7czyKAPG4TmuQf0xa2BYQWoRNL4Prp6o8sTQ+xc2kAwiLPXNoJ7clrVZbmu2s9kuaRK1SYEHZIx
xW4I1SVkKNscpjoiuBi3zARwre3cfHPdlWt6ABaU/PNnx/qokD0sMvdZ//6Auo2gVIpOb5YX7CVG
GloaVK7EIPfpGT8HsHbtJXWzwdff86W/zRBBE24lqDiv/W+wGKQRJceK/vaT5IpPsOtq5AidwEDZ
I8gxzGouVr0JLqm6gAp3EkcoPEVjvxZKg/dI+nIKM+PknvgV9qtYaDhOOgjtMkl144ROdsF3vE9B
s7ayNlvzDJospyWhj1PjM2b5PoG3s/HkglGrm3nGTy0xVEfcXpYy17omknjUgUVwnCPY8ViP679p
7f3w6Hnj3x3ILAEbh+Jhh8kZ98q6XcmcrXKzr0btydDmmIiqTC7muzMekgC9ugKOqy5eoOmxDbOx
B8w4wtHkAvTP3XcepxgHpuy6jTacBtLs3B3VcYZI1F5hfItYhn3Zsgqsm/xWF/5OMbqt5QoGenif
JVBhrJ5ShmYzoQ8yYpunBuIHyyftmKytN2j5kQ2I7inHCUdTUyX6CSjJxI9bggLgA76sa2OwRSTf
GM3VTtGSboolUXCPXh9L0OoAnxNNwhf7PBwtw4J9u7RC2yLTsTcGHp38bb4AGAJR4VfVrIRYYwWo
YhsrCuGlTB1kQGSUu36Mqc/OK4w3QgUEg+ywqrGCmpwaOENd8JmhaD0kyY+Jmn8CnTP4LXzkNn8D
TnpzbYT+AaQunTByJYn9RnAohRijxjm9CJLGtAK1O7PJNMhUeyCiXqJHtwRZWREJZvljgiH4rsQE
STPJRxtM3aMUk2HlhgsswpIAXmKuK6BjddmGHbknzGPv+IUZn50MEy4/Vzd2DweNIXYWsfJQ3Ryw
kwnU1Ff+fKIyaMKqTyEEBFoMx/SGmHRn2J2cdHtW7RAdQkOzb7DPmtbSewzZ8tg+Ci/B8bvdyzmQ
+rp2Pr4V84wj8Iu20Xaml2uKejkX+nNuOPhb6zTDQMm08blW6OpMpQjirxZLwksBqVFv9SxmSN6o
0+lvgLGv08juP71fHlJof0fPhXMiyt/dACEcKArJyRtaETrmAhoxJU7Lxw/1Urxc1nRoN6aTqQCc
WRwull/l7ATFIxppt6gAVUNlth45BpkcIE4gH41YD7bPFPlhPid8F3XCt/YjHU6TIE/YU6ERGNKi
YvVgH19wTVNX+FIIPC84+JcYl6tmee6WThIyeg8XyoNFlpjbZwS9PjD92OVOgV6Z4QLGSRo3YU15
OklBU8xM2hF/bWAsfmiPrlmbyyhVd8QC4T23a5S2pYyz2d0Yw+grXOPs4ktCTP2sIT/UjbFGdkDI
jlzBNxHtK42NpwTsuu0ANpAAJupXpzlyjNgi+9Bm8wCTjTCWMd4u44rbCKcwzerTp5N7G2rlIfR7
rmCg1SHLLRLVz77FlV8iW2Jkftj/izl3HguRBojX6gNszbfqPuxfMPHB62mL6YlJbqdU+PCR8c5X
tMkdNlY4TTOHQKYy1Fv/Ss5c5Ky6+BVDuMt3rCAQfFTl8dQXISvttLHZlFLJekzTJw632sHzRCnd
w3UEGwIauDOTrsK5A+jv0RgDZJlCkcvf9TQmNEhjg61TSY2+eyOOUUUtiE0+DwCqT/MWCyl8+AY9
fAArMqIbJZ7tIY3iHTwRAsdqeHZrpngbUDp+Ltp4gptAL9tJ8jIOW5XeJjDz/26MoVqwAhoetOOn
vzyIhpDaTCkEPzgLRPhu6VCUeTv6zY0ssSDWardlh0vT4UnGKlz8vXSxQswwOCoxXNapq63N3GiS
r+KWRxccEdvrCe0z0hx3euNuxRjlUyABPH9vN7sCyZvWomt8QEpYqCvks9Cf/4z0q6jN9H02lFJu
k8GUTgJhaCC7ne1z510HcxcrcJ/A7v9g/HQ+WddNtPy6qpMbmC26dVX2SjDML4U8z7GYaOoyqJSC
oQkWHuxHOEf6DMmHNibbIWBGGI/rauC6HbX3+62oMgIqtWvVBi/HJZ9hnwedgIF3OgDsJpn4MFDX
YVSlcFCMQ4FUwZzbePhq/8svlzS1602kqPAQUVJaha6OrN74rSSPsblnpyvuT+0YDK7yFb8tmQIx
hlIxxxzes1YPuqdPqCWYnpQzHJkMH25Q52Dxv0wCV6k7+3xKTqpbUjqlPbndoEM3Bq44KfCOwKwe
agI7CBybjcuqcQiLbME3JxP8kduHb8vqMHD0tUFukYjaG9ho7qol63vUjCOkPRUJ0HxSPUXZ1e70
V+OUiaw0s6IFoHOyia3BGZmwP2WIBVHsPp77xCRpqkTcTSyzDqbIs+GHj6bT09aQvzeZR9bZSpz8
clKl8pvnBpG+ko+b9R/kqXKtnbpL0IU0fsgLG1i3PjdQgIL2+an/KUIEbaW4R6XwZ+ju5Y+mzXn/
XCYOEcNXSTPLfECcii7smbKfjXoigip4JpSNQU11L+MaSL0B6aUCnBC0LuZnmjGEpmslhMaAUzwS
+EFahCvRWIeHuWhnEgxLuMikS1ZiqWbdF1RS+scUFzrJkTRxdbGxX19B+Xt9otk0pWY3fpG4joVO
suaw8YefMjMCHvElWuHrruMOgdPXkT4A+nkSTIqaCCJrYcA6nKd/fZ+RgfWLUunRQogQ3BEabuhJ
ohGxk2GvneDRKNQ1rTsaAmoVjdRNlGs+WyJ0o2bNlIL2DR0/XrIB6M6t6HYggUu2nKgmJAv2XGjS
SNxA/5kTY+F/9Gh74dTw8ZbkVNG76GpNDgPUaUQnkJpMV2OGLvY5C0nWE7SmBXIW+OekqO5trrmA
wX1hldctYuCeFkcWFnaH1skTTxxw5drMDetRgSI68H2+KoDFm0pr4EKy5OBA68BaRy5f4XLkIar5
kpHUpCPn6oSp5bQlxsIQTtr2h2eY9Lp8eJ53QFR49uqBOsb0EanhMKd3q4cyVyfeEuA0ihgsFWHj
JsN0TTgkxYps0yvFQJBNyOuB2ySZMC7p0pVmp13DHNN1s73AEBN7DiQ7359TIuoAltNDUZg1jMXO
zQVDmTx1o/K+H8wxdge5wnjHAfz87+wKKGmwgD4g++au64JI47zxD5nn8vylKY0Ie53YCpSqbMAH
t+/6re50IlBFwtyj9+TCGFxCGQ6/CCHc/xGrKjYSujDVxhLaEc/rUuoCEVCCbrYvcGUYP4sgIq+X
zmzlUdTF9PCC+CAH0ZeFrZLA2v1ws5fviXg3pNt2Ek1yqfxEh4kIcrIgv23oH3gszT9yxtZsB6hv
UrHIUsy5Syb42PBFPuLwYHA0AWksALGfDcRX5j/yjEZX3f6fbPK21biIYKc9cR52wh30c9Jmvpio
lAeCnjFw4qbbmueZZ9tCWSYlldaTyo5adx6zoJE5OtBQyZk4W0ufUOyB2zNPDJlpCuGD7u79yU7p
IgbNdBI6MbgGmdnBdPkOBuPtAsMKPgIgA70xzwuS/dk88ZzJ/N3tqRAYhQkPW68fga70GscZrsc0
y0q1q4e0Kec1rxjDZ4qS/0MLZCPzwiXrK1uoM8Y5LY3kNkbx11SbmPV81IPrNeDrEYFOwRvcJjMf
deCdTDo97GOv/l6hlEkc31+wqoJ+H7nS6r8wnITtP/agk8VHjYrkPdun6ACL0S41hddKRsXAa5kP
u9OZkEIR1sr6wxdZC07stJVA43cy7w6spjeuS+GoePhQ2kwFyPgIp8qufGGEkiWQB6nQ4sAV3Mcf
dCiA0CGz4v6XmFyxC8EeYdmx5GEWKw1z2kri9IG6eZhe1qYI4FnMOLciA6JgmNsP4ivq+wIx5Dyh
KJWCMzXsRFJHzkfjA358A2AOIArT1HKRF8M+pHr4VXZ7N7d6aJsgjkZS6fB5q3ZOamO3XW8hpi7s
3aq7mHyLYCiUPSv68RkBtM/1ZnFCkYgX0H1mBiJ8iNhhiDPYSBPvkNF5NhimMx1icb5KGCVuce5H
VvukCLVYseMDbAN1BZBu0Hj6YYjCksY/iKJ7z9TKqnE/uUselWNnqxfleHrcn9g2gJ1ejPn0ZI7L
Z2OWynEDTihDbTm0sLXdTRfHb091nlgObdbRufvcVbrtKYuwbTnFmdN18LwcUS59rlZUQcPyn8sW
xQIVOhQWYikFvyLeEr9hlswh+3nK8FjXDmRE+PTkFSIKOwh6JzRlZ0TLC0IdnKNiDnPfFHfh/hvi
YIgPAFgSCgFIjb3Yn1JLLVbASw8nxKkwjci4n7b59pgGVkKlUIaF15GIzmOV9iMimRM/JYWOH4eW
/WcV6kjyGtn4fyEhUA7hoTiDxT92buHjIUKIQA1S4LPQecKBlVj6Hj5Uu9pm4m6+SVApJIwgvnMG
kow0sRdsIp+35x1KBkmXmQ66Hrp3wJTlLFdVq5L3oUhs7z+uKFW+Rk8jdJ/+WaD3BDEmLGIvA1vl
4ZIjwZAM1HNpcL3ZnA6rCIahwc8fE3W0SJoWIo60F/TRWBcNQe66niR5RBdk0kjz0fgCdr2lY3DX
Uvg3ovMZgRq16c3DDxBt2jhxb6/HjBvfjRhNUB1ciVLdXupyAQVAroXzrZLpZ+9DOMvaYyUxQuu4
t5QlhZLY2qkEf6fEt/uszKpYHcC5EKbs031KzPLwGclDTezuio5VILv78pmhcK0tzcZvHfJJPq35
pmmFGEWcw7CBJr6un2ZIg5T0GNKpUl/TAzUQXP5LvNJF02LOG703pJhtsz4ffPCuPsawHH0YH9AG
dHvx6Yl8wPlldSKCjgqXuyyt0C854Zw48/iAfPXK6+g0GV7C+S6CJrmBkqIehF643eE5q+9aU5Zz
cxpFsMmDS6F6k2vs8d61xQ/I3p6uEnes9eUR0qmmA/b8ge/I26b56fEac0WStSgDlZroSMIzBpN5
7NeVRrbA8QSd3ikr7rWALVMv2Oj5d0UfEqO6DNAiiVsfLMHkoBbhcfLIM768zXzZG2M3XYMPDyPc
binBeTrvesV0qoM+Jbz692DETIUub4ieAvbgjdRTL5ocxJ83EH1EgICGDBJRGXhGiSfDkLaTawpq
IwHzuV6zSmGZBymPJ1qUOClvmq7LzbjqvmGYBSlFFngwNwcqNS0jZgooqTumUsCq0ohachCTbEhf
dhcILLIrq++3heYIKBYUd4Tj6ypDJW4wXpPAhEMLAl0D07HRfvENQEr0ahRWSeCxjX+9aO6uHO1G
8hxiY+O2lrgAAmy+7nyTN/3/W3d68VLBABLBvTkApdASgXnNx44KiW4pjOLWsnpd+R1QrSchL4a6
T5W20F75azJruk4R015rtRel+RWX5x8oZBpM3qZ3/ZWQtGX3RuT/Mtnhu+exVUpyUoWMHfloLelk
qcAgZ/JIHSmwNfZSHk+eWI8Aav/JIm7K5t1t2WPq+5B+edV0YDFT4TQfVEeKztzfbPYOcdtH6hRb
45GCngRjU5RqG9cHzLOxoWa2fdCh0/jOba38MHDc0GEQ+LUYmuP5hPC5Ag13dwQyTxIEx7oPfl4F
9w3ymAS6fLr8XHG17hmhSSVTnwXpGAJkGkViVmRWK5zW0Gg0fe/+eMlb2If8NtDoe1i8PBLBAeGT
nJIkGkPKDEWg5aS8K+kgo+6b88qLbdHaGLlEQTFi5NumSGT55x+XWaUUYWwTRXwI9Heq+aquy54J
O5msmS6ARNplkrYgDn5CHpt0tTuLbw/ZfxyBwcGo8rfKoq4Nh6IjE2UhiGsoriDI4/7ayb4kg8hB
OgcyFGJ5GZ9XomsAYv8czrUsmouoM/GvIf9WpzW/k3FcQ8BiRsZnC5eCGvqR8UJKXUjD5KopAI/I
l0hVKr7JuSe5FqlXc+MGob6c612mFRzW1UGo8WlPdFd+gf4w269v+Q/jQGspsyn04BeV1R/eBZtJ
FPHYOFF75r4ZO6bxJ5V97bbD/PeE6F+qpQoqX+kSnTCNVqE5Ff7YQls/LEZ8IQb0QS6Yzg3cWQpz
4Y9uEkVu7QBLY1JJsFsBGsl7o7RnG8a8qYG7jEUQ6y5vOowhHKcn1+eJ7hR9O1KZPPWtUx8S/gJ4
QvvSyThxNppviMUY0kjqRRf93U4aQ2DoTUILVYr/R8zL8KVVQTw5pSVcq0KVy/vptZYhiXBTPf1f
zaLR2dDNsZaYHceYwPDz0WQHJ0ITsY7brGlekT2cAzSNFgvPwRxwwIIiSO911K9uq7WGOALhu8iZ
PTVHevbrBeUVw/OoAK3OJbLBjL01ff86fXkrxIYk1nfae4vha4iAWSSWqdVy0BiWESTWSJhYBXFv
Jpwphdz5YsjFgTF2rLVQQrECwabN5On4SYsCaD+CZ+Q11jI4d0ndqeMSbw7Al1xrz8NNsY1Cahyw
z8UD+lPaTldqzrnqDhtwug4h/cVYgWmd8HA2GTB33EqXpzWnxSM602HQ+VCEBN8p/3fM8jziQU4f
1sbU3wfGBKA8Bg5ECA7Hudp+NdJ78vbbHJ9mneokluegT7z0e/gbK3wbZ5gjpYZ13r+nNVf9nzaN
rBP0qvZqKEu234Ird6YpaIPSYpmdPlWx8jQqQ4QtLNaDtdJ5RaWV8uQY1snuJZHLX57ljvD4TLs7
Wy55uSqrJQyzNcjf5mdO0EUjHyleo0VFeEPzYzQPPAmhrv9rJ3mDV4KZicf8TDfj/+vr9WAjJgqz
zBCfrLthyEVG5vb/VRPsnTS8feDQcw879KhGJG935QcFezY7OvkBLVTWr87V6btze1Z1YCkzI0VV
+JToftiFfhxykb+ivbCK5hv74WIyu/t3C37nSirlKPard95HDcfwjLzsAMbDQ6vp8aZCIbTgUHMJ
hJMFF0KM4cDSqgqCkchWc5wYhvu+NPU6XQ+9uBNYP8BfC7WjVUOs8e1ZcSWe0I+O1hvL3huZzOZA
wOP2GKnopJQdWGDETzsoORQAc9BbAjfZ+ApLjYKxMFN+3yp3ltT6v/CVrIGNYdtTNgLOq0SJQp+c
73PuioUrMlnI2XEKrjUgBCr80LbdDHfgy4OV2jVl2sgtIFpTdNxe2DRwfPeXDpM8+zwwbEg/RfKa
J69BhMJ4H9vkPK4UVTdYl5ILqDoBhNy92Qpm+E9UI46dvU/nXP1/HqkVQiD9Yh/HNCR6EGFCRDRh
uXmtsggzWREF/P7cDeE34k8SAJKmEHfhNMAg0yakBm0vw/9aVlkOUzfzoWVfDXvG67/cYAS0srO5
iELp+YcKd4z0pBfZTKFYn199K72oLXo7824q9Wz97RaU6zuS8y1OPzoBdCeLApoEKLgrWl/7dE2H
G/4WDR0gYlU3aM4c37DL58rCMScAGu+wh4efVAsWHXoCMPPZCr9aTldVR7WMT6g3+ZJT1QdW5Gyc
TtVmWya6jNqYEmQgzQHUbuIrYniRH+GqCnlalmpPdDoHvIXuWPAdPldtPRUdqI5jy32bpJd5syk4
KFYo/WBDjMyuMTHiGTT4dQZRNoxYELSyqac/Mks0cvcM9myvDVGDvOitl2q8P+9E5pHQbeeAEF0x
C/899kT9yC1KQHpDrpcO4bH/qGBYLpVKcB4F/XnnSoqW0EjPbhsnVb2C52IEJVtbH6NtNYv6HDcH
xt0ujhwRFZTpRXglevev6NsDK9h9DjmwDUjl6rqhoJdS+zEtvmGA4DDL+FS5Z4+u+KpTfUmD19nB
TEg9EJNWJAZTsZk7dBomHuoA7HUdTokF4WvX+a5R3moqDL6KvZFCExmeg2/z7BKvGYubcO7J53aQ
Ji9jo311rmT3zq0ekx1DGlpSBzIHUQyI0xPODwHdq/+Z4RrB60QGRlB4a7u19msZ7yqQ6sw5S0eh
GTOr/lxQAR0LTB3gfCqSVrUn5NHP4l/agtPXMzzfvOyNHix0uCgtPA75ZokNeLK1LJvy0c21yX1R
IzsKBJxoGPcj0Ba32R7IMpyrcmMHWx0uU3siT8DE6fyL+XoeGS98Fecd9ZIgKhEKbs+Cq7H3U27x
yYjw11AnNlmauk8UFKAaeF4FvDbkt1eGP2Qgtn0ueiDjJ4Og5BRX3DVOpTOYPVAPq5Eaxxs4J6tP
4Z9wD1LsE1OKpcxi26lw4f5YLR6/f7350ANAw8jbe9qqRlzX1NlXs4kZWcRlIrGrR/wQqE9RU1R1
kC7HeryB+EbmGKrmyXF7leegWCvE4EO/Ks8Y0Qn1Zo4Dfa05VckYjOg8q3of92POktxoNyMa4WgD
YbMgTnri6QhC6PKxCICljtUrMveklUs5RS3m2cGnJl0OLbZavu3I6ChvthKYABXjZKOoUy70KfDJ
qctaB7NvgZ/kix3GooXwBdQoXOU+O27duvpXpiHyp+cDUeJLQE+v4BQek9w52U+d/DkBcbp5vHzU
F0MAQYuqVctmPKWZAFzxtcAKz+On35G4wzM5qSC3OCWuTx/GR50ASFMDheKx3VSksxfBsS3WyR4N
Unll6b4TPfOnSSIjsUS+d43OutFSBcn9u/hJs4+YkDfmdjsPLzj4KFIbpB1b6+RaV1fvxRmlGFQ6
RUUHluIfHfVyXEHupa5KP95T3us7RKDTnzbCixkTZrEzDyuZCNYCGptj+ObAjCPOaTfU46a7rcL/
nUPhUl0b07d5unhST1/hQ6Tstv4pCNUKdd62CfWAenepKmxWpSkwlMHnB492PNADp4fHr9EGD/Ai
bYB+dyHxNDmMlq4nza8CENtkq5oqieYolnDAHr6T1Vl8jFutrEXhCsOinRTaZYNMPGUVTepw8oSt
cV6V5bZMKEdyzXUhhljXN9Fo6yfBmE2FWq/OeJyh+GsMNiDoLPEADLQzYS4f9kzKUUhe0mcMx/h5
CIV56N2ejgrayGtctgK9rJxHQ9m/8dHAVnM6i974FsyPv77iu7y8UgdAqZVtJyx2WuHbqa5eB6cH
aigQQQUU/hGURyDQD8VwjwMKTeEnOijmsUZIzEqRgd6Q6nzbX3EWHxNvLmohsJV8F232W7kxJb1u
f5RlD34DorOolT+dOTdSdx67rX/2PtAei7zh6NL/l7ZPgqm9+HWX3+8UNVHFzR+rEhhBrZsrImyw
sGKwwtxqkVbV24kq4V5CB0woUy5UdiRBqhJMYeRIrMguqrndgI1T7WYfPh41Olqb7dk7AN/GyFQZ
sSqX66rX+rVhH4AMGPRXxAXdkdCnS/hAmGFvsSBW8mfzJc+310R9hwj6NP9YlXzk1HD/TiGW7bhA
DJxcJEMQNDNqMYary20/GbvoHivxgpH3KpyrQ1RkdyTD7jiDG0c0f72Ygy6tt4iz/GoYWywXTMbk
CFp1hhmkBLNj+eJ4xrmQLMIGyPfIjTXp6HwTCKXHKg4Hiym8dnEwznBhYyf+qC4gRtvB8O2xAivs
uOtUrd47gz1sLQwKgdtccckbhrAcMSXjjDgkCIH3ZbPvrbE8+0EUtJc0fIEv/x2d10DDlHvH91eR
P88Vf+5ATgAQM86HGZ50v7CBimuI/eO3nelmBAso4l/GWJrnA0WH/gutiM/ZhUHgE0Nqc3gWCMwI
vsvEGdhyXfhr2ZtWn1wgmgXv94snmtO7xxeCdUFSzmEn+NDciSt5GbiFJaRRiGwjqmU/ww/THUI8
OpsguLDHWqNXH1ZWeKEZuRhehcd885wZgvIFID1hFsPRfGvkFQPrF9r7fa4tua9e7jQvF/Zlig1n
HwGY7NvtKCL1bAsN2SxgvniiDdCBz009cpVctAOWfLIOEngCINOIC8XB8TU6N7O8uT6Z96wa9YYO
oaRQohiz2AdUKi3Kws1yoDLwUUlQuUAftIHIb8WXjcOC+/YoXfcwu4EWdz6Szo0+O3NlEs1Vd39e
Dr6KwyXwbMBwQHvIfFGKhXWTyaWdAbAmmYlKPxp1Oi80ccojHbKQjQb3gOIUBGWxHkWbAyEeq/j2
xEommKWHZNFlyL3tAW0DU5JrzCTaGzXJv2usAP8TvVdOwx+R9PT1NWj6RleknfmS64nN47UQ9ptg
RDTFM8X6q+8txUDbtS7lnQlmFlA+HLoZQ8ojq6q8egwJd7LFNbJkOja+jFoU1InsExcba2jQ/vHM
c5Idblob+Fc+JQv8y7qU9Ods00ztfBn85pDk5AQdvd+9hnB2Lf2/4J8ErxMrgMUMV+WzUgGr+J4t
2sBxQxPOpY8dKKgT+RHWRXG4Q8l2Es8QmV+mubkXzZKw+z6cuSinRoXV5k0YZ3tzPTH7YTdw0mtn
vMvEsb7qkOa1gmZTXnnI4woe0yD0fouH4sQnXlcrmoKCsMDK+gFzYa2yW/z7YBjreGke0/0m6Wrz
jHdVgi4XpbG9bSlAljrk4r+U1+RNKYOnSLsfjMtwHb8Eb2+0hLnwer6pXgBr94PmGY97oIKeMIHs
+wuzN9+sg4fHoHhkyze9cjNxx39NQYtkMx1X14fF0rKuTyf9YVeEbfvQM/rTkPUmzc0aGKT00MLy
hy9QLo4gh0xlCDOGBGtQxDc3IRfD+X5HyQf0jcWwxD7aiEs8LOYUBYZJuvkb8/fJCqYBL+TNjUzu
QdGcwIi+kXsM8kVWE5mGlN+8UrXXA7R2EvsIpJhBnTykLpwgG3EHctArX8D+i/lb4VW7hcVlwRtP
yBYuEqIcaF+YXPfJ0xLw+1scfeHujqg+LZkVtmdE7pjSXXZiS6YLBToDfecyb2zjtsc8yVH1wLEQ
Kf0BejuKq36aeLqmNMudc0MDmYqtUUCrBigiazMujgKN3593ZY+DaXCaCkkND5q2EZ6Y5NA9p/JW
KXRXnRtw4FlkVCV+UaTC/1a4hbXvl3GXYZu9khxLl2d5HjO6s3DS0MVna6OjJJ223ppnrEVV4m6Y
ztG+s2FWvYO4idOqqsDSQNjUV8t+yk5KEI/YwfL1hwswBZwJValRCcVO2cLUK6I/DLXAUnL8yVnp
ADyh9xL7o9H36UFYQFra6etNuM6Z/ACvf1BOZrKHBh3GDYoXYctVW6vWN7iK6mh6TQnQzMSE6UBh
98nY5YwBJq3WbvGGkpbdjfl+IndAKI8G/TNlLs2ExAni3cG5gSpz3kszxGXxzlnaFwLZBGEK63G0
vmDRjFESLEa38a4q0VzEUza94hYnmaWXU96mfI1S9Y9COnghXNKoIB4HEBwN5e+f1qAV4f6gEzwO
DghdGDYuKGsa6a0jyNVth++g5sNyKbv4qxtumJFlKHby4wo45U/1SFyqZ0O2jP2rmNrSQPF9mwRi
W6XsvJr295cQuR8tqgwtYdy+jUv3FSZeiEKnckIIqq6+Ly7UYy54eE5Y105ecprU1LuLB1uDDbsE
bSXImnYUgEBATq2hx1QcnmJoR46H0n4raYh3x5J3dDUC5NatKu42rGHC7dtNnFwidjtjA1VYEV1G
mLmCTASMHsBmPynj8OMFAXn+d2Oqn4nA0xRuvOEa7rQo6/NZ5Xrn28TDZN723NjmVE2dDwsalIk5
zZr7v3NSJ3sSocAJlGtjKbAerSanWhfgCY8H16AWZxXtCGuaD66+CzqOkgjIsV90NVXZu5lDm2Qv
0tgOMGiOUBXcxgIadOb7a+UYWbv2fIbzkArcewomsDBi4azDk2l6jY3v0Z+WyA9A01TBvBryk8ec
yc9bM80DXkn/8AwmfvkLJOdMs0lcWd9O15wv1i791fdDUg1+rHiw8xHw5N9PslARJMaCmY/PB/tu
rmNt/SvalpqGEMRkdy3BlA3rIkVAYXjXQ5MbDryALc3DP/fPHDKRcQIfBlFR1vNgetkQLkTXo/D0
984cEGcB/GV06qaedY4tzQ0EfxnqHgV0A0wLqobIo/ri1RlOiBuMOLCRo0OebGpe+cHA3rBQrzH5
fTQ8Pv9lEIbEeZJR/Ai9JTRHr2QtGrEzmm36RcXJkOF7TNDkY/xBhglIiLTjX2rT1Avf1QRNFK4K
xZ2YqQo2wM4wj++owjJ+X6VTRylZ6OPVag11Ai6llZNjKzEyW7s0ZbZaqSkMmGUY5517Y/4Uti/r
IzfSg+BDifMT82qYPjtgA2xN4TRpECeDQshSTvpOLZCG4t57Sf6C1dCRCRSCj5Sh+lxS1TTVxpXF
kYgm1zm3qC037P79ikYJn44OmIyJG+nbLkhSAcEw0vRodaMWNje9xTIQrcqb+FYZ+lSPaLuI9zRk
pDwxp6LvRqV6dzSjo2yPpk4LGpyOOiL04bG9nH0Yj5hRl/7aE5RObhNsH4DY+EG2B3e5/vNKQ+wv
qc8aJ+VhlqOBlTQrIbqXLXPXoeWrP/Vj25gcG0veZaeUYBvLHQfcWfCvOaIK3ODATwK7GlyfiApa
Pr6EXhr6Yfch8catGAhV9qTQQs+kbp5JS0sj8bHwXf/vHkFTM7xVFe7k1OYNRyQZWR2q+N4mI+xn
5KpQUPm9GyxHZPp2/WoXo4Ho+ju8LeLDXBc2iNFQYwV9ADTe8ENzJY9bS+7LVd+LAUu0ZlgPOWTa
wQ+cgiQ6Mv9yx8jLYp+bM54wt3Wr4/pKwuJsjCg2z+skHWFvZh+bijSRsIghBcDS6ebAqY9KAyFG
gqwH6RS/9LcDATwvdMZMPA8kN+p9gJ1OTA1taicei95U3CM+KS6K180Q0DWA3enZarryNFu7kJ1s
dS7cfulvlaicSz4LjRLDV909P8QlcWoBFaGcvaj8NMvdBZAROj9TMwEXUKjkjCAJ11TRn6CC8+D3
Bua0C5qwE1gP30O1Vugk2YIFMlQR5GGlS5jbE/RQGHgvw0CNPYer1AVdXKVKgvKaEdI+cZgs10NT
uczxbCpXsZD2lk97xS+hUadp6TJxlAmSZs75Te/n3uX8hOGgeaHqU2j00n9XZ5lotN8UZm7fYSFD
wSKcZEi5ANlO4CHSBWKhNYp18hF40Kz+mtkr4pW7c1mmdqV8vZOu0e1ZXIGCVRpf9nM8bJRYclIy
YtKWz0ZrsBDkBV3QbSZHl1ye3iHqwIFljmNZ23zTVA0ufrRSsCpTgNN5lU2wvslnk1Xtx2oSXgEl
jDzRc20KV2RbL8OqV6quNfzdcB4IBLY5yWQ1hh2755WXPRuHUtJGivU44jIplCeiuUiccLV7IYZp
Sne8iiPOpIncI80n45IXdofckEpbg1CVc0cft3yFPiCsqZpQAj9sANiuyanf64wKc18XUUtm01o7
EcyIwp5TQDNqy87NV+hmO4kW3oeQ47aNJq5mpuFMCK1xGLbO18MWEtKx+favytEIJmmobvREuIDF
02onBHfZNgF4a1IJDyHm56jH607GxQOOardG0GGXl2aOUVuydep+czfwyMU6NcdT2iTSmZbVkXMg
uTXipskRRMNdeN6X6wyf7jvQjgt1PEvPZVCnou2rpBAkdLCsUScfsNJXC+BSycwqFAax53dhRNY8
KpjIzHwdB8FKnXW9F+YgaBHXM6lDWp9QSbV99dOaG9HqpZjiTLjAiORVRgKElql9uGfo7GvE4LWU
HTUi+ESaQ7pZIOt7nrg8EnrTOsxI7Hi+chnkavnG6jQtNxxS/Fm39Mj5efvVHKifqEcGMYwi25tS
qbLr6N45yfwMgkQkRrpZeK2Ua2EcKOSE7jIP+v+oZUaP+/vhYaiH58qhnxQiYm1pfh48VK+9Vkol
PAbqtr0y1Py9SOpLcjaUDDm4Xpt/HjjVSl1HqmHdKs77vSisEW1x8HI2YqjNVZ6WXpakI1+1RJUs
VU9GIq9UIMLJozCS8AOB1JgskI1esY/jifm2lExFszdFd5qJN/VqeK2jwdQv6rg72oLlmmG35f6p
az6SHHU6ImuFTHuhz9dy1/+8RzVU20NNxfu0Zt09XgGfTGd3ztXVaefwcjG+1A5+LOLYcAfuhPJC
XzIomnYGbWhyuLvK2ZXwXWLbLruAxWlZruOiOdQ9UB/stprm2C9ovnVn7PEfqYajnapOYnnCGKXi
zhtY3nW6FYiljlgfvBNSBgZ2jvaKG90JwANkrMnUmrf8L6vIEjgN+skqXeoaqzos8264xhT8gMXr
rlSvSvBFQ12EYQEuf9Z4uf+YtN8+mYBTGnnpkOwOUjB8SlLPJG4O9+lr9Nj3/fGwHfK1tDaVuL4B
iF4xzdzEGIdV6J7GPo81yKDef5x2NxgIZMA0W7n7ilPxJaNE7vzidqBAjP4BpB4G+XmOhlEJfHV/
ZnMtdNBW9T83zTaTlaQtmIjsBAxjhUEItE32hAbsWd+KuwEH34Gx0vZyMdsoZc/5tHKzPEI4vjHO
ImE+JyOs7q6pMziY5WM3/rgP1O/9ktREvj7hlnw3mz76aQgSfThp/i7FtGajj3/QHBKpy1eC5HQG
bi6X4xSLdAY1F5rggqTtdY9dqaf5cU6/QhDmR9OkfTRwj6uBFTGLFo/J3gP7r09mQLfZuYu76Nhu
qs1STSj+bdYvS8+52o6GmEHw/I1w3JOgvhI0iVHOal36Jc57YzssDSbNu1F0lVqIGUSi/f3YvhEn
6QkU1wOvZPlSbi6t839n0bM/LRMzqBGkh2KrPBWEg6hFUAlkVgHLSQW2Bp8DEfeu3/w7CHqko2z9
oKgF20iQ42mRUgzQXhvkAAFUa3UFsyzE82V2VqFm69yBJUHtzlBwfaewY355AXMkZe6s7Lhk83r4
xYtih2wDnuxy1yKpOSrQ8XewKY1dFdg2xseXW7wPpjyEtlS8mrH1RqKopOgtu2Sh6egDZCsIownJ
6o31+6zNCVmxDCQ+a4NQTtNGnGHaewXQxJZM0aH9rmeNz0XYX+9JVuMTllCtLG5Pom8UgsPniU95
xuRoxrQPporcpC/9EOtJWZ28EXg2RQl/HfOPi0+UxhR7QbMB4KLecxoHNR9izZvOddHs894Mqu1p
s8U+Xf5RCz5sOHxAOSGcOe6h5/2fdYl24WPwcm+YyckZmw3baCNJzDIRXx6elxxmUtgBSGGL5o6T
SJPvHW8RRBtn31h/jwiNTfmAVfEQheTA3Au9mO42fjLeD6CC84q9AeUdIJLEvlTotOfbZ+4IMGtX
Qpp5iGTZyDKmzN+sPXRjZPZYvb32mVz91PkuiNt1xH6iycp8mVyh4OKb+1L8VgTScN6ewe9TpHWu
iWVLGAH5D+8pIbxkOLLjLaTwpcszs6LdFl0fbcldyVgcHsaEuqYZGm+2tBYsFwgut6WzLggfh9Pv
SA9Wvg78k18J/WJytaGIJLOUoWwUSvyqFHhZMINHOOMxWZI175fQ9vlucY2c3Q96s58zw9yFxDWA
kVjKx3TgurTZlAx+mI5tmfjJJAemVxRilAeZi6CWx7hnDUESt3ETgXvuAlPRrpvoMUVFjNTkuAvf
NKTz5GLWS0Ag+p7H0b9OKgCaw03U+euLrqyaQUi3XJd9//kv6IP+hW0nPLOzuAe2+Ee62wHRxUvj
Gmqar/9cFjI9XE2UcTZbmQMJ7mR3CkwoT7PkdRWxUa6tbnuRQQp9UUn1qbjM39iLDgU3YlJvIyQb
WzVl8MFaVFcOa2u3N9G9m/gu+ZB9Cc3QtWJVas87I4qWXsY+VO0418hz1QUAca8IHVHOb1bFTmDu
IgKa3DLo2L7Ql3uh+MuRwoJHMrR5fDQGhsKIL2a3fMxyQfueIidpqGiSShT2yLSaqOFyloUUnKsG
cv1ca4emu3khFBDB9GEmXNarAv31geedG0yYSlhvDablUUdjAM0TLjKwhhKO6FfCZKGB11Tp5xRm
UUQhwBIkNfUCVO1Qp24UWcAEYsGvLY9gzpWHw7ceHSbRUB4o0H4flEjJxmtNuCo9wxM7oS5sDeU2
C0KoI6F80kvgC7IeCDxkRTtRtNC1s6+fLvKP/2G4LzW1NmztepuPueVk4DSh98uSzb1vtq3+WbXI
iIfpdWHm0Qr83LVd0uX2C09Xt0kEAq/mFPSiidohi8hE4y+Z03sq1NK8Uajk+N3NJL3SH2GjA2zi
VNEfyuSaFNmq2TIq20T+WgXwvBJ2g19NHb3ftct5JwG4IB5zYFcWcTJhQh9wtMNfVRq3+Zv+ELqQ
5/GO6s1GzQt78p2dVpEt/Smkl9SRi4JAZiu1ezN86n74UMZZlg12UD//awwSyfep8QPEmg2LFHcf
C502VljmLptzxLIN1a601dmdTONi6+8hVRaoygoqdi+xJCgmKBKlV8ufLBCgOhatK0+KRHIxDYam
SDMrAFk4IY+oEfMEelskh6pvT6o4YJy2Sn7s8yjPBhyNeZfPAM9yxw9KoOwNp9K1V+RpYjIC7xB6
W5GqolFPyXYT9Bj/CjhWGqJB2lTks8F4xlcI3fDzjMgKfQZDmTmNYBmf/gnwcNbudIH+OwVmrh0A
o+av3i2XpE0HCkazOYwksE7WeyK0nBquJqMsfOHRHKrHoiS4Le38RcD3HrtGJHoU4W9//ztgf5GE
PdEHjjJ3pZcUUrB/U8JVJVBT+5V1Oi9F7cIVZ5MY3cSd08ZURfqpp7rRsZv5voYETKIFKaJNETTF
nLr76PSTnTShWEb4p5IE1cxfvMdIsvK2xV3RmQgsUzdzXDs+EqZ9cr7ZxU0JxV9ldFoYxqM0SoT5
ZbZdbz29bbeTxzZ4p3yKlMRE9kTsftwsW5aEtyVOXxbK6UhphmAEDPhhKimp94u4d/XkZdf8U9tF
9/7bsLxKfTaGFzpcRGRVXV6xZuHnycKjlurdxbhYWWKvAUFkCKlz+Fq+Pz9VDyA8iTNCiTrmJZHn
anY+1PJfM+VYzoaZVPQzaOU0kBTYd78Og+29Bm8x0imM1xEhxVo2wqidNtAeeV6J01oNfH4JC3Xq
TJ3Gww/SP3egkTw2hbzOpu06b61FLlX5fnZi/P87AlP1bz3LXjvnT2TW8q5vaczIaBX0SlIbIh7T
fo2NicyQ0Rt+c/iCeGaqjLYE4BKBNviEbvesl2vMXapCjA3KCGboizmL994xUkN6RguSUbYn/OMK
dmki+UVKpbCERZBtACBShlleOL4Ml/2lDPeIucjJf4CcUB1BpJhfLQRmjbsPZEiq3M0mVGROjvlm
16zGK5Y7S/SEXzqH0ieLsIUVrGMweIxpNkEw0CpF2jMl9evN+VmP2Gief31zOKb1g7GRVnZXA51/
7X3CBqNd5Jcv/6CX8hlQ6+AAbc1YIdcUfySepqwADh0StzYMPA/hQZhzBFfLJs74Pn43Ed1tb3Ci
Q64x354WptsYmiAqSgKE96sWIT6ANUeXy1KFX520eJhZSf60uLAz+f4vBjXgn0A6Teu0TykdvE9L
y8US1ZZZE+wJRbKubR6frrBXmB1iX3pW0Z79giNO3TNRCWVZ7BAjC11tD7M09XB9ddZSz7M3fUXK
3Yr/dnAzzZCAV6kz3iZEfF4+GdjPVMX5DQoVGNI1g/lZTrRge/dX+PrjbB6v6dgxlEFg7LIIoz2+
aOLQmI9zg6OQsGm+a864VcwI4yV6IoV85TNyQ+k5NF7YHjlMDZZtSnqoD51EbRAtISmRSCypADGX
00KnLhM3oVrXaA5hN6iBV8Iz9Or0c1IcDx1xEXL2X74dx4z4hophcw4T9ewEejHSv0tKN9Gxy7ND
V2PqDkdc0mXr8Rr4B6o/ddHP5J5tWuG5hSOzqv82h/bJQYeDHLeqMeVZ+XoNUfHl9nIS5XMv0C1O
TdpnPXeRKNLA8zuiU94HK6ZOrP+lhMV/1qezf740caOKllqV46hsAAhLELpfGW1jOv4fDfkZJyky
uhDmiUMrd6xSsjmKUd1l3vpohb7q3BkR2kjbOY4mrC8+qIl13lP2PjGLHJk1spAbfRIHlfqTKeum
oA2v3izi8nCSkyhMCG2ZVy168C79NmuAwcqN+1ZIEM7f9d2dpW45O1rx+blcxYW47NWlHxEftAw4
g3QHe+C0b1kvL7j16CwqiYv0WA4u3jn+hWoA5gcliV1KqRQq9XC1u+d465vqTnapaQvGtmVxgelA
/3RyS/Ay8Xbvt8Zw6CyaxbtyhcLOXLeQYBagi1bUIqQaqRlvCN0rAPSBWnqVxTqilkAgxEJN4TGc
M+mn0GHNdgumICESrYQ+UWjbDO7cXyADPavH66wZdwQp4rc2ubl+jHAYVpFTZFPEjESk0sUIYMDd
BKdgOaNpVn2Ay+6UzZMgvdPihQ//sONWjDitKFEzrLZR3ICd+f7w+4MRJEM8GwTqRq8L7b2ENYrz
z/Lga1enYH9bM+Td44FGKq9DwbQmHKW7BEx2tNttLZ7A/9771NA6kkJ3PKKPp1XwU066aL3Okwt1
rUyWZA6hMECYOr/VQ2GzQbtY1BX/Py80rbdTIr9cKyWDP0oLzoch1yVm6tS5bwqrHm+Z3rLpn6x3
78aAMN9JxldBwTNZM09QW6OfrWVWrvL7RGY798fHwgab+ZiDtd1C88zolPyxoVxCbmUaliUNGX+b
8Btge8eRW8/g/y+iXO4CJzFXSajzggeaTNiM0kHDyBH13FOqmxcVihv/EnQrdaa590k/FUkyyeL4
F4sgwzXtKzEVwIrMkWIMa71Ujdl1xXL3ryGXusQQ8cN+3e3/K4TxU1G324ocUe+9dOOOwNG6oiRN
n6Y5qlHVokfd51ST+rLMiB1l4vl3U1CwHe5QtSAec/1Ut/QhJ0D6e1VrFmnRiSouGKe6Ewb1BUWr
JHSlHJKsoIL6OM27Uhl0jfy4IRmcaNduSZDF4RlHJOqKsZ5iY376Uo7JNmNPJkj6VLB1mUcmRsKA
53mnTzySKyytKdUX+q52cokKHnmz2p/6zgL7ODPiMhzN1uK61Rk1T0e9tqclfseWv6Kt5muDlCp6
DST51cKCEdFcRw71c1vxXxP3P6IB7k0PWZGNAd3EgvEEl0bmAkpOy07tO4k2tRItIExZEEbV+lfC
9txXIs5qfRIqhQca+ygtxA17EnbEqpUbmQEjGlweCADfYRDbqdSYKkK85FiGnrpaLx7GHOfPKn0u
H0G4QjGKTaIzJ6xrU+dNDbqnkQacXCvuUlI+vi7XGGAA3ALpI07EbVn1JvbTXCX/jExhMyjRrTJE
85+XBTlUYkK5/x5zc2Xfi2ecjNYj8T7+yuxCTSk0ZO+ODrdelZXGQB02/vbFOdbf/xb4jeRtSuY5
Fr0/vDGej/EizueCd82Icre2NevqPjWrl8JhhOBoslorNTfuwJA6Rrh4YJpPWsqEdnPE9wnBXY5C
4hoDLt6jIKwPBBxl/bcOTj/QS+GG9n4JXJVHIWcVOKaGYj6VPrvAHRqFGqthqZvCLPX0Vsj3rELt
B3spKr/1EeiQFsnDPCID0VfEgpyMcQ5t9sUiX6pVJBpR68a24QAtdSKwWIGExrdfo2yV07p3gD2t
wzK2o+a3Xyv2Gu8FKXzG6ogsNrQ/bkP3m+n81k3JCF48LSIQpDSd+mcY8sBJaoATQbuMLykgI3Pl
rmTc769//J1mxJCTJhBnH3JhOwhAwVleYRLgnZWAw/JGTsVgM/FHlLG+I13plS7td4plS7IXxlvW
hJv58OTeiwqk7NnTJTRZrkJjo84j9fSP+ucdi5NQ2coAN1vcC1NN5dLFAUJ+ZyK1lvFeiYa1jbQH
ej8EKBc71IReMbK/G06T6RBHaX/oE2E25gSGOHIzZgqgWMukWlXGgTpQVMyAxKjC5ceybUOxgdwZ
4JYwFHLPrYBYudX5iwBUfiJhQQQLbALrUeOGs6eMothYUpQjhIhKKvMITmQAcysA63HQ55oaeCHm
igMYCyipOk+kCpgORpDKbdY1dkTFinnkUScmSF1NKFAFDh7kWAhuVSQ9RlVdJvF/yxzeqAusnk9a
Ww6rPOcxg/BX5b5Co1+vLc81MD1Jv/gHoI9gRkhDFBIaaEMXGFGmKZ90lK6A9AOTa0g9qImotTfy
n/TLzmloLF/VV0HqDbz1eIoj+0wA6/aNrYfmFonzSLFveSQc4M3fSFFvsXicgFsRYuqnOxA6PIz4
bChiKqVNq+4Jv3fpwFc/nxisyUXBXF5+qk0dgoL2AO7DpeBump5j71sOEtp6ggOKqTRxujbfupNu
Fz2en9HAUG+j2RrCMwmyKXKW7eivUal0A9UpUO69CoZZBk1dKr3Q8eOwWrzqNaQkUMxin9S1B3n0
Aww6TEPG8a03K93rKYy551icBoBoTvGjKtL9ZJuUd3P5ohFDwo0Lg3esZR+HynVb3f2VoNMBJWw1
MB+FoMTWdGE4w9oaXw9WdZaIKZJx9hp56AIqNIlTupsZmw6m/ZN7f0PLfarTqjpBJXwMX4Z4/v2z
qQ269AgsnxPtaTFHgP4yBshvlbicsJFUcPvJTgy2rRZpb1kDMWNbNP9ilYe7yZr1/8tDsbrtJpQn
Ut0F98XmzNqs+VieRPZ6xEXxUKawOFsHYpkVTUK2+sZHe/N8lthVHhY3qv5FTgaspIO+FEasq1JZ
3UPmfN/kkuCbDHQgKi8zw+xCBd3OHNXKhWarOeFJ2ghAcN6nqTpQCm5ULH3NbDnWKVx6OzDSqHQx
W9pd4xGdanludqtUo+RmQuLJLbO9rFAmBM5928J8bH6gLsYnBFMIxcfDXFJNIAEPhhMfQ53+UOu7
7Edx4ZYtdlJTdx3ILT1uE8KdmOvmYwszpD2Dr4CXF38VAeZctG1KX0zZUcRPPA3sUwzRJd6aNzt4
YYthb7m4DyK+FJlBOVi9MzmsjNiuvQMSCzyqUAaNP8hWwE0aewIDM2KZefcQi0arExlLPFk/IZVI
LDQOGoCtPu2Fs+yJLpo9/yxO4i51Mdk7pGe/ECCVALtTdcAtftRyK0Pt8t67i7hsGfCy0HUPLM9Z
5ykJV1gPjre9jRb01DiYauDx/LsjRtsSDLPvKPzAXNzFap93iUxlIcbMjmTZYuRRZvYEMWSuVXfK
sVC4IZ/p7OgZzqpZMcUjJi5UuyU/DgT/cKmi3fwRApUrzMpTjDn9KKaSOCQrNuzHesnaFjF3nKO7
8titBHeHe2+h5nL75FpN0Nmng2GBsDpYbMwJ0V2SU/BAOe8mWFD9TU3fMUw3Tx1vEkQOcTapVKvF
8AV2in5mKvI1Y/hKZL01/oJn36CFEGF3bQZi5W/+ki7qyVQTfafG/84MXvbuaZnQyYh2BvFWPbBh
LMuyKchkA2gJTIpDj5RrDyjiDKxixBj18kePtFqhQvllbsxlbR1xi8eFO8gTnTD+0bLaHUwXSjjK
Uc9Avu4sOSht5cwLfmOwNlwIMqD4hbx9X3iAPZBLyQr6HE0wJw4dRWZlYeS7kfl/bXqEF3KCAaIm
FiR/zXOjGpL/kGojerxsHlxqFymOmp6rHn6PSOZmEZV7yQaFB0sbjDA97KIoBLQ8BSyVLS2KUhzP
kfKJ/aY+F5G8zm/n696CgZLPvISXEYs1uPCekxDB5nJzEQ2tcfw2k5gX4KQEx/0y6pWF5OFr5eOT
MutStAA3wgJk0COZ6CS5db8plTBz9NMz1bWnOjZtXvp0xz+/Z7JkpnDS69KNjXKG3OFh4yCtrfSh
GJrPww4coL2JcvnRIggoAXJCAvaYK+NzkstV7D9KHEFlmjF3Pu85t3A/dE/rXxQFX2RQ1xfqNKyT
OXugoS3pS438tiA1nfEAJgCn8eqkCU3yHsu1+Adlp8Frd2B9pe4ROJBfkYIGMRfIvU6ABkeyF2YP
ANUwp4zS9pYnOUA9x76XmGZmUfIm8WBAb8NCejKIwvb1mHkWZ5CSlXzQmF/CyZkzZLOq3erx0B7U
w5A38kqjOqgAQUGz1G1dO9nGlAz0Qkes8C43o8K9PnrIo2igSwNZP55RSw+ZqM6qvIzQ7KbgCpDO
EhsnDTDHt13warranmj9TkJ5gvDvX1yyUWoojLgma3zG5aAhla6IOvZtEeuNJiBJSUS89rOBxaJS
7W9SwQ1UC7ZlOyuf0wWeSDvS2s3y/q685oWEqry+zWwG38B5E5EOHPhmjDuqhGy7HmcOxEDMH6jJ
nyETEMcc8ErVJDfrwXjk4IrggCAhB4cDqfTw1xKFl2K3cjHGuzynWxx0eSTzEVgeNWFTTg5JAdrO
6rRIaywd2DzrIIWm17Wuqun35h+rhuQfzqq4yS9fvG2yYXXEvEnqItfbaU+rryJpnwWxLLOsivve
GXU8WmJASjE32bL3hoB1EPdksrvckMu2GQV2JrxVkyA2KKI0/TruM3iefaWUlwVdLvTPsPq4ehas
23hRT70zZ1PmBZZd/K1FkSWP+Zgd3TIrTrrXdk/Gfa+bPP1eBt1mO6iOgfY/0ehX/elu+qMB10Er
uB+m90mCyI32O+7fEnI44XSRMNPhp1gCDlpg1rnRacDjP027s0aSeIBqozk5n9ri/UHDhlJWVChu
WiOsNKMCzeP9yZy6cggpxcDvy0uSjzqkSS/l/JcYudg5aaT/+CjWfmNxwz9bD1pvgOAVBx0dqi85
Bf0xbVdCvPkNzc5Za1Ihau8HQUItna2jbZvxM2SVPgIlE3Hyt/Ulilr/wvIZwxjYPmCuexvcj8Hr
V9cX+Rhad/HAAWIdpkFZtoinMDCKOBB5dTq2J+EjNkfNJLjN2xWaT3BHuxm2rdjhcaJ1KPlXAwgd
Q3QlNMWmECjwpC7fhqHSu6XOYQidl0iuxE1cDBzOhwJdp7Zh4n6eWRUOtON2BZOM0ADWJ7J9Loyv
XyGwsNSdN8os8BH3mnaMK3CKw719fBj21BYD1QJStl7uxdTlGQp3a1rxxoaeUHbD6eGtQ07ewoQ3
35rWTTALEjOKpqQLYk/N07d5bbRm0s5ZU9TzTijp5huSMV2bGoj85JrLa7tbVv5t9BSMijKiRdk9
+Pft9AFScboUVgD+3Z2TNLcglyMYYznpUQho1FX9rjrjR1WOGeI2Lay5rt8ITC+Leizmvw1pw+Ja
y8iCrutGw9CxzRG/FbE08YBZ5juAzu4BgjOHtrIhpgJuYbgS6aT0l7fqJqADWdYlCwvtsE2nguHs
ULjxnV4AgmObTNQFOKfv5iYF3meXriHBO5OxA5JpTE0S4fMllKRFxAM2hGzYaNv+c/JGG2gWwgQx
Crsw8s13PKRQzVKl3Ndi5AKyTajTjsGUY1uFwDjO2VLx0k2yhcUL3carPX14mPnkd7fWTi/N/qE4
26X+U7M8MrZ+++3X1h88UmO1l+/iwKPf1XudIX/4XiWwNlqGbaoLlwNn7B5LEtSc9GK3mpAiZt5Z
LjoenMY2kZZNb0yTmSLemvB2R0Fke0s9ML8TLV5AUYd0ZcL1l0AdIQVz2Ax+75QDxrOiSDDM7f6d
kJ4OJk0A670O8d6M9/sK5GrdUFlWheJU218HLacJX88Wc4DXtJ0hfQGDXldJZePixl5vlBdSkYhX
qMylX47ZroNK1Hy3TnsrvEKi+VAfUqNutZ6E/2+DJRR4WsrZFp4RUIMTgfEnNMyehs+7qJ0BY4Qd
HoDczcATsW0iAnm4VYCGmqsIaIOSK4U7ZGlE7uOA7k9vOGyYZIghkIf6yokfFPdkCwPFQXSBq0Tl
wawAPXWMzM4tQwm8vXI1WriNp3bUOi13hfwrBu2TafdqabpD21mqiqh6LTO60Q1f3AJebfh7VEDw
IxsdfTggVv6WPD9O36q9s7e+z/5MLwEsW18o7ewYDuyvuAN2Dhl5N/Db5G91xQlpw1PMXIkjHq4r
G5SrRUepooQnSizUI4spsYNO+AQChQqNdCx+mwTywWh6XHVx2HOWB65AP3qYzkw4zzo265Cd6Gzl
KMFXONMRo7TmDgp73WviGOwzdqEmU0yB6CN0QYVnpSdmK1tHpdNEDXsefq3esDfYQgREMdoY9w9B
dschgLzp+y+OhIKBuXQtNHwQEWIapvFLGWEI9wwOLkRLJJQzRopgYEOnQ1bpk18cij2KA5bXa7eq
OmIdfkYNbgetgQYW2sr8ZnXsKpgA8arW1hNOSyB0pJZeuTsdPwE3mfKznCkfTBw0G6RqQkdon15k
BKJ1GBff2TTqBi3ftYrTxF2DieHxr33JyLI4ctddJzakpRE0mPhr+Iil8NyAJ74WzEeefpraS68T
lBB+JC6mnht8glvV+lBvjAHmhtLQNH9040tnylHrWJ0KNMXxmT6OGUc77dWgCKN5QePigpPNZzh1
o0aUTPv472duX4MDx4zmWrndRas27UDlNC18JnVx98wkt+mm8ymIjjTizaeaLpeTwgDo9H6SufzH
oqpSYrEu0cK//BcPqroP+2wEmbtEC1WFLkrjgnxJY7a/aIjZWEl2Gn22AxeTTShyDJD4Nk94ixbi
uP5tjPahbISmnuXeM6C8hLxPRIUH7+jfzT/JGCwwwZ0kB7hCh6IULWDBiFYRyxkUhBIfdqw3HYFQ
yd8spbpQQd774FC6L/Nhte9z/IQwkWKDaxNAbwY3YuvnmMhlWWGYKKHyZhu29eKiDKgysPS85r/t
7bZD8yz4JUQtH14mml1m/WM+0Vji6etbeJ3YzX6ONiLBJs9jDjpKoyrhAx3Ee7GLEhrE6h6nIDyp
I1QsvmGm2JBVcpgROi0gHh91nEoOTIpZB4Y4c6vVZEZreFIpetu7waqh0UO8lfC7bx1lgc9ACwFH
STjOcZmyAaprQobvbNMPEx/lGdXMpjem15Jl2jhmdZLhRm0VzqLw3NtI4gXc4vn8i2yi60Wd/OCv
R2Mi+/pm7GYab0PVmx/o7mHfOXOxNMfjPePuH1U8bLUymce98yH94HQf83MRRkMlLMtFr8IoxkYh
EU51r4VuHNDBxm6CGEw0i2pzhjcxFbXCeBGQjoaSavoAGuV9L23CeYswwUXpEnAgCUPwfq5zNFBX
KEaVNSMbeSQ/JP0UxCTImbD8XeD4MzmwEj3HStgqstCYYhHO/msqsijuD7NTBg8TsVRAP9o2P5HG
ZrnieOn6BjQGjODz1uWBPRX1hnhLpm1Wy2Kx4D8QmFlaQYvAJ3XqAmKqdDDpeRpNucw+63w5WNyq
fuLHC6EPZp6HMcbLjUwVI/6XvDP5mAiguApDcxh5UnxUolvSyRa8Xiwxf4cQEagkqiWQYgOfOC//
KlsIuCtVvGGLSnthTC+Gb3Dr8nhpexKhkT6Ibn+4NTM17lN30WpiZHIHC8txv/P76tivb31zdmia
WcwbKvGCeZHdgXa2Uj1iWnuNiRRDIRZ41+GPU0vln1qdW2qxMdWOJIkDtxnIl/cUlqgHZgPCydrB
qPVP/0axR5ZptiUpYYF4RtxPoVlt6hGbJaY9Hp6CLs4EmXzihsZzSgLljMr/jdjqzc4hyi5xqRWJ
m2AlOKKAha2Y85T+HPfkIxJZ2efoF7b8djsR/YhLa/q51E3OOdSuqEltUDxOzGzCfYRYg0NJil5s
eJ23wyLGx5vG062sbs1Skx25tl6Ru1jER2HVng5hcHs1zWat3A6W9LN9Eko5bb0hGy72vGK1pUmu
/Bna2PZspyttxJ7MixjV44wV4UPL/ni5iJ3rt4uMAQF6fm4VFMnA1o7OT+l25Pr4F3wXBhEpo35A
Kyq8WQWKxx+uYTZEpxHCsHa+50ton9hcfEOMeGpKMNaxlxp455kWsi4icg8n/ZzJcPGQFbbdsn7r
8rVDl5C0EttJ6bjY8gw8QI7d+fed66EgPZAzj68VhSvsSPfvEOtRmW/1YQPvs6JtJAyWjUaEk4i1
8tqZYoelpiGXNbEtSzS050a3o2Q2pZKQxdb+6SQbeA6IevOWn7jxaNjYIFAEkZqZRj09yLaDPFMM
oHG3O9BSIUWG9BNiYxWD+gbW16+r7us9z9Cf55H0BrT+jlrligi4+44jamSKnD8yoKyiukr+Qa+n
UTmdfLRKGfgyUnQaCYo+/NHqWY5x1ffIj1szjZbQuqQ4oHqCikAcJs/84z0q7PYsvHfi8cCwJ/Xn
PLy0/xv9YfAGsvC1K07JwoZjet8ahKGmMD7vLJ5ne4+cT+jQCKa+AZEPI6H3zHXn5eAFMzRj7ryI
52kI48gQ7vAbKj6inK1w4JSl2HvaM0TRyULfWTMWt5l+Yq7/iqWTsflVXrNPp58Jm1l82soeIYaJ
8pWil+hx9KNp9IC59LSqHq+mlyjoJy3ab1YT916/TPQjj2R9u3jqepHzO6L05i2NSOGtyv2/SFxB
ZNwOf3Un/maFlxGjjbbfEt74p283L+MZOCycI1FN9KMeafK9iCBxRHln4gHHH2jowp4mb/rWB4fQ
Fxuedr4JpVtse1NGk1yFVMergdwksy/5njNs6cJvTtbdPQkbL1j+JogAxtgrfIXdfk2m2FzFenqu
IA3Gp72pgIZTHHeODPzzJ0DemwVsxa1rdECeS8vng9I1EuwffLzpNWjlksRYO5mJHQtI18apn1cC
7fA0F0D6M3eCA0UsiPUo11pqobJTRRsfguJ3zOUCNE7SNmvOEXwAfKJsxAlJeGzVwlWtAa8f+ojF
2BnnZwaT4C7QO039G7ib4s2wJ0Fwvspamyc/P9vH8QriXhg+u9fdb/xEiiE1DH0TAfndIauurafU
Y2W4l4FTjh8HPBe7W4K1db+XVTy+ajUgAZDBIjmYT7ZP53zXZkmyrIK8woQuY42GDrQMBy/wN2K2
A08Lx3ahZ8svEHUOmovujb1L8OT+C/9WIiQAew8/8IytXcPtSq5HLlgwRPRxJq7ikmOG/pqzaR+p
w4QX6Ztv8rOKxFbHs/QyBtCIOj58vHPnjFIjnmI4Lim5spDckBISh0GCCBI/57NJvfPglir0s8LY
7EM3j2SBQSEBZGlaMnjGukBo9sc5cEkmdlq2Fmijg7YULlPQj3mpJrKQfVOGO5STA/Bzc6Do6Juf
Tv/a4z4TLMAODAPsnP8iLYx9mWBG2qPMgSeh16MvyDjy3tBI4AryjOFGEJC5ABWjPwZRBVygD20j
ztroabbHG3oUbfnbfLPp4mFVxvglG4EoJV/spklvP7wbujaieHaSrkcOI46ZTbGF1cqBiWjQ4PJp
yGPoFkF+JwwsAdfbCcW+iPBOhXQ9/n2+K4THlcnAP8Y0lHQcD6M6umTwDnVp6fcdSBKoFnTkI7fC
Y6SbKowKyQAphOZeOpzT/wPYWZgOCRX1+Odm8hh0XvsZCkoIVuIDn/xUO2stqECMk18m1aEfl0o0
5nNWzaJT0CSdDZYyA3TYkUxZmMm3xuS+Sc/vUJs1yJ8nAOwXDfdy4zlk6ftfe3uHRyzw2Tewc848
j+GfTOWWqxoGzdYw+coLXYgtBnYHv3n7ByfqqQb856WWM0wb5jPPws6IARnbQ1//uC5rjdI0dsDI
HZA7c7g9ItjFnRmPApbyqM/PZl0UxBl6I4UMNI8XELqwG4Aw5IUBfs5VoycJI+uE6/FRoI/snbys
i+IpDDnnS3gOeUfT7WjnkOwqNV+3vQ7+YClew82Kaoghs5Z0oVdRAw3hTuT9GmULbIlq1jbdEVFw
pA/KB2Fb4H9y4ncvUkUqufLlbqhPOFnYrsDjpiPQJj8zfrOiGkO2+rpQUXaZ2fS1MT7sjKm2wVlK
qJdrH98Skzgz6dwLLrlRY+yAh29J+V2N6dP/pJdX64jZQlH/9tj8Xi70S8SWjSKSZ+IMS/Qwdvyk
8/xSXHvDlRo2jfnjjEtmyL5Jk2rZ4Aryk1fdzRFvL0p953un2lE8CEq+O8k988TCPs8pj+BvcQmf
UhpfpxtFfsa/nxvgA23hPvdyoXFDRpznEg5gC/UnohjLeCaane/j+Jff6X6DTYZB58wJHetJ2jbj
3Hr4crnYMD2DO3Qr7Xu4hMWJ/8y4g0DS10+dU7h9tkgYxgsHLGfy1f4v8vkbSJ0nFO43B2NeuBi3
/gz2/kPHUUKCOcrIi9/eBqQFiB38WDuLckunNG1dH2kj13cTkzAdBuNsb+qkY4Zz8llmoXR6orVw
NBtSoBW6oa9JkKYMqEqwWWio7CWzmg0L/pwfdOrsxDy96QQ8bGKHSXfpWNVmr/hc/s1AP4AGz+Am
tKt9xARaBWMWGqaMEwQULrlZNpTKyA/LTyJ3aIYq+8rpEiLd7t9OD0xW5Xx6OQfuLgKuQCeCZgF2
cdrIhfh8BRSo1YFgGuBEJgxc3jBp8pCm5ziK2+AnpEkI8bf2FkVdslHHfjdebEq+r8o5OvOKvBIz
T80Hb4hJTdhUyKDfxM/k3tazfO16CfKarp9tj/qxDHjzZ2njNX82AChPopDL/KYGmOCprJdE5TG8
7JDVtt1xzrsl3I+RpqSWheq4Cw5upoVX9fr8oPH0kAHpaf7GhaLcWXLgI5Oa32m1emYwbW0d3MG6
aHneFMCMXLMtPsWcLSYvUv++8dWkCXJyg0F/dfCjbhKGT3MmytpFgom5ovLUy+F7sHse2lqRbnSt
+Mny2jmWNCBA+Uy1Zop5AGTJ2vw30S+25A6lNYCbrKebA/ZMpB6aRmQ7zkdwT29mdQNbrNDMTAp2
SWCs8CGPuljjEpxo9WB2tO5CEmj41MiZMupImmeFZNmAJiTQXJ9nRTFW2f8j1SPHnkTDlzYd3tNf
Btk4ZneFjsJCOEF1SxZxwDTsLHcSgGeNMBFrOfPk8+VtfXOTivPC3ZGQgwkpJgcgZnga36SxAunM
PSEfpUhwpnRCeVirpYWbVUuGQl+oNIVXqDHUzw31wx5zmiyaN3ewNNP4ZtKgPtqeBiGTikn1fZDR
weqKsL+Ui/emu/mExOMaqIP6I0ktQBP3hqtSc83StPJ+Ec4ncKdN5QQnYRl26sF2B4768RBSmVR2
vmUyF8u6LLICP8M1t3l8VWoUuIwz4nwgNhf6YycpK5qRRYnU79x6l6pydKRJZG8XElZtXU2VgxCO
xIoHWkABEUXsocHI9JDB+zL8IvjATlUoOy7uN2ytY87F5L60MMBMc4g8xg+PPzLSecLIiz9jUy8T
J5bE5DYD1If0wVQbIeWq2bnhgYV4eIEXnsuZmSwFObK7kh7a3tHswOqE8CoZY7hzwtt350JdwXCK
o3e+m8Fj+HBzkEA32IDfAcdJNm+p7ZpXDThdO6XuJ6InKvC/CfrjYYH92a5jkx4pE2N8jbtb4qT2
un4aRLJnx8HMqGn0t9QBU9CW14clYdJJcisFh0BqaEXa8qEeMyw8A0pNVDmhJ1T1rl/p4wn/jzkM
qvCF5XeRutV1ZKO6rnBWPsM7OY0XpYzNMfWuf8s6n6rFlmTg3v0YElx9WHp8PpnIWsLUlZoTH+Ji
TwzWPJNJoiEhtFuHYxIeQaK4ee4OzX/MbZsU1azeSO5FgvatorGvlzoONnTVFGoR9+M4DPhQBIVY
vXfNkkUshBnEjejA7tV/aQgsoqj5F4MWpZhyCLMgncH0K1Kbz33+dGPgZRWLJmzbG+uLmOQnkxR/
W7w1OUHl+WJmxpQfv8bT8QxNTH1+FXVCvUm4IMEQPAufwMLmVOCNw9DY/YSjGgLrMRjocuFOjYYT
7K2O7djHQxUbHb5I8CnjAMNf2PmY9ISKtuWFiiR8StK7tZeiG/HEfciqct2cumCmaU/B7Z2t3NYi
JOCQ1uhw0TeEFMfnk3Rd3s1cp/kvTyahRcwoYcpNeZuFJOtYn+20IaZbRrvxum8YQUpWVJSBLw21
KlSyE1qOVVum+UTX8sRqHIE65TGxO5ndDhfy0qqjOjODo2aOUKaDD2OjAKN3KCC9JyggeWa22Mlj
hquXN3IWrAclTzdJ3x/+QWn5+Rfn2re0ColI3Q+WC0X+CshG8suJDFixqd62SvHsf5xjiP3fuFcD
TPvKfslumA+vgqf4cqhOcDcJVZyxYWIXkCah+aBvjkr7178PcEoGur22NqsBXkq1wxVllTVCSxVW
O+ZU6Z/aqwbpqQ1aZ9l8SPV4i4X6ehUqyXdK2FXuGTEEfPz7kgMbsXQ+trZOBSx8gxlosydzG+Or
WOPmEqEE7jZBCV+po8pN87o/TI6TwMGvYUxuC3yFxaTO3doTwEC2vzrHc/wgexGwFB7LqgbYf6Gs
7jFnWGW+hKHUoQEpKkEcG/r8KaSQf66qQpQaGe3pxexswEOGVUFqMCT9bmzDPUQu7wbzn2XR9aPr
ShbhkKkfUKXjIvRaiRJH95QohpLfuQf+KXnHksWIL9DFiyxZcga+LJsXqpdOa+17MJ0ZqFdZJe3n
rFbxcmBw5TW/lAeMevNPeLQDUbfs8N1g9dxNkFH0yt6MpHv6MiZ9oVEzloev6uQJj0hDPuSRNy16
MKln7v/G92vl8USMhYSM9SbpOyIff+rUddVORPE8MZC79rZALyoOFKmOI9DDk+/Ht3K/6tY6pNwr
uyYrPLTMJ491SaYifmgfIcFrzu435TdoRLU/bUIlKdihu4LHl5ipATzAYtJ8SSj2od6h/vOHDU6n
9xQKaekKgHykMRTzISHlnljf+0m1+ZH9h2RaqXBXEjZG+bEnk6UGs5WtK743/aootw1EL6JP+h+I
DdugZ9EV7EWgq4ucvr0AGtL5K2kgz+JDFdBMkYT3Z+wlROV0pQqDNMT4OqIDYcIPdiFX6iNe5BVC
yuCGdyW5pQmp5DTGJYNfZ3/EDDNq/8wjUtWDigVhO8dJ+tCOQPvLMymQOzsQuNzD33yf3PW8zan3
FsGsgnZbSto6Y6bG1bRxMFo53KJzKLbEqDzEX67qVAdMqYFMJ4pw9XKpyAS6iEA633wtAD8UWnYi
I/sVoVdCPBZaZK6VFXOXmi6uBk46Sdu3i59FqJX4CN7dr+C0XVm7u5r6RpcqcnvA3jCDesU2tZdT
ZZyWfFWJapCjvQKt4cePYJZQa9GCatXHYV1WD8cDs9Ez1XvDp0AD/zhZHUKYXO5RsGavp9K0gMc3
WAwjmjco0dSkGLKz5EGal/0MKI+cGzS5urv6H4EvrFCuYaxoya1hM3LRj/SFPfLtynRSm3+cOeh0
dGOE2mgl+TVtIZ/R3Tf+MKWx5ZdZzE/CY+bu2pN8y1QPH1na23YgjnQYTsWrPnl2zy5HfEJFJ8LQ
umlKmU3UZPKgNLwj8vO0lJE+bmt3XHCvLW2cXImWkxrdtr3EK+t0oyu8QQQvhvTVFCGaUvJJIkyy
D785XXewTPQqI+XbkydVp0WGIQ7o/qAZiCucAH5fnAMbKdQfCdk66os5UfNdsNXKSbon93nS9aAA
qC87RGDwFxLKh9PCv2t4zhmM1gwwXspZobJAOkVqx6xGlCCj35VetpQCkbGLq0F5COcjB8O4r8jH
LB43VjgZtExiYShGD9SU8acfjHir8TGwCL2Tmcu3Htgz/k8fGGO/yvs1YehkhN3C91PVh/WQHpXX
bdgVPiQTEOaYM6HyW5uO+Vu4B7MfVZEIXpE+QOaiL+fnxUgxzSF7Fmj1USrZz70Ii4hvWzTBP7VZ
9AUGsCNiLqJpgKG+UOJTDZ871DM1JJSi7TtZcPgXY0OivM2pgLQgZSFnK0xVWpHvvlDIk8+pY8lb
BgTMT4BgwRyTOEG+fSzuHOaU78yokY5w7hQk2baU3oKRM3Az7JfpTmk902ANwMl6+Fh4OXxJVuw/
ywMVYDMuIm2RjIjpHWYsq8XIIBrxZS0IvAcsxCK0wEtoO/+LUFXO5L5VhwQV+NN/mM2qVtB2ISc7
d+K6Uo6g9uWxoMWjT+gvAxhoP6zYFjr9u6rbWF2dClZsDr8m/eFx8llsKulFFVAlzc1BJOEqyMqn
NobEkQQsWa9uDAqUXgwAZ+52sJ+2N4QdOosUa+g8OsGitw502SE1TqrgsDanK0bWHtb7QB+VYLqc
8l3aZ82rS8CzaMD1a7tlCfrHQHJ7XsR3XS0AeL7lGWPNAl8XYBwagFPH3XjbkoJYajB3mxPwdU69
5w4Pqp/gLVV0/Bl9H05HYPN1KRcDXP1+vA/2Vwid29PUbJKr2kVAsQppz7qCN7FDfOU1/Y9myfbF
KINyspkEN0AwAhz0yR4AnvPamrxj90CZQ5JfFc9uJE94k75GIVezvaFZC9YDIfgKCcjwKmt80aFb
eihD1UDZTRKeOlxpTHXZ2HxvaoP8DZfbN/Pw7TuChFWWrc/gZGu9K5ZFMFGAIybN9teXVKsdupLS
KDa+4PogOVsBbkHvglaEGh0wkIrCZ8JJ4EjyTpnIfctE4t9ttFbWNpLnNlXqux7aJe5548oEvgTD
WsvJpS/RhL7KowYn6tYxIRMY2Ju04KtBMWuBeom64yG69ADcoqupeqp+WWONvapg4d76bK3/KDZA
Z+T9bNul1CKhA9/zPuAiCrmJXACUHaVGBOwo0ODgCV3Hk6WL8H9fCancxP17NQHWaPVeRAq5SLxg
AixW47xwv7RyslPNmwvSCICT0LuMIekTIu31ytpAAlWzlTdMFSAiL254xVxinMt3+7FuXkR4YNsm
Rgc1oMUW5ZkoqdWqjAdUCzId6z7XsFy5vOpXgI3zwcWfdSgyinuJXYHh2u9V0UhNOUXKWo29Lqhv
aj2272iWtQ4bbvywakxYqzAroY/OeyltXLUi4jpk5mwCwqObG72R6HsHaKiAdW6OtQgdB8vMHYAo
TtUssBGYK3avuUyqN+tJiyIiLGfC32b7Yii0YwSeap7Xb1CWCSKve33+lk1iDFvqnT+iIckk4+B8
6qHzcLVIpH/yMDdGqLeHJQumnj7RiuKL0U1OJP9OLQMwvBeCGbPYwbLJF0cpUXRyszmuJBV3EZfe
PBOU5zQia9h1xChwKMnqZ+wbJ/my3koQ0nE2/KDpchURPvYEmaEEmACAiCjBsvhG5lK3g/IZXaNh
Dq36ALfZxuC/1Oms3tduz41ZoBX3yUnwxKwd3e2/xgHfliyhQoS0baRP8tex0ewh3YNn5xcwXrbn
vD7dGyYTvqho/iyQGCjX47nWsyXE/bAlvwj6tmcstoiq5eVGt0JeuldrOVXd/KowkJUeV7gIwuSt
NMT7YqtIiQBEhsmUvIGOpIDuhq3dheN8OQDNkS1jY3pcWsJ8NxG4gfpaRNbLsbqF5k6NKSLSAMcX
QHE90yYoFpwPuLGTyfiM+mb/3XxUL/j9jhvVjC/H7F0KsX2DJAxxtUa9Ozu3c3lQisKD8N5cuDC9
RWphu4BdT6hlzcAfHN7HNlZFtcmnYL2MYEs74SckxaUXOLnG1uXMbxH9ZAnEP/XOlWU08WL1wOn3
fmxdAWgxksyOFoMxGVCjn4xwVYFmL837mIQc545HRXF6HlFMjnymIKhRuUFbCyJPPMmha8xQcmrX
DTGT+U1/HRBKzmweOugDIyknvRh10Ek5HabSZrijO/0Qc4MIhgvhEWEfx0szO10ZVfKekR89c501
SQ1yCoRWkjJAemDKUwqHr9gTEmxEJu6q2pEWSuUpZyyeaMoKCL62QC5OhsBNYfS1zdHmKgXjcAKX
1uPJlMNZ/WlM8g1+2mEhPvNfEdRhmWVKYOPcIkhJqJqR8spNXImIL4oO/tvEqFVTre7FmBZee4gA
810sv0McbCjjA1kC0tqlFG/4p1nTvuL+LePa7dnSBPXvZmTvdvCUbyRHRV/u5O9YJwEyPq5td9l1
Jk9XORxPLR/rQCYRaSo+r9SmyfZDDw2rHZ7Mn7tiDAjQU/70YWUbwNtUw0GxqnjU6364sMLgKFrw
ZllMhi+fj2kzgzOg0WLYClD/5VzppDs6IinXM27AOUDcEDew3swRAmMgbkOT5ZysRZ3167RPHXR2
TExo2XjGNh41Xr8vjAIE/ESn7qozaoa54lqA2w48Qz6Bbc/cb1/r82UQWF21IpR9pvi0ucsFYJBx
tk3iPKW4TfUhmUpfPnbZwKGbHrAlVa1EwNpKTDfcLnLTV9DK+whccvwlhHB60f8+BZOPtbal+Lss
PdQSPTJJpnJkyAqkKOQHeiWsulm17ntJv9iWBm61LNwR/g9KNw+FH7twtqtrzi2C5SM7CcNGxXrC
VleHiGePbTT8XYv3TJmsVlvhejMdv4DB8xDy15nPmGmmf6j4UWIRm1p3tzGI3UcatUvIecKgWkcz
zRAegpB8idb+c3pJOh076k1DEbSVJf08chgOGE1cybu96c99+LkVr+WH2mZPlut9/7g6wDB+ItIN
wsHy+6HxWI+trNVaub999ofGVgPdKOvm3vYEQLYVmwORt7fwVuJe+EcWvPoBMavVWRVkKWrx8SVN
QgR13DND1Vo6Whr8FewKq9F4l0TgODxtrJbyljg+ijI1Mje/EtiHs9zGMyh1ACVg3Qd3lJSczQRo
5+LfarLACBI9BNwtJIz4XiZnfpPK9YNNgavHl7SBbAZghXZyMwhT++pY0s+4DOL+nzXWa/Ls+N/E
tLtWfFT7sAPJ1Tt5vt6S831YsFAlv+EUE8T+Sjt3kuCh/r0hsRLn9BZ4MsIyoPDuIIyNZtXeOf85
iQ601epSiYKvSbzzeGV53vAQLxisg2mjpBto8qnFxnMT5/qxugc9TG+iYFPR9PMi/31xJes42cyc
01ARLo4guBmNHy8Dk/dSOPKyb81gNH42bVdXyyLoV9rErgtPeRcNDIjSKGtRmiQSJ88TwYmT8Oro
CpFojm9m1nFuK2k2egTzehmHC1x6m98Un+QeXWGonjtGg21paCr9RSzknm8SxWPoz9LXYomx5s4P
3N4i34SK1eovOAjYOMnwEHRZxnEvhCT1GkD7CEODBCd52evqF1CH+yW/wltpakHPPIzFLoIpwDYY
tCTs3EEUx+OkpF/9n8nVXuie202PRSuE1OLTvLtXpUtmHU0bVVkXwg/3Mq7aRoUz5Z4fZKlcal6z
w/8ARX3ziXfQakrN883uPFjWSDn4mirlHLeLxlNFq2yaYyQIYLFytpLjRM92wKsJbc4GVe94ROox
ZYlLDstFIeiDgMYam23DPWW4i7T1VRgzSproRlxK4a9u9ilzU4csvY5OFy3PqXuibMP47ndDAYHX
ElZgc2vK9u5HLd4J/71Uo8Hdp7gN3+A32Q7K0jszP5KNdtILq2iWhiCfH9zh588/w8yNqFTiqWj4
T/6xIGMepXWJgrJgsMWPRFF/pJPjdjfVj6s8BgxA/y3heeFQnICqInUiZoRu5p5Q66HqTVkvE/+h
ndwfGmwcH59OEStd8crFQGZhY9fr9wynrvr16TODTEuDT3fygtgWk42X5QM66JqqozgmX1deRnlt
+D/0x7TC/9NIfrkSRZAusCTIl8fpizha5NDd+OEpTesh6QT24ZLgZCoR54nsXg+WVsts8k0vfsEr
0s7iz8ZyIpinPqPUfFF7mL+c/LLZT/xMG8nhkrLPUq4iebcNQP5FYBWmv2V0nSnuHZ7xVv0X3UmB
s/Fw4fe+eej159ptw81DZDUcvhg42kYwaGt5wOopLVaKTcj7+ie5IoOj4Lz6LUu07VAmqpbFaflM
t6TQ/Oj7H+Z47cxGC0u7S9jHNc0BmLY9seTtjAW4gBSez8fE2OZpyIizA45lYvAMcwoe5GeYQl1v
IuJ/yb8dkAsZ2IKx8btqh5fuy4K/MKrvMVAnKFVRvSgP/yterYR4I4qTS+p7Vs55R13TPjbqASTx
LmnODoX1oFQvvkv8zkZvY3WmMyejjCH/bWMoz7PyVmU504DmVn947LN/uQhzeeVG3OcD4r4VQF4k
OXtXgsUJuuRGSPYzBKFKWnO+CPqbYoIR0wciSC1OTD1FJP1hTYif/rQYXfEPKt3vLL16blwSII8T
FbMGC3rlSst1+LtkPNS/xVDdhsd+AHoJTxoHr+YIkY8AHKhkljE2pZtaj9L7qV9Zt/7UfxOKqZs8
R3ncB9+rIjAF46eg6DkV6j3C9j1e6MimBCQs0x3SLpORJzvOLSEbsmqtbuXkvZ4AJg7rjlDdfHHv
T5Qm8kgQ8BGyr7KhfqGJhlP6GEsb5izNOIb18mupiVXSnoPg53TxwD/7HkOCGekP5UP4d0bDFi/L
QBGDERaLZ4f0Wcunz+iDK39R6P9dloBia4FglOKDfbJSJxlgS00ylNzKxLj+WlKz1swwbN9zt26Z
cht+TCj1wozpo/HLhuiHs93qEgbvI4Rn3FB4zFA9VvOPxKTBZUl2idhFNZaSgYuzBpoYbypc/rpa
Exv7fStRKF1lZMTXzx8Z0TL5l1eyp4LVr312EL0PvP2VqOWDWFuslyAAEPh4pzTKikUF6Zf2Dv0M
TEUMr6UOXTLXqM4tTwILtnd9kx58ycQBXt7Iwwqs38UIMk+LjNYu1R888HOV9hXonGB3G3oKFeRH
Eoidyuy7ALd0XqEZ/o7WON1+5PrcJheNXdX9m2oNgYztkSEpEHJdU3mzxPVtBLGJ4Ibmxu4WyVM2
9y+lpcyenPnfsfAOaOC67uK8LwmcoSe3+DBIA1oQlvajBYSnD+jtsjtTmCSzbfDR+es2ZyrRYMrC
WOgkll4/pfwSyGEi/hHoAMuu1/weY5BFSoriFZKzJnhJPbfKbuHaXtOVAK5/R3GXdeED+GbnpCfX
MKfeiPbDvk5yw60ZZGWvMS3N2IihSXqhtVAWHgRdYjq+iLqL9rr8CsbX2dp9Ck7tfZDcj3UMnXpf
sCrrNxTwQ226p5pjnLHpArZ4Zn5YI2npdJUa3ebmnnCosmX47xb1DXulFa6UeMrC6PURNdOwoZ6/
i9NS0olrmTKeE3zA9aYiw/zCOy2PsnsApLS31jFOp4nquM7/VXmFyI3iqrLrrrpC47fHkeIoX5Xm
rscBrm+Vg/IrPsI1mQM+RbgVMdeawdnlJGqJU0HXfkx2Xwg/oCKLl7gi2aeivXxGTGD03/pBqnAs
Pbw3l74pWsjWIIXtJSP6C8xg1IWxK6sUXVwXVfjC9Kbxzaof+1kErlAnksNcOGCx+CriHq4qtL94
LM58Yp2zAhygS/pcJUi89xyy7z07XL/w0yqi2CPwkN2hKExk/355l14AUMeqOaGfeUONZjDs1a3o
srG/UlwluE3zD9NGJNfVvwYFKAxNpfNlgYnQz4ERNorCGEcs58ZqaVNB2v+b/G45N/D+xgLQDlKi
vzw+lok7f4P+XMPgBq4rs5hz+TPMF3OyEp7aHo3R9iC9x0EeF0ONYLFTT/bu/34e1WMsHFsqW29d
p+OZ4BvpQfe9J5FyMCrrFmB+ZZvuSiF+Oo3TCn77YaG+a7BTzd6yVnt9vcnNBhHIO441+y2sDJJh
pkI7ySr77BIxO3eJ/wbBLRZDm5Vvf3CkKvT1uYyPPgsiZqbT1eW+PzXgcNSPN0ZJfVwsRtdNEs76
F83Dm6xL2NQgiL3KYQs6btwuDxIlUD2cXRxnd6aztaOX68KCWDffsmamEeBIOc6jT+UMB+wYKekw
KNv3GVSy5wGOuG9/yhViHDzSBT2m5XbE7Mwi4y7G2Zx2fM91ypG+xgWkax9VzvhO5qCSsh3FfMO9
xRWRAiXgqP969GDRMIc1O9P+rLHToxToONMKya3scT+WMgP9KI7c2UndGdluSxqGLogQ3jwfKgq9
fHjMT4L+0Y3GKfkVm3MnN2V0qmgOilLqALpLfTLECxkCzf45m4sCuYB1LTpwr7tkT4ywAgt/nqDO
SOzeU7mO6XZN/+XSoJEYAOZLD5yFun4LRPcx6ST+p8yAf2LvvIAN0InpP9tg1Fq0qZNg5hbFwv8D
xaEmiMp1uQb+ymxRzMC5GgXjTkhn2YiJeWnLdcdSGUw3D9iqswf2WoKVjZOPUAEgYpLoZc+cb/Pu
QVDwSGbQDX2TRXnctck5zblC/tghDyajKBWZ3NFbLNEH42ue24xJ8CgzXO+ALGMoWug2sW0mpzuI
csXHAJqC0FbOQIF6tcrwdjbYIdjmZQu0oh/q4HkXtEmEHfR8AvV0zu9EHyfzB5+z9U+tB0criYTD
8D31/MvKOFWEEkJjMxINaSBQt1/9JhFXaZ4OzV8+WF3quVA6yj92myEQGs4YmPZIHItsujZCSwme
YMIVHepaZGJO3wilLNcNq9w5pr71q/bgtoSU+aABBphQ54wY0RTl0rQUJHgA0ApLoGNHr7A5QN4E
QIthYnvz7goWCSP/3IPrDUZS41wJicNA5Uua8Pw0QFxwb1zSYlWWd1+58dzfYAbz/kDfgwq+l8Bd
ycPnvcvMXn8vGqZHQqEIobiO8lGyN+8LeZcLuBatNmh68n4H1cMwOHBDtXPUvjW/LiBvzlQvcJ2h
KgD+82tXOiE02UUFGyfkXshZ1rfdxqHUI7fcSSlr2qUY/ptQbVmBKcEtd8QEzfaNyIbNMfKgzdPn
MqxHuHaYh67k2F4r//1bVaWRj+zpEZ0bQwp6+cJ4dFxoXGUnszbCD7o08ziZtSFnRist7bipCJv4
1EQ27nP3eA3od9q4/zKFUcO/NOU+jICuKfeaNo9D/zWtE6sROlpWtBh+NeRIdkf5+kazGXyHg2b3
b3Iw+3+Zvz0GwdumuyGaDZhgDOeHfGCHa7XUbzX1UH8WYbHtQzhOlmuclrfJjP0EmutNN8H4wgE9
1I/u6HTJAmgqiJJ8UsS9uKpVjr+eZLvgoHkB/JfscG4pCp3w67CjVC4DwldMbNsgmCjyexXP88O8
+OC+394efj+ygOU2t3yNql5tOp3CnkPQo+yQO2G7QZVuUqsXjrVXbrJ8RhZ//AJRnNE+NdEFdRbS
zQN68uC9PhabFkRLRBumvhzOho6jeQmiVOQ1ThschrWKZcX0xN+9c1E4NOjhNlfTlVO98XKkBFlv
Sqb1u/CFYBauwklQs+KE1AENyq/TRKX9YI99KLzwNImSKptoYCUIbBhhDljb6hiatyLG9QZ7ffMp
iFxZanmfOPSsRNagO/uJG6bgFng8pzjr25+LD47FyggocDsFb0h23ftlO1tMh6yoz6GIdKgy1vOr
es53nYNrGoiTy/OzcpsF0uiZmH6g6MGV+hFD4+XMMrxMvxflmVdadSPNXYlNYM7mbtso2dQsPC7w
riDXgOmewKNgC+/ZrlBp08BCKr15t4NRDCS4akrYVXELHBDxlx2CPDoZJFH3awseDgt3N/95/ll7
1R1Pyah97MABk1+r1B02/a+5+OjO+l5bZk+JhLyxcv24v5rayhmCYwX8Wm0c2utsHxxuDE0663ie
jWFMIHcYv1+fTQNwmTdi/igQS4tfLI2PMQ86mV8E5bw3aX+4KwUieYK4UPoBpv7qjSDlaJ4YdzfI
GKCRilE26tWljmIoqdDwD10TiXkqfOPrZy8e4lblAM9rqePLHWDlZpstIdfJYsgWBN9CMi7IBKrm
2LhU7cnAPtER9NRwtrjUPfPI/r2kTdbKlSvacjFBkBQqSiDNCT7+yY8t7Vnj0CDYUwbqZUuBpm13
P0HrQIOLvHfDSKv1CabAagTD+Z+AeSa6Dj9q+M2h7jRvOXCELFpd1XHviOp+/3HGNtZWIRJ+G9K5
FDdjibEXX9ojDmOK1VQQdoGYu9GfW2H3EOklXnFxqSOwnSZmtUFZqSHotj2HHmtaL2tTyZ+TQDzE
8W3qgdtsspYSwguH0k5JnR+JCyYa3m2fCDYRIuQWO2GUhgD1B/YZI2lNMYHGyGd5pkpkkOxkda2l
kxMMzS8nJ+4lIKa7J/zc8HpxkSBJb1W3x5Im/7+v3NIan0nNQL5TWfGYHUvE2nE8Cui/158vg/bw
JcODiJrGPgYwLfKRsOhsD4Bz4dTK5Rd1ShokUpPPM3mkLy2JrRS4fWg1PlOl3rFN79iLYrk4y4iA
H6x2FKJ3zlmYyc4oynQjY7WCMduDuNWAXMhpDLEYY4/gTgf0iQdygNFZF5GE1kjwh2Eb3Xem98jJ
sbzTBAinxGcjvP19P4XhinvtSkQt9BGmmAw1sNpmNaaO11KfsWBL4Rg75vxDUfwIlG2tNK96t9zb
Jk7zO3pIpeiPb/pLa/uU8SgCVQSngEcqb5lht7SKqyUT6RwLYWWbl0tqCn1HysFzFj5KYyrVyP72
m0fbFPs9gPX3B1uFuj2tLwnTK4dpBscgVBal1G3Spckjh2Ml/xJmezWc2VsDrT2Mr/HcY4UPPw6V
zRE0anLQ2K/oAozTzIERlWOeuTG2VtoZOT8m2zlqlrdZgs/e2bJkOfb1xPLXx39ygFbgy1bGFkPh
0bzCsWm9bytYmvuUy3ZVft4vcSWDAX+7WPO7ekwfrhBcu/qGrCt/2Q7AHr/CQVV1HOaBLYjl+S8E
xVNfECgB8NcDLpncZrNnK2RjR0+VxlVk5R5+8GUKI7Q1fx+REN/wxtfkPpmsqeB93NdpnOXOPwlm
saINCUnek2xVmkvVo+2D+p84F02v2tb0TLBbJyG+BT3Ehgc3UGcjQn3i9W1hTexpy/iUpDi5WPSs
PxAr7S9u/0iGv8mCDC46doL1Iv3pxkNAncTv546j640FWlNMLq6wQkfLw9Tpvqip4ovWVcoxkChD
YTSL8IMEIGG9wneCxtGgjSgDfcTor2j+QH3JZbbnVkONUfziOCOgR45Z9D6A1RNvkHLJJBfRhdoF
3shkZcJ4Ye1Wvy1stxKWwseNFjgMKayR2DzOl2BGykXuR742dadwaJAJPIKDCZFeruzRhENnzp89
6DH2sKNsA3du7RvkoqVfgfiJG4DseOM7gm6tjgdLiZP/o+QRMqHbWG4wQYfVXc6MHrByRboae0FK
7E7KbtpNPSZkqEyDcBmuwmuF2h3zq2a8n8wx6Kzt+tcw1txAQDewKNN+2ZTfv2pZpe59BVfSxjYi
bGfufAE3imuEFqM3i7wiFnKmcBm2TcD1rn3WLN4uM3rpVtXKKjOobb0HrmVNlGJEB59eQvTJEogr
h1esEPChvTs37Y9gohjI9gXnC5YePdQIr9SDLHxGHYOwlCz9n9ckB5N5aLBvO1WtBFOsHQqAlz/K
pWDLzV7h4pKvFLExtXOTLih7RZPfM4qWAXRAWEfgEpG57GlFU+mYP+Tb/0jNU7uok7TSi5Ufe8hO
cMqLAoCeKBpEjTnutaMdri5cpGPf2+KIzzFosrxf8xNHoEmgkfcODqKJMM9LC+gwtpOjKHB4sYK9
lINYtgNN3AjeTX/9k51rd+/2RnKqMnblsgCLuQkXH0tnJJ7KVt4f57XEYc2Jkr897atiwJqeAqR2
IgEshd9N5v/JqJmT/jU6YoycKjmdHpff8j3HTYFlFbuDrj7tJdxFOyv4YPFgh4a1Fh5OQhKyLtWz
71s7KEc68pYO7n+KA6DX1xDLnE9xOHaZDt9+evBfwhXRCFEvSazTjKO1uKBJuzEQFNlFiS9BbX0e
lS1n3r31AJtedAnKyQalEeT4SzBzGz2wwAudyQQ/vOlecXqRpriiharjbjIk5DMynRGpTz1UiOrO
RKnp5kc5OH8smjbHs0YHFBbruChYjE9uoZNYWGYQnAIy8JTu0PRY+Ot1B3ISCxPNkNMJCGWpy6z1
eqNq2eq9FV03sKT5MS5EoC3/mKl3YopXvgbv0MkQK0VIv5DqVnQDTvsdZftbbBDk0ff3cFmt46W3
g/CWZRFmDmQjxdD2mL4CDZL3g6WnfacjSBmhTRdeYlrvP0O5RSJuiw5Dh2MzVHGNBUaLBzr1FxYX
iEnsyd28fH+93ieaJl2+3ggJoBon0Q4WdXplLKbb+LSLfSNYgfnzwSHLLBb4HZTukeAA4Airb86F
oOIFvsluSbUTPciZ67ez6OLePFjxcirnmJGfmSA07dwXWyOR3yzFwTqq3P6FX6Swv/BY4q64jrEV
A4oMkIv9a+0JahVthQtcQgx+sD9M747w+/fAqDxlFnGMEZgdzNIE6CBiV6U5AMRHruLs7AhyCm2S
FjRYEOiGxPOSSV55cUkunaJIXrjouVl8SA2B6Sek6n4BMn1mLqdqe789bvPTunJl5mM5oVeSGbiz
cN+BzIYcY1PxAwwR38EHhqaRNE5wX5YAoacRlQOf3pBH5WMVBg69BqKJLwLOqYmHxi0Ha5jcRBTU
qriw+nl2KHXnvtCfoF5BZ6fsXYhllBhANcrfeS8FynXDyxZ4loHZtKsosjx3f8E9UoXkm9sa02xq
PHmAH/8+QY5egYrgs16OZARywmr6juKp4ppLtriNovFuO1OjoOfoSXFJppbb4IQFhSNSqoprdKLa
/re5Z0Z3BQHJwuxawL40QK8cbgIkX17XjpR0Y+h2pt9wOFYY51B3UqCVKiOJJihfUC9QcIQxGfqJ
fccIfVLIl5d+k+3fUBTAf5+y0RQI3T8r2fu6Je/5F/Ho/RkS4D1fudFQEzjJSJv0KM8alTX+g+AR
7W1xQ74jAKMf4cVUMTo0LxrekkRzLjq4arQiHZ2MEFdd1KQYAA15K+nitmmsdqwqQFD4/DojRo7g
myuH4gnSC5lNkp5/kXp6eKU8rWdtRqdMhIsMtX253L8vWFTWfnakTY7q9A+dv5mB5cljBy83q1Xm
cE++aybMW8pTzU1A4nNnHX3B4wylJ7trieYNcCP7QjuVfLi8ZByW8ozV33p53o0DQ4j99/QVkLLA
X980KAbNQO79wiBdlY4bcVEKc8d/h4MAsPXxuTUYWE7F/Uno/QZYHZpx2lu2sBZu0BIoNA5lifp6
q5GPJw/bzbpDXznXrIa41kdhrdpaDY3+2G6E+sM7m5MoVjJXO8j93oL+Y47eb2P7XlO0BY1hjZZi
gQQjlYCigFX+DUCAENLU4VpE3P28kAQzma9wD4GPlKuwpCBHVA+qeu2NNXOmXEQgfRfg1hyrSRXF
BEo9Sc29bUTARYa7pRGpKxDeyPNa/P47vHv6ElnTptqPMDkyNWLKN5UkjxbMrYL5+DVqooiI0vxS
JZlREAVckJQZMNERxCRPAyjst4AGZkIoX42CiCDSVTglU8XdJ3KrxI0rC8F8dTHsM75Th5TAVCf0
NpBalHn6PfC6DEbiY7FBqM6d89etK0+5kDX5J+H5zRJLXQsTZjOXe2X6qAuwQ7cAzSZjNCeH1kec
G0D2pdb03FwqyFlwjmV5+PzrhTxTBzdGF+QO7yA6Dez50IxDMFfSdWzor9j6I8nep920R8VQXpPF
YSa/cHQAjd134XgI5m2O1dEj99O6yq1OBX/bjs/YOwKW4F32WXxnhAEsYoNoE7SvuEoyCoE4NgSe
C5IyaYLNLwDCM5mpMaTFhRaM1X5Vz+XOV3wnTWCMxV28hHYInG36+JWJjKkdA7KXZnmBlR4FbxG3
cm8wLDAsogFUm3MSDLxGPVNo08WHQbbrnXmc+Sd/V/2MTxHmWL+3BVgZPMgwHExG7ETLMdQqXY44
voE6Mu1wV9EGuHOmr1K5Ps4tRLPuKaGwvqZMmSDWrH/2NxBurGj88gdpDBi+SJDQw/RpKjWkFkFi
QLqBf35et08lUfhTkMApBGMgs7UnlStV/RXW+jTm8ucvM/XBlrSm9kKTbz7UmJX8sLC87nfGYrEW
lxPSLiirkTPNeEut8sGPgCPTj0U7qnnJdt4OZchRRgW8DUxNfi2oKJ8jSfwm7rMimSy2XKLbAxzP
xf6x06/lT6KPfL7f9XX4n9wLpy/fKyNseGw+sr+2oQ3hSwcQzl+EWs/LnbcqkX6ZURcfUN6vCgLT
SeKVTCTnbQi/a+iU0ZEI+lEabvh+krJVD6n9lsOS5uCZrIK5gmtBiDl3J6DKl6cT68NEwTb6RLTX
FbpE9OmnWygHh9N8XiRuR+omrk2/ornjl4FLlA2AfWBstZPgUXXaQtKZkn+tPqpNltuxAmlt7xy3
R9nMoZ5KcCW7eJhii9iopSrYdalTq/nSBHy3XAhhKwjCcsnzfRcaA4Ii2uiuXncJ61Byr2NKQWjV
pmxF/RcNCPTuTcYTC0Xpl3rlr4Gt2ym2UXPhHGQRL8jjPToUy8HJbpt5CBYmQ8I6GSIEuyyDMzJH
b9E4sX/hXOqHV+TA89LDWQbJdT4VS+qbMEbVw8yGFGmkDxVrYA0Yp16CttoEA0z5EMBlwVCSIBMr
9Czf4nI/UG8mqE26znx6V/5h11nboFEjC5cNkBHfQ5cXXxT7fNKo0cIy5ydWi9NAf+z25H6xFwJ6
iAWlnK+9IRZN8CZxMFgrJY85PToQGk0yWKvkvLOBdvxi0bZGUHxWgWkVY940CtWzdU9PZaojbs/B
V2WwaKDT5JTuM/bAwzwkWRvf0hR7Ty2UWJ731CtPOicwG5/qh90+rxQTBi3Xvnfrb82MU3//WaFB
9WvxjFyzYx6E+wVqv+ZywH8LXmwP8SRz9vlrYUP56tXh750YsgHIM/UodMtogh0hdacZi3s3Xyao
ox/oL3+hkTTf6ypJc2SRfq8QwgQQHEMAVet4qdODba++SqOogpn808C4Riv6S7t7Ytte6hZxtuCC
ePqLw8ArvtVVNugejkoOvQHX3rAHkziUmhS8MFDwjHNrw3+chq9gSkZJhD1CYz6U/sYidpe9LZfL
aaD44zrtGbQlY8jXit3KLrIv/DYJFzy26dFhjyYG5N3OPP4c8fvCK7hkWcUaem0XGp77JqYjXgSn
X8gp/5WpVb4sdHOOrXmJS+zGGJ8oMCoMENRNMJJ0fojbcpgC0vsPk5gUy+/SvS+rvyBZI7xharMP
T20fVkwhp8Lcn9vT0fP2ZYS2twX4JTM+eqYtpfXO9f4i6nXcaULvsmAyWiE+/S7b/h3VXmJ41foI
kMTjojS92yX5nO+PDJFGHuYwrk9CR6W8w/Ts4xQATbIMA76w6urmOA5X3HWqNQxRdBOfjee6bZCW
1IaRFH/6p5LpjOQp8OfLBtodDuz1hwwY+RmBdghG4gX69yQPla/0bE20xpOQY0lab+/qxL8T9409
ATza6S4C4xhtFmLYM/51BpnFrwuODP1sFFT/M6gXWzjFo1cXFKXkYG+HF1SwciqaYeR8Rq6Vv8YU
hSdDV2yse7ccfMl39BLcGBzxGUER02hBooV5hXYW9D03zSgb6poirBZXoyXDhpg7bf+sYZAOBrbA
Fhq0PwLZ/oflTpwPZmUNlLYysF94l7MZvOrx2ciSvSzHMlah3IiwCxF6O1mx9MLkYJzHCtlx0vdZ
ESI/Gx0rpguIN1gDToQLMiisvM93y/VpM32hlgcMtghsoRoxLlNxdHPYgW/Sq5gDi2zkLetgTc12
aL1hGtEfsykKzVX9AwPo+kt0P6LYGoRLRl1+jACWe5OWEbMjtN6LgxkDHtbHZLxzEc9QiDyx2Vvz
uczoBUJLLJ15XYl/TWjzfMmyO7X9Pn43Lv/yghKOm41BRPhyXcMXkcKn4IctDTTtihob95A3dPXw
LMNzIYblcEdddqX8bN4gYaTEZjKwdpHugDeRGN7x0aQO7xPOr5s5+Ml2IprChGGkpYP7ei/NVvW5
BIFcYmlLmi/jLBpNgnFVL4AoD8U7/Sr/TUghGWz0New9Z6EJB8aFrhvXPAVZxSOYjrNbWepuj8ZQ
77puxUkzIJiW//8adZNeQge6fko4VXNdwfpNQxmpaLg3k9o1CPxiMAkzaTQCpAYEU6UpMnVAWhSA
3X1UUHzeZJxTBVcBUOHg9bP64kLD2tPPwe2ra+okTSuxn/1zHG6d07XysPHwyhZXVpOMsADVdDID
cBLcFv1vVisDC7bqjGCC3mCDsjI7UFfLTuKjrwodNT7n0PJ3cueq3I2sr64wC5t2mpdbjnNXsCjF
Vw+/DMy1x7RJL5JLH0htG7YpFwZ+AKq+4GjQruzuN1NB6EQhimayf8tpgQ0yU0EK9b01ndAuX7WY
jctqIR36rjf9iVF1ZVqt7kGrf7VBBqE8sZKuQkY8dkf0ZjRm7rngIYSqsIYhSt867GC7TJx7ZG51
O1fONlMNDRoNW8G5OvKIG+9rHcAqys2yNonaMDDpVlM+pvz6G4MjJgQkuZyRjOElZ9bMWpvaXmkl
2JRgF6YcNdM9HE1fGBedN/NvjwVXPTaOWuCzQa6EFXegY8OSPgiD0xoJ5lg0b578r6giDsZYoFOu
lRCFBYeY7UVAz6FPfd78nqsWp8CCaz20gaFKMIHTQP6LlEMZ/qZsqNbZgSUe9dAbRkBK15iBakkF
apj86jBGLo9n6u0DrEJ09JfTwAqPIIVEfuAEMIdmDYxwhcp/BPjeGS+xuDTxV/wV6t03WOjENT/w
tK96SqRkm8GR4HlrW4VflMieAgiI18vq2Kg2f7GelQ9v2gbRUyJE1Hm8dc33fHccskAKRdFPLabG
V/G6fbyHjGul6WJo4xMHrBSKco6U4SXgDXfiECCcc/SpYMUWDOjMvoN8BSa1PFzgqDrPdiPgmgB+
Fyt61zxElqQw/tSXqrfCFraV8VMHJFJ6mLBl9PAgJu3kvmfujGXmVCl1EHV2R+MixjbjnE1AS2i0
T79qFOBIcTqxCtUgE1QuepZta34woeDa2I+FVUXES+OMl4LkVyl/NIzHZp1FyGA+dlJ8gfqkjlg3
By5Ka3YrHAjFomxuSFwMJbvBkxjCATl271WLIWXrE49oT6qWkri4zsqzN2OjbEbHvdkyH8KH9Xb4
I7XVU07Wl7p2LTVtEQQ4qGET46fVGerSgPYT71ay9Yf7ggB2Qm0bO6dYA4shocmOBbSPpNbb5nDW
uaSQ6oOyC3znTaO5jmt6J9WRDx4JW7Fp3J1pPG7eF371j7F8htd8YD/FIxj27cKT93C8+Rbxcdgq
wFHfsy1QApLe0rEZfULDDLMUUAYyhP38cRiNSJB58DexhyrI3pxfcJzWRn5rKMtlSFLpkj9dz4VS
JHFH+HvysgHke+1qU6xxyeC9QBm7opX71nisfX0ft3/d5CbGSHGn7RzZ2LtHzLXnddCCeAkiEdvD
tmwOgb8BdSH0SgpLlKRQp11occMjYVEU/Hzm6SPDPh++8P1VbAoZPvDDjdgcG7S3CkoO/HKk5CIh
gwZR+adG2k3xHw04LNzzSwbvN+L2u3gMrwR1zYzQWsMjIz0BW8g96y+B/SyxgxsNwwTQpVaIQvSs
Gz3qbg9sSwwzheYl9hGGciz5a/BgWzniGHrcbDR8lxUVkI3wTs8hW0/yRMSkGV+cFyyG/HXawdLy
RNRh3pMyG2geDmHhV3N+2MCOZ3iEniKfWGZ2HvDmprFT8Y6M++kVSqRX3EN+shW5TqleLwnHLTey
t12VGebKt5lAXBwk1LTu9fkUwh7VsYu/J3vnt1Dhn2LL3gWM3M25Ftoa+QxmHcwj5IuDr4alafQC
ZS3qYPsBTE3FLPX3bSO4CA8hGpLcYFYfD7mvjEoo+Ek95pGt8xfRG+JCKxOOiul84IAKQ8Frnuhb
RESUXSRXLXb3IQumPs/j/yujAX7qTOZkMBdWDxMjPbmoHvEIzipNsCBEWMluOteHMRLWilkXTW5s
C6QtFdhHYSGl53PFD5nCbToeL3IFUgYLV9RruQ5UWL3oxotX2sHzVh4gZRLWSRNks9f6dcn4QBTd
g3eppYsqxmv3ZbM2V3Tyv/NmmJiMrHhFBzcQYkj3nda/Y7jivM/pucEdGimQbEiAx0F4hFrO+OrY
UDr7Msx2YtkwODITQte6WMm6T7lPYRBejI7ykfeXdmfex7rWMSzcNsIf9PPNiNE1T4xS5iSp+Hea
0+qex8ijrGwJUIsg07kceT9IdKT3jFSisCf984Td2GDXRLsH1oaoKkuHTMEteSGX1yU7BAzdr5dh
ETjy50hyZtZxC1e0gQhy8J+T3GjOQZgfS+5mBlyDv4Xntk94n89lvGMQybc1xCgTWQ4MMtgUvV0f
zW1Gi0o1y0mmISXEEo6wJSOU2NTpDAmLaHADOgHj9v98VTyEC1BfW56/HhAZ6lwbNcMpGtgFG5Ts
cMKk2GTpw8cXioFOFbGVyx+MpbiVhLs/Yg1W94XUuKLyAXBPgamnM76t2f+G30VIghNlPBvqq5Ke
5tI+Cq9ZPt7tuo62e+uKj5uEawsxbc+2YlzoJU8fiQ/bPj6yXfP5y9lqKZaFHyqFIBFPK0PmahnA
LjtEQ3M69Dz4AUB8mZ4Bk/HrN9RkcpEwKLaaEnYWJFJ/NyJuNCDJxPc9lK5p9+QEKPBWIUmR1gP+
s1R/BaRRCZ3CGuXZ8/gB9/OJVijxBZ4DbKiAu3cMK//bPRKwqyJmWAEMSaTNFnowLAFolPKlunSK
m2ezMQkS/vFC9ik+e/Ci2/twWXGncomJAboStCYaYxTpRyV9rlkJdW0AbsuAOxllrev4PzP3GLEO
QDmQPMvtj0uii3FiY2tW4ye0EgL/nbqjaIjB5HuHT60BCDVZq1pbngwO6INJwAgZYcpLw0McxkRQ
n0xTI17GzG5LCEjoDIIU0UUl8vsPgpAKk7Ns8pHLht0DwC5dYaI+TZI8Xh1uMvZ+fOvto58TRKb+
rQoH59bbVYpovvihYYkDy44MJ0Yafur2Qwx2ow3aJ3rxA6vpGuDAaqln+SvcSjWJ6P1bch/d/DTe
0v6q0SrU2KnxRtFsOIH1MXr/XfeYWOoxZskLT9XPrzcgoQADUd5fE2wAt7KPnYWmmL0G/CnvmNs3
kbqEs/AqkQX2uqtfsJK4SMpr9oF19q3siA3R4GNRUEN7ngQTZ274tJMR/OY0eqdWxrs3mNaSEEm1
6M8lT+pO+SzuQj/IXPnV4xrhU5UqneAXqBQCWKX5y5ELdoViAvH9MhskNsVWisf+fwkVSiiX2QUw
JwCikEwvljc6gRijNKywkN28XZyzLYJFjDC75eGkFbx2a8LZ9y+airLHl/mZnw4erDTPcX9frOXM
bcOgaxQwBGnhmbRuxlomDPez/mMv8M/908ZT1RSG8VjxXz20p4l7RsQ5cW3/w7kNtNxd0iclnzCp
uDfYj+IlOc/lsi3/PIO6xxjPoiH1GzvLxBcJBBNaInXO/Vd4TBT8Tn82RrnIyr/GdinmCQ4OIuXJ
fr5bI5jifytNwqSqCthuGyHppYVNp8eP4zOO4yDRa4Lm50vxdEniIpzqsUxem8IvZ1KHoFio+cyv
jvR3b04F6ObEu+0A21JcriWE0/3rz7UJVt00uGC/hfrYFE7vcnaNr6uDHv+SUr21VVKqJesFSI5T
ZofaiYpcojOxprMMEuvmvFVjcj/g7BAwrMV+TOg9hJ9c3BR3hfi/cGjt5Uq2BUr6r9nQbGnVJ1lK
VdEsPqtt+vYw47NQuGB4i7AxEtAnPCnZPe8nak8SKflLNy1jHwbZc6VFHa2dZCUW2PKneZzVZdAk
Gru94/J6hU/XPU/06NcL76JpHM0/3FQVjG+I19GI+/1nf5b1jNgBH0/U5rAgocnmD0/Pw9eTX9nI
Sivr2uWbnVZ7B7m70Z0qUpxKCphMZAJsUeNXS6Jy9kJAhsLGuNRAzHQveFoQi3m0NAaoo9Cjt5S+
SumbWDiS3UFDXNJC4FkQdD5NXU5KPdftpYH4HXIKjAw6SVHT1AD/md1fZf/t/mVxEpJruzSMDcG+
Lu84uVqG+oyF8Eqb965/kOjoZQpBLpjUXArLdKxDyxHMky7jqk4eRfxEwBPq5IwFL9LgrtuE9Yi4
WkYgHUKIuadp8Bepf0JteBg7v9qcA1CTY7kmQkAloHp37ft35j9RSJHobDXkgxxMBNp+cDblk8m1
GrBYY2a2xLT1UrYbW9kppm4tq0ifufEmuKWAmc7mOE0tsbBB5Pw9uR1hpHp3RQMovDsdPxd2SZDy
05rhGYitrNHespFUzrpZ5pu211/GBAWEI5+mRQZREtU/SvesTb32a849zNdDHU4q8UA7qCIUu8QO
tzpfuBC5kbk7kZEuhD17kNmILipvj/qG+4+5amuQP3QEUlHEkH5j9QGK5OXBZ2F2GMj8Y6YffsfR
afSjtg2YSsGfWWjgsSd6NCRGexIpd2jt5eOlkKqjCyo3YWip8JL9Uk3CTiq8tgDopmvBdbKZE74e
q0vMXviaqdx6rU2/ElTcrm7Jzf07AGMBr4GhgyuDk6nisOkpWVUQiIx7ai21E0suLjqg6EHptCQJ
mMB9cRk+cqa9pNWAjtgDl8HAgeQKiIFpLLfTvUKO8w1as0aBIYmGwrnPjYTdc5JYrWiEv7GY6zxv
k3BOBvZnKr3QsVkYj4quY5YpIvIEDm6iLeiH93PY8kieMuO2yj04AB4iImuLF9dltXEcjL2dTkgY
aT5A2ArhXOHCUR/zKKwpnDOqMursWeIfvfUQ7mfm7tk4TuLZ5PVEZgT5MIJpEKh+PGKaoIy95qMU
iaJm6g4MXsq0WmlfiM6TBQa52RfQbQy+K0X+KBPkRU988UmH3mh+1cFzoE0eYwOpHL3FjLc/BSwD
quskN0nXA7S+VRyfbWSgqtcIQi3GBphR/8QwAyuZujTr2sNtaNi3uFx69n93jANcLteCuc+WTjqg
GBYngFXX7ne8TKs01G2JeQBBhwhxvXYkrlXuSFlSlXDno26wOhGx29ZOLv3XVkgFtUX1GxxJzD7l
2F8815Qub2dCaFBh64wQKK/ZABlpU5F0StJWtCm0jrzoAn/Fbxxii5hY9YZ42pf70FNwhpU8XHHQ
7VLpXpmhEJXE813LeCEKwvT7Q8172QLspQwFu/VveF0Tz1SMmn57CGyEJeSsC1xCJlECV9iuIQWb
pafrNZfFci+0+fC+/9/gEx9ONtgB9r5ccIbg4rGngm1XBaza/sTCEpww+++skTkpITtP/v1hxict
++olKh/w0A1D5/rnQpSPJbzoVsov9pfkoD9LOkQn1nSYkrUcIMvF0oYb8xtHZaAOGMjR7ajJM0//
433iPB4IeUQKEZiYljdrcc0DX7bMAARJRayGQZXmIzMGetJ3TOm4kgvMyAYd9iVBCGZSaMrPd87Y
CLfSNWHZWTsyLJnNvze4lSJ4OjNwRIKWomlMGrYNYp0SL0Wcu3uND0qg8J4MqWWQMvkBAjsYf/B4
0k9kpsf+QXBI4EgmM5iD9XZUCG1m+nrSdBrAhZ9elsMY0LE3YCTidWG9vdas3xf0AOgYmSVmiWDe
6nyMfSASUO7nJRKyt/Kx3dDAReHs3DjqOIeUCbEUR+jY3O/SDyC4oKGylQEV7ZNUJXmJVSvd+T/N
zvoKBmrAxfKrccy5VrOyA4QWiWz72BlZ4b1N3d3QZ9/bBy82y5jcZDFHpcPUa/xL2fa2U/1cCwhZ
agMtsGBGIQtmoFcR+2IE/MswskmQK61Ru4IF2JIvHRIgrE+wQrKG+k0BkY2hyxgBvhYiyUncSPfg
xL8hgAdJ+jNa2TXwz9kPuZF6vJknS6NSBgO2t2zI0dsajA3E4keqgA70kOYn6ByEhNr/T4VthmTg
2mvjU933gG7cShV8NZIL7W2EccGfnYueE/OP3xQ81YDVSNg76YpXP8XSpYjHG0RDrx3/LqCe9+fq
LbBDt12yNLmobflE5J3sQnzCV/NZ80+5Mh47aFwmUYVcF1QLEyQiBIkSMoYm0IK5p/RNdI+K5526
XJocDuLoRBLfyb7vWvD1PEdfRfgU86VTi1kxK5R5LVNEBBQxTT9OEaJlSq0o0ghaise88XMmc3Ye
/bXFvYSGEs9JYnA2tpB0gqCnjkOAKZRjB07BHYFG8A7JgJz7v85IrpBfDqfMNdkcD3ZvDsJt8iNE
QTjuws0qT4evY2MtNpNm1XycLiRNcli3lk4BYNo62wSh8PU44yy2cjdUmdNCHk0PYTbqEszwtKBM
yCbPDFwdgNnTyk/eKnrOE8g2YMoTPxVQtO4v0PvnV4nt5bSXoY6o1dLj2GDXai71d/W5VKhvg0MA
cxaZGqsULo18T9kJhQBwv5J1NwIls1uqH9AxrRYX/vdUDF9UEGBPbeTP0PekcERtU4Vb9ixvqLeo
sdk8SuxSkwcLTi1sSJSjDfC8OHskrcLDw/R+Bx4QmIPUa0077URSajZG3YjqJjckkF7Sb2IKF3QJ
1+SlG920eiVib5MbOQUDlUnIQQLPiSK3Dh4ECh9YSK5vpe7FJl56bqFmWuGOvZbApydp+Nz8cq/O
xzd5Ev8FVKRCChQypnopGEiZs/1+QAOIt+7P0CCTKvZC0+oG3tJnxjRZtEgJmkUf6Poijo8n9fBv
gvgBDP9/WDtWa6ZeoFKFBtHeFQa6IHGlUq4FciLrrkMKs+B+wU+d07x+2ZeBbAyUzJcKN1aojurf
WoFSgseJoHA8HcAClbJzQzZAIEPFSMZOQosAJ/C5l4bTO7dHfYgFHF/OVi07UADfz6soPGa8lz1p
v0jAmxO+rObwT/XSAbRtNrzpyIzvD6/vuVtfLhV18zM/reolbNzwRX8EguDvyrmeGtcnNOSXJvej
pFpd5JXHn+j2O4ksAmVYaEqUwhB/tw5/iwW8QexCr8rezglEpQH9Vaa7Lxl0dShpRYsmP/KArrdW
aOpHKn6ZG5to02/v4yQCaUJCIuupeOt70roSbi1VCJ5xWmCSr5uTldPY4EQ24SN3heIGoBXgZnCZ
DReRmLPR0t9ipDV3Mu+/aDSHCW87azYbBMlibFVFaLs7FZ81el2EpAtUgWlJAR3ZYIGmxWcqwosH
rAN7ypclM4YUgzs2Hcuyx/1/S/ZhZAUzbhxrMh+ndzBG6fn9ZyWYs3Lu7QRIGMbK61syoKxTm2jS
oje39gmAbGin9KM5JoIpzjV5jCz+229tRmqM4En9a94YMmRxeiw/FRxxoypx1HhL8qlu5UI40VXC
CMHy+7ekK+kpgWISIqXUCP/GbRRd63RZYG3XdVubqAoCR0XbNpoUHOlvrxMqxloCer4HaFX6QH+m
PsnhxRND/yLa5S3hEXRc9lkcrsdDuKzSq4+GJEGlN/XfpW9xlt4sPk+gQyKC4ooWyvZwKJ8gqFS1
wGRrJBVXXLoEtfCmFV1QcuNzeGIRxFnF/XQmYP/XTbBhrQLzWnDY3zyEzHsjDspIENeaQ9BBEfVo
1QU6iVpJxGauAQCc9Pg3ZX7+XV8C2k8RK2Lgvm9OFojmauKpOVQ95CFqlsubQh03w8hdy3xh1DSY
yO1EQn3YZdsIdxoRZ67gOOflZ+GEPNYmFytO9XwRUgblYMoDXC6rJiOQdXRwyfTITaP32OjLKY6h
5RuAl/Mb4kqxuVSwQx7pkLQqrIYAjkz2cJWU6IhNnEUji87+wpR++5KZMQbkCFxZK3bzOHzJ7/KM
SMhHNnNtvPF6MCBYfHljVc4U63SkLcAZcIFNm8TSJjOdYQrTI/z4erz+uKQgIXRdtO66EZxjNUt9
8hpCHvIYlJ4OQ9QjdMqli0XXygPIBec4uhOAqZj67E/MZ3Z763yEpnQ23JCyEEzZxHQ4voXYs88d
H7J/PAsJQRVSclffsfBXeFSCecuXFdIpr5fP+CO7jihSPZ7ecvXSQmuFFO3BIfrhm+gekZnSvqKQ
5FUkfkdZM086d+VSKhfxjahm+0UXFXJD5TVEgzzMoYRmO9rDWaUHTrv3AcqKHrOGdhuh1fuNndvK
/aTc13WhAvC2ZPy7tJ137fH0vVFcduWKZFwYMIJ0y/29qfM8CxxqM9m/bc13i8PfHkJmGNRKm9E5
1JNe2yYNf4IDn1ciYiCkEPYlgYewDv4LDzNoJLvzCK1y3UN3+oyQkxqwJv9b5+DVdnFQ3qhPrXz7
ETwZw+hr5EDiRBRrJe2iBKYLSrzYEW1JLV5iRXVQS1aXuANQiP+0sa8v5xna3DYiGPdIdqqcHZu2
qb2OgN13Ffqb1DbdshvxnWA9lzfuEaYGbxIUQZVb08FRqTKZQazqaVBiGBoyN50ftFMAm0yD7NsY
5jXApoAidMB29YUsukrmFI80PlzDVBR+Xi/wRSacSzA6XPTfWePXYpdgF/3k+vWtyBJnLwDuknaw
cCmTSjWtqZWNtuarQedOQU6zaGMhawWAv7QLnI94zNbwQLZsqfI9mf46lCkPRtTk1mXnFXhpBdZd
FOOgY66gtstqN5nkskza24PIpC0yD17zjVxOcFUgrIKRZ8EhXSPnEhvE4Kt+3y+iMAKw2Vrk1wGl
R/LsD76v7M3Kqe88v96PY04c7F6lFcHvkRpHvxYj4A3ZfCuYawTpSWlvLizNm0ovu/s9DU468UEI
Q7j0dojyL3wa95SKHEtj6VZ2IOTvokiXxsfNqK4wwDT+jRVg5nrAMejVqSYxGT6sax2+ZduhDbBQ
7ZOcgDC9l2zFrxvcrcdpZZZmUtxsD+TmWEm73sdxo/UW13UseSNk8UL8j/vsqkI5pMRiKU5erDlP
fimNeC+3Zwmce/0FCoUFJPKk+WSDbWeaSyv9cczefP5qVY+pZjbym2wY7JQUPBjtRs9rtpAE798Q
+aFRzv9LM/UNc1DkjejurYoNAOnBd0mKP3fdvd+6MHY4Nebv0XUKOdDoqkjyiF61WVFgTj0DJx9V
FFx8F1fgvBaJpaO7urrHb8PPUI+wP1EGoCF8d6+g8R+i+C0w9Z+mhgv4WaPhMuJcN7emwuR08BbI
zuV8ShRHy+6nIivJ654krBjTQ1dXBpHwxKfkaPWgN110x+jH/lHwR0pE1BaCBIIy0u/MkUz5GusA
R6lz/oOjjuyiu6/cT3bK4HQMJJF8SeTJjgiKLn/XYs5FFJHIrEtXT89Ws5l9UVZ0tg3Ccy37gNAZ
CXIWQzoA+lKfDw9A23qQWgpaU2GF21qLtwQkWsb08hPbUi3sRRUq5B18qLv+yH/SPvbKk/nR+NqN
mNaxUBVZDje/jgXiPXTnWQEiv8kUKDO8sz9mutakJm8EV/tVJ2sqxiV+YXIjKrq+YUXpUz98bREF
ZjnO+J8oh28rSsIi+ElhX5Sr5zs2DqPUkcrLh6u81SUyYjrlTkPWY6f2hR1nuTWVyGdXvc1ilUkH
r8VRCz4rkj3NZwLcCfp7qdKyKkgZjtbyZ75BCGnorbqhPpkoB/FO9Z8CsaXjL4wRloiLfDrCiyiZ
n7nek/1koGk4vNOXu3xM4UuyWJaLm4G5nSeIuOysJk8E6Mw+EjyCGruC+eJnSOh0L66pfjAmUisC
+sgt3hjCQZh7o2+wzZTN86E1FeU+kH767YwS6Vv8juzLAD6guUsJLu+4ucFTW8zJ2RRsaWHAcBlv
XZnI+URCdLf2SBnfSSQ+GCXDSrVVO5jQXC4LTezijfYIETot+tLkTUXc0dvCi9j4w4HdaPCSCqwa
1AEtTQTfcIfuGnkefZPX5OMfI+12mpr4QL93qim225RrYa1TfPSTJxL0kFWRhOwqW8veDYULFUKj
25E27n83xFs3IFEFq1LB4nKJ13Romke80EyV1w1AwS7CxIdFTjSVsTxLT/IcXypDgcOFrGNmQM/4
w7VCHyiZNcwuynJ3tgFFlv5iQ1Z+Wox2qwSlX1bE/bnXk426wXE7qfysZ3OFGcvdF/LQZ/FaBL3x
KSDvc/ZVg9bd3xaPREo6B6UXxBrnpG00tlgI9kwpcvnUter3lKEev3KBmuEQNMJzypQ/u4ypOzER
EjMFbFhL1b/TV9JU0W6rGbv/mBANPGKFVetrz96AjaQQP8sBR1jGH35CSXsjpfggNX+M0B/AnlNF
6UoXFFgLRwd/v5ZSVgbHM7/w7V04SF0V2PjAnVQz3QmsDDtPe7zNP68eGQRzZuNWAofaQdbCbPBk
OAmxsJ1qGa1r9LjJ/sguEEuxqE23odw7dkn2rAZPhqa/2v6hQTcLIvjyzNzsptlfDoxpmvqtz96k
dslMM+YOLTnuk9OK23ckxPdjlYx6mbem8u8/0eB0wrpuHFZZqaFVc48/uRtu/64fw+fwui9XpqOV
Oh9XL+iNZhNio7vgaIJIByXpaELi5nSBiS/GpARNjo2COS2h1uQgrm5UMAOqRZRAnUoSJiDXnZyq
N/ahhOoFc9OjZnNz9805gcP341p93YL+LbBJRrtkPJK2UUy5QhvFE6rTM+1NPfVrL3JAJFIvDybq
8km8cRJ1qAP0P/oKrtyopjWyehmq1WWX88Uy+uq2wXhOu5Ru7k9HkpLV2elSepzGvnF1pPWVfyp9
0G/T+4v/aIRkfu0wwS6rYQbJ7at5FS7jVBnPA9OCcr9xLCX5v8Bh1+R1QhZdJDrKAIK9EM1KgP5o
VwHlSzMDUH9uJrPZ+vHcE+jE2NqcqGQb3/ywKagMvc0PqkJOiwndAyu6zjNzYUW2KfRSkT8WwqZb
hFRswB+uRsC5fXCa/qdtP+rpb/Jx5sV62VEcO8aC1BJ8KvT8adO0ZGSts7lb/wobZ0peB/F9UlMg
g5VVAKhgoZZxZIq5K+44J4F4l0yy0tIT1z0ZSYPU/vYy0hWX3uQUCMTawZKH3R37VqYPn5yCuRsN
BTcvaTOjmXEnKbjbwlQPncFZU6iNLGBsHJDO6QGVWIWz2mKkg+BmT88SxcNrdB1e8Z6sJHUqjJnD
xRsLVIIWaq0udU/fcR+d9wA2XO+vLfXl1Zzdmdi6a4Lqydmq54nozFjCjGFcxBH19Ed54+orXIqu
hwMZ8hvPY/pEk+y3w/igheC5My4eYc5Zvmk0TAWe0P4UVVfv0Ol6QLyOuVp7ZDfz+Nc3hFG4cgCN
r+qXq7JJYO78Deq9UJ9xjM5pqWsSwzoCAJddo772tpHUPHihuPlji8/hRZ4jS7d+3rl4MD8Ess4d
TwC0eAjgEODkldubFEEcaievRjCCkhNIndQeoKBs55uYc6niej4zW6wkMj/RyejYL0qa91MPGow7
1+PKbbm7zmZgVVItTrVU6YUOUWJhXbeHPjuKcc4JimoUyna0/xny/B5ADdpSrm6YiTUqU0c01vlF
fwwYkVX5yppkAOmgkGk0HhFB+u1WWElqdXexciQLOwlUIDvA4tOeNwv9WFKMUZUwjyjoxyHSOoYV
matPh4m7kHK/7rcAxR982Iqz232EuAqjU+OqARtS4tHwnI3ZGDp4Rf6k0sQ7SKsBx9FAJjqu4JIA
R8/7Guy3SUMYKfyx/hFcBZvYMZfAI38atwNfhxcEf2DtoS6m4Ijd9tW1Fb5F9lIrhAmV2CXHtp1P
TwQQAylvrywqXeEBy7Nr4colPNHNGy3dcusBokIQYpb9tuHEnEatLLNAlO7nhsj8yL6d7q/gmhZI
L5ZHHxk9EQZDpW2dFvYMFVRqnQ+uf3mdAmOLP9zxKzeW9jy/dJDQxYUxH3CPVgxlTpwDdTU5t53L
I8Otmo/fOXOVWgux5HsxVjQrtqsLAuYnDoY1STYvGdGflhUEetr9Lp5gsx5lwhArNXNJ6ofU0Dkt
ZvLvaCm/AIan5CzF4Oualy3TxT9n/slQk12i6yXDSKuEw+cqrmAUG1IuxklxmovRNkBf2IijpXv9
SYFLgdTsK7hVH9ZR0SW393Lq6JG7nAGdFRLBJp3JmaxwOAt1cGPSt/fXy2HfaWujHyIG5PjHCkza
UE9UqHCziMeWT2yoOpWo2iRpUKTbvhwcgmqZkoZy8i2ucJ8TowXxboV+YBPff2e6FzuZCXVnJvGh
K0YGVWhvXrOSh/+lywLFAas0egpfDz1zkk503XWOz9dkdxJsMOCUwU2gsU4xzMm6EdRv1mDd421k
PNe8PQcHRf7T19AQJGYo411a2frV6XV4Le+a71ESdt9GhOCQDV4xgnS32Vdbq0RIBLL5Ka/I6Wz9
8UqAWHUGCs1ceTMp530IIjF5Q8PHmCFaTILOnhlgYsZ9h3Ax1WGt2RBqxqeZoqahhigJiswKd2Ch
fhGWztAtwT4AWYN20BVSXF9TPoaDwV/iEQwbyu+qm2EK6bsqTdV4fQCfADWGg9O99J37F607CTGJ
+ylpLhscxtnbLtC55QrDZMXdce3WbYXfvEfp4maFdlVu6LsD6MBKWVvgAz7Rxvg/A2NnZa7oH2+Q
E5FjVL0jYMMES0EDPRjqpt7nXySnmUDXVnKlxDftwduL6QgjRbu7ZreirTQxY2ZuN+6KSx6xSc8c
KfyRyXvQkGMSL2bqxegT9TtdaGcAeXSpYtyBcb72wZbmUzf5G5WnvI0/6Sjvbs4oykVvDt4k5X97
UbJmMUmoiCjmpWwpXHfU+6wtApZ9XUc89cg+YrpzGjkhljyuKl/oYSz4tkPBn/RkpKWYffj16Oxe
W7BChoCS8CFygP/afgMk0QQjLIO0CQxI15k4XSMaRnQJuwT5/O9eBrF3A1KCe1JaCoyNhxL/kZkW
7pgUtgdJJxQiuPXLRNoNYj2Q5IHyXBCvJJ4I4ZEN6cT+tBuRHSGnOPeL1jba1JY4mjy4/gDqKw/P
WXsmenF4zSDDuOVfx3xLlpfcrLs1AORdlRNWxe4jL0wQZpuX0e218balBwwlza9YZw75lesQ+Oaa
EjWK4pBwo1VBgQC93Pyi+se1J2nPUdgh9zd6n8IPjMpzZipFPW4kc5gnREolDFD4dUCCIBRR3F3L
T5acdlDWQstFf1cD1Q9cQ/9H9GaZBheI73Bk7hTUgbi2XHMeipA06p52PRtUHC052YbcmgUBBJxX
AAWohpUSr5zvfJlEgbF0QX2VQGHYLWhyNoA6zAQO87hokCZ7jRNf5lxmP0Z+eNMNSULsvsSYAclh
OhrLs4XoAABDjC5D+rxhFY8Ec+iFoj2z1FBIPYjDYKbo1Bu9mxeBS1uJi9qyCbHUDTyzLzHROA/H
GsDIg/4aQg4GzdOHzEpSqB2Ty035ZZ7fHcVphdl8AOqtOo0DLqpjqN5Bs8fzLUnQ0IpMk9XnFakn
bgRaF+XnB+t9Z+OF/FV1WcZnlDrlt/b/FrLRzeHovmwwmdOd7CktvlgZAuU4QTh1ugYGS4KT3C/y
y3CLlSEJJa7x6HwZhUAWBNsKQoXNNOzzFX2yacgSNYYNuJ3fWtKybc6rRvGeFsxQJ3npR7PRywOI
jUzSz5yNeZDZzqtfG1LlmLKXjGJF3mmooy0qiGJZe+GD4Lm/Y7uazEQ9DdKbU/AEESrZf5eVvW/e
kOH/z1a43uz5mQoFjwQfSnOEu6HBt5xVEy1M0SpkUNAQEgaal6rdOdOS0nIxcHtfCBCR8vObvgko
+MrabmQ6IvNX3PLj75z7ikumyba1Gv1KXl492Td7Xa2NpVHsQoW1wNcfXNz8qjaby5QHMgMi3HOh
ql3eKflEC2YVyB0UilB9xlCSABcCCMbf7ZYDEkh1by3fhv5pyWFcgkdHSWdrk9X9sU0ye+g0ytTE
y1gAa32nNAf/aKWj7JM89fQL8OmTdEeP5vjCpvASt9ySuynb2SpLgt/Y/iFvkcQKNBhjuM8ag4qv
1HhXPDNgTRkZhbwS4YEQS937gCIQC80p46j7H/mBOm3ONorVvpupQ/kiBI+N/0TNIkQdQbi2xkkn
quJhCtZ+USnCH6zjtW4wy/WKwF6Udpp3xubfiRNgp+QbDAhMQt+nEsbYeO/HwjargkOcg6zLMZWq
EkJSJbUIw0dhFKEEKfh3cqb/dIePuTIqXTRoi/3vFvJuwtZtEV1m+BvA353eE5QsO4NyoYreZQvz
On/P3FFKiKl0JyQdShlJFi9uxQE+9FlEuDr6LABgsX28mQDJCe2S6WOQw70AgX6jlX2YGmwjLuCy
xQgqdvw0jy4mgXTayPmcK0lGRpAX9/ws9ap1xk/lftVo+Wj1FhErOqygAcisrPSl7nbS8MKEssfR
bC6mrPXqn9PizFG0Oz3KDSCDWqdkLZVT2PVQKTPryE1lTrb4MryQiwnGnMKbLIrI6+QRjg1FlcUd
m++9HS5sc4+O1aEL6otVO5WkvNuzYQBBtWX1xvoCeZxYB5BOzeCfj/hvhSnJzOALA4lu9HNKfn2P
zF8xZaUTuKGiKVi9V2WT5MxdC42cbHzysAnT7yN/VHp+KZvN+wjR0ScRSxKn2h7TMpwfVg56S5N2
vmql9S+CxA1TLJiC2VWgjPIb4LqLBvEJE19NWjQ1P8AWwDR7UtwsYVR4TJ1WcLCAu+1CGIxMzivh
FjYmOR4hu74DLRWdjz5+xOSPH1Md8TgNhejMJ2r4FuzTi2uw51qaY5WLX1cDNTNaRH1Nh4Pm5CKI
qjz7Syn+MsZgyadsRvTM9YEzezM/q2tR7BTvjyFTTNRtNmObYo1A8JtrV4MVoK3Nto2KhuyuCaqr
YYy6o14iDS25Q3F4q2Zj6TViGiUK6WRg3N9+QQDaCZ/cDjGP9D4IgS01DrD3SJkfBk58MO/Qa7u+
RdekmLzvBccl6Mz5+yfTkc7jPwJTrXi40UZiO/ZG/yhkw+RKBezWw3m3x8PuYzYv6/HK0cIKLP/x
lppXmKapRHioczM3vsw/gnmX/fh9Ky0bGKMdNKXgaHGJX4oOqcj/+48UR/dNp4AVAsHMENYkF0/9
kXVRUgm6Fk3upIbS32Pci5Yq/RNiyl2+Lr+Fa4eIwgHfg8RTEoa2xuoax/L+h2aESISJ+3jSEaqr
TnAOPycqLer2TdIoxMWte2HHIaqA9qBhr4qJOvWEatadPeNYlwk3AfQkLpR0g1aNLFyxNltxlwmw
Yf8CXAymKRWAPtYyXHx/aIuWVB47nFZZMEkbAVeZRW1Qo06v3JXlhdMmqKkIuwzlcVn2Ryo8S9nc
PqCAztIx7Lrm8dGAFEXNtc9PWGCIKAedWV3rhx51aY955YJlkg9Nc5Cw3YyJfEVyyGKJ+TOb6yhe
CTgX1A4u33S/hzCtfhj7JFm6rc2KSrImSntDqimGGxibdo4rFTQa6kAo82wffs9oMBOwVhz0eRjG
Qxghygymp+n8fWUNLSQBrBvVJ8V8Drx6128/ZaAmx2PenZdBxUy517IYXK/hjnMafaX8RtIx1SjX
NDK3ew1og/oi9xY85uHiN2co/K961/0wTvoqUNmDAM04wJPT/6SOAknW/+wJYvJgbt9ms8znuLpZ
j8WdrFc9WhpV0kh32/mp51+ipVWo1hRd1TAYZ+StGMaS753DgL0Vn157oAyYnFAvOg29e4RLiEv+
GJFTFekZW+jNAmMNq6tcVhvbG94+qBL+PpH+qBzkrrGzYfnMMSNU83b702V5MSmEJzVE8Sv0zAwK
upT2ZrL0NsBDeFGFAVgwvWIYLQV5YIfIpsauzaiZgJJR/z1ngknIjvfZk4Oh3ynh11FcwZSeOICz
NOps8/197jtn8cobYJ5Um2/HHsaetbZnFmFIvxPI9O58ami6LJGrWHJwoCv+Se1vMBbIa6PROTqV
bhsQb7x2f6EoeCa6p8ROm3Qp89o+9xUm5u9m/dTpi/9MFZJUZIaBRwQYiDAzo2AFHTnxZxFvuibS
59PPmSL4P17SSo0H7M3jgxZ0ikI6s6OlrPpdynqQfpZQEjf6+3W8aA1Jx1NTUL29TGlVWJJsujjc
xKQ7JWm0byIQtyQWH1kZVlZ530enhYdsSgNcuEZsynfqpQubOpEdUJWM8B1fOkbRk3zDACodJ7Iz
jvfl+NHrnhrwldhbBvWiVm9MzY6si0F0KvHLMb7Azl5ZwCwhkKVTooe3wYJhFAjzpn43eLcBHLEI
klV6ELUgY3gy3claR7R8cg6Ovs939+1RUYor3V3TK8Mh2lejgSwXqviJcZ7P4th2Er50bOv2p/Oi
Uv4i/GvdKiWrA8lJQBOwbtkqaCdT8HHf3uLKG4aECtIYBNrI+kmnx6rLvRH8aCzhoFiPrCJjr0fs
pBqtyOi+ZScktCF9hth6ko68nQoTpyTi5QCUdMQW/p7KumN8kxYXtprqCDv7lhvcyfDUFmp0hIa5
0DVtUAFW8rvC8zo8jfnHdeN8hBrTZbIiDB84Wpu+GgQcddD9EXvwe1ZfSxWEcRoZSw955CpbQxYF
KOyEMhDR5EclFCsDljh+ntxfrwV7FFBPGpWMKmbAgFYyC/MVvH3itfwhXmwTMFGKRUDampy8Wn4W
qpJ8B5OVa95NX5FDu30SyDGRMoyzrfciQ2GmM78GXVN94bv5qiRj7ktmt9aMZdMPfepiARdIUDSn
0SgZXimRTyhf6JQVJFDkaKLev6DwKbBp1StSxsW/j/aEjMWn50Tubm4AFxJ5G6oiq2jC6GHNg4km
ldbTYwgrxaDpRSvhAorWjBmTtOgS+zLRZaiZZTx+yrJiK31aR2o7D2bS12rOO6paP6sv7+d4kD41
3W/Cb3IN4hKwxTCdC8MD1MRlokgQnIz2oakKmRqCLKmjiH725oWhIbshZolDbkmBq9Pfb0+r0+Hx
VycLRIhIc6DgY8RhnYEaC7TelbvQMMnigtgZj/wtA4Fnmxk8GaLi1X8B3vBG7RmwOVPWqjCeud12
0eXdeVVkzC5ti3Sz0UQw7CCPuZq6VV4pvhENOM0uX0x4bMoxqfKAqTOETR7h7ySozLCpRlNm0Gwu
6t2TxqY3G8cf/tUg05pnaF5DGrZXcYv6M+42FI3ybMOSRZXJaN/Kpd9G+N1UaG00QosOXHt0e7H8
b6YGjxzI81+fPHrtP+M8UjW98EC4KlT9CZ69/vxA3qMRYcFk07wL1kfXGSCVJSGYSXJPZEkkdgSG
CJ7VOfkq628RoyhQEiQErrrZ9t1m5PbAkCnnIVZ8cXZlTkm5ypRBFeZFAlwd7a5dH1T2F8ECcUcp
MOdoZZCnsbqAvgG0KK8NagjZX3dfArOZLze/13ML6xThOxBEy7Tz7QTYPCeu7isWL3/CjoKWdHve
GL5f0mOO+rcyUUgpu4lnGfoFz0fTv9gkupnEar6GnDp+1v//HLITZhALTnOZFJM2D1dH6zJqvUWg
+bJNjTS2Sq0T5n3eBXM8rWhS/jJ8ZfG4s+CPqDoH3y5BlyKb0M/QOIIkH5iBtawSjUtlyDQBpvT/
IU185zwUcAzs2ld83Yrl4AwMpYXAWPuxBniK7N1VSSbqc8hWUPoMoacSD1kZP3mxfGD5F/bkveay
DOe+DGDQD9jSdNLRAfJGoGOA58uxkzZxVL5SIoQ4c1ImIClHqtXcoUA429CqVAl81TQYEC0cwcIx
ZtrVH475e2rUZ+SevdPo2ycVdPtWiyE6MYnSS2s/zF/N3JnOq1LOA6vhsgbiO+F6SdJxsn0yi/Xl
6wW1uxG4svIjjTkQ5qzbXImg2Jyi/QIfN13O/NwzLzCQO26OYeBYcFJdl9eSiNzHPuQ7vQiJoayg
x6aJnISNnCgu5ZeUPbpcpsnQOD1gxo/2DJLQMYQMLBA2vROPjpA/3FB/OeRYyvYpyCz+8SddpqdZ
Mysy8MroqghcwG5PqZj0RMQrB8qhcDSJ9MZ4bO+6f+2fZWrMcJ+bIjl46xVl5YXBjFtJKKbjhOQ1
XHzwu2uLru9rnEfPwVUn1hGVyOKNAoRS4Ti84Qt2FQ6gux7Guk5S+/kRgFk15yeUSFUvs/f64I1Q
5Jj1GwZJWr7EpHWhijedIhJ9gtIfD8SuloWEa1A+3BfXgsJWca10WbLuirERfyMjiDYHfiVpK2Oo
t/gU3tV5YJCx6e+VcdkTRqBxmOp4QPcTl06YObRNE25ZRcvaWAIXB1N3xhBxJeeGInoU56CmJeBX
t83XDU7wmmHH/IlIuFSw+uYCjNvx5MAJAZBv1jxyGNew4SpefZuCXrwqGQ4BX8/xsIgsAZ+hCXlb
fyoz5RSf2nxKcCVTqsiYKH2dEWK20w0Uj/leynzWIk3Hb5Rp2tEcR2x2b5ccCREuLb9fOXcEm5Pb
v05d4dsFxgXHH3P4dltLSTi7Y+lyq0FFevMeoyHRJGjDDec0Jx/wAIYN2Cu8v2VI6VgKfEFMxQgG
5p5qXuCx93UzJvwd+6BYcJA8qsvJggM8hRlCWbUkUzbifutQIejlAHXEelWelWrZaGFQTe3vFY/5
432P20URhRCVAchBySTqildDE2n9gisbOFEkbA12ebib5OPLjCVx5iYZcqJst5HRPbqy5wv2qdMC
9FzrCm113bWS3AbPPHPUcr4pCTL2dSUaPxDoSJJmdM3Fr8bcTAHSPvRqj9HzlTUpXUlTPy4AOofC
PYQYDQIxcFhXgVG3AgF41fqHmwnGMVd49JgIyNDTizxOixslQfT09VaOc5PSpDDbg0H+emBmyMZn
ejXN9eZAgjlSbNGXPMfbPEKSQQx9zZ/4niNYY8EyYdaAvn3SDWZ2mq1frwNeAw7e7/V4iez0gUkP
Vh6fDpWbqfSGG6QBloJOi2pCeBS55gwqIFdVQuIa/J/WnPfKcuoX+DiMKHNm6XIc3R3jDkasjP7Z
fcALKt3tOZjQ8pXakGfTf4uGfVFcXtxJEiXKUpmy/2vBpaBCToou+wce0LPyvbaUhS3XWZ2TZsTm
ucm/yq1YCLuPH6bKDNsgHu2QVm3cKz7T0wUCEVxjuVMqujZ+jEbjvZO/s6Z7sJgJrowh74LPp0tx
rLBlrXOmXj0aKr1W4dyZ95rqvKFVzZatODE862X7I3JAtU9zHhdfalJUobRNa+O1AmjaFJeLOuZO
MyL5C4ip48626KBfwoNC3zSWb6ddY8C2QQNiq3AY4yMcbHR9SizZP86MQ3svwGg5JpbcHD2Y2Yli
se2XF+CydhsSJqRkpE2dE6XBQgQ5+V48UEgJbc9TYP58BAMlRQOpU/rY1OejEYNpPCrlTzHCcO+C
pj0CVpzII18KARzWmXoOswwKXfc3D0OCNuD5+BUwXCisy+T6xgQDJdPy+8rp4etq2/gZFCkZzVAY
F6ntwv4p6TfJc1MTgK95Q4fc9IqibWSUCAiMwybEX6FtKGv/5k8VuSiFEc0IaTnRBr7ZVswHmxoj
1sb/8esOhXdMtGgE3wa1O7UANt7TaAw0lqCU9PC3MaCJk1nLUtIc9Gx7JJ+r2A4iEA+yKDuF6MJH
wXpVNr7vUTLtiWFaFcagzGwDQS21m/+eEsbgku3HU+jZdzn6aCUtRxPXIbunbRcoCP1l7QzkV/Yv
g2Mt+IRSqxMi2Ve2twJ/404wbdamfSc/EH0doCpZIdmP8/xyChstigCxrcbGNbPlr92BsGoiVrDO
CBg1nwvnbj2YTaafbH9bmIqzHbeWDBjxKBpzXcTRlEqUVqE8N6FfWpAImu91BaQqqs4TiNFYttb2
/S3qForZRf+4N5O1ybFOyJw0Un4FyUZEiMLYPZkT8dEMvchd/XQ7aUlfqH7IQ+4ZdI4/iW7XsVcj
S6BY8rAzfPe6/zYacIMgINeMu6nL4eP34vxWNSk18oLNFN4MyPf+M5f0qEiS8TqfezhC97n4Sgpa
OsgDJ0VfWmcB0jFvLkN2Dh1JlZkpTmKCb46YXAZrY17O95zUob70zmlC2Mu+RvJtLEkIIU1rRabw
hj4jAdnFvCGLXTLE+HpXsy9p3L8asOIYlpdeeLerER5bi2vgEF0cGEVaeeXNbjUlYdC+S4nNp5Ge
NXd5g1Tu3E0dwiEEO2e1hAuq+Nlb1cG4j4hvu6J3rMTdCj/Xc5I10TLooRsgPC6MRfQ4tj9+BUCj
US5jCzUnxiw+JRMdN2xD8p+gvbSor/5I0TmpPUDRjh4Gtr4kmSY6n8ZXjwHj/ut5t8PAR2M0LsF5
sdcP9pEY+n7pUKnfKdzGT9iZ4TMa9avqgxtWih3uXdP+APwFq7Dn/r/0mcre/czlHWhsF5h/rGZT
uIA8rwMfPpbU8eOmSV8Ir20OHZTrPhZuuFIVA0ScUFRdgj6IQEIgyOtmI62WRa1gMTDb2z24dYSe
FjT4dsqsqr/nsD/S9/6LsrTr22OXi8b44XnMwALOxRlnDgFwJlbv5JLvDE/uvIowZBWDFuNIbl/U
h/X/dk3YtdbEY4puB886CKZ5yl+HDtoAB5j2RDOzskLObh6Aik8XH8gL+oUSZN0Db6yK96sbIBHm
+4oheMdHmMAZKAmQ0MTA+xDWotxaNwU7nkS5/5IQ8d1dHBqxGYXaknN38rTxA/C55tVK7QCJFkwk
uiciuAUUAWQ4qvPyyhUHhumvAD6toovczyvfM4KiDIJWmXen3WcCIYrsFgSINdJrlHc5FKmRgeY1
P445UuOk+lEhLkBvbGGtTr5fuVpmtatzz/nYdkFow5Gc3895uGtBR5nVVi10Cp0l3OiWjTVsyo/1
t+GdAAWXPnNKXJ1OoJC0vNGAqSGnOSfNUSg1lDFbaI5gOrimAHRQqVBucadQANY3ex/tz6Isca3d
qlwtqT0ZKw1OWvnjtmJMSgGM12yRPqWJcK3zn01JJgASIXsb2fGEzxsiTLbfTEz6G0EyOMWRa6hV
6Ey4lfGPk+QEFGHc85tZwgxUuZc2A3VMkCz+Q+BheLU8Qx3xPszDR6ocnbV2GYXM8sjYHkd7nckA
2P+YYVXwM4ZyiVtxUhL2MEWW4oxn/ArCNJmDF8M98fl3DIcH9EyWjyDAWNVziKMG7ajFNOaN+DVr
x7+aF19kkSBZNEEGup/aA7TfP3soJL5K3zN3EJzrQ0xaUP6QL0Yb/+n2JTzpUetk++xRCxoLANML
FEdETZDk3nQJfMBVwq6EqwsctVVnB/2VSWk9eKbe5rwXmC16wFiq8Z92C8yRDHzan9XuEHLuAeXQ
IssItzb3duG45KmcbaeYQTX+UvJYNftzr1oYaRalUZcXt2sqGUPsGjbmgX78WOdsKPA9rUD0QO5V
Cnqu6yTQeRtUvYGZYF7miVx8Ho1SR0WMPFacvNWvPTBzxoRZvOVrIIQVm96LKGsteIOxfafmlIu4
L7NvPwjGxobefAJZ1FxGYIovTUZX2OYgZcbcZqMaLPccXBpR5iFFbpMGXNfn2V5QpAkicWAUvzIh
O3OM7QvROrpsH2csCF5JUz8auByNRkX/cw5EnY2eK9fl5OPKWiaue8bkGU+HuavNXsvVY1ShhkNt
clXcINDdGFk4w3rJzu4NnhcZ3IqpOCgmlyDbSBB6sV56EBm4Av0S1xyYFg0TN41MWjWs2kV4kZr9
Fu5spUwnv0VQVRcw2rRU5Bup0SBeeMmzj76isT77cOpo01YkM7bnbXLTLrvVYgQ30DRC3DFFP5N5
MIe6jd9PuTLqL7DIXt3brczlN3U9LvH4LW3RSTdP73wP+xPtWZc+CmXzUYeRIH717lBE4yhGR9Lk
WsKGeloPNHJhJWm6Mao7FFjwvkEGKP2WNuotdU9o/ASZRmK1rVZ7IUsZsyTQCSu6du3DfZANQgT8
zTmW72MwRZyw8YO8j7dO0w/wcivHvloLJakmmMwmJ2HZG7JKC0KYYHMyNA13xk6lGxLunM+FLltt
5hf8TamQdDr3K6oXAg58dufU94xlTUMk+VOMpLXFGOpjSp0vFKLsr7At78RnRYpDvGATjN3xlBTw
1uhBeGJdUHg99QQ92jrR4mue3q4csoernCPP1giTq9TBk5a65GovfGMTBMwitGihMjLal4MAD5Cd
wgSXPkzSAsBDFz6xjGffDV2cU5pkqCxOOKuA4mQg6Zo/r624cB7XFUpmwqeVhVFEsYerWTnyQrwi
ezIC+yfSNkaYU9v3xHLviP4aCtlBqP1ZsTEhHotBPGAke8gRuj5s+EUHxGsRcI+sNI7Jy/ICgO8C
NFUMZ0f4INX43rOLY/bizu6wd5trR07hZp3tt3rXcKsDQbQnHvWCTY7CtmsxsU/N/qg06LuqXZQj
U1JS48LeBkH2XeL1X6HvZjjrwgSZZV4rtSawfWyZz/qF+wJjoI0FenoM9ry90Iei6kXdVX1CY1A5
j/1I68q7VTlkNNP+pZzGUI4oymauFzVxP7/oIWfiFvpZQQxrDbX+QHtDEu1e/W52wPWeRtz7c17S
5STfSToT2wFZCoKyqy14Ez4Y/J0LEMoKjYcB+9Fur447RrvlNK/3B3emvMufKW91/6X+rVughzmq
NHOo5DOMpmD8W5ZawUjxTPJquwPGwwkMfBW4+UPTJcf4xFVgOUgYxHg9nTwi0dAz+W+Yi7crw+Wl
J96q+od1poIEhRhVvLN88l/lSdpLFd03flKyUp8J5/ZWuxpzZB97mpPD7wWZbhwPXbYqXpo/LViQ
9cifwgzfNuZD5Slh8IiBz9arLeh0YZVOfHYy/NN5cIQHh87Axm9vVMCwz/JYUApQRygLVv+7zfSo
j8JFl8LY2eF/m1bkRfM7wX70i/nEPbgQZds7GSmJIPEMb8UgioOWt/ytEQTUJD7r6u5kj/YZyUoh
jzr/Y1ikJ4qfc/bSXMzcFJBYlzmNNBUiQj0StaVZC0/fO2IZd9S1ovHfXL43Wu9jMElCkDsln2LQ
slMFVUzgVfG54yf8FcpHqZ/18zf9LAz37oLozzLgCpKNs3oUSEnEtMNZPqQgKwlfpYN45jYRAexG
KABMH9Zt25wMbWEsZdBMwmMGDEUtUeN6qw3XBlFzDVhTDbYJfGsc4bFWSCUCorR81/yJjW8WMd8M
PITcZm7jYvFr+IWZSEnquFFEIBoNzvfV+uEOYyMauE84uB1R6P8+qkD8MJVQtjQvwXrFCuMxSP/M
n4QEohzyMkTWggTScYWH1hdQJCJtGv3tzRJaXmGEyfufa3XXB4uDXGvHL5YRNSnUpL/wxwrzk4N7
ZIxXvF8Dc7GfVJlZ5Ed6rEstuzRkEjY2oZp4jo1RzFLscehr63MuM9MnVLxzGuazWzj8ixjLu5V1
AbIUXFQ/wBUC/bvu+ht6NLL71ur71Pgfbj5A3p9QgiNpYNNYsrsOJDG4UbmQVlUMVBj9INkwk92w
gj6MLPbpvgBcyAd7OYJPlnw4TBfVZnwUJgiglOnrH8N1Sy4tsiwgtdqRfbHQBYPmdAnpUPdDJRkS
ZGbhJM37d022s6le4/J6vGnzaliX85+qkxwUJE8CRUzAoRCfGF6aD8xBZqttZ9xSB0GvL5AYzeJF
ndG1ZtKpaeCj+WNkYMVFgbzZPCxKMfalwuRvG7QxI7R9u4eVmkRtXo6XlSY/hPIH6zjzCiuS2Bho
Cl8Qj01d3wL5L0Kg41zJuaPtjb3imlX4+Qa3rA0W9GfscfrbZ1d+j9xw1jGjUpzrGSZrTKo/sdG8
gd1xfkcaaaH2aIqxpOxpW/eS6kYeVXl/F5wE/G/aQvcjiMLHgzCNF7Jc9p1nefPYWTpdUqr+j5LC
LVWKpP4E0euvQG9DmRfMOlECveFWDPg0hIf35VWUoEMEOF2deT4d4qvXJuex1K4HHJYojGcxdAMJ
XTh438rpLxMxH3XIAtihZ+iHvr+nzdQ5rW2+fwl2fUbxmx6yCU4QSfBX/p3WVVBBrniw9xFvdB0f
P3/VorXT9iayFQTAzLrcESAZ5XLRdjXIyVlo4Hz8sxAhzrXe0BVeRqrMWg1JoAlW2sEWnFq/tLWl
7CxbONl9Zev6z+OXTQXB6hGD+CBC9MNGeDP+XrEzdIicaUBL4wKZ4yCtvEUuZ3Qzlb5c17ta+839
b1XC7qAquCqdZlO3pmrkI3RfRr74Qz4bnsd/TFps5pbmJuhtURICJnx0Qxj+JwIjJQS7OqB4p800
O8q1HVEqg889S7Ex0BjzXsfzfk8/zEX5RoY4ZDMkBk1nPZTBohgpzoQyoQ2fu2EXPC0vJetqy9tr
KDX3MxXxKVsly0hlt1pkSvMIpHHZ+niI4rUio27jy3j9UuEr1iZa/igt6fm1TB9fRJofs9D6ipwt
L2JLeWOFmBikCZdexxOOFyJmFBECI78jwkNXo+ZiYEnn/NkR2xUNJ/aWkFPDQNxfHQF8aAWWC7y3
9P82oZOpdkIjhKTNl+aukR4NpHDskjS255nYix9VDrcEUNfdL/OCbi2zmlx8cwlkNS61PgxcOvpr
3GYLU4MTP611xYKzzCFB6MQyJi5Jz6p9OxpWAAbh4IWGJgyvdp707BRF4HwuqcEGi6qH8F5l+IgF
dZcpyYwdW+jrRbeMI5iNcO46gDfsMISNb1mqgiz64cP86OUVLRFff6gHHjNNCyBLnT0ZqB+HW712
XdP3C+8XMOJhfzLaDxuRVzbVK0sdXLuN+6kxbC5VEn+2kkXSOEPWKIddqoEWVwcEE7gv67hrafgq
VgwXcW8hV8IAp1y37BFFXAEa9YzmDWOmezqOsZ4lfYN5ZtK6nG2SUK7c5WTJmhvRRaeMD122XthY
RbCWVRcf/9kBTTRdte+oh/umMXanZp7jq6VyT0tyx+5OvCQ0HJZJGE7/scIIE5CeU1gA6IC44nmK
7//qnJ/hHJao4D1qgPVI2e7qhiI6g50rLYpnbzyPQqgOHKfAL2+fNSFMncEG9KZ1IVbEeYYQQbD9
9t9cdSHvgy/TmGMfwaeIkSrsVYBammUfv6mtQhkx0FX0btIMyVyuJsotF7ebE/DN2oEqeT/hvrHd
4Ymqt43tZPHA4IRS8hM8eXNju/BfEgDloC3HbK8MNt9euSywwQStbD3fFqLIvyeukb51U2S8s3Kx
SGBUpEMk5XaWC3ty0K2Mv16cKHiZwbTAXPWM52UaOXsItFOvHLmp9fhZlpign7ae8GCJsS8/893X
gGcR1BSXiUCPLOk1aeJChafhJY5OXiUQuXaHUr/wGk32SVMP7lSTQZOtuZHUqk20JQ7Y13Lm2olw
23dvDTVU9Y0644bSdi/CE/LPlLyv5HjlMCu76YCDk3Rz4jyPfQ0O9F37jXMIL4rsaNl2qsWC4HVL
CCMYfpEs20LfasS3AMvLJJe+OCGXzpTRNJKCNK73uN+AwxEyIeDnZzwhcxQFqAUZP1orSWd8ACci
Ow9WW/Kkg8qpTsnorzX4Wc9PPvyMMs3ZO03xtZPSa/YbLFfLZMakGi9VgUSGT39P2ld7yDoqQ1Jm
uSOM6+N4f6zU5EW9c+cMTsaRpeskrVBgeDGZC/D+LCugc6agT5L+5I3yYWNCX2/u/rFVylf/MqHh
55BH5nrzkCHefhGNzOOFwTzz4V6jBE7PQ/oaynxsuF0D3cya4GaYW3FygvReYD6h5OUVdSpGhQrt
Y6n43gzvaJzyyfodHZCndKkjOwBawnV9SN7DqD88uNyZIGgFw7ycwi2X0LwX90dyxfVQcH9Hewc+
m4okr71DYdudApcjKC8jrZP84j3TCah0Md7CzV7yXIeIPd5wQI/MR8Rg7N/RH0t4vRuS0aVHJJ52
PclaSh4BE7v5K+vmN5urM8PEU/KBSSI4o7ZpwJNCv840Zp0rffXmy1jNoHNbAhuzLf/vcdmB9+JJ
YBTQs1PBXCKlpWcENAINU2+tWdRmolcb3KKvM30bvWej4pjpN8mxBBijT2+phagHNxPR1tof41/a
9JDlhdgBjWgpULavhmdryZzvcdFqLFtN8F8YU1ViJ/VWTdDeY4VkfVj1oybzFeOmyviCTkAp4+Ds
io00gLQMPA32idsLX+q52WdIIdqeGvc+7GiX+emH/5zpwE3BYi4fskRANGKBujf/UOfj+WH0X9MM
EUZChpxQJhub3Ga/LgglltH0KwD0g/AnFiuYbwzhW0w+VsRB/6shpSvPi7xwH4w0fy6RBdO5xVwn
ocgprbxLQ45827KvXWnLk0xj/rL0ZftwiOn/r0jywOyn8jCK0weGzwVMnhyhjD4BQWdTh/UDXPV6
wc55N4efkdXfNg4G9sXbNcLMuCL/r33xF9nsG0fMjn/Ip6BxZTEEewdLlAD+x+xBI2U8h2IB1aeO
fBKO8N0Zo9HoU/9qPhFMuGkNUuApmYpNb011n3cC/ekvMLX/qj+mdbWVgR+0aMdL/n2ETLFAwNGf
fTJ1wcxmanp63AUcBswAPxuWCqZIYp73884zZVsgpwsnslnJUsjWl6niwBP0l2bXChx07K6E6lEW
hsT3QEjRiG9rN2X+BdjqWgtjLm7+grEUJkmhVGD+HSkIHYEX+7N5Ejq/4JHHkbB2zFN7CnNM/4YU
zWHfgAo6WT2ZQ4i3hZVDaN518kXuwKAgzHEHNqNM9zUaIyzKwbg2imOGaSWE9tnLJQtRKceji7Ig
wzkkAvecvOmCKyBlVp4TwWSGTCCCt/bWdO0UuAoJtpL5sT2CbNUH0L210aXCrA0VRSVUGF6E9tK3
BCNHogZvGwdJIPYBEp5wvHEr/9CBYT8p6u5L/v2/9x+rFhvieNXw5gxXNZ4hdSjP4NaGNigo4b5K
LhSKK/yBZ5ncboK4bJCrPOeXoGjYW77gxvB4lcoaHYwtzm1+QIN5f+fEmBrFoKwT+i4DJDv3X/IY
1tq9Zkem4tDHqxy2zO39Jzj7AVutIXt2/QIVNk3rrZfyPvRfTf5qDyPqyU5Zt6nsH5LW3L0rPkjS
U1DymojKj2p5cQX17OnfCdavE0GJCLTbXOkmo4qdhcr6ONVCMfxj1nCcmOy0sQhPtFG1I0nnHZRL
aeLV4pkv4nghGsgHkmdyXm8PE0/WRUmJvoiHhyCyEdGIBE3g9rt2HyeCZBPE1wEoeI3BaI/QAOJ1
NhqWi+bOUgE1M+KmmE5xpNm1DYzV16hHbF/fnvnOIPB12bMk2UAOefiXL/w8w3xlKcT9u8iowTgX
DTUgekhMY/dANUPamzTNCvKruvouwAgwUnqPRxxs0iReutwJTlwSsztdvpLly4AWXfFK9GrmSL6O
3YPqK+ktGSjcTE1WTrVQCMcN7pjXx10igDVG3oj5eSkKiFDqRnockXkgh01c/iIozlyFRXpe/uS2
5N5SCmE3QGs3TesW7U/TgDpRwazIhWXqMOHKpYHoLEXVauQD62UtSjNjuhl0HwnI9aRT4fUBVNHx
tlFBFnzYkm/SpLE4TODPZelaCPOCutddHWbAe6u50yD0+MxGlhhdw/nYeKm3F1FVxHHwGuWpgzDI
pRZ9tnU5pmtjq1xwEnj5lmlv56RSkU5ybuEJbgRXpwCt07MwdFcxT29WiMwUpFk96xi4X9gcw6Lj
5Zx0ZLhIAGAFF0p4JQFzITLpjOXaI7FoUnq3rJUkt+RA8RDIpjDuMtgsU/p39qmIPVNq0raGmerU
sbYj+szXF86jcxOq/elfp0VLIHUoar4+wwBMKoEQSqQGH4wBqzDlMRg+uilge5jETem757Bw9edk
Hpfu/h624tHxjJ/0Pn3/ITKR5URuyaXRBHfOkauwH6WEsP87kzMjY+LMKXtFDUYfdmwm0AuhaGDW
XXkhTU8ZhAu+GklB882VDJXCFgy1yUHLTUQaMLF/zpinVn4dKj99v7lpWwYVXs//VcAvG0yezowP
wRqT/8tJbFDN38OOmvc98Z2y5V6hxJ5zOGpKcktB7xuP9XM+qD2+XSbb2HsFspI/M0ZyhbB6xNqy
Uv9NtfpdAQt5Z5xCDRylIHyZd25B6+0pmXb1nd7uN8U22OkKvEiLVu+GlQNs7UnFlBPz1Fc6m6n8
0fjA3Q1vnj6IA5Bl3AeoM9CkhxYw6BicRkaFLV3K59yil5I5wy+ypkYltLIA0VATOflApbziTxbB
JvmfGebP0AOkZG7c/AWXZC7TGwZO2YCyGYaQX0cgkUoY276JkPw+bWjetPJ9Wwm8OsiJ+Q4Kcgo7
i1rIbNqdiVcduB2aHyll2MG5wEhuGxtPweNUiyZgRqK6e73+nGQYgHLPZQVeuWXXiQ1htI7xIYe0
mxKP1Hj0k/ZW18/NT20ZKZL0zFrW4lroIgXp6k5azMIiaE9tbhSJPgkOdTR2sUxei/lGyrLw9lfj
xsvXQ9867q+lNx7wbw45rbYC9UYeSVg2lwD/yzUuvD0zVYWuuy0byEGoWGZsygxHIY0Fz7iwhkwc
m443OU3kGfJD2pCgeJcfMjPFP8Pu+61T6wj+B/RCTwIyUs1OyVY1HfY+Sh9WDJOp19Lb4suMwRuZ
uJKpJLvBsR8LtzqqnpEWCCahZMzxSisQNi8pQlrAXdl98+lSdSgErRrsVr+gzffo2VZ/iri3v5xi
Nb7tlb3j8c1/FS4zDwqGqk7Jv8+0CkWgmBN8OTPlEEoz7qX5FfX65F4B4MEXFpSqgfPTowNy+2RI
wjYoWGn2bh+ChT/cw9ZXtnqyRZNwvh5JHWz3TslGaBvIWyfmcBs+te5ptXarchwhGdihsESRm1md
/Xego1QmsZrV+8zS4C5mCARGaeNYxE9XeecKYlk9DcXGJ/sBrWfsjClAfI486JsuoLSMR3Aui+5x
LzFZ52GcWzSMcYtVIcZHZ9oP/8I00uMVW3Y0lkTqG0QLGlwaB0Fv4uu74vV+oDpFbrbCmWI4yIMS
Ocd8aS58pRK+u9b0k+sAqyuwKXNPHurud6GdQyN+ZIJN4tLkLG9YjNyZnShPet0hE5AmuYX7KAdq
PjE5xqNRhI0chwLHVrteQuiP2HPFilWwaBQl5AoPWvsmyl9iOX18MqF93QeqWZ/3ez6Vjsddf5h1
pGbafg3dwBCnSS7NWQhyzbdOLNeSPjv2lj/4sU2fKRun1d4gRTarPTtRbF9tuqV8bcedRksDSBF/
kgj7llGSXGVOYxq+3eS9yVjOSHlyBaqxgTDbdEHbAcIj3cNY18Ag97r9WqaN0r4m4iie9SpTc9tu
qh9yMvOPJNgkc6b6KoS3uI4PBRGFc3s0Uqv1+ZuXS/l+7ULcvRVsfh8RaTQGIG8Lyj/ks1ihEHck
X5kPV+TKGE+IHRY9C6NIBSdoIpIktQtKV4Czac+Y6ViwnhYCeV+33CGoMTI48KJWDs7bZOYy4LKO
RIKoatX6U2gJ9hXCFTFIzal9Sss8rlF9hcCF8cUrXK0CW1Y7xA31gj7ug+l+VWTvZVv4AJPbOIQJ
uY/NbPNdCFsdFTKgjAilJRZMmEoahKWOjGnD3/Vqt+Fgys3bpjA2efmDambWjomumpY+/WaA47hy
/gSz7e4alFUN+LtnSD8KkxH2pZQHlrIsfFcuGaP8hL0mVHcZoNagdq/FvKpeawh58WG1VGFftUz9
qHP+HgDl4ruInV3lkWGSOueRXXSPMRfWqp1vjRUBi6V/NCIgk9Gtq3q+eM34hL7+uEv8P+2/O6Hd
hWOGmTkh3BVK/Pp/TRmn2QB2kC1+2lDFEx2Pzd+NCeD0rXc4ttrV/CTmYP2fHwUSXA5szj4cH94F
Q7uy3yAFHZ9OzR9qnR3f0IgfY4Up93e7RxsOFGtWMj5iD5PeL9b8yOHqT8okMMGQ671+FUZEUptB
cXuoRdmDeuhh6X68zb6cKVmrbl4kxt/hes2NR+1kWuky0nAoWDw0XCy7S+5nCuTrjbiVcScmaEkk
6LfBn3ffOz9Vh0BrcnJ9TbqItogMxpOKORd4lpx4laU7rvdM4UP0YhYWHfX21bZSaNO48F1M758h
NeRNKsiJdvQDGxt5eYUH6FI85UuTYI6A9TYWg3iTx08gpk17s+DHPW23YF6qjSKZRubIGz9G/QH/
vGeQHYvILJoYgKRThc1PDEcnKXMQVVI5W9TSBTYUHt5CeftjyRx+wTvNny+E2cPwr50nzxeG1iCO
oypqYf1r01nHjoyC95cNUEsZI36VCtqlBHONOpQWinItAarlTZ61gvUEYCIiqJapwKqwfsdKy+pF
iWUXmdQZoY/axdLaU6Zzl5SAo3kkFyxkZw7wHzt/dapRRVnm7/kxDhHetai1nNCJYZ6ZxGs/Nv0d
HMS7Yq2GK8Rz4qHRpRAyP3GTdKXNBG0K5furIOxTnBzTF6qN26QpCSNPtW8bbeNiYu4Mr/4DpbgS
1EoKO/0KmtlhK7HUORCCHOPGk/0XlQ7JnXfzL8FzImuEKhoSD+HCTR2zkEuM5SGNSfFrXB3lxvQz
U5hhdjVQeBFKIsd6oLNfdcjvmWr/R7AWmbEYlg9JltekR8+xc8/tygx62dg1ZrN8k8HOwh7J0Nri
/1CGe+nZF4fjgAXMofYmXvj6+cIypI9MyeKslmJwySbe86/s/rgd1WOhxFuXYoFtvTxztAKpHOD8
W0wdTnfoguTaobAI+ZcCe36jefFn4UbOUce0CcNUgrJ9Y8tJXs+PYMNBzGIREwuxD3lwd6LbT0tI
uYmdYrmQAVovcgdI4Z7xmGcNnoA9R+uZtEOt44aLWZh0cVaJqw38mHChFANtDgcbGMgamKaVkkMk
cD8+tcrrqpOZlPxiVhlq+2a5Dn1qghblwcJ404+mHkq4GHtOTK0TlM2tB0lmPL5BxQbMfpdbBFXb
FyYvEPsIk0OZzqCotH+a9owZHnLbgHnAyOBnU9WkOo3dFMKd3HRu1T3QBVw8TsnY1R4nqcmztuIB
OPtSOBhp86tVvd+DnvRAhQo6/MIRKNonfKWXxu9rxiQHjPO0HDzM5Q+c8GG1zHFe/WOq/U7K+SNE
s0y73cFxZNdGKchqwNEjBVxMu252RzHxLCuxtML2aYWuH4McZcMQ+4Cn6L7U4WAxfvOQCibX5g7o
k87d18yTlyJerm4uXaKN2E2N802BwXQikcdKNeTT8f+Z9wk8yNirIpDZE0BXi8441g5/84tGP9Ml
swPdZism/8SJSxKheHHOGlCVL7uwf2uWPWL+N+YtxJL6ypkVj1ayQlCoj/ZAMEljbkl3XtE4y9t6
bx5slPQUcaN4h4KyPRTD6sRtTLNliUfirzMZiMZrMvYNRxCox3irbcWNi8B+/1pCFwQOmb5Da3hB
M5DFznMhr9NRHBSQnQhljIgSOf5PnImSww/cY36X+HshHCOUqem2imdzzAE3nLRdHYk0QFFfyzt5
UPG4PZgg3rrC+1X6Nz3qFW74QuNBVma+5Q3MxCCRJGQ8n17rGRAFs7tZYTLEn0Rj3ewE7iIgF9Cs
lk2ETUe1lGH29pysNHoTdo4Nb/aKMbXbVEsarcdwwGXdKwE54x2c6FTvZCt1lsug5U4P3EUmaBQ1
SsH3oq/Cp23s6Mi/e26wm6hpchjPu7rPoWWU6UXYFbi5Wm/i7rUg2ACUGrUy1CU8zOelq0cZHtMv
ipzUYterQ395IprPvCtfhcOivQEr2n0YAYQaZZzpaWex/vHk+6uRPXGkXy+whEEPBSlv3r9iLbVE
aGegCalZDUzFqKFxUCvVM2qnY8U4j+V6Xzjrryimp16b/6Q9ob2PGmOaheKe1X8KHw0NDm+gaFwq
kok6uRPxrBKkIeVtmITXYcC6Kny6xNiYJYbdIaqWSKHRLnPqJYQrbYhDqU9y+N8YHzbNE6NRQtTd
Lcvu2BUAo/byMJHbQHDjqZgzR+nHV4TBskW3kOC/1q56BF25cl5Ctab/W2bn8TVB8PS3xs4Xv7gC
8QAghOfWzG1GqkGa+WVSZCPe7nWQnt9FW+IYysUSJ9aFixtZuT4RtYBp+4s4m54OV63YuULYB6EA
53g/sh4ncKYGbqslEMx1kNhkoLa+fYpwV7Sa6/42thz/cgzMnSiCfiW3x+CrLr/cu6dAjLX3UT6h
t0q1e7K9A99fmcVNyGGkfs8YS2wondc7MgOz4Ek1iR9vJm/gDloD3skTepMQiVR6Cq/6K+qcGDbf
43zLFux/evnWu1YM5E9hgslQRItZNJVzx8bnU/xSxjpo3j1f96NXHqtal1RyCkUQSAj7EoLp0cIm
w3TD4eFy8XNE7wjBNnooVoP5kuCm4O4TR2sH8JGNAtfaeLVW3PG79e4cS8fDnWI+Roi8xxRLxdmt
Y79LpTAnsrhzwSq4GbcL0UaZJzGVgPK+NziFdd+v6MCVBWbC0BueVZrit37PVVtDhBQ44bCdNo2V
VFvT8/pWGehzkM0YRlLnC2pFLtt88oIsDwYeH9JmRxxnHQJX69KhkQq6xZH8Lsm7ye8mvb5yOjDT
4CTdPMdlclxgr0yaVFFLW1n57viDaaTblkb913ZOmPWW3/5wJ9m8P3VNucJnE/jr/vE/eOV6h4rP
jKfOANcA/2/im3sfvKovxaKBpNx/CsMWhtuPYMYQbtrr6cusUFGS0Qe32uU204eK0P5IfJyZxfwx
BAAM5VY+aUec9WK7CtLfzl9P373PbsJe08Yzqo7MMUZNfnsDE7ghR6GDrEl7e0VkNfezyiJwtviX
/kjXKMkcFxwdA+OxUpfWx6wx07ECsk/VgbyTORVkxEclqb9k6RV4+7J4mymQy+rS2EUdT0FFJ9Cm
JEqJiJO3CsYKJolOD1Nco3zb5Y1fxRLGRlrWcR2zIT/AEl7dyDHb1PKY68bba4e4Y+69iuJNkEDo
NSRPjWp7u2QjdURP/JLkotzXKIYmg6q9QksLG27YK4stmvC/+s1sKIBYGZQCIVNirsGk1KS78uhR
66g+3/PTcVpdHh7mm0D8QcAb8fE/DiC4PVxvvQdERkQejOII2kbsj3P4znPyXnXPSwTeYJjl3lB9
B6g2mu0+YgukDEsJRNjPd/WkWgPawkIVwA2qy9OMyjh91M5PZDWhTacvEv7FjjZacoKwMRO84VWy
NRiXLasonSiNhAkJBvMuxYRYcycmW4f0GitQDg02aMTmBC2lDVWT3KAhYvFVNfB8HgRGfeiSfVXo
h+K2Bfhmcdc4q1byXYu1uj24hAf3e3A5ZW9olliEHTL9+tSmvchWXAK0+CMUFS6hz2YXk2J+yHCO
HTGeqETtrnwx3oighflieigjeNx1PIRCYbS+OPcIw+3CYrBK9Wa2eI5oHGAF3WdR/hmJB1poGVro
9V6ACt/n6Ih9a2o0EL14QQpjmVJiFM8W6pWBKCLjjw+lIrqXOi20YqVXYLPx30mXonaCgutVLbht
nQc3+cSnnkNMVhUo49G5y3a3KrzjD7THOnb4qATRZJGgT5BhZ0x7LZhlqsZoOKk5XJmMscNRxdw7
UwX2VOsyTxlp3Jr0HO1RY48+mZFC9pbA4oc2rd7/2IHnYD8EvxgSrcI4iOkjNrLh78dOV4nw5abi
qegDuWEaaDyBOVjhzBy65SJ8yolCnFiO2fEbp4Z5ZqXIfabOE/+3oGfUxhRgfL6riGktYGBQfh9I
zFrOpu01ojSQW+O7/5UyhZEeJQHNrIaqsGiknXVpYvtsYIrCFajYq/DeExzIh0BBQ7MhhsfLg9a4
Mn2ldvrOWEMFfMyCeXLV10egB95PDPlRc07YPH8VyUNLFI5aC4Inu/yzFLdfJDXePes+Mkuw73AS
AMRKPykE127/kdkwsMSQHAiiDBgrSDIwWnH3XUbrG/EvVQgkBKWSTmpRpMGuSn1d91SkJWkXZ7MI
SUkcxfQWef68XXvK8GGqh7YtQf6OcjXVJaLRqgz05/EUIdjVkz6jWSwvVMTKOpZO7KNgF8tP016N
pYGCfICIdlCp2zgqwP5lbljWwOPnqfin19FdvxvKkGxexCGxbU6fU+f2PLBujNJLj/AEBEgj/bxi
gx34rU0Ygdyr1rFfK0+dknBqOt0UExwj6NTjwwY7jD7hjZrouIZXDoVLYJdLVqw/j3Je5wT7FtP/
j1aIcJiRjETYfrsxquT5s2g6QMqEXF8/Ll6V8YchXOy7Y0arfwACNPd9K6QeZo77If7LdQ5vnMCF
VW4wlNkhiX3G0vYNYbON/2tJV/R+Oz2k7uIaSOC0RHkRtNa95IUkjxsNonJtzuabIT1JK4jRJspd
X9S5u/CjIkzgNtiWSEm7e2SylQEJ5eScieUWfT/o0w7YrptIvbKP/jfl8RyqQJdsTve0Jgq/BwAM
bOvHc/tbC2A+b0cKWujC+JzFP+3ThUEComskr1yekc29hd8Cf76jSVoDLP7qHRvee/X7Z5ogEX5w
OlxPMWvNxZ6fBQJfRCId5bG49iuBAFt0z72IbzUUckBe6UPoyVgfuWld24jil+ZeKtJOpdtL3WJf
zuQeJ1zvF7zLPVh3lACGarQpGdLKWyP3XAe9skZ7LC/h6CaLn4OLDYfTFvikV1bWUZZ+f+6W1gC5
4Wb9dFdS/W4XYJrPwQioe03XBD91aFiMlnxRMY5s0q3EYaro4J3l4ZhhK+G6nsMiIpGedG2K+luN
xV7fZKec9keASmv1HGBPhaCSRXOhYF1q5dxfen6m7UpzYEzwWNJQdCpeJFlz/0TmWXDtSioo+kMz
28J7PEZ079XOKqkMt3R81ny6pe3GgjB+BdOSx9JdzO15RMwu93QeSIzEizDYbk0wDKi2KpUbD07X
IFimuu27IeDH2AXTKVnnBUTqudi/tpjxrrXfcF5kGmi6FE9KChtnilfw0T80sZsjMaGsvIp6rAVw
2MMjKoRSzOUyC9jEWOABcJ0p1SdIa9fBaHDb0cGtzK2nzLNBhmZg2Z+wWXiiw6PP4DhsySvfjyUG
0a6IrzGP/TH5ZDKdzEyPPmPfBDEQXRQtyMi/Kju1pjvMclX+oi+a/RpIo4Ro1GKpAoV1tAIAgbM6
J2kvKtP14ls7f+lqh9J5k4zLsvP/Oj9OtvJe5jDXwahoML8TRwy4X6WvLTxBg9S7ps3DvhwKQWZi
HXDDL2Ghx8aeDEIl3TIiVhuWYcMHFwkt5UfCcFAou5WhorMSEFUN4kBSfNZ3fm0lQiwIZILr61Q0
rXY4v835LasCsrr2MZx0RJpgnhv44iGncaTlyfber8RN31b1JvLB8UkNnCStm8K4j/h+AJ6a/+38
coYXWOojf7YNl7PJPrwn20uWecfuEEmd9ARiuY0QFQUV1h2ygreGp5fQ/tFbGvIGUT/7fZhhFu6L
EyEl61KE+apw+U/76JlCVeFWr4TV2GQUvJiN1ygAWHZrwyrDTqRq0MiERmUKpRLVhOZyfXO57XJ8
Y0TIx/Vjn5Ls/SPLN1xa9EBRhN1rQYYUCwa3mkPmaxTcBPui/lgNQqcAkwYfGt4Vm/GzHQZdv2OP
wHTuA81rBE7cyzDT9/i/lz9ES6jDCm8Cw8E8EO0AaRiFMZVF1wH7sbpD2PbWseojuFIM2VP1Nn+u
FIlfQlJ55ravshizH3Bnya2HKM/lD3JO1MRLJCbPjmQ1HkdlMEdCOB42+o9U8E7nsaL+EaooKDxg
Ld0a/pjpL0Uxa+pvukvDNlQxJvMo2hSFPDKyQDCsYoWTKSHGwhcI819aB6/7QQnGEQx2JXmgOluJ
0wLMVeFqBkeYQxQeRuo+CKu8cE39uUI9itGivoGSndNq+pOtVI3Kk8p1bDwA6d61LCs4GwUx11Va
piIy37Wh4ppMPUrfLmETjZwkqZ6RBaU+Bk8NlHXpsAESY1bL+r8NqXUlc6uYwGc0YZrsVjryjR9c
nwgYAJs8xG1Op5lvpBZOFl/I7C4b4gT/XeGnUdCun4ilGol9qzfvS51MWTm8pIIjnRRY0fXzTUBh
nz/wv8qeNCkSXHWrw88rHJlvCZ4d6yNvT4piZVCrQQoEi6rf8u/iCp+E4+FZt77IU1cb58SCGYma
BuvWoaxKiqGrGM0vWBPCLwYmvL6F4VmIruHpH+empiJXfmcT2xvkpbydxYgYINorocA7QurXd4kQ
6H4dVvutkPhJlDGAsLRBZ0pgPykPNXbQ2o26MOkGjXE/3WG5DHyXJpUsgMXxLY113y9l5J05HkHM
+/A/khxSgMLQLST5G6J2gpi25gh3dCb81IQhT2PoiZcIRY1t62EFxKzVFeYIk937MkMUpL0Y3w75
LsAbhwwY/5wVh6L0esFZ6GEHJJ3+3Jf/C+WqJdSQW5Alr/4FCrwRg3vgfDoLvoirlND1vL57rFF1
3vj1MA9nGPlRAy5TSq36JgVmFm4HDy5EKi+68JAUf7K3XF/ktT3FGyqzHLluMLI4AgmKiKukxebu
ZRoK0mPecvFaKpo735H+odvPqtS5DT2v3R+RrH1XZZYosXunsj2lsRbdeE/rpaBM8sHnYekKsJAX
VmSB1SEvMqJmNHD7OHNpjzZpOz682ELhk91umQFLDutVAYS3GOhru3VOVqWiDebVMCSqcmRdHekd
tFR7bFxVna7ioM30tObIILDts5twUHT83YsEb6V4vVdapQGkBNbspLrNtpIWNPQ+lNymLuIYwW/Q
l2oPVdHJ8MOlMTpJd50ItcloCJQiEjdd7ogbCukBVKr4mHeW5U1VSgSATBYi5kvoTKgpZf/esgfc
YILa/bY16M4n1jvYOpbjOGVDSW/en153IugBDJdIkEPBU+N3UOAhLM1g2XIIsMyfJzn5GbEDGUHo
kL0sZZYtBrfzoWobqmxIXjazZ3oH9B8wgTcmscLYwBBhqWdTGIfr3/wbFSI4ipMArGk6cBecmZPW
ImF7zTyA4te0N6Mxw+KJHlSwcykmlH1e54t7QlTaebSbCtwBPGXEFfs0qe0HaSO8mo5fjEmOrJZa
9oTNn92shXWj4TiSgQYDEQZrGejUgBYmu9kO+EDlnVof0zdectATSF/wtISuztrcQj+tAJbOi1Gl
7Uo6+EjFkJoqGJhJCNhB5SCM3O9EncGPPZ6H6nOW6TzauoMFGpqU9tOeY+10ALi8/1EgaznpQXXy
xI++VwtRE1jXNr4EfC2RD+LlC6MLEvb/uvZ4/3BvzvXwK8fBjO3IH7tWHfwIDBU7Yt5W/ZBnr6Cs
RjXGZrEuxqoru40oY6cMUsi3y/HGyyFhI4zNf7bTBSGkAr/xbMY+zoOYpnu6NuNxPjc9J4upnnwZ
+BOlnffjjvyGmE2s/oZj3Hcx1hE04gcBlJNRiq9a4shn0m3d+exIk3Lo9qfADjDV1HAWcQR6UPGK
djn0vApazQOrZFrnp2vILNENgFztLGsWABNIxrenqx/rqEog7IU/Lb04nsHhOBoCkPMHfJCMWIbq
7u+oAvA2O4ylPSyUuW+Ae6nWI44iT2UsXfOR0MeXmdBS37lMRhVDf6fi+TCNR/le+dNxzqlW0Ef/
gMIF7+HCLqFxvzt4O4NmYnTQOI3M259tyQVaiNT1qOxz4rz3vslebZbAe5NaIWFMDaLRAaK12NkJ
hwFB2w8njnidijrZG0nlSXeK5+nxkiXDk7X9zxlexRx/azUdSEllDIG79StWmHiDwHVcoO2xKxOl
Y2bkJS0KKaHpE4cOF7noWUbbGYrEj5eKQE/5JtpYTtA31k1rosHSh54TBSwc9YE+PXvbaXgE67mf
XRDV/PFsNWOnM4UDs3DjtE3nYpAk0vnEBlsk+58FKPks+feeHcSAhkAUe15+tJrpwwejVcZLRYFc
lzjfVXApZbT/RhEQ9ASjV3lJfk1OxxE619ktRVX2ASZRWnGqv5FiGDyyWl5Nj1LfykDeGDietvRZ
zWLwoxReUAoSD4cDKR+w9fB3mSjsct3vPi0+FmzyLIkvaJDbjZZuNefeolPtqodzp0gyp5/Hn7nv
C3QxpGZSCdJmLwys/dq/yCmPhKr+5y6pl0UzMFjoDvnTBvwMaNlawVP0DG0qELScpFlJgPajmKPX
3NKfD4n02rM395ZaYnoy3dQMt4APVHf0oNpvCxf738fTjaJd94brBi/yhOKsFkZqPySUsQ2RqoRU
e5I8yBv68oWxy/SZjCfxfN+hmZaCCD7DS4BW4C7/w3fNTI8dBJERMCXFcclsxSWAQhZwhy8le0ao
LzkmD5SYspdQOA5fMFDcs6v/MRmTWJavws98NIFEDEqlZJcPf5mxCXnbisONeSqEr5ZzPV/hjmdK
4a6xg1rj4j7B5wo7QtRTE1s47qiQJTVhCGcSf7/KF59YBarF8U+hZD3cd1TaFan96QPVRiwOonzm
4xkrRGxGxiCKIsDLk+yjksXO7eHBkPCQhjGN+9+oeMHyE3Va+lcTqJRHAcC7+O8AzP900hV5k7aV
MDaMdByVxsaLK1n5SYSjvo2yHfVysgkurPN98Q+pb+T3vzk6DZ2rHSYjAS4WdWj0mbk0lyebV99/
hB6q/f0R70Ke+HKS9nLfiKhrwopsFjIVYo0OXl+g75zSH5yoRwwOgIwDpYShXskNyHUHmgBaTLkO
z2zcipwylqpKnouQYQEDl84qQq8SSYhXCDl57FDd7535R7ph8L5HJl01FIAC9iOES16fNRkJHyr0
lDTQfaV/TKabHTpPTRkhBej9oqaw7zW5vRbWbkJgzYm/aHfQCEK3yoCihVOL/FkbSQ+dCtSz4GhW
A9vFPFatzbdu7NbBqIGsnQa9dev9kiPU06LfXQ4W9XVqhjuw8G0R9ITzLz2bqdfbD5yyNUuB55mM
t0lR/uem6q1MDWb9/cc78z9ZrcdktF90qz/wOkhPsnMX+IuOMm6IQg6SOWQmopnu7ixb6wVwZH1A
RhxVJzj+ZH2qBimOy1bpEk3CEOoFL28gIWQ5OW9LI9NbhpmoO5+wP0vWv4u9WAGLJ+fk+intq6a3
7D30TXbC2kCAonodpGjBLtA8XI/P8QFBo3vUmc+02lACiwoY6gV4xghgwrZ7ql3c7wLxR9MXmkMT
+5xLFhVOzomDyyCc+XfA0wc1mpFMdLYnEdraqQFOgyoyWBzOTxLWnczesOI8+hbcQFf1e8KAhDJk
OVyCmMpFNi7dZikH32hPdSL0Hnf1e0h87R7kwRDUShEkXuXmdGyo1YpV/Sk6w22xCkybLyjWyymN
P4xY92Zf9dDiJ9k2Y8Vc6jUqsQwQmA+fOGLXumwMRbR7FbKOWQ5DB5ii8b8dO8EUBjO5R7FXIDNE
xEKgchLczXpr4ejsR0awfq/EH8g4x4rBBbar0lN90tyET1sm3BGSucXQ2McY8FK/poG59yCjFoFS
h7XNhWoqPQ2qbz3Vr9vwshWMBVOG/XffGv89hzzPQLeHMap5IKjSs3ncerNXNNNlQ7/fGg84/6qz
Z56sWoSVh6YcNX1uC0aLdawiZOF383eiFs+2MdYdWklVNWRbhk3X8ISa88xub0QG0Ert/eDzINN3
ZbLBeW0DHnPBV0WUilhFJPbmdN5Pm0Tak/fvE3trO10KrmIKg+Yg8M6O5bB7F6r/n2TM/TU/qKle
ROSCgJ9M4YwbUpEiq4WxJP4czXJHhQfFADonC+edo6jU9lwRVDd3+Vpxdo2kORS/DVDSlfB6Og1T
vNcRRdFc8mV5TB6BQWp4ikzmyduO5/FBkxJYpS3SkrssCJiZFGGinSLWpJvRPgtPWSLFw1NJwePR
4UHMtgtsWhrQlRZlZClSCF01NlDqXmRWC6hMr5evqgsTBYEhjGstxwvLy2skB7LFe3RW0o1PrKrb
e7AOKOKVuF00Lv3Y2NonyJrpuT1wR0QFbTYgejC5b/PZu6eruDlhwnm9pdPqWXcAzl/7djlSuM2i
lbi11UJTFYG6KmgSmHUhVWMdBwRLv5czXPBZ9fmrRoVEEtlw3OKvwYBN6cqnkffNb+u/DkotZBn6
P4vEHNDKZ+t7aVKc6jezFa/RrFHHWG8dzOAWTrzDpYeGwlSbsVIr9c+l5yhwGFij+YcOV4Ra0Dq4
7xu4BX8I418n35H6xcET7xK5CyY+p05mlE6HHS311lV/SIyp3ohDTeyOlXHGQjWVq+SuSZya4kxS
bnjjCzEAN7qoNkvGDGjeRPlbK8pIvo7d9vHsse61E0GmY94wMz+0Anelh7gc9CC2CSX8RpDir/KP
rMMEzR9hYI8U6lGFcqM9+BfjAnKvbLVbMUJF3iAE/K1JGVI5sBKQg7aQiUX27lYO/BrM9O9p2TzN
gODx3TD5Iyo9znqdmco74dUwX1uEi/E726n5+AqsHWKqKuJo8y5IIxHlOPitsUtrAvmYZqokANwE
8J+Ktp5PMmy7V2jk3RSYC/6+Apke591uurMKlN7N9jbn8qmkOWm1RnJBS26wyYp6W3Sr+PUQbAOs
w6AxNe1wjpO6JZ6cZUAGCdCb/6AmgXccmAxs4FrHxMl9TZNEWmMjZpYyN2GUex8sP/fCz3LucfpC
fRG9FZ+lJ5GqXdhFG1Lh/tyi0DzzxnY8fVsHgFabVszjJz8p3lfGl6hvucV15tqiJg94UUeJcRR7
RdpoUjjrYlAtvg4IMP7A6ztWEfjcjSOi+FqCnYwozH7496o4WOvjM8f2E+Rs3rHQaYgv7+lQp0VO
kj3Y+3JrkeVmLMsBhsZqjRjgMpA7S+qOVa/1uWh/zERM8Kup2V9VuuZRNqQoEo6kUJcoKFen1fzD
2mV0HPhhDIBqXCU8XEGYHrP6zLIqzK193hXl4eLgWKk5OttTN9ZM+oyqEDJPZJ3TBQMKPX13frza
Zy77BztjpBYHwd+hmvk9S5xf2hYrKLk49q9PZ857Tg0VerpuNm+NGht2BwMohr7ZzxtAfCp4N58j
Ndqzv60bR5YGJ8N4LoS/+7tcMxjd8K0FkCoqrqE+VfvTtLbi/KX5sbbw2202P4EgHsq/+scfD9yn
J6yXO8EmtPSN9QuQ+PPdIr0QtLPQiXR/ijy8GUZVdYAN9A8Iso78BSQl+jy787tHtmokRrFyLkVs
AUx75JD4rmJi5wrl3J0gL0Z96UM/gbSRyVBqqI9Q80M+66LGFWrnO64HhTIhwqOO5/402iEKFInz
breA9qkWTxzfk8SJOVwwgOD0BrAOC28XN37c3BR9Dv/VSqCXqPviD0QOtwhRZiPhFdu+xIC7WHHK
9DHwRGTUUh0ro13+wvouifGvxF24vEbop/mMF0hoNiTKIS4UMfAtH+gSIjbriYpB0xxJuRf8dFrf
roZWLLw7U/bvBfSatcqpS4bXw8hv2iQHzUu23w/SolIvCL8rbC4/mhEoFZCwY79uTlwO4LyYDwbb
UzIvBhi7k+drP35hG2qRWlFpzXZzeUc9MABVF3517amdDXd8S7fraItVvFZ/GVInRWdFniGbZC8l
xbJnreaAY5DWppJDNtD/7q6LIPmJyRvPCkNUf+QLm+B5dU1T+TyeFLG6kWm8wSeaVrAvw9KtAPpX
2wVGKxq/Bpzl1X9K+0XsAc6kDGTbqe3IPpfuhKvPwdJ6g2wTK3f/W+c1ArnY6QWmwdKyIU5kX/Ub
A9XB9PbCpPVprbGOzmHaiRHOss9pmLFE8V/1GwyvzxIzH+nOyDQFyhgjbRskFa2QGeatK0beC/XQ
B6chAAnbt+0sr0ByOVUv4IuJ8Q+KjtPkKjoWZvSYm6j/GI+6CB6xZp/rGAknjf0+/lIkQu+qbFS+
64QBuhrl9nthrfLRXM0iSaUxWK+MRkdwIg8FRFGot9/r7ctQz9T4tz+eStO2tW9stbmRXtiRminN
G1Ov5FrXRALMzEZeiy1mN2xzRRJZztZYrKjsYkjIkT9Kkw9uDbGzsM4X5daMZJBU8UY0cJbZzBdN
7UtgNbWgfSuh7uAfUVxvfrX93I6o8VXlYW+t7Wc7+MflEGc0DcmWWHhJRqUtBG4/9pDet22gCnJs
jaX22C9MoW+N6s4oq5E+jiexJC+NnLOvpcx1LEPBZomqv2ReTmo+0i7AK8WBu2vMM7K9gndcjVXL
K2BuP57MfFBsrO7TKtCAK3HrXf2GDiygKuZTo3u7QUgCaT0tV5+zwJ5QS/nO7qpokcKADaASRyTQ
R8AHd1febjSlvzzOOOSBh59OqDJ6a0ut9jV1tPtV7EojrK34lL8ufrXdyjzr0ecDQtfy5b3colfh
8s9jh6vloInMmX7XQA3NYAsFLy4xUxsGWr4njM9SWlpfDN8PsW32DLApR+HRdYW/eigyZ3z6K3jL
TSOLEET8ARKlDTWKEgD02uXJbQVaGZNhBAipiQ0qCmeSEBA6JYafuLY5jBNicTiI2ZEiNYObf5k6
asqL3+wRjCA0DBjaPqkba+8gsDq37iOxPmd2UJ9V8lmcMC++HpyTwb4w+wlRzuKw53CalhUq2Hfv
RgxV2MqVjs1Fakq8XiGvsS7TXwqQgPiGYP61FrPA4iq7IoXS4ws7ShcOJYVYg112+B2+XucoJQ/4
eTDi1PHmMm0iG6Q6VAXZtyz7LLeQutAfcBXfQOyTfsRtWdWN7MY/ka1chHXkPaUlxWFkd9WZYrEd
/niERH4hKILKxHufFl44vIkJIl1YaYkxF0SeCWkoq8+DnpIBC7jV0sZ/g9KF8oyqQleFj2WaNu80
CFzliY1LnIeiIbWGyFwGGS1uZIQ8m1WyYdaZvefq6w9PHaqOeYCN3rWGj1Cwaty65/81foeolxHn
+9iB4n19bqr4n/ndMemm0qpGGm+0NDv7+dw2FRo1QfdTd+UffAR8CvbBphMyjNMCz+o5ipsyTRaQ
y/GDCMowL63xnMy7lx/QqH11pibEgsU6hoUrB7v+FuthnRFaqaUc8T5h9YgVX9UISzfoTtKwi4C4
gO7/YSfh06RRze/H9aFRG0L/V7i8bbNu5oksOGwr97ufBUxBlM0n2dWfBqEyVDQ4k6eJtd2s+gyd
3axp3AesekGmXacCeAA0c6dir9FXe9XPqdvYj85Xm/mFmZLoZIt6Wm6a9iTgvJ8HbmHcQjn0G6EN
bt2/ewzj5BDhIhOQSXogtzXQhzSU7yAZxsAc/vWeu3wTE/7FtwZzRq0PWVu4wrI3BvUrUDCAqrLl
LiS8RdZ1vzwPSzNtQTKJdFQ6AUr82gg8soWqobVmzoGI6i1FL60JycJo8WaDdpvn+N7bzgDmxizO
FcSgE8quJzvnBP9S1bKNP/LkSFMY1JLwCA2bTVo5jPJFChuLWRW7ffrfRWrDE5Mf+bzztnBP/OUS
h1usiiS2hUAW4iTb+cOM8vQFIOsq44cCFvSXM75T8QeeyLlED1cimmtpTFiHyPVUBqn2/sXtpeGy
9TgiBz8acrUGxRw14mORCvx6RWjJgitGJ4/UbeFp6RUbUtFrU92PvRJktTjMQH8zcNO7sgCeRI4K
3Z2TmHG+eD871qxXLYxFBYZJiak8yMG57OEfmWI3HyGqmfUutzjfasvN6ZphBDpTQvts4R4L5nr5
+XXglnz4ZM7neDzSW8VfSEEz5pkKoWncQyZUXetsL8hYVpOS8k1TORPCyHhRT8wsDiI0Q8IPHfZz
OHp1tAy/kXiHY0eGRTefbqCWbxQooKpB1mloBV7Mntd3+81DVoaAr1UttfbPSSxqPHp/quTZbQAG
8k9p2dfT2pWeAD0CTolq9tEH8/P4o7+iaY7Ut/WXCSxyjmGvBVd/q0IlKjOmvtIQgMl1RaYyOa+B
sId8msnz4585VEEO+ZqEtyL8OaJapEJobvCsZalYesbSw+BtXNL3Yz99xnDCk9hLt7dC2ybEuKCz
qqlO4bPWSN0mwEf4tjBmlvrWzuz9ny+M2qUl8vYNpVnf29HK7nGRfBUO128o8+O/cqAXXRqCZoBZ
uZEWGs+RwEkr48Plt6c5vmHBTu005ZsnReoFsXpLAwcaQTvy1U3AfvcXxUI3dY8F/5tqeocTbR2l
jCK0PTUL2K8U+/whJ2m5cPOCvVMsLSyT3sgzlIL1LqVfmlVMQik0TgyV6WGiJgGd0JDF2TYVY+QJ
RFAepao4Vzj/6ZwsRlwW53VCSLlGBrex2/bAAs8TVK4HCD7x3MnDYWthwLSJtNz6hVYRwYLBYICj
v4hk1wFzVQZ5AAuEXT/qevbmcs4A1kz0SGzrjdXb/fzEqqCk28n9RIsn7f+pTqOSmKuIWx6kDeoo
ItblbPcoPXXxicqqMvFDVxnIvUZJsTAjGDRc4e7axzhUy/yepXtupDtS9aqThPO17fez23sij5fM
I8oATtWMDsvK+Q+ixLWMBibF0dJgmyZ2MnifhTeoD64WK6IBlJ9dwTLqgDasRnngvCwfjH3/3MJ8
YbwkBerzSOKkIAdPbgW8+lGdIGNvXLknwqxZyljVDMIv8nH9BGHyUvVfFvclRrdAlckC44VV1NBJ
9S6lxk9HaQjffUQgpiQLR+7ATpOCBbOOrbG8oKiPrRynCZgQB0D/j7kpskMkaGZVfT2t49VyLWeo
JG8YoF7TwmMCdizrnAwxNuy5rZvlU0KAmVBl2lgYISE8lYNi5WxSNzP4l3BSjZNTgcp5ZIaGN4ux
Iq3g00YiFtIsfm1pCrMccx+EbhMD5itg4Vn/ZzsGnxxOLSOuwwrx1UtxAAiXbSxPhoCTF9obnMhv
cevpXs1aBtJ/iAyjnah6F0yoqGho/btr8JAjUu9anSHtgo1SNyvDBGkJbRRivuwaBsFV/m2OBp9m
Zz9MJqFhGsaTVMDLkmNgCMu6RmCpnrYdiEWsSWuopZMH3q7mR+RGFcuOoSx9aHVkYuJcyGF49JBZ
WQJmBdGRwkedDdg6ZTeZ9YXhsAa37df22ix0XqXQiU5qpdqKZZNzppuhrc4QmeYOxcZDSpL7s82o
UT4bBUd7+BT35UC+aIxTVioTu5nyuP1rRM8X3LWWI6qsXyXQsRogvGoSWMKhS0avba+wK5vCGl0Z
VQYUZVs69TcR8F/ISj3LOO3Ykjdjuo+iDZhIyJTZ/F42JJ29KSvGmAkMrS/qJFgfVSta9ZTdJzyd
iFFCqaj3F8M+gaERlkOPvw6/3OLy04qizBjFv/1A6rGO7Ad+tAmyPeZ4kw6O1eBLZAZpeQqGok3S
QmpxMO6lksL7r+rhzeA6HrkACSMoLeQfsc0l38JbmtW9t5dDJVViFXqPuL7rcjLMqARXH05X2cNq
JoKTfg8gYpRigIr6GdxO9kAeTeTARiq38ywZk6nc55U+Sa9XCe4jwstNRPyU56NiZ1I0XdI0XfSR
VrXmhRHdB0K6bWxC9TaLyFDBlnVysspLVlMRoGulslN+2sUXTzYZ5R5y4Y41nWN61N0SouEm1NfX
XDfQ0Ij08HI/+bJXXIzB8UAdVwTm/CNXAbXkweTNvxnq8QDCazHOVdmFAHwJUx6wDHiG82Vns0j/
6Yuyn3vAAdx3gFLcrNYi2C3UZ4uytzg66Kk4N8jwGir8bAr5z2KNMAS1SM++oDQBivrJlhPj9f/x
3Zav4AECLyk4QU7Oah11d5ZPphlaYOesWRBPdXPKaiY5NjtkFEBQwGu5nSpzIh5wtE6fHecSaydY
ooiEHJ+ObzRhQNUcuPOAF9D13BMLhD6go+3iP56ZAHWvhFqFh04V7MzCF95cjLudZfbAIHbu7fpB
SFMWDau7EGDu1yVUJjWeut41PtOUJoEuGuTuaRHktLEjjKCnhHG5vQmtbkM1BtKH0QhKrMOQnchC
kxNjORo3map87z1prxPMHsByHW50ZTmfHwuFq0x+051VzkJ4pmsL1IDU7ZCk3BotjMYqpl0og2Ua
rsB5iMYLApnVP1Ure6XkHtS6f+3zsLZSyCu2nA4chrBT31e8tA6C6OqwDGSTFvHJU87hmefZpnlj
CgPVHd957nUWGEsoR+67hCTS3ph0CuoqDaVd+D5KvGA5u7pllSYGIpghR98KmBg7umO/Y0Tg8AkQ
d6fBm8nXxbVfR4AaQqB8uZ6Xscq/YsKVD/4YDu/uOgUsjXMd3EmMiIsYkJJFKQXK7Hpta6pSmuVR
muwj2BUsd62bTAsnkTsb5IW4aBUmUYyO5SHyB5DvE0UdBElaWfpFoYF2y8INVW1LpJSDFaksHEBN
23x5lg/tnialkrKPwr4BemxOYqn6tYideC2ZOfYmasLk7eqheGgXR2Vjgjg+G7/kv4nSfalOetfP
gMhuhlmC+dIthxFYXffjsGaH7g7IHz3sqeEI66PX3RfjY7X9l4DULL27A134/Sgy3fnYI1H/zZGm
ZkyikuuT2YS02d/y7E/0Um4IPtawguU87kYeat0EVA6uVATjJdu/p4yyxMD0nEiXcu+abWe2qz2c
0rJEwJJIV6GqHfpBtWojLbjKTxFbasUvHZB0rc+IANcFuX+nQT998Ys54pXdj3jQYtgJIayfZLUz
u7Ow8YCqXF2SxeyBidqimfdnRjfeqwU6JyFgydAM7VkhyUvu4SrWftV6NgeVuq2nVKZ+nWycNpOW
eMcsk1eR/LyragEeGI4kvN1Xs2AWorY6FnmCM+ZP96anWfELoPz5XWxf3elYMEuOr4MX7HN7sfq2
18bd9IweX2xtUx1HJpcSndbtJCOnKryQKbICpGGBxi+83KkAt2049CSFq+CtNhll5tuxuo+Ge5OW
48Aj6HYpsEcJdw9yiEhjGvTbq7OCKBQ5yCBXfzL+zqTB4lBrycXYjgh5+mN+8qXFwlk0T+KRFh/X
36eeIXrHEZ1NEjoIcKEqT1YCc9albSAlsREKKrbiEBx44pvjPJc94DWNik8YonmEPfd/69vm1oNB
/7Ng4KDHrvvyKYnaJx/DtPCSJkoAERb5p2tqNYsceLDEngvURbM5/ye4kMZMTC5fipQynHEY7NHu
oJWX75NNNiNbWXdODbxia0tzhXD3d6Wmf+9i6DF/QDmewhQ16rxKPBfCyZH5tP/tQnK57F+9qn8h
s3QUj3DKN9BaUlWZqKsNybV4C7KtAV/mBViJzVlFCRwbW50EFrvsA9P8pQ+WUOPN3B6FAvEC5WU1
oscQATcbi+RmnLue3SzKeAPs3VBjadHwdY2uCSTXmxSlsXPD1+sybUJkLgyisAoLtsyARR4nc/xv
LzZ/71bc0VDk+1nb0gSZ2/VLtV1VBxJMSg68rN6F5awGLPIArPygoadFEFwsMes2CAh1g8XcF3cx
Bro2bNoqb6L448yyAbPzPsP8t7h9p2fu0jl19QeUuT3aaNi4CGqwRQhyofKc6NxOLMV/yRdb42pB
sEmpuWaMb4loB3f32TMmEuNpT+8hJqqvr9ZK2WezgE7wRliTeUo62j8cwGqagTyjr+O7B6VeupPc
RxrwQalkJs8nSONExnBSkiQxCJ+tMKRWvFkCxmg5yo6IF5t/YsshLcH17iXgVuTDXN9lsi33Ts+d
1nYI6EGJ0amRDZWT17lslJLNHZ+1FVVhQrADxkFt94ROfM7sXH4wjaKAdn1m1BoQKzlacnpWgJ1m
chgBNXWZY2IOm3xwThBSaDVQoBy0G12HmJfxAUMwJjwpnrQsFnbo1bH04pgjnooKcia+dNDhy+8D
z/+ucPxMMqkF/CYk5QWf0Z1vPGoz58Zfk9BPP+l21hvizF9nb+R6an25KfI0+XFRUublhhXJDaUD
UUw4TnuoRKv7MLPzY644bYt5sCfjelyjcWw/FLXk9Gqy0D1wMumJVmCR8HCRl/bjhABQT1648aLM
EvVwNakL1/GGlyid0p1W6Uyb4UDfyxnqznk+fA41wWNWlCalHnu+4uiZACjn1rev8etb3RTMlswN
Ms9arBxBuLCGnI+TCi+hl8h9kaujFAFhczwpI/GQdfkFb5MMuFEMOi3GIcj/98QUoEU5k0+odvrF
42Yz0UMNXyVB4c7xRK8Ad5pyMZtkDjU0LwcsnpUoZ3o5jPZef4jAnY4QLNszFCk965ooI1Am58LQ
fbzgewQvd2zn0I9UONi3rb/nVx84bJlALej2bAc5rHlkW58onXFlm20hWVAOe8dAxXbJbV9WYqSi
tUx3zl0Ph6M6j7Q5Z0BYspnaeIa+npQ3/14ulB9ybll1m8xtDgmICJl/rwZndPjmdbxh8ENmrBO9
sUR5lxq41T3FCQyaRarostc0AnLHlTFhhrcwRspX+bsZB13FwEEH5fHOL3ePjHaFnnD8PmF2Kbfd
nT476+hH+1fjAH1/91lSsnl1H+qZT/fJyYzEeV6bt3qB3Le6adLWE7kHZj1r2aT3GAGmgjuhcS2+
/6faEaxGpldIppdOSvT4N7otI9QAuywUAQPP7L11+KrynXNvlDuerJkdQ5HijYvkNfKoWwfXuP+I
67Oh/DxgJtlqP8BUDUCZrBeQFVBIlNAefpNE8uHyvuPGtxVJpPs9uzjdju3/YCpMH9uFRCzNQunG
vXHagRAAPrqgUdN7XUw8L8WgqwvDXxIXjg81es4IZmTAzQlXfHioCDyfQEx3Ahp88hq0Cho39MAP
KEYXARA+BOVJK9kt8axwVVb9DMgZgmQ/4Qc06NqU1XMasvZaRiXGJ5BtGOupDNwp1d4jfXpZ1y6B
Xt2bvV8O3KiF+JYZnVkBXBf4mUEjsH7Z1KN/bokc7N2aJlGpBnP/iGaCNesSvCS7FtthXYfUhaKo
rbzP1osN5LAT8lJadeWQdCubIkhQYulOvQMMsGZA9FzCYGkLuKdn4nzBE/a3Gy/6WQ831nk94QQK
3/0WXjfstL4FimjiYlKTo1QSME2BwukxqniyIWS0yfF/ecDZKdcLz+WfZDN+f1RivzeYxfwYz3gz
ilc+S+Ya49qoHSc94XPuhxUJ0EGEVQ2CuK6eR2dVqG9bE+6JdcuTbDm0N9dw8ie1YwdPJTVekk9b
MRZGkzRWyWVbDOfW+UCqwRatYQNwf+PwvUhZz+6eAJ1BBDMcRqtQvS4X370vTYxnVl2TIEHOBiPW
U2oa8XJwOkCdABgXZ/QcKpw4hh5BkD1iHTUUtPt+d9Kfi9FFTRMbC/s3Qzh2aLLTQMekHlVpBCVp
/EVtsGILHAMiGDr/E0DuoqSGPN74vK12Gh1aeop6oTX4UXLvT0/NWXNzOJf1Z6j67MD8ljMA3D2p
7sE//83Yui8+ZeWwKSXZzmHSwK1bDHd/iLEdWTa9KlRK5QVoHG1eFyICpHae+eXrjI8LS0fj34CH
9wRqea94c6JdZuoZbxo85OeuLKFrnCJlYFBFJHPmTBr6fUAKSLw/CH372I8+yanzPaD440L4j68P
SM0Cva9tcJsgD25KLQGZLV0Mc6wS6MOCSV9wePWyH5h2VGrjwtyQ3ZVwL6qn+QNCyKy94n+Oeqek
gwU8eItTytOq9Q34MobkJpAoSEEYaXCR2YDoZK+t2agh5sxZfxNYjXSfd2/R8+k8DMoxKqgok6el
bCGfI37qhq8dEYOoSoNvcJ1qwQtFoBTUEBzXXquWX7iXsA9qYuLfF58exnKXfkUie/Ljx80Ox/H8
H6Iq3Kepmfxg4T7J7Ycd8Ub0YtLDsJAPQsZKah5Wvo1T+2o7MrxyKb8EyEM1Q8vfePIa4/lqM5bG
73iEhvUuTdIYq9knAAG4PPmfYHAhY5lpplsNSC0B+qsKQ7j8MEd5rYF87q9fJ1sY9KQTVHwJXsDV
3fGqRI0Sp6NmFKF5SEnWlWGRLwSk7hXVG2xyj9/QFEVqfq5MA+VjeanoFSa/VILVTK082xcxZgbk
3sVAs/RgxGNWe7ALvOkGdYOWxjw/p80ZQeTUbKLN3nhsCyWTDQj91umJ19h5q6pEvgh9rdcirUjF
bF/6NCyGmHfqLFkZSc0RneqqARseakutBAanxrdSn41lP6+iHoLZ2z/nzUOT5T+6H9dF4vib3kpf
RPhq5dW0JgHkdsgATJk1coNJAa2IbAlUvOwHG+wHEk33H3X41bcHL4QHiXp2sJL48nQIG+r3Cy+4
3RcEpYaISCY8EqEQAqZ5jFFjpX6g6hrehtaJ4IwtLJwPeG+R9hFqrSU6SxhxWaBw7lArXY7g/mAm
tQCTJ1iJStoFaSKxX/5NpEHrOY6VaMD9wMG2aCnnOqOrXLJEUKie+P4L1hK+b3GRjA9v9PxprgH+
VI0FtLkLoXN9WsJk+VgVRWVyLK8xub/DGuOBkQyVhhvdsyD151YEXU90H03dvfJyEYqum0upxvZK
YwZ+0z/nCb8OBo8gNZhNVQ474lFGgWjP4r/h5edvhhz4BT/HtIy21OSaaWVYJWFAKcpOwd20Pg6l
sQ8euGB1nJZk6+8yOe/Ir1WXMi1u1Usn7JmwxeDIACvs9D4OvUZ5lvD64nwqvRx4tPkESwLnNFHZ
3mLGSSs7OcrPSrN4qYzmRF/Gz3ceXC1bQQaQIrWG5XFZizrbq/SwC1vMfWG10oJTGwY2x9cy+PCL
Uw00U1q9KbKguA60gLEynTYkqtGph4wouDTYbfpLlsV8x+Zk6vGt60q/KwzmXvT4du3tVoINNXa2
eylzHPvhi41T2eH8KvTIk9sUbv681YnFJHs0Ye9yzxm0ArUBFS/gp4KajjMc6ekRkzsMFvWxnNd8
7J0iDzzrgS9hbhJr2OzPCsLIzjFNUWpXbLDgaraYb21qAIkqewEgoLw3UHkUWlCepLFTJiips8Y2
yEhdXQ0/wyfEfHC2/f4sY04cM6RXQN4e/h2RgbSwKVDLxc4qlPEmQj35wwP/qW9TDprRF4R2C6ZT
bK2dkugQdHgvMUPcHHkf2Aibp7O5Yc1g+RhAbzq8ARWL78R5XXnyiT2flrJs1NL0aIBt128YsjeT
t4l9b5C6/ZC22MA5ngS+M/AvBbgmyNk8ijwuqueMniMTjP90HhwNLcCBWaD2mWBsTTB+0M90Gshh
85OSJnlROVBAIku4qvVAJDxLLI4Jw9vE155IP7TLWKEonPi3bPd12m8IlGbH83cAKCZQ82IZhyGJ
6RftE3uBQFbk+QyilA/YO7zHS9skIh29b0+fPnO1K8MUFrHB+yrBTRHB5NEHGDRafAB0gD0y8OOd
SAvTkZx4Q+/YPvLGOEfIX0lelTxQwYTmKozoQi168Bg1TcCyVcatOUcnB3vRZEe+BPzmFdbiKxT6
0KUhRzQNt6CacdMTzvunvFjcb2/a77BWqR64KBX/mUsWKIcc+dza81cIoivDncbptWM6Rj37JtlQ
vwaX99OkiWv0G4tyvHSqjM/P8uuX6IiSqoJ2Escy+qy/8OIsrkSdn4WpUUzNuha3SYNYIBDwWz/J
m3nk8bDRj1IdLkGRyRISDEmT34g14MZZZ9xEFLs59cKigLbbjGWlNW12P79brQbLu72TJ9KRKGM9
JfPNDqM9ZIO7K4/lrhEXlejJKfcO6AP2zfAUx7AE1BXYi6sXfw3AJiEQs3Y4TTo5u/4wWBxnWu4/
fZsSL2hJcpLzyTopsmQ62QQarDKQcG+C+z4VY0wqCNkPyuxC95GYTFbX0ohPwhBQfEQfaWu1AWnn
fkfOE3S6r0UaDQLFG/dDhlJY/c9bwTadXv9ccWD3ym7ZeM7B2HR/sbhEssVA9rZkGqqj31JtXxiN
NNWv0AAqF7SS4/0KtRoOnT9FmWcSLeP+ns/l1pjc8z9ZlzBGXrYdsk2OEZSsre9fdlTaruVGeoi2
RtOf6jxsDReONEDPvLam9Ztxpu3+CX5mi4EvoxSIcXKAsym+297zXK/5aWsLxfuNSPrgcqT5vNoP
AkV8zjmY4atQlNaEmxFcGUeyEyN9TZQSaDKvLfVn24L6as5VBrysqX36Jee7f8dR/vyb6J67XMHN
+bRZ36q5Fzq8AqTx8sTwPF2lXPJC9AFARfvBtx0e9jIL1JSnTaZYagUnN+sRE41EZIl9DFIsgh8y
Uo1d95LkRXjKKMHKbD8Hg536xHd/Gbl8Y7ML8cAv390ccHHYz1IHcsiITfYFfCTylTwAcx2C4u8X
lRqC6PMfE5fu7zTCAQl4jq97e/vNBBXi4Kf6xPu1ops/B2Q/cZiO7FipRhHYokisma8iqWtJlSNm
p9mTmxp/MFKqM8ararwPHc2hlRf3De2NrRFMFIikB8fzhruXHZCeUz0zuXuxWpOSNdc9/FEE59Na
h1FDlc8L/lRvB2Qp4Bv64d7+YSGWt+wpdED8HGQgZrUVaL4mFArwEWNydUuVsLDsqQCszwBUL6u5
XlpNz2qBPYernBeoM9KtrqlyTRUM3rHRgndUpyS6wvKV5/OLs3Qn7PRBNs69OdaCgnTKr+rjo1Vx
6vb37VnyWN5rqKXmkGiKubjcvztvWTZrh4OnQ1cabLSFPm602g+6PgG5Tq0ZrJFZwU9wudczXu1B
wWm2spkU+6GO2VFfU0eD4s88pWalD2SyhroXcvLc2a9u1sQZgVeE61op/gLEz1J4oRGZj/QuAhyP
+sUzWinGAkIAYpeomyhjL9UayqTC9mzF56Ow0KvQ2zyzR2yfFs7r0pdPlz/7KW57U+E65mponm5G
PHGJKzEe5Tl4h9X5lyIO9mS9QcMU4QJ1U/4SYchURMvgd1h9PQ/lKS4iNzB6HxcynuNWLn2dgY6g
hY3Pzhr3ZB/FH1Yl73NuUacshmaIDFldVk1d1oVMAXzobR79XiKvH9hv95Rn4KcaQgOvu1z6dGKz
V1erXZDxZcelD8hTshERN8+GZuL4QhU3VK2cWrIfFcChdx0/Kx5aCcjIRXI6p0OponS/dCkz6Va2
w0rGQdSleHybDNh6c4GDk/r/aUvghcyV1BR/hJPsz5nSipAw7Zs6gVkIhsPW6tT1P+rpCUwEtvfL
Al6ZSxwe8tWVD52MFa5y8r3ijBDX1LaxhkhA0GJytuV9tk1wVQKVnV2I/qzobMVmiw7a+do0FPw/
VE2tU/9TKrDlJb2HVyVLWnvvqbIkiPP06VuK520NZybe7eT+qoljVgvayI1joQ23yApnVrxaUFLP
Wc2jW6Ca4sqTMEJ07fw/ep56qEV4WGID7GfbrqqwHFXjBR1YBpPWQxLrrHvLJuZDp2xo08t8shJa
9VShrllJ0S671RGPH3bgjT6oHQ5U7l6TkZPlgOqCsH+QlHmpM+okLGTp0OapwdojPC0Ppb3CnTKC
fFj6lAeYMk4r4b5N8fGsJvJ8+Ok6CeTQ89tsEym94EAiVV7wFVJoju0Gx8rBAqHutJbhhh1BKDTg
wSL+D6i1jZpKEVbSN1oK7RROAXyU/8japWpaWO05kA1QM+6r6Mlf1yAmfcdwEr1YsxwARusAeWDP
WRC91q5DnnkKNqsG7fQkARXMDBfNoAyH5yzZzh0HCUsosPAgrsCm2OiUomV7NIbj9anSNr1EdFUw
1ReLZrMKJR05w/XnJ9z64uhL1Gy4mQJnPMzbibKvU0la6sO1dfYX3SxWg9eW+YmqcydcMiLfZTpu
QwcETzunChVO3F6jyOpuqvPezE16nA+pG8sXQd5gkqIigA/Y9hTuaHXhlspuwVZRPihccM5DYXVS
YoI8MrmM1f4WdNWmvs9KZkvyryvr3L2egEPCuYMeH93xpshUX8aeL1PgCU5epsJccLv8KIVa0oLx
P09qvjhACLEq/GyySvTZhCKNjU+EXWtxfiBOvATxlshwO1EGqNeWeY8cVWWot1xf7/ps0/0LCIcS
h6C0uOO1f3+gG2a/YeGlR7P7k3DmAqbXuXV7IqUzYZV2kmQHzuM5VJFp5WPPRsxw7Hp9NQbquJif
/GjlyPqK6UopAnMgWyN4S1yECY+6hDRjRtPCCZyEgnju2kX9VlwIn7J7q+rLCVb2RSizlS/ACdtv
qppSWaBYvcN2R65FDdAM4QM0uRTk37TRVssw3e4xKUVT8AKhdI6+hQ1cRAQYh2f3HMRM6CSRK/zR
zHngBWLbCIwBu5vUTPyOMU7DE99PPQLM51Hie+GXqiPjPw6UVHI3cgpKY32sJQiTjhuuH+Mz1SzG
1+VYXS309k1BA7Z/UCUffCdwh1wuvWMNlvDcirI7fOnSSbadWiKnd4rBqosDrXgdbsLgpd23w3oV
bztf/mpSdv45eY0yCL9e3CxEbcMnI+T8dQAowF46O20U4krkEqUkafdvPBIvSLLKyYgI/Eb7QdOH
3OWiPchxKSwmjForfOIIQaf81Z2nLsinK8SF+c2c6Nmrfih0r+A3rGZrWLnmKBydOngq2f3r1eLb
+yhth43vsU7JnNW0mZSao3qu4S7KO8QzYIsX6y9zpejFrFUgcsKWt3BJhj+UT+rdXTL9tXUD86t8
PPZ0pxu4XOMZNzG195eeB2rNvjTK79A9iejg7hc+/wK2DstcjjQam7fFqhUgIIOIpBkwtGgs2/ah
WthHLRLxmW1DKbcM8Zkq9rV1uvWRtlb1Qnr7JA25oK9exl23oaaAlrwD0rJGnxRSlgFdCjmGKB/H
+4BMKSl8GUVjJ1kZjbFLKVWgH868n5GCY354ax19LnyDAH6N8Pn0rgkMbaK8YLWeFrw8iP7roe8R
8bzKOiXC8XN/8R/PFvZyjw0miVU6OEya2elhkU2Qg75PnjLsuOMqQfhTt6YzSkfOwZ181PGPeV7s
lmhW8m63fMOEV41giaJ+lNdP8tajXvn2rU1Beqkc4A0He/9IWlqtRA6IC3/t2VlpckmS5fW0cSd5
cvTuW2fo0tzerJL4U+VRj4kqsi4OkP3+w83AKoBNbLTmB2DmSv2B5CVv5uM9D6SnGPquNc+MDw60
JPIkEapSCpMuudph200OcRlERKhY3TNH2fsLWiqOKeo8WKg35eIQE+kl9xJnPU49ajYQS+syvgKY
1ytKIqHNhQdL7TJT5W5+vANeAufqjm/bhxE/FjCMFqVR0E2NF1CEytS0avody7T6kR0evGbxXA/e
uNIzLziW0UalTDleS3FpMnN8dQeERd9qfHSchdiP0h09N0tlSDGJkby3+qhBRadrkesPKnVA1Gyx
DeiEHx2a3Noyt7mkZIcHRKzNDEz3bHxO729H8376K1fJAdlAJ0Ka22xPZZk2qtKCJ26zHVTyrT9+
gfYTE99eQze4P42v7fZRS0yMDoX3bVwuRIT1qH5oAj2mHkXHjD4crDHWtSqQJPqKQmrGNFffYgI7
Mn5vxQDebGyDmAUiG74QOO5rHjF4pcUIQo68k6kCo5GCyyDhAZTpyLM/wwc2WBrUC7+A8XGuDehu
z2k1wvkcik6HSzoo5QoHe8RCFVdxsg2eOybi6rIQHWx6rgixBKiu4jUSz+n2WvuxTE07y+MQ6dc5
tI2Il9J3yTGLZMAYXGJpXls2pNjG1qHuWaq8aNFxJfjRtTlfLhBMet9D+sS3Vj9auKAjdT12+hIp
uhI8ftWwF44GQA+WHr2eQMMZriwQUuMNLYR8+cRwW18Qs2CSPQsDvGWWZlUqN+fIy1ml49QL3GFw
ik60lI62cqJKWwA9mcGwP1BTYg3MtQR3kgrnmk6zYRtk2vTfNExXefCQoHQGZxE4xMpDDfoAdiew
2onplP7ypl4m4rKGRmcdEc+ukaCtk5fevnWdkEPVg1aQWlWNyjsJuHHZ5SSdaUYlV5nqSMHM+YHY
54ncF31WfK8V+gzXOfdNVGbjMZvsSEn++CufvZL2wZ+nQVtC0k413au0OuBGvJcufz9wWXLCPPxr
RwJjLtXgW29sta1Kt8iqoOfgkMYunjzZtQdjpkLuEwvV7xX70rpJN4RdyYNOuUmzQ2VZbQhOr548
8/XBBLmb9GYQICNJoPeyxOjpa3Y0G8uS5fQtTvfbe56FgWC2+4LZfWdzBrdCl720PNt+sK7mJlwu
h2DaGEFNLqMl+8Qnbp6AAEOZaBP/Bfh4R2YQFXSQ9bxD3vi1TvHdZrto5UNZBtM64qHNCiDdel3k
4742Rdk8/EBJME2qzgebG+G12aEF+kXSLd4AsCzYqCu1KBetoctCBS3jUGT7G+TQhW4d2TSyTfRd
zCmXO93dEdo/YwIxNor6FKEva3D6fpVwRJL5RXMklcCfBEYGyQdqwuNN0P2BJwaeBBkImIoXds49
7Xv5q8unnRIO2EqEec0++yKtxKSUMVhr1ctvgNw6raS335TEfU3UnfFwZWCC3vG/VnduD0VGt0tE
WoOuTM5knZ/9dxW85a//+TW1GmJZLNhL8W+lHxC9isjraNcq3KPQY6ufeBeKLeiOjYt72eud+d5g
c2czPZ1jk13h7Vo5RkoRzbohKjkrF1sl1DKwATIBAidUbCrsdqrhqvmizNQFUk3dZeGW6kcVjKiz
EPeqwWciInSYUH1IIz+mjPjPfK1eMruEo7IYXwojCOXR34dwenN9vVhdC91bTmKehcYzFA//6loR
aXptfeeekdy/MUcXVi4lsY3doToU+ybJKmVaBFbOZs57xPPNAa23o2hbqqcBs7udbCaDL7mbzjVL
MIcfHri6w6KfiztHYVXj/2DcLD09WHqOVkBFUe27cLPTMJjj5gI9KwcroTsRL7ylAJu2EinHkhfu
DzWPdXCB7PeMdvDbBf9VLsnyqkKSDEjL2GlExqKucQe078ckeWrdABO9uykbveMNiu/nK5XZ4ws2
jYS82Pm5HZzpVheKHzmz9a8eHfemxojAyHXBXRYNy1FqgH0K1W30g5mkdLYBA7VgLcV7IyfHzgdK
n+KmRGtDVWrAGkfVHLwSL2HBhxKFFp3PVVQNftklREH+oc0xEYk68l/2KG3emy8Y8LUTLC5pEAse
Z6oLnzAbQgmxIBYyOs3YnjZZzpXa/86qFj7kMrWdFZkhFH4VG5MdMxL1Se7TlslCGWv0jPm+aIdn
9375VcbbuCSBKUosc7jqJw0etC6SyP6L4p/YDWoDZVQtU0wVRc3FiaFfS1d5xYbQW0t9lUspDd/A
1ei5VT+2pUDU9AXzMMft1xyY6jPLaVrdtveaGrvGCKhfzN4UlMgjFeTcxBsVlqG3ECLIAlIN2/Y6
JULcqDZ/H/iZOO+wXb6rQOePB3tp/fOFZiBEyhT0biDBv2uX139Qq0zTICyNRo8u4JuEjbEjuAtf
NL7hDUHLNcOq3h9FvJrsse6CXlHhy50qTVnjJ4WpuS9rG/1T5tgYNCAZnT+JbMy/gt+aqY9yYmKt
mCz8gAgq7nroql7QvDJthMtqkBCx4M3SQxr+/55Ls/zBZXA9pHLWlee+wmoCR9OXzYUqA7y8lbkY
ixuoL9FnpGFGZpe5/d0IFbbM0kpDf/xR3/FRVT3qFqgYgWnTyvKhQkTiNokvmxo+OC9j5LIZ5KJH
MIV/l9MxeUtD1KatiV9vQmZcfo6/+QBka1H0OJ4uX7rzn94+lLnpG9/NvQ6+hH1axiqD9M77/5LG
SdOKDvs7NHRAnXhnXokm1VoIFLw7XnYzKkfciPXrkxuruR1QVCKB2pqXZljcaCoxPoFVAIKVgOMs
olFbx165n+Dch0elRvOo+d/XwAnbjIcdVYkPEflp9cooP8ug/9OXGdrdfDr7DxmZkfEYlLef+cKt
sH+sekk2tyEa3Mj8Te51Cy3LeluJHHVJb2gvQnmqXqYCsl4I3Hki4NI8/x2kJO717L7yGRT9115i
j1kwOZW407IkyIGSPayHPmAGihbCQMz9e9BSOAzoWp1sp7PAPIki8dKv1SRJIdqS+OquNJ/ID/ir
YcL8hQPwdifEFLYRxnlWBgqrxvT1uyb+US3VGMa8rGoeSY9Tnz7neZxogJ3zwbT5BFtJV0HyShTH
TgmrP04+lIbwxnl4kHkASUJUmC81eWKksBFJ+mvNXuavrIbbDtIhIeMYnd94ZQ7f6EvNsSnqmGIT
VEe/PPZgJlw0HLG/371yB58OxZxv4UVZEWL74rr9VjbjqJufi+ND5EhnFCnVpk3/X15CihDcKppP
q5IfBgg5T46jVv+GHcYdTBZK6e5UUEgA+w2Ce/5uE6YE8j6vxFenviwqwByZh2iNMhzhPzGXMGHm
pohNNg+7yzXkajhdsxWim4TJYcLmMpFE1zwZ5OLwn3Aut3uZQG8cOFx05/KOnXoT5GpVdWkJxvvb
U3gfG8t8Ps4X+040OQEkflVBZk0+oZzWvxgeBpsF7k7d14Jgho8Lwk4YdR4ErU8++bU1KO6Tsfsv
YYKWMwQv2UZy6G/VBKu7JoI548Kt7KfJGhFGWPj3MGpMTiaQgZJGsHchnNR9x4FSpDLNUHm2hV6f
NRrPWmdh8DdWGp7olWy62dB5q/aAkI2vuKI6KKNKljsa0ZtZhecaUva5yoZNDHfNd19R5hpNmJDW
Q0RnVNWObS9qMM8frnWlmZPV7jQUKDQ4GS73XrY0pF0nqWOAGOwbkpol9aG4lEZvowAPXBkHvF/w
E1cKEB/N866IzkpCyUk2P5TmgL/13RlU1z6soGKB3mEqtatQt9nok5xrvfwmCWTk/gKhNiLt3M3K
XFLFHNdQHWNWQDNbMfM5081NESLLBnmwjTJb+RVViYv9WQInO4EB/gYEqAVhwtEC6au9mwS3WO/x
C//B/NG+dlB0j9OBJW/64wQGqCqAXkeY7UxObc4uWNXUcWrUk+/VyP5Vl9oxooRQ+UCUZFLA1BcF
g4eqfmGYl3mq2qolMskt8+M17dFJeMejin3HYH5SxcjRtS8vASyWW8JDwjzzCrSNHwE5Qh0Ej+Fy
QTLZR2+cwolfT8e7S52+Sc6OXsrDnBPft+y9rwzqxQb6vx1NvEGdwPvN8rzcd9PMhyViFElrZDQi
Bbi81xD3D2IpQbFtMIfahQGK/IovAn5kJSU53ZKlwiKsTYrLgtgaWustJmZAXm6Xd8OVC+VFAJ7L
hKNIdNN0D7WfhPjge3NiPI8eH+tkPjb5sjqrq2H88EKMa4gXNdSL5XB7z2HBtpbo5OggKbACRjNE
JEqgLrZW5K2WGlo6kzqQMLTBlidDEgZ2G8Ukqvvrs/arInvRbDaQCSKGJ7oMPE9Hijt9spNkqeuS
J4p0KQcy6zp8BSEJjaJwAMlx8a3zKsdePnCPsvR1+iwyeNyL0OTtZEDBS24odhXVztlwugEKAMHD
zouN9nU4Jyp5CbkKJddTqsEu91yHP/70QjBGUIgoAxsda5iIrQapJ8j//IhW/sAiX/iQxZfnm26P
a72paw2Ik+5ke0r2p/h5668wdu/S7e+BFyjTocdn4Dq+icwF+ixgP+LfNp7fl1yRIhpyJU5z4VcC
lVJu/IXYaQx7fBalihPal/0Vv7l/Xza4VplivbmRnGELcYTmZS4mU9IB3Ql3cSinX31f7lCbRidH
kICwIMR38QiC9/ZiblgJP21WwfUSMBXImTEtB5iTRjvP3mSlGYKm6PDj2LKAyL4O3rfIDoy+IS+i
Rpu25xFr2e86wQxLvKJp1RkcNv0Ab1ngh1XrUgOBRGKV+rGSS5kLarSTPYyrzI6CwfgdtGZr89gS
ZJdYd/t+Tu9agdOo51thEZ5vz3q80p6tQA5CkTRuLwKIgsw0IeGCDLO0759oYDWg86EvSe3eds6C
/LNXtKQKIHPBmBZKfGPdYwEsopc/sG3X12VoiKHJ+ZXFB14B1iJO2lXf2FjQCGBPgIImwexpotY4
YugDL2CXb+q0Obyag2j4Pkwz7vGUJDW6lDx2Atn+WOrZsbQXZLeJe8pp7iLatmJ+wInxWjjQcS6L
OCvQqW51MOOhSRNKFqhmu1anyv2Z1CyNIrTv5yV3j+fVqCANplM7sOcxJDRMoJBRgP8x5IDo+LA1
RdlNJGT0X2Gj9wP4LJLLFjUmXdoThhPy3/8eY7kcZW7XY4Trk5nfgYaIHaiWhkbXNHOCSyDw0Jtl
1Ekc3PT293lDnbRwuJcMhhjsYipv0+fJBQtiAlxDjQ9LWWreS+aid5oS3vwjUcBIEej5G1OXXsb7
V/yCnOhuPe3ooArXe9RVKWqnkZ2F84f8DX2LXc3WzER3WqLEYdCupUwCbXOnB78XSI52wehgnVEA
e1GBv1nffPySBsU2nqkfp4V0M0KkTSIDDKswcG1XKcOjetAUZmuExruylBIcPxriPg9hlFDxZZbt
GkiZ6Fvu0Bg9PvzINCpOvyOmLXVdt8Xd9I8em6voclEIXQIvp1+ezyB3BaKo3HC+t6bCDxD9xkms
9Gx62KNSElXwOyL4loJzMWb3xgAJ4TgqXiRgPveWRfoiQrd82LCtpqZ5+qrC2kFUU3xRu/dQ76Tk
6fPNkZ6Ufzc51JFcdMv6zTenk91t/wRPUQb1oXKvQJl+E8gFTtxwuggNxgLTDIuhjgx3An24fpO8
W25JJ/q6ogAEO8m7CCnMTwdJyLU/v/PesZK0R8y/DoaEtroq/xIW7Uz3DAJC0x61g8zGkpzx/sOQ
LXW1703cPSZEj9xqKs1un7tPdTdy39S0VFMFU0uIFTLFoKkk1wxedno2scs9egQulyTbNynq/ZBU
9OxPBy9u9Sex4GwV/+snvj1l75CFKjS6rK9y+qwHjJWZrVkwQ9Vy9ppHnTspFa7crFCIJV5E5h/Y
16Q/LRWNm49hiOvoqEWe+Go3CwZ718mb59skVrv9WyxZfCgf8EzXk5ZB1ng/7sWhI3bXdagvch+7
PtG/e2XbKmKuzs3T18sT1kYoLsKga53Czi1QmJoX9MZWRuSnslAOCriHyKz53eQLFTzKXX5+O6IP
shGoRvDknBB1GCiXN+/OCNEw2KrmwGnfWLLbX7DIRArM+NtKgpne1+EAyqKUBzxM0hYds+IFroEm
e3WXYwBkXJKw1XHO9TBeEMYi3QyAdDPTmDFaHDtGXfKyQUEIEW0AV5FOVY+5/5fio7Qm7cYwbUUN
1ouTvObatQ6+mUSmLj4ubyCDk0rXzhvrlCGUgR9TBrYEPVdwo50/Z28q3iAwQ/JWIBWGedUvy2ib
0akdm/c2zki7qGBsyNijKt0rlHd7v7eM1OhnUtsgS2sUGMyWBKyNgPDEAVZ/Kjhdb1Q0w2Jsr/hE
yAfoT7CVLcliafhMPseK0cAky7ziArWIRRA8Qo7jsDqA7nkv/62tnGL3fpm2jRovOHPptmuoniEq
7iM6fZHqpv9BpMLz1jhna77p0hIWxaZAUNXrJsVOUlzHJVe/rY1VawsSWaqhtAMYEOIUpEP2nxTh
imSvPwjsBqB4kiAjX6UNTI0TNnVETSlea99WtCzEhyfU7WLa+nUZPDUdVKKaktW41UgyVlBTRfEm
mDhr8s2yK7W2rkB7+80363px15qeU40oP4q6UOUHB5ukuT++AN8+NlZWZgj1Dq1tKb/uSf9h811h
T9sbJAzq6zkHG/13m2vrGs7Ol1LNA6n1uwU12n0eU/e8M/rYGCCVdmPa6aVzFUhcu5Y8rKZUW8Mw
f4W+cQ5huCG5aey8AT7wLVqqWjEmJeejmo/+Tq4RXABZCIOYjguqYHuljaqkbHDgG0IMhojgg9X1
mnhKFX2luBF5zTFJ8GvPbpuhR6cRXYuf36ZUJQAzPv6OHiFXHdxgLe/kM592ROx6643S1Y7ZQz6q
uT1FAUR0E2IEcNnHT/wl0dGQ0rBkyvGHgVPaXWrWcHTSS9QVQz/B5Uf3YrbDGs7WxI/ek4OCC4Lq
SkxKvvDmNec7z2RhSAQ4ASjYuVwlt0CKbl5m6Il4cjQmkNDtBdDrPbiMCeToG53YOdcpfydrhnVn
LgLMweUcmCFpIVS+c0osP9D3tMXH2zLW0mXyvpLqR+EgKAsW2kmNe5w/+JWBmcZLexFQgZ9jZboP
1KUyEumnC9S1GeAOvp5ssEEeuUMr/sk3P2WSpKpYlv8220HDBRf2pRv3ajIOp05FiP6K3LZBDdYi
2x/mrA0E5jWI8sKu5oheKM9ATlLdM25bjDM5eWqBecl7bfJE9toTGLs2RWU1GU8AXP1WbcL2Pmdw
Qz1py+wWH606qN4F2cs8aNsUERahrxDgndidGUjxXd7Do2MMeXHN0E8+XTEAa/PqTzmiXVuLSa6X
I5i3nNpC+eQpK0lLCed9IXOvCgKLVA2itqmx3gMSE5mIFbGTWjA2T2e9doPSXo8YZDnJuqQN2vtC
lDiqCbnQtFszpHlcG/P6PTO5XN358cw20kv6bcb+a1JdLtq7Hd4jjJi0eWi+JMoazv+KkaDH8vk/
6tjpqHSLixHpHpp8mnl17UwNXEj2h8AltzkoHbSQScbKEdlRHBLRsk+rdezCSg2PtKITodgB6IYd
GPSJv6MZed0QTOo1167jpJPnb8D4LD8O9xIo6AjXPnDvnqwNA7TCH54KxyE+celUWbCE2JkfHVN+
pgVDkrrfKhbtXdi+5L7goOWRiPaqx/b1srjVxE8fyKTEEvLK3xwxFynR6Vg6LJIw4NUGqnXT+6SR
2r5kuIf8qfr/TpurLcHPqeDjQN1slVg50AjAXiJ1h+5DaiKGbOQ/JaJ99JV9pDOpOt0z9IGoDMk7
0oN7vhJMGqYrms5a31v1vrU75iXNPpDHFOYpPDa5LnBB0vYeRUCRDMRBwdLX0h+pE/8okdBL0uw2
Oi1UqjH2cyDbMMbiGSVjfC1U2fGsYE2Z9cbV8a3oqCWX3SkV4f463MRpC/S1m5yVcWrIq9q64jRG
huCTe4sSsrfHJTHCve/Vo5qBzS3b/Vr5avZmILI+kL81YjpWCEdlyFBSdGUtVf1XUSZE3KhjMbC3
RHUSx7sle5oaPFgZVzvVmn8CRqW65cTWOfIpTI/Vdlb+uTMtggFB8ScAvvZM1NLW1yaPSympVKKI
st6MxrLP59Tu6gHuqpsMAsh1DaeojPDA3VoV0VND/3g9odTmcKRjXSLEf0IROI3wK8pqAonUkuS1
fhV2hEQ4/mNN7GMxxgnBreCJxctwPpSGuCAhoTM+nOsUfBu7zmcz8J8AoePvhihDPQJunPt5UVL4
VfrDby60DcaF4HzDcl1aXwYDrUT5fExJhzZrxWeEbKhnn0nkaIfGFOoMOx6oiD2q3xesRpevBa7e
VDX1uN/BwET/WJgncg6NZTsIWuWLRIpF8wIQgxSuVutzwQ+UxM2NeK3wXkfEAHxoU/trwtykPVgx
S1Dm78PFCVtfB52YCHIDGVDlszuM8zSAPSnJypP6M9oKptb1vJ0efN5CUv/G0pIRaE7FaFm6hojN
H24iHsOQo3kA9/kD7jABXG/LMEtPax02NZh0PonYfq0RwnrBlziHxazJAjyQ4DF6EiXvs+cPQHje
jole+n4lRbiv4ZkCmNpK6S5Zc1uB2uBu46uyyBC0WaszqBM1lXg0lAi5KgQoi0h6BInWaT+7Z/52
4D4/10/ypXxw06EgkB/6rgs29ehp8uPz3XHaqsn43cu+/Rw52xxJVAadgrnY/5o78d+FLQRd4l61
fkMMQOLGedOAHHhX5/KConpM4JVobVZU9hLKK0d/89ZWh1zombWggQX6S8Qhau1kVDtVhxfQwTE9
ui/fm3Nf/eOBTQWLZ6xp4meysiRl9j6LQwcZMIfLjjHFaBg/Yk/zSYzW6uH37VEqmhisDZ6D30nf
LFWEd7RDOkTHA9ifQ9N0O+xsIO1gUo5EoypuLUAu24yTgx0Rl1eR4MnnEcFess7XOG2Ccn/r8QQw
VV0c5VAFpGMHMnSG9+1IRpoq40wO4HXbQmRIFwEpH8ECvcWh+julBt352v46ClwLp+nInlHXbKQd
b6ucutPE059+LY9EmkGoBh1cQfpsA55pzNFAicupF6na+QLEjv6XRKcqI5Us2ADY/7QeCK7pbw0A
xs5IxDNXdj2rfm0+VdZGlfPSaXeJw9jC4ZQKjk17RyVEQ1hOYYzdQ9NTSlqwm68Anb0ffYUzJOTO
xgSwlOA1i+84rLBjmLVGtyGMXRKodyItIMlRp/xQh7ubfTBYAevRNbq1Q0p114VdicLAFTSWfrPq
cdZg3dFGWY0aN2mudcjPJ0L32ERwoJN4Fr49DgUGApjRrmkljCjNhWtX0XaYR6dERNvZVslnzZEo
rZyseQaZEa4Kviwfx3ArmkpoKsm5lRTkl41AfYKfRQTrcH2FG83P0WJd0PCEkpw+bOBEuWEhqZK9
C2xCDlxrpjETQWFmeaDweNr09BYOoLrT4Z1+hDV+fLY51nV4YjF1iwmgWaXEiTFGu44p9IdzRnbK
H/TQNtFC1YKOk2sYbSK31BQEb75OhgAlbTSAKyQuaoWe+ggEzF3Mp6UFs6f7/fkjGPhlzF2P/ahO
AWKam9uD7YQ206sTLVXGahBpyXoNID4q3x4tjnCBy7AwLXtuaj4HYvXxVlCHH8DaR9TZf8HBpr0L
dWxVZxdW1i/UnvrhxMc9GMgTHutf71AX061t5ZxJ7KIMNy/y4RZpBp5Dh/Nl11fifm0USLbM7748
b9+tGjWz3LKYASQsd8cF9ZZtL2yri7n4zqjqrQqAcfwgtE92ivLA1oszVn5C82hqJzNOl9yMlaDu
Cbjyq5QdT9yax4GcpNkims+2C8UfGEDdME9Kh7kxcdWKvVUmLpzOkN65g5QUqyA4fHqnVkrtmlkm
T4gh7Nz7KOAzanCBJcYszsTpgXCuwnxSMJCQSx8oAhqS/GYdZ+t9+3cS/IEbkQMZc2xUa3gg7CXb
YY1FatVvCiGgqtVMBlL2erA2yV/6u/KGc4B4F+1mUTdNoGd86cxrjbVX+RVWTY/y3J9pf0nzBR82
hvzq/9aDrH2J651NgnRvxzdDrYVO6zV1iBomo50DkrGvHqDQUPVVofuUk8JJKTgkk4Oy+pTx7OTd
j0Mrq3ppcp7jL2YEP73hWluPfKDkDae+WE/rkeOxirCPQYDw21eEOSLyr+tB6qLQ8QAnqnyNdb0L
8nNI+3B07JTjscfFXEJS5ooSJqpPmvCBrBRGjuq0Yg4Sm5pvFUJ1G+zSpKcjp2eTADuC6ydRoJ/G
c7gYxdAwrEKD27m/T3ZNwqTuznE2wFnl3vJEs41wS3pNoJTvm/omd3n8KupJNN1AdBAydZ2kjdQ+
HUhrLKTBHR0LI6u7h8UNOMDHcmE9vnVdfLtK1LypNL1OJQzuvc/s1iiYjZuQrKoNJyCLVLD3olcr
xhWd72EEsn3CQ39BIZO+xYRqgmN5r9tT7iFlVTVfpPx+/1YPCvmSUY3ZeSKWDc5OPiq0UFjxFylq
B5coU8A+Nq682KvzcMoXCZ7qeeliMRBmYgqBZUqsT9gPUUvWmfKPXNulJjSdTbSMmwdtUtNyEViD
A9yy/xRQP4NrDXWeknptIJCqdW6+cFRMMRtuKjuF5DWsvCOWkCSkEdlLtvK1lBlLgM+PQSjJpsJZ
qEITHVSBZSqYI6rM/HPwnY9oULN+Vivc1bGyoFCPHV0/igY62/xMAf0E5HIsQ26qNJOsfhOoYG4x
6wbVE3JpWzhpIa7mKajPRsaq2y+klkwXt4DvZvJsRVlo88d8/lXGgJHdbFVggb767rzWoaF4bgR5
NkLVr98+h544FclYvMJ24v2XE2AowouK5EawlSQ5sLlxTRj7bNwXG0L3G3IHqskpddA+Ix/8Pvve
zlJ3eFDuy5l9yLpGw5BRZjQF1SAaaf7JIvkdCKrcK+m8txKPZrIwoRnwT1vobuFntpnpZc3+h+2B
xD+G4IV2R/b2zyvFEvGoQxSwFd+ux638UqDnuWC+LFvOaQY1wHMH6VkEcx9OKQjHlXEBBvY+8Sk5
Eh5vZuJ7yQ62q6KmdPrt5KEqvOcOoWeOSMSMVs0HjHoCcth8C0YvaO328FuqvsrZr6akPYlsLO/y
+7tlZTyOg7OSf1146w0U6qIBKJyIcFrvmVZI0J8xa4nustYy+1py2cYBtHW5iKSlOrogeiIYr3u7
FoaeVYfRSW7gNzbwMZB6Z0vaz7PIRupcSqFKFuW1YwhRGeV0245q6x/AnvdtLzmfnwgjA75UgDsv
xXbRrkp3iIeeFHDksJeUGwOL22yzxcJwYEk9urnw+NJLkyVp4H6U1jfkSIASsSNXgf1qxNL7fOKY
DECEJd5S/0O7WTS0DFBPB8TEAuGbA/ezG+IPOtGi8+Mf3nA2+6Gqn0xmiqEVgAENOQW8MOrBUtU8
7ht0M0WyaWf+6KdZzNqLTYiR2qPnL287TgAUc/aJAsl1GBF5T8OYQke3m9wQj+hGxlftg0p546uh
EQEOkULOAKX17izDXgQ32mYD31sQRiJMnjaM8DddOfLI9kWLuq4KsZU9Q8BzVd1zMq3qcqe4i1Om
vjxlRdHwedsV89VWGNwQlYJrgtDzT6ZLCddd3a0mIPWcpAS6fISW5cRhSUYnEdFQkYAdzH27fn5v
Pt3KnBdORLB7yvgpSs9Kt5fAy/hd4aHC/5yST30YYZJ4VaxCFYvCaj7mdIosVdtQyVxPmEkDSF9M
TS9PlEgeJsOi/H5JybVn8wNJiUFP+EgiRJUk5nXmVaqxFFHankjcH1NH5C8mtHUyaghpWaFivRiD
tDKjUoaRigh99+eRUNTq7I/VyJHVXiUbTJ4DKJsOvXpY5XH1iKx1m5XKuL+cPAYVGlqoMAkJvHUw
/6dVeXBjPpJumF9CqAm+hJrpN1/qf6eaypKZkNZ08MP1wJsAXjyh1+lbzbt16OEeN2XTHMbrR+CO
uKIlSpalknDyGcj/14sqbNL9Z7ippNfPBE74Mx3xw+C7XK/J0TXnbY5CSq/QRR9RYn0NwSallqct
TMm2MURVQL4/Zdthm2Jixkd/QeJbUG6h5k3Xudf7MPzlVw+t+/3z8JV7yqosZ8nWn0qtJDRKnN3C
0tp72L0tvYAvXpECXa9LZdAAgOC8KpD5K0DYcPMlINuids5uxrwWKdxd0fyu+w44iULSxB80yWXg
kXamJM7J+36hHUUtVQwejDk2pKWyAAQyAzMZWPhejKPIbWccOO7EuJ5DSzMOZIL56nNc1IZuBJZb
DnqJS6XGAEw5tREaAaBN8iF0dj2ZUAFwe2HcRGR4M/ojgBiWJK/7sMe/L4znWapXJ/w5z8b44EfF
4864thDItzLAZaIUNoBJmYQAfSCEbqtF0s/SWXfCsiOZQMqu90oJiE0e2PBtpedbY9T2Uh8Nhf96
kVbnS+vTK90BWcwGJBLTZke1njLZhare+/liW8hWF+1Pcv2fk/wyi7Yjwi2OjeWmrEF4Y00ikrjX
VJkePZ5b88aaRgt14PXhEHB6uq4CA5Z7ASp3DsM6KtHzSa62nXy0gcxPx7W2sqLMDo43XzUOQv6z
x/++p48ipgfA/EWUEPLFO5VlNNPAs3f8VNekFXAstu0utZvXPUH6qHDs8bsCDsIZLlFeuA9wCsID
FR5Q8XCTVXsL1U4gCVoXotnLQKGHG6htVZB0Na8h+9344gd7OC/B19OSuxSk8g0XCcVMHv1EprIL
nHgboCVxsyS0A/a1rhcbYDQAJceTeY5ii9HjT/XXclV+JVTKwhiDtcQLGEYKZsmMjYwaRrJc9lGA
TlNd5GKw8828vOi64MxPni+0M5nBrZclayOYTfcdhi4lDgC56OVenr8L+7PIqFv0N9MuVlKZ8snD
GIHtgnLSqQil7mDdKcLJEQ6gzI0n6h8TMwJ/x6QlQP6rgS6FoSO64XWVjNbpMVnMYp9xRWtkP7Wv
owYImKTA+fljXq5P0auSgTkiyyaYYESl15g/mpJEwBprOL+KnnwsUa+aPJeRwFEMEbSKEGX7d+fi
9U6W/QKY1o+/01syCNYW0KmXTPknsdr7dBM/co7eX4/0bvQHcf/meEHwaOjv4QUTlallHEChqTag
1eghCH1kL5RGxUvfU/eUestaXQD+DZmjltuwDeg/SgrYRghfE6dATLShS2KWy74977xgON07RwGk
BPF8EYcYAwAmuGM15MLgPlL1E4rE8vcgZ+JCCQLi7hR1NwnB515lPC3hDboVFEp3KUBu6FJQR/nh
4XPRnsClCM4P7plUjROHKKXO1/2rzjCNQ1icvHJLqprzeXP7WP/suTD+dd/3C5pkmSONQmWyxuxF
/mdn1tEmzp3fQd4I8x8Vn5Js6FTSAT+uPBTvDJX5g2QqAIOE4ZJyNZa20V8Bv9TX15xHSqLQx5rL
TH53MULJTTcou04VJab9rY0+ki132/csK/wVx08MRZ4+Js7ef5MoCnrMS2r+VmuZtyiKA8pgm5yJ
jZd7MOFCIhrzoJUxc0jOfOwfavDZPTTLo1+UWy4I2GDRIeAJw8/BmN8VhMyfHkUBkB0hAY6/1slv
AHLF8+q3AvmJTw+LuFEc+jBnt29NfjovWiAQDQ2AHeP8teMtW8wVggkASmvJy1wh/yPjQcmPqtG0
QwtXYzfP1bGAUDIvU3bVWto8Pwk1+tXeS3fbSYYaFsOwKL7c78Lgyndh6R321e1GD/nto9x7lnZ6
a3vG3i2Q1XhY8+osJSa32Y10ybR3XXT8sJiB18oTZCoLyKCQjAdvRoCSZUXnf2qsn4NBv5RlS88w
2MN2BmPocSoGq2Z1rwzDEFpnIYMkJ3TPfKmbSmygQUTxxlZ90FjL281ru1zHI9rd489F+PtzhdRg
jrPFm0n+UdK4vj6fRU34erFp2jVVvdNvbzxCMWmnfRCVnHGQdSTPE+8r/Jmhixi8eJ/2bW1HO+v3
yWDk7smtU2eiJNFQctn2tfzY0Lr9jUmvolfBtbv2YAsu7j30L2H7tTFJX/KoL3VyjHzR92/bSYe1
2km/foTGRo1ynS9naxyibwex91uYyTOKqtanGIPhzbXTYKkVdRVnbP75j0L6U9FKkMOUrSSV41qk
9ojhezca15fZieHE4qH0eAPV4f0140kBKobDgGTev8raZA/XHRWrrR72W+Syh7/LpD7R1gmO/b+e
FT4Dq6vAJ+SQyuf3/xD4f9Lns8L2bmOFRUljQS9wgTm//hXHXMtLrSx2dH44U5wcKVMh8GACBstD
4FW4OA0kPXNA4nTr4M4SLEqwA62zXAJf5ZTxLaVPO3SYwMlKOdEk8r/rhqoMekOccFDQK1nerT9g
NPZyIGPzGY/D7873N/yiYOc7lL7zYo87demUo3fkIq17z6L6vmCRRP59hLV7acLhZnvifi5RwKSD
93dTpljCsFIbtDkaGma8Z972SBsLu4hWn5XWgOeKYgHrq8EcyavCL5Ed1Lw/P42pLbr/p92bWxdS
AR7jXSgxVFXoDNEPYpsw9yyEwTxjjFGMZT/AuJWf9eoUTONxRVkAdNAOLYQCwkGDLQs6SpB58EBo
phyQ8jA02To1/OiWMVL9QiDZNioyPD57kVXmAFKsMBDtneyDPgBvv6CLsGlElvVebRKwoTAZqHCp
ZB1va15QnWVqNV7lTtrPAGc5tUkNzCxq7BR3wHrstxf8ex1tSB0ewHc7ykMwf52dTKS6KCpHJE94
USqn4cSX9VvdxssQNnRhwcgZUL5TC7RBSqZBPAoqVpCds22RcfOqeLCXAu6CP+A6WfsNw7Fgu3QA
ktEbswAmrrZ/w2Evv6YFImlvI+39Ds9Npy9VRPhYbu9/cns/Y35CXtCl8+UjEJHTDg6oVDsME2Vp
otVydl3wujsZy/IuVju1NgRaGTYlboslPKQsm7m0n91B42Lraf/rP0Xqo12y6ZVnvsBKWCNy8Q3+
Epk7hxuP5mOyoHCnU6MlWjZg4hdCc0gcCV3iYC6h1ekHj8eB23yB3hLl2cPW2/B+sKbn4OJg+twW
gTtJPVJc9f3D5YEEeBfxJkRST3PUzRYTie3Zoj1pwwKCan+mPzgJfjd0d15MhhtF1VBZaniz5Yqq
quvwN0MO6PKR4eIm9I1UWUnmumFi5ZU7lLLJpmDYo5VSxVYiGHk79OhSSJ+uRi2GbKKmflq+3YG5
hcRPriEMB0ZnpnKTigH6fIv6t5RrZW0azkKTs8Ivrcn1lebhHnRkHa6tLGlEt/t77FWV29QsVC35
d7yiNVixorft+l9lFQf9R8E7exECKMGn+WJDh8d1q3GPRhOonIVms9HtcTZYY85qgrRNQ2+IjLKZ
dtE5QrDz8oeZjP53CQru7o9rw1nUXJNkzC+Yd7Z/Gqcfpx5OTLNct43V3QKbirFxV8/BWlwz6HQj
YCXfYTBwmIc3GtLvLfeQ0eqslTqZuXNsBBsx30xFoYxEilskfsbT94eJCg/mYZ/+57Usz91QgqCM
q8+wN7B43uZCnX3Pxf0FdDuNj2MVdTfTQXW35Ana+2l/j5sUPylTFv0XPmu+C5YxlaIi+qdjrSpW
fGkAE8B5WBsqjXRC1VzS/V/8FArJLqBZ/K1x9y2q2x8N1VczinGVDdeGu0U4Jvw2fXOlakKOClZc
XJ4ZuykwRNIz5KjS7brOVAcEyQ+AM1016NwkFVXENJCAVHV1UJUlyw4Cgec1x950LAu0iwmfHHVG
Nb+rucEYPyzGcRW8hfRINw7ejGeIk/VyyMpsHvYGtdcLaDSYgp7nKe85ZLG2zjl2e9rD5GY4vX/y
/bibf2/CkJo9gnX5Jtn2h/ilTr7KRVqvx5/BQ8NYn7dGjaLUrGTqu2z+9tE9z7771YFUxG+DIyhy
DE5jtXEALHE6LnmlyHgXLo4V0XULSW1tDNfaWGs0Rz0oBr9iR17tc/xKz8xTx1IH0dfOuE4/akGG
zs+zOiMbpyuP2EU4v3hr2vhj89QkqXgE1HHX23RQORElnyXUdXJFpNHZMGnr7z18vpSqCFrxoN/Y
b6bLv5bUyR8GVpN/KDkyp0v8tzCaDmiWk6tBhb4v96Nm43ik0T+CzyeVh8GSJREqIYO3H1QAbqsV
EDkDi8vp9Hgk/2Its+RPstNasmfSQaSY9Cf8MZG9YITwVRMbyr+jlFNCNrXyvGkrsjb/n8KeieLl
AggswS+/2hj0YSvMyaYUs605fNXqBnKDXeODN2kuOJd7+dbUQT/V9zEZoyvyqMAD8FBlBHukbQa1
eELPuDB7hpN/jq21MBePYpe108UoTWfjY5LqTqJ9NwNi2kobYVm/pQzRD7TI+Qt1Mqf5G0Tblpl5
AJ417w8/WpYqZXxjoUBebSZC+/q/pni9PgJLXd+bu+fPjXVTNjKZ8BN9MyS/oghzYVnq+eQlWp9V
fBrO6t0Y4ySxeQANHIxGs3FIQRJ6PsqZom05RvZteGmXuidUSBhGx99I1PthBsI2cO9zzLKqzmlp
rJhCPK5hYlTceNoeX4GgrOC9kl5uW3Jjga4ZIB6WvY8LPUiKpK7sIhcdZG5zvEdvEbckmCIgw3hQ
1GC8M2J1DDq0pz/VYi0opb7SZFPlA8CnN11MQS4iTpEYeYrc0LZRn+dGdCCuOCX1Kms/5qku0Qgw
nqawy70OCm47NAdwyjcZWJHzpp+Wc7t1eb1ror63feVeKvhTRu5kvLsI5RyftVIymhM1+hNfMKIJ
hiCZTggqwA2J2aMT2HWovVqQtMmEsiGbOn5Yk1nOwspocWW81Kb6T1OVzuqkojoI12dDOTmmaJUe
lV1Tgc5bJ6pixXFm7luz/RuRb5XG3yL20/FNV7UCfreUGX5hvr6eAIdZFmZloNJHcwBbldUk0cxN
GRV7zMR7Qrn+KXY3I/PRhDGdScNIGSHuU/ygKMM9GItc9j0v3VoNC6C61Wuy3ECQ81XVxUlRi0R7
SqqjW3Ut26+QcJYWLBIbGV5+9vH6MBZwK2s5nyAUl2Yu07di1jbGXMMiPoNZj59Llmx/Q0n8N1WS
6Bf0yn1HitQAwnhTUU5fjlKj9qrQ2BLK2ept8GJZhP31CDfP09J9sXGsGpse2Mfo8VuaCnV64ZYP
zB6iiQpO21D+V08PBwcXXtlCjGowTX21rUFDsslxsy7RjMyVDoEPSed7pvkAc/2DdHVtOWB2vfEu
/D6w9yZCQKHKuF+qy3QgIoH10vQ3MGQiC+j67x8a89G4dilaFEMhH9ydzWidA9KoZa2CYgWCIhgn
nCFMd4MMil9pPnJWpFnvGqJSJI+hsBxB3YH82fn7lvJtqS8XJOj5cflpm/s4JEZNDkXQ9W8l7y/3
3N5lPBm8D4Ff3iZAb2JmSmhl4sBsdmqZDERJy6gDF9zK3Fthpy1zLiKKkuFCkZvD0KkzZBpGXNty
xvoDrLXOnZM3gV1SEtP8EiG5Jt2FNkXOhjvhgF3DREiWkKy55QTSJhUpJ2zhWF8/9bv2WDxoNJsx
rkeqxvFYov4CyJof0EEBIkNc5pSHJgi924z1wLrDzam4ODjKpy/r4KBotqCMupmWjXd7QJga8GDO
yQuYXQdyea8xuvcYpJnlBTW25bLwza9YvmDA8xc6/1ia9o4PZFuCQPDp0i3+8v1SFm4BevY8GcZX
hykYMXaPVvp7T5BDactirP2GmKr8/FkhIOb+D7rEQ31mjrIx6c9dYr1lyqulT8ATKNh+uf5oZgc0
BbWbI3/HLuSSWkchJGW/WWmb4J48ieEKIotrxU5c4O9AQ91Bc4qL0zHS92Vlay7FT14kYwmcyeHX
OusD4DArNRDFXRPLBTAuiNSOXXb60lU7ViFo1xhL945+2mCabPOcQOIGsoGczs+51iz51kWAfQ9H
3i93dwsxk/g/flFUAQUBMVojRHbzMQVGWN7rR/5Pmt7ClV56Y54+eHB09/XYuuced27UyvsWUyDQ
NRR8fSBSZUpJYCCy6nVGjGItZHqTKcMJBE+fiFMBCRAuh61mmMCvrm05yaR112+CpOinenFi5S1b
30ZpzbkNfUKwOWtmqUVMt/Wq4uRzBqQefLNHrbY80VDEy4nx+NrT990ohdyCHctXjnaZhukw2UEM
d7wBiXLFV4e+1zHc/L94LZJSIs0xp6G6gu9V52sRdUT56bkt+nxw4wiiDfbBCtuMVtnzmkT0Eeib
+VM/g6NWdiSHiufpbIX5O50KOI2N2T/jGKFOSxrfJJvIXsJdVNjxsk4W34GCqSKihiVjFbqH4Coj
/Q3GmNA5P/6dluLuXp7t1VIOuxbPrQSzoZjCTDxEG45iygm1NLLestc89SSl+x2WVloTiPoljsD6
Zgk9EXaay21d64ZQ1jgWkJBDD0eJvVhA6nF2by16/6Vmt4tzMgrCWvh/5b+UVmj8TR2X9843uZNK
RiRIpPLP+FD8IIdZcWEGruiTnVRO0ltoWzPgizbM5Bk7cU43pBYe2xQWpWFAIB+/5y5aAJ0GBycn
h7yWekmBTQbeQ3CByRvaazqdsZdW45rwDiiRs+UNM0cPPhHQy75TqK+3SQEpC2UixhjLbhxbNz1B
ggK8Bx9NEBMU4WXC5+TQNcCUe37KQFjQDMeUrBI8IeQ7t7TugbG0x/DzN++lsT73p8EW55ACboc+
lh5s2VCsFcgKXggUEY+7Ng0RfjQKj0POWBcIkm3f0uLKPdgCj5Ll272vvNARD7z7FIJYRavc1lP8
mWLeqhZoVTL3+r3SOvmRAWlsWBhKjd3LJkEI+9vitA4RyU0dTr7S9Cjkj4+iFBL2xQCFBZl2Z2zB
RgvRMInBKL6s9Wg3Idb3PZ4TZlia4yKfOqYGRIawLrMSxLLNuKivJ6Qa5D90FVp49+U65VWkzfde
6DPbpFvEEoefg7jlQPAi+AoGQCBeIMztcVxCvidpgMDFn8+lSaSvWAyC1ETQ7HI69sBEmSvfKNE4
utDbjjk+jdApYshDSE3msDenQvQA+xPezeVaKezSMRO4AI6bgKXHOxfWMEzy3vLWe3rW5qa3FhQM
O6bpb6ImKBS63Zoj/1b6R/j8UrJpXiDArtSx0Yngq6qFLX11g6bx8K7DzYnAXd5dAxmQEWLroww2
toIQpup7MqaQMmNwk5MQcnDEOLjsMeGc67uuRL4wixIB43q0u1nD4s2crVbeRPfS8pHZQZ2dg5pJ
N9XdYQG125V93yuo+mvXMsUFufaTy01MNLlCWURSswwfb9bUJqo7BEssSlMLNa0Q2IiuRO0wYHF6
8S4stYZvzLdjXNSDi+o86Qu4R4pHiT2KZL67DeJrh7ZGrNap0BOyoFi0jWqsbOuTgb0fIjxHLKJx
iVDGVCeEGUeXqr4QEdtQl/9FHrU7mrO3ZD+1yEmzr+/FTmpxPnMo3oSaWiv+R1wW+JvElQ/0qBbO
jH/HlTLaEbokn2/iGOx1n0aTZdC29vws5kAt4Ir99XC5tRs25NZmcsjMBrJ9C74zcd/moDcao9jy
k/TmaoMakZeR6Jsccy/hTK9cyjuZLyy0NPw+dHVRT6wn9KvSJamno1ZeZkY4uL71gt5LLNNece98
ua65b04N+65ZsEolQqVCn6xNDuntp2Wzo6VYfemRDf2Yzw7TNc7H9KWwrvUFdmPnJjtu6PtJrpg4
KHnX0m6WT01vy9/KMA/Uo1SCm1lEDvLHkMT0phd1ZjmC93Hodq3/1OjC7q7CafVjsidgZ0lYiMeo
rVIMYSPWB8WhFe/40kve93xuFJhdu9ka2f+77Hh3PvTvOiKKCMVNFVbZ5/lNmDXf8eC+Y4jpUEVa
eywZCfDFtKG9ILJLqpse8+5LBElpE0hueHmgosSwUPmsqMCVVKkhc+XeNrrPQIBNdRCQZq0CeRee
fmSARI4aT0HuZ8HgJS12JA4+3j5no89Rltct/BXpsB6h7vHdghgNKc48n+Sc++uS5XoC+Y9P6yrU
y5QD+m3t2YFkw3cUOwLFL2wwS89iza8e//y29n4494sF+3uUxYJmtk06jDxURqYk0eAuBXA6O2Bo
sTCTHqN5IxQsKK7Wm+Tr1QluN5oKgMZX1diR1KNI58c3SysAs4CM/Iz9H2gtMo+zopCnFtoyesGs
WEXB1/hX+LaJJJ7Gy4iPdcUTVAeAip2+9gQVVT3GFLYho7T4Q7Za0Z93Wq0HMMbeM9LIEGAdmOmo
Ux4WPeha4Br++eyM8vcjf7oOD+NeHkTzlSJhnte0xzbLEww59ijC/OnXqoYW8jfqiVwf/lLqGvqZ
XkDh8dHE+pBi4Bvq2LPWF+iWPeH1Sqrzap5jpE5upqaSksjZht5F//4Hr5DE5gA1VCq1n/8rNkFd
pk+r2sOYwHKF4wpAnHaOlxu/20A5AlGBbEqN6G3YALYfTjSDtpqB9UDctdyeux1rnpSs0p3HZPvv
Z7TvHU3n8CpOa1pR6l2IP0gxL98G5pmZbjEJbSbHon7CkRNyfBwaU6ac6rhe4iTN5EKZCEwrLpLF
VvBVUMEMy2a8vi1aY7LcqC8Q6T51NSQFJwaUQDhCzrJyazR55GmmUTKLKxQqOjXnl2Z24IelkHWd
QkH+jcy4VN/K83h4hmbJik4vOhGZoaREYx+flE/A4O3/egh8/N+c/rQ8RhPIzLlrHxptus3n/mBg
NZNeuOmVL6d9qvktLEeoTfqFCkeTbRndNI8k+jiYxU/c4pNEoNBCkVZ0wgBoHnE9oqH8oac5Qav7
6B1r1ohT9/R+QcpsWwkk3XiuJro8fyk2zQVNI608BVD4ch4M9UpigMKnbeGPMHgLw0lWlLHs1SPU
QRAtTKiTHzcnVRpavNI43oMzuyr+EreV7KVgslDCNO1pL339UWjgtUrI/GaZrnkN42IfA37v/smT
3gWl2+PZkBpwwnei29KHxJIOgbWFHHLxs3OW17L92x6okvVs3IPbXk2IKHdDybvcZs3kOdC5tZHQ
jRGsqqrbiqnjdSehL+nnNYwaF7tRDDn7qaS264Sea7xzAqd2yJg1uCcS3CYqAu7hmcgpC1gQlrk3
Ba7v/rtev7pKZtiF8qy5MOM/rCQeUINn2N30M6zQgiPLd39fF+iE6NcXarnvES9BAKQQJJwBeyCK
Sy6myaG9/Jh98PZwpp/WvZmo4LVMD1JG6Od5l+86djhu0uwaXi6X/bUXsQuarxFGCfb983Fx4mpO
eOxPTPztVCCM94S7w+R+jEf0oTJUtALmJwkLL6nRg3pgAi4tsNzfpCO1kQ5jiGZaRhreMngU51ol
7qngJ83Of8aV6TJHHIjKKW7xrILFJoN2klMyiKfv5P34b2emVEIoD8JYkdrDNtDI4eI+w3F3l6kD
HMvTy8JMkqnG+HuXvIqA8156hhIad84RyO9y9ByRvejLJWqZRcHm/Neb3duI/+wq9t5TsLS97Drs
wS1qrSmaEHjxPgPr5dnJqZnyPtEIGeeE5Axk5hHxDnM+/bw6Pw+JMWOqeDlcX4Kd+wTG28Ca4L1R
KHofTXbdwq3VCnJQNLz+Yg0iGvhOhrfcGSFQQup4R7TraCEr1rUjyJlSxiGrrASB6VTyMx8Fisat
0rPpibBffCHuD/QizoTWJ31W9ApeAQcJeQbnZbrYoovabwzptfbOy9One0ycmMbeSihMC36NmD1a
DB58t/BGhAL8lGQ7m05KawmtprX4BIIJrASQTzm5ezlYgMugI1BGt0TtmzZzZQB6x/R9sH1cLqCM
5aIXWSjQ5kqg2ahTUbIwMvaTBNqeOBJWearqUmR7SXov2UF3pRdXxMVn1cbkF5Jd9iDB92gLHjiP
k4CH7bIS4a7mkeEMb10D9gpTyX9xkBlgRzkS2gd5pCPA7TzbJGPF8Ju9y1Q4HpFtlsm9ZLRzfM9f
xsL9PcRL74mrayy0TeNpfmxXsIB59lTjLQXoDmOyE3+gotBBpfMHmNcY118dh2+c0yU/L84svGyK
Jd15/OTnkvPIINND+QOWmBLJ4Af3LvYI+b324uAbaXrS7JiDI2ohXupp9cJuvtDfhcL4tQFtdPi4
iuhY8eNOeQ/N8ngWJDSlSFmJE9wXKmXW2xfXtDFv0AlHqmqibrXOrP52eInZrpe9js7DLqHUtXS7
6ydKzUNjK+2z8pPozEmpY6QhqMryA9ucSgaC2xdYJXUP0tH1xuQqwZM1p62FgYLUIsQ6BZhEj766
Y3eEI2d2O7Hd8rt8tKhAXTFqlsqFwBteMvwJ56XeCfXvFNe3mmlC4nZOEPXH6MqFXSg6sbcKYcib
eNYNTGk84krSw30WoTUCQHzaWpmjP9tuesw9Fpd0KTRtdGTOoTp+npscj85NLZDxf2Yq2shkHKr+
qwem2kYR+0NQViqZ536BX2atfIYKAeuaugYnywKY6qguMQmmx9qEqxx82m/xlSUM94uNXKTS5knA
NYklPglkus5hqYguTKiXZOWSEcw11s8kCFJYBBKzbeEy5P7gPcoKzvPd8NRTgLWuXXFp5ZYRCK02
VX4fxNT4zSdV6u6gIwsxi8yCXnKDSb/DwuB4astqPaBIdbiMxDGi7pSbAbMq9RMWe5ZiAVYrizlG
JIZMk2kCO/TeywiQuQlFUJo8FL6eRuJGiEIcAvUaVq51vsmTgLnnXeP1vH93g7XP25Z1XyI+GN4Z
TM5a2AS4KJ+DsPYCDatKyV9PIGBbOEzlpiJ/d5uVsaMNVJ6ZUXGx0VwIbD3I/BVW8PdW26Ig2OH5
e+/cJgNAAoN7BSTJTtgOychqKfb3V3YGjjuOQLIbnt3CstLRsJPwpIDhiMU1BqqJPDVePLlaiJur
Tt0sP7CgY9bwDlMJDB9JEl5DVR46czhEovEHKGN0ahDshlrRxWhWerRbnVoMrAmjHMsgBKtuEmZK
BBypswrd1vavxeNmOX43gKdkOF7zXLIXQbM5Qj7e7V2w9nNjDX+k756oRWPlD3ad82TieGkgEDK3
4JtRZ38hKnoxIGpzMctGmy/UTvA5i2VI1ExsILWUZH+WsgGlzLuRNr9T5rfT9GuK7QpmVtxiCU+a
Vse++wWFCeH8DYkPjqvPUfnl9FZRFizCHXrgofOfzd7NKcgfz0kPw+xXbL0MihIveTSXDXQuItWc
4OovJ1b42WezJhAPjZoHaaVbXMQkxMEwJeXiJ7uDT7Xrw1TRjiH6Py/S2+CeX6j3sQp54XGycQMI
tqYqopBlXokFF+2mGvBBMZPYA3onSfOyNnZlM0s0lCeBO928cUzQJmBy9Y00f/k07y8e/2gTu43V
pYz7UbsGyWIw/26V2mnvu/8nm3RDZ7ngiw9wdOAEYHiGjXD9O+y9EDxF+SvlCvxqr6BFo7+Tk2R5
EyNVXlRgrtZfN2mRBd7T0KMQcej94iNrX0Poj/4QFG4qOI496w30tVKGa8a1HmbVsXyZms4uH0mQ
QYZLn2P7hmC6Xz8mXFQwO1kcL2gTo78w6pSZ1Ud0BlIZXYfi+TJbNimMBo3+oydz5FZ/w97c1Aec
hVOsmqJwbCZmS2PNGDU5kH4f/VL52rFnCDrid3Gry612jfncJ4IYtYkWphbsN8uAS/bPoTAeenvp
YOTA3c+RaA+UNvRok+wogYQeQ6EMzkaL/yQM6kihY/by9yjRqSJqwEcw/4rl5Jucjs0ljrrZmtDe
idYd8qYVlYdA3APTr4BI6xICiEc7vEB4aMMCDn9I2FN5knI+1UErYRYYW6tTw9pp6sO6vOHNKCUk
P9Cga0d/1cjkfu9bfGrjzzBl7x8wQ9kIlFc96HsHDqcT4xK08Nrt3oCnJRp5x5SHiWiIPI+jBYP1
2AHPtAgFIy04OJMvaeOgdbETsOfugfGYq9lEooh8sa6y1PuGCd4lHhck8svLa4arz626QsK1pksm
isL8UQGRj/g0vy+vX9gzSBMoahV1+fc7QXXFxiMoIb+ZwpDoLMKgn2zUosTln4Cq8P1WWUwTGrAF
keyv4Ht+VKbkZsElyCcmBC8vBfWw1dTA9ye0J8YqEXWPnWLd2a3Ob8Ra/lIv0zKpoihMLDL8s+aV
oZ4qcPMCouMd/Lq41wNGAxFBGr+olBKqCacTriSCppjNYK7EnMNJDTe7h2pksOjmWVaFvoXXjZDQ
AUjWcBKazTuYJyx9LVLMOycyJEG2fovXDiGz1mrcGlTtJ08CqZFwbKalPvdG3bKFr+aIAF5U3jkE
KWEFxr1+QprTnNUyBTS+vRk7daiR01RHaozKwNZbgf8Mxge6oJIkhIxmWDmRo6ZMx8JuNB6dPL7k
Pvzv6L+R91TzGbelYqAqsupoDb7+MlN2itfirCGBu++CSQPnVq7TcKkqlQPPdpDDPAZpfuDYNpVe
DlJjCxf+ASkH/2wsXVG/Dy+SGGXsCMbfmqh8Ayr7/bCpkqTvjfciBLWSjLVJrs/V68n1ajViopfu
SEoa2ZNBZ6UMeVY6HW6EF60zTF51tI4D4MNqHZun8mjJ6UG6PiMxrY3Mms/UHv6sulU0s2jLfQBz
QEH7f5JGDpXmwGSpq9bWruTCCvHUECwtFJc7w8ZcKVxH0j9pGHt3dsBO04FRnVH9q62p0w3YjcES
uO8AKbZCm9eUYNBiqgA9neIKceOS1r5kxeMy2aPBy1YOVJzypjg4J3UsmyeBlyipaZT7Cu2EZlk7
bnpxGYccn+Z78nQzUuODQDCnYTGy6q3QhpY61h+t5rj9QpwUjLvVlBqEssH6+k95xHXDSZUl1z8f
7Xn26tizPJ23khdZuOaz3T0jWEihHAOrnCntywNfZ8pehliPT2xXogOMFG7MlO1m9p0BGBzX0T8H
OQWsp9pUvw0KcR4s0PvdUMVykFNfJGw8AofJKEaSyXJJa5m32MTV4bh7nhzJC9OwRBvC8i4nvV5E
TAlBJ2BGEl5FaUojA7/KQVtWXAB6v6NOiDatoggLpn35sPfP+Nk9GvVd9atVNf00cFKdfzm0nniq
8opyHO0tho/Vk7ui96iut5Z8kOj1RMuZiJZpIS6PxjHpbtZb6i+Kmsl9XcLmuaD+biu1U3Qfx9+h
XlhP3WnX035mKrpqdNS/yN6ep11rnvVnJtej/R9tF2sNYmyfUp3iXq+9fSy05aHBX+7wg5IyXWGL
uV10WWh9qKS/0ygSFPz/o4VUoISSbFPyAT1vEXOLd8I/+u2aYzypMBC6S5nIKgBuQniWAVBNzYVV
MVGCjYVu7XJtTabIaVmEHg60BwYfM8Rv0d4rKjvyTrNCWucWuC6Rcd60PvJXPM8jLjiL7rllW08H
bXSdgH2e691Uwz+E+t14qwfBbqTmQHFseqnUMv9ZRmHEa3yVofgPFLPkAxBqG13aJ5kDi+SAzAP+
3eFBBkKRIShsR260SW4eMa2nT3eWVj42SwMwZwhHtEhrzWXaK/mSoLBo4D8bs22PZuUCwRE8w5LC
eMCpKXhxaFbN5mNwZNHnwtLu8EALWXGWSVSYZ0mpjQYGj4IlZ4oGuxR0xm0RG2ryWIYPSYi3zbP2
1w5bjnuHGkHxZ7875lyXr3m0c8qQI7tUuNETqw2+cZ+4r5hlcDV7wzU6z3mwv8lqq08UFe668/iX
FxS2s2eI/ELw4P+6pgIeZFoFJ/7Q765ElrAm7PEWIb2FZD/lzhyT1BjuwyGS5VRxtyDAt8zwC1GO
YEKCDSqfp399SyqimsYgNUTZtUYT0nly2DhYWbagjnF1Sf5PmQxB4S+tqlLOz07gGmHWVGwi3Ocy
pFGyaZxP/azBVI/Yr1/dlZuk1ZQFFpf9fpoZ9yl1v3yuT2zsdcxtFgn7SmRiL8swP7KbuYzguSRH
/P9lTYEvbUOaFG+03LU3sAT9gdFepyWl9+X9KS+4Okb5F+jeiWJb2wE1EaUtJQSiClCSWr4i3iol
q5sQ+rh2nktB+iD8riVoWaQLQIliqzoOg/twfFtFmxrYx1otoj+eS5LgREBuheYFj+xX5SyrK4lH
k0Kuyy+169gH5Z42BcPBHQDLjdGkWx2hiyvhI4TGxcLftZWtUMr6WO5FS05SelEfmk449uvxmBDi
auNliAh5we5+e91sF7RAm8YYwk6IsOHQy2AoS0ti7kNcX96VmSX2ykHiEgf7/toc0q06M/Fo+NB3
aBvAbS3wL+m8yFWaL3uaPVw56KoWPOasgz8lphJe8OVqudrAA1e6B9pefUFYDiD0WDJ693dBmAp8
98kp/NZq1t4ySBLyF6mMvI2H8h0EsluYPi/95Q4vcHqO+tHkNVFCGbUe2TKQfnK4b15dZYFtap2I
aHmJUIwldLdq+VbRpTOYJkDFnCJVu83eZwi4InjYv2/phvu8Sm95Nb71f8Z6NB0STdj61jHmRbQ5
GWugaYxwnwOfwJ2QEr9Hr+RP2k57+qPlNLPYlnYMes+sCryxJN5yG5VGSDpQ9ANRFKpykq3vazhD
b4xqNZ4xZj5fDSLRcBBlTl66xeZpLzLqEar2EDaiWwcynNwRNYSUoa1yKd9TUtRq5RgLUlVKXwKg
oCO5ejUqlG4Dgi1Rsn9BfgWtO5l1gq6h6XeO7ZPdGbNTl9Kh/jQNo6t+jFnFT7qdXqd5fSmvW2fp
BSdr0u2GM/mToG2TbLvtCKMOq8XEMeywxQit8xUQYhtWuirjqXKTeUJu+KuYgcs+lmlV4L4CLhg/
bMlDYdG3rN2fk/mW0R6n6672ZMUXjAkCPtTAXWwPlg+qGaem1x9S5gMVjGtV2PVIaymkyRzzteEX
gyPPiLoi5Kyhep5DjF73xnhEydhSA77Pk8nP+enKsqaSghTBokvosCum5yxunr4nwq0wMyMWNDlt
Zb+gr89AcMAJ0KRzP0voHXkzNK2XlR8Aeje/SIpR4LaqkDPK4tu+QjEgjam+8Ia1Mt8MkiPiv43x
Bv4Do39+ghBgsd7SgeoLB1MbOeyQiVgsVLLS4PzAaWrI4X6lpXGxbroPCB+hpOjr0/2ipdqW1D3I
gpcivc+M1eWr0RUc2MMwM5WLdKxy/GKmrZGUyw/L5Zb01Ss2F0H/Eo3GpaAQBkmPCUiUh5B/hRPr
fiKTrnfHa5hgSF6QAqXbQ+jMVWfjTz6G+TZivLGic3Fmx9ABAqe8wJ+b2EGV0CM0Q88Y0km+MGLG
1bzFANo8prC8lv2o3hNQ+Cpa7sTrWIp2lnuCwWGv77ejBelTv7ImJ0aeDHVvL/27DnvBvoFMFfFp
iaAfFowUpN0w5sMkA+v0yKrDjqk4mHA2PynKSa7GmJi8AFf1SoNTXrT7jKoMlXZ5vvnxjiVrXfgI
Cbyr3m1RsTieycaTcJWDpammNohEchOsa4yN0hhtVLILCKbXu72C43qsV4KADL6X5ykugLJpeTj8
zz8BrWLi3MtxBQDk5FrMCwOQ+8aVdvvtCkNFdZWMwD9p20Q2nwP7GGM7t7GCo2QZV6VGctu8xhvb
amJ5v9gzfNivEnoigO06haJBdRmrD000icp9x7RKVZM18VCnG8tZ5peSySuAfSBm3EsTRbD7VdZU
sN0Krax8IK9BouuaUAI4x4ng18RtgGIVsffkMmaecQef4lzwhzQUx4L+vrI3tWxUSxHhbKng4EUw
rBGbCkbq1XZc3cCReRsdfCFkPwb9MvsMXwVkYLNjwsDhnlycq80YV9ymbpvnr5kWv583RPHoCdpb
tUGsNLRVNevFCcgFDurorEfVDmhu3+/Ju9kNHGy+/Qov9NRfgEk1zr3qfLL1tr9J9B/78cLKklw3
LTaXynC4wC4D9xoU/KI4ujqUVutn0g3PQmevLkXVfWIQY2C/4gMLNFhzvdTejYv6pWchvgyeo0m8
PehMpJ1aV+GououWURGJhowlJqy920+H5muJ6ePDyRhMubfixkVicKHuCIrG2lTdtWK5a+lTR1uZ
QxxudooQ+Kum/BbCVfD/bJh/NZjGqhUxzp5iHwSdRYkYP3q9qhGIIj49BfZ+uyh0RsW0UElmLfEN
ppDuliezSMuGE9EgGWgJHJ+aofgY4rGvlgudxkVfa7fzZ82J2ZGgGFTt2pF8elPiRReaTsZrmPnL
sAIqgF217ldUDSdl079acDOrRhhF5l8A333onz4SQWuv4lK+07CA9SDpE6W3OdEjIYhFDvLQgWoD
9Mjxb5BdpI2ArOlXt70XIaLSApLXB9tkH9z/luPfGxC3EfiafQpnA1wvjr4Nbqp5+RZlI4hoH6ft
7wJJvfeF7KvOwuyu0hB4IyJRB8dxrJARdO/Mb9aFA2ADR3IGZOA3dWAa4C/t5FvDmBSp8VLbSfIa
zp0lpymV751a5TP1jN/G4QUEsspgCW8w/4Hyeb1MxhLqWc1Qd/NQR7aEQUHaBFwXozF/oEd3Sxs3
eAv9xStsYU/ZujqfjXpYdU54rhbsQfky6CDZyCaZEscNOH611rf/VIO0E/AAllRY8j0A4xZzmNa6
g8Y5KPA+SboYbWaSvaDdzeE004mhK/xShnqIwPYMVc2sJGnmODmnbYQMqngcJ217mjvytXyJxq97
PwpVoBkepdzl6Lr1jPJ2VymMBduyh6r7R9GmUhSeKX7VsVVLn2yS76m3YDIZz5si88rhjp60Sk4K
faij43W78IDrUpW2nKIR+oD9On2K8j3W7DmAdFFb37IKAnjWl6m81/ReGzhc59fIWVpt7WkGLRPr
a7epypJ1dP2EksMmilMFHb3kPzfiGYvsi5fVMMdNVV2ZehbItOhNB5nQ7RjQ+czmAGSosy5V5wRG
Kt4La5AG5pbbEWSBJ0sxAxalgYVnElaTsuwDcg3/JnMSmNILc3slB36SnbuAyvt5m7M2PJPT3vLY
wpaSWLtR7/7Q2m3DXeHGIpn7V0uE0xEWSOhw+ACodUxKluyOKMR3HgTZoCzLmNAkVLctBdKMV2pJ
/Nn9+0/pZyoHaV5lvnz2odOrBIbreV2aA8LOlnTN1+5ouYrU7qQ9NGgBhUboGM6o/eKhDjTmaD/C
+g7oUyCsyI6A0dxn/6QKPGD/GGOvFb/nX8M9KyemsIy2WbLFxEowGNXomQZnbTrC0V2P/OI9TFXd
sKppouewat+ST/q8GeYXEPhVTGagTjaFRmd4qJfUxY+fWEeHNFN/H4LFqFV0zO9IHDGNRGHTY+NR
EXd4Oqrfq/IXXewAygxFQw3SqH/DqhCAgti3nNmnhohJmUfth8f98lj73++TscJIid3SJ4eV+ozO
tGci8UF14bdtb3N5ARmticf0GxLQtKJGVvY1PrQnGX+sl8R67Mjw423+B4Ue5a2LtHFh27j2YblQ
O3DETJUfEoEX3Nd9Jky5Z4QWJqh62Nge+yLX7ANzmvoFRY+gQfnbBGHzPdKpQy+0NZsHz5vHsfmz
Bs0fo/i0eNzhqAdvAI6bhBYrYro5oG7TKZJWWCx5eXPVwTKqzcv349D1EsONkYK92hqNgJcvekqR
W81Pa+4ACcGWVOoQyiTMXvekq3/INvdTRo7I9kwxitXm0CSPhPnJ2uIWQHzVM9QHaU05/7Vws0Fc
fry258wkilrLBIIet5rE9ARgxoTtWt3HwZ4osDAcY/hlkC1OAlrwnSX2x8cn5ZDYd1dwpUDdQBQO
RhKJ/NyOS6EHPlfrQ8uy2EateQGyRMdDhtoaXkpwINN5yHYRzqgvBzPQyE3UE/SDvytECzsdWROL
A3fC7djH85QrXR4kc7izAPoU9uO8XNKzWqnrTFpiiLn7kpNfe02LYpHIbQvlU2k6jXryk8fpFORg
Vduf4H9fQlTvmRvMpsW2h8XWi/+BPrk/Cc1ONqQ9twhMCRF8476ltGmGWXWiChh1B3OXNWnhyc42
CiW4oOinT8ieyD1x4lOBcNJE2S3ZRUoZtP2D1mK+h4p/T890PNHN+DKK2Ueau8VQ69KYnL0H54dB
QWqMp6Hgf8TfnMPVQFNdUMndGx3+musBrZ+PRmq1xI2lVwJI68k+P3/j0xtlwCq3+LS/Q58uns0P
T6H1N6BWi9or1UQxnsfjTSItOzOfQjya8olpsBRtT57vG/hqc8lv64VZPieS4nbVNvtivA65t2/O
L4Wo+l0mRdX3MeDKE780YFZGtKsphG3DrZwxi+q2Xiz3luk9VI7MnGpmTaIMPk3bBGFkZuH8J7/3
QQYFH+7A0BAPztVYMv00qc2EDNPO9rYsUgNMqDhF0ig0WVN5nflG1Sl6Duv2eWlp7+RhKTWZ5mDC
sCvt5vFVcn9rpiquaDZdjQmlVp1bwpyEc0MmHfGXChMlSvKI4wBxUkhaxJtrfoc6jpSIwd4Eppaj
SGT0nHMrLNoTeEeKAizsBWdKEdNBoqdp1sFYjP5BmnMFRcBqFUfbmzSClB6IM7Niuv9UH5rsEcjY
DzpluaG3LTbz+aYDxSls1cA43DpJP3n9FNHPwgLCxEhsYegdgqw21UqPGbtHtFPQunqLcln2P+4k
oYUkYI/KjLINRVDeIP0Eg600lvErhy19X5zNYjmP/Hl5iouxYw9c2zLGB/0P9Qr4UcAbrUfrAB+Z
Bvy/7fZvBhgoTbtZop6NtTo4T+HxRHCEEJZIQB7ciJxA/ghsIgYcMqbZrEyaS7HKpqp1rBnaPEiO
Pz3CbXGXck8RANXfQt4n1LyOnU8/CTpcL5SIjZWqqZeL8eifqF4MR1spxL0f8UuWzDZ9W0y33l6y
z4lD4t+PUoO5kqLX/P/R9WKG0BTURbkAOSgRvMV8z4ihpGTy9129EdsV/70lVd1h67drZVatoiAQ
qFlQKDFnOMH8or9RyIQuNYrAvHVkkcSyM5NQAqQuNanUj/Uy0d7dpTxTycbx+KUEQ5IUKBI5ZfkE
aj1K2twZrZiM+5FoXRD8uLZX7FITIST2D3BIY20Lgdj3gPci6t+kE5YBZhX8PhKF+06lnzBnUETd
opk8FQkoL15HwE/giVwgz/TDFe+FZbr5aZKXUQajKpePDx5qDL0Cxh37xTTgVpY+sXMF7QX7UeFR
vLP9RqgYH/YzUGk+2ZS2M/LLWfSsfYI3If+/wo1Yk3pMs0Y3GOtuqmm1iIWJdMd9GzsenG9rmbb0
c8I+8+HAkE80krlpHKMEr+C70mQ6F9a8dHdny4auG4GYxlY5WtwDApr6XLOsybKxU31AH5XHU5ww
25gm0D0G697p/mv/wxPhfr63tOQK6Kvka/EZAMCwPWkCl015y2gPBjuJVbnXhIQmu6LmRo9l2JP3
/etCEmoKNr+dQLvHs+Dcq8flQ0nM7GKx09pjyxvfpgGowauCERAbaXQYTuGtiqL2CnEPDhNxjDZ9
/qFV1u76q9yLA6QN6mn9SrLQKTneoxcYGTjs4GUMm7ovV4GLzhb/s+XpNrRoxMtrv2umVm+jZZod
3CPCHDyXEzzdyoPesNWdXRtOaOLs31EBCYZHXV6n5wOsJrFYo9+PrBJ9yzUTm1AQIT7YauURvlgR
p3dS8pkG+Zr1KCJ2aG37I1FXYXZ9hI/1eufEWrIqtLna9z2+HBJ0S5d4IEiyOooKDj2ZytWwEBH9
pjvCKAv748wELPr6QRR2SnorppUtriQ9NyLeJZYSxJ8YpcZxll7qLMWhLv44ieCi1yk0UOdxWy0m
xPVxdp357exYTETby5xV4G2hrxkxVSNS4dq0soCufRrSYIbhOeHtZ4ptlKhZowzeHxMAfvHY86xi
EI5yl2aic+MHMETasCgqlrR++pROZVwkXfvhWpGIIq+gY9vIsHWvpgUGdNk6XqLxPEeMqjUbJ0x+
R9uS4DXHFhy1lNagbRDPVUBzGo+XkETmERFmymFzLCzCRxfHOee1qhQd5M39GC6MTWjOyGqZa8Ge
2bJZdvKoeQuNp4WwVu5IR/BL14zXpIeUI6HH6vFexuJ7gxnW9rMpH8P5cRxaWtKeiRFeDry+5z6h
7/j0/e2EpwAQJ6WpnwxWXDZr/38cM0vUzUStLZjGKThJjtyzkzvWM/d6T+66iZ1cOw3QfR2NHt5e
57QMbTwUH0OPUsCYQi9z5jWgrrXbWCPhk29/u8QzWHEV/l5IMFhscpEFFGwCpSkU4r9Sm/+KwfQP
QleqyoJCL9N9H6J/qHJPerknWJxX9DF+sVDtDkLpXFbHXWysQ9fB7tJB9paMefiR6+bJ5zNP2pt7
LBApp+Q+fn7HXe+nr+IbnIWc1uKPxTggziyxiN5dCsjhUUNPLyKuZZ35W8huacTeNFkYet9TGUnT
X+n3O4Ulg/EpxDTx1s1vCBUP0zcchPZE4Y4PHTpkAHz+ZItiy73u9ZkAvc93MUG5Qe1gi9vnLvXb
TrG5gqktKrZ6gZ/k+5ZaXrPWqUCi4vYDb4O5rXoFKqvBp3TTdePSvjk+DUNF6PDvTHyaHfC+q5gE
dikpD6qxMYZCpzOPDhPYTurAalvd45RH5MexGj5NefZ5OiRhCrD7A2qu71ymNaKO7PKPR6/AGyQ/
ikPCIXVz4KPVrY2avEl/uSmAU6K2PeDgDlYmJBa0BYg+OVT1wS0Lqi5jmrdMP2aH2nx9xv/CWtec
/KWKoro22aoOIiKvTrNfwDj+3SRiJDKYqv9Qh7VKMStdMH2ZkLFxCBlJ6fu2kFP0b/89r2phZ1xg
vjDUxqJ7LeWLECbjur7x6Emy8OvFfLHEXIHg0YiVXVmpE73NDhrUbh3c3r6TAl9vvkMG5mjJREOm
jFPw67+E27XHJ1cVHs2eT4qKXtRa1Gjll2jU0u2XIEvHmXx4IV53sM0X9/lT3KMJ3NAz+VeBy8fy
bMEbtwmiUI8UKbq5xkpHtYqs/iZ1wN0VoZsbvdOrEMO4NlMCLWlg1jcu8Yg7ROxTn7birexbwSUc
Fh2WrnQTaNpVy49ZKHI+dW/1tzwgwLsyRLT9xM/tZpACqaGQo7hX0cI9BoRyR+gLRdRS4Zai7UiP
xzCaHi24gYx8CZVfkgG2OclVWQgAGSeTeQ2VuD1M5FS6OHTUq66cLwy2gmkQBT3cja6OBYU1Hc5J
fDsxSMIpdHK5vMJBlWIey+d4NMmjXq18QyfFD1NuvX3pqxhYe26qLoZKRM/Z2J15XnjkN6nZ1Stt
u+eOUmb/+7OWRv1KSzvZe+sxh5JLUVeilZIicrLbEWrwAgLpPyWWrBWx5L2c0J5B5jt+vMpQWtce
5rtqf8YdLD21GffubLIOQXGU9SD7srj5cmAz3oKU6W+BnSAVm6h/GWU+w6HCMKDU8kZE+e39/RG3
KMnYc81W2OSgxAWnc9sUbL+L8SroUEudLR2XpyTTxuqhXK3PwURoBOiaeUhBLRhPE/Fz65egO5gi
/W8+21zeQQzZ+CTg3gNvqdzn6S21aBmN2qdnYkfineNI4cYMIvJY46qidr/x6+wKhAYgdGrLiln0
qjW6wRF7ubb9db+wCV0HJHzmR+OMMvDpjUygmmdXiNvJN8wMxJp3CFX7/vkNeLMVdjIYpcjr0hkh
8EFn/q4nIJmLqQ/IuY7W6FRFqCHi1QSlq+qzznsUSqI4O1sfEJSePCPwhjIBkVSdFxymN+sa2LV+
spyW5/xGuANlWyciTh2aBUCLu6k4wxgH5QYNSnGVRsdfTHTbT3pyDp88ATvpqmGUKDLkHYKjOrty
GlEpfL/cnZuvydHIle311XtoBqo41w4k2LIc+ouamWvY+7/Qf9VsgqDU1DuXmsZiXmv6ytTmz4oY
MCJfXzh8GvNBSAzO30BiPLe8lvhu5v4ALjhIga+saqZGEsUEesfnEFZo/6dOjPRkuek295KuXIzQ
ECmCSCPOoh5FQrUFZRer9NgYWUZDMAFzuf39odOelUJTQ9K8Unq8sAA5PzcJZ2E4wuJSBQ/rvGHN
Gs/Ygi+adDP4ncu/M5GRrcxGQcmORV/Dhvpqfv2cEZKC/XSBpWUJk1OwOdBee9BFVnXVI++W3IE/
u3332dbfopNIJHOo1Kv+UWbiCDqeabPy9OOKffMgdNeuhE+4/NZxCOv4+0sAkdtsSIfvBKHPbz9q
h9iPnawljg3KS6d9UGIZTJ7LmK3KZQAy5Kl+3NKcYcujYe3Gus1UVv8yP4VmTIcuxTOmEZMsPkBC
VMKrcVOec1WJMU8lsOKvXI2iNAGU35X4HYsrc3iT7lx0KWv2yjTDLfKWlLhuHY+qG399HwTIbQYY
gIZ99AlXkTxocRLjfwwuPtyrstRieIGsVj+ShxHJcvht0dtSVpQgjyF5RUCXmwiHqkCPK835rB5E
4dbplqd7U9HzA8/ySXrHd4rg3Esf8f9UUXEd+VLJo8ZvX4WVAK9R99o6JnE6yn8AKnv9Qjq+Bpb4
ffmi0IQt5ttJgVgIJi04YqB6/3V8z17+zuFnoGV6OFNTsw6gPN0klAh0zBTrB9y3bsGaIpwY1l3G
irIEB5LK9Yi77ROnttsA1estqBmQl2Zo27luWoD0C3zYEFYj50m8/v8tYvMvRqL41rOBipd7I08I
kRBzEw+RzR8CY/Y/YQDKfpSP+mO4mkwzq+npjx9Kx4QyQd7l0nLDqqjojlK9jRZ10njeCORBjwQ5
Rrg/hI+3an/W8nhnTi9ceCoO3y0qftxpfl4nsldMrU2AKKNP7HiHt6Voi0Ls7KT8w/LobOB5+Jru
JWMcPekWZd7f334iKcwMYJFeU1cHSIZWSlWCg+do52IQmQF4OaaXmPKjEosqsaknFFwFQ4mGT5KB
ppT+XamJxjAJrzP9vOAaKOyIshLvII357mpeIBaL2QX1CX6ITGB4lnmWVMPwwNb17XRCA1p8bHcg
sitpFKjXKvrgGAoedtJQcMWsiUToaeIQB2+Owi8wIVbA5YE175Lsk2dmhgvaE3UagFYGbtqrMisr
uFC0IeT7OFyZMfTUDFzcsjcL24/rs9EHQSTUtI3goZx1/ytjwWbZe7qcXonXVK0tgh7oatj+DM+k
xyti0ctEC6FJhn4afPOkF17i6jV8cOqtQVcHpwFx0JNu56YKTAHy5solAzHUg2HhhKvFBJ5Fluvk
hdeNHeivU6o7GfJL08Dp/Hy4IY2RMDd6PrXcDqBsbi/VXU8NqllcQrMQL5sYGu+RinKyFE9gl0+v
NfMqhpkFTLJcCgBfB6PNsZFsSFtwPP2J6vXShh7hEg3KDfDEH6HGy7mRMnRi2qVKX8k56ps3Uq9D
UgyJbMHTdSKmxYPVuuNLWMThWyhhMW/FZolpIPP6DnFNOvgb+CbLkUDwPQRJhLJCW37zuzoKz+eC
H6I3W/ah732GYmbNjwe/ICu7A5ny3jMYb63VBJqFuV2DYWx6F/VcjeJxGF3x9hme3ksfeciOzWi+
ZHYNSDNm2uz46gGFgj2xrTWvSBiwZw4CWwy1R0m35nfjo2md2NOFsUEG6iMEP4d+b/9Ph9MmD7H1
L3ggyQolRWiDr9T118XFODwn5UlN8/UjfOZQ9EwZ0CezOKwRN2GEUc7JlceLWok5vkclZ/xaA6Ym
S6kIhSrU2BsRnYlF4y3WC3Zv/6qxCrUFxvIuS/bH7uOORl9kUwCnHa6NC2zTJsucKVL3ByweLRqm
f4w9UNjk8q+x5rf8FcTgr9KZozAXK1awlnOJHZ5ok29gPOfs5NVIrg1im66HiHzFMYPUUv9hxb/o
xREQZUymDDSoztenIw7eAGWHaGBvwTtfTRTs3a7vWwi8sm9XBNSWVU4tqLzBc547n07Ji/Sh6s8Q
6F5g8fElJrHrZWTnfONzu2kZWr+RztLGkKpFwcjYA9gdLQY0e8oJUK8dAaWJkJQNurpybfwwvQrI
K5RMQ05rJrZ+M/cueeerCqbLyU+lEZIZlX0B/DxJhGdh8aBPL9qVb69oRKQnaJhicVn5tPpDE+eL
T6JhNFioFwjvvd+YXg1eRNx8d92hArqeo8C9onmsJmjsVf3VZtvRzWacJoZhWAHNmGm7tVXxFgY2
OvtHo6ArLFW3pTUvzHQE8QzSaRitOR4wGZxlf8V3bRD/O9sV4D0mJ3HXz67PctOoAlm16VdyZDVm
x82cowKVYxUV8kfHNHkbLf0dlF7klxjm+z2bsDl6vNwraX/8Z82eQx79Ia4pcG+5Vsfh3DPKiQY4
1quG0OFGcLexBnlcPIvrpXTe8OXIKh3AQaG7QiFBQtEArFLfxM98fzFjbSR0mzTshs/EPsZxpFUB
i4FnDrjzcjqOh/16yePugAriNdHNKykFO6696MbJL+0Wct+rkAuIM1sNgQ9JlfVugEffawhwic/W
Yqmqtiq4C199jCEZA/BS0ADHAfeq/X1Y8t/tIzPHx6sMgAxRfLNvIEk02jl7qCkdU7ZYW+ufzD5i
YfAqWPSmvb8+zw7b+OGJ3s/sYidPz93waGBGtzmh/JybUxkBrjE/kQS3+m/TqmV9VZtQfdP+3m8j
dzHLWpvVDtInKwK1GY/Xfsm9E+rsgriolLdmJDk+2hMsJjwj2cF2bnyUa1gyaHTiiEG5d5aXY5Hy
HUzSc5c20RZC9gBhwiPelXIzThq24OVWMWQpojhV9LufQtuyEq5ui1o4dpC+8DJ56ExlH30WLJak
wJRU0jrNkcRsPE7A5vVqjhDstdi+C5qKQ1q/Mk984Em8B62ojbW60wfppihd/hqEiOiRT4sZIzpi
yrXKmL+o+mlVtDGNHP7PXTXIOOtlFZK6mLKvX1NwKmS+5cR111iNrV9X1qg4/aBXFYjnrUBrrKK0
sDQAqfRoFNL0npCq8oYleD02W7+QLZxBbdYeVcC4iuhHIkM9STvZ2qvyVSHjNTicFbAnRfa6eGJy
QW62AHFmV4Cj7fBQLsnGtCFulS7NvenSrmJ5DSN+kN3y+vxjDY4xccoQkbtWQqjNvz3U4AqQlv3s
zmefw9oAklq3s/pjdArnFI4n27m2WJ0y1S1lBoBE0NciohFBLyREyQXD1L2G6syD0W9H+ls2kAJz
fZVacJwFVxy6L8b1ZGcwalS7lcUVfZRFBnBUfG0Ta4lztUZ9ny9tERLb10g31xVTVq9dvK1eklGv
fbbSa51qdL1La1yTMnJqs95xfztfxAHGGACgyGg4OekRdJ9EhjHC6OuHI88xK5XEhgZL+50zRKVR
Xu4+qO3PLgHt2m399YiyC4YytwFpTnPIFhlYotZgca44b86TpJJ+NIZPIw+DMhsc5pddWwcV1pdP
RUPoW8H33OYkIjxL6axr1FdMbwLFpFKEVaLz1mpKrjFM0IvtGSfNW3BfpuOLgKo1wprJ2bteGoYc
cRCbPUd/doAABj8mQOTTS+H9ehnPunY7xzGa/m305b55KlF3zxDZwZsfviBsqoO5XA4jpAIZoYgP
+fBG26D7JBlk1uALH+kJdRNSyGmcbA7brPecCk9iNG6J0/Ein1GHNg/rObPOUPSQ2SozoB9pYtQx
xqAquFKxhAY/gG6snzsDceQ0vWuQ42m+BM4HecdONvSUs5L4LeO7zEgV0SyTN+qN3/v+rcO6+hmk
Yp/hRhdHPkcmEAmI6sEjyolI676AN8Rf4s7Y8dYXNtnfg2dM3NP7X0rM1BQIG6mqF3ZYG8isBFxk
fDUw3w7mmd2Fsdlk70yeL/neoaR42H+RaN+Km8QDMAgy6xPXksXj39OaigcI2NZyE0qplLtJBoxU
t1xKjcDRMchLD5ItGI5uxCSD3zwAIFw0YbTlKC4MHfztheimqkMUiYPzxMG6OodaVIi9xKZmlv2f
TpcIFpDyrJy8oIJTPIl9+SmtgDtAY5pkNFebwzY1Ho2EnvIAj8Awy7bO2DCqDvdvgv9G/tFDVSTc
Q9SzL5YkdLlnCfwc2GaofGE7+P9VrZs9P6hHCyvBkfXSflrRvJSxAqlfUlDwZxjgN/e9ub69TV3Z
wcxMpjBdi8valpoqkAdFkSM1oVqRT3QIiGcxTFLgwR6EKlq04ST4dmJAHMEPx8s/OjFq+aMRgVRp
6hcX0tA3pKu+XwOqBYMd6jCFzUfAA+YWamyY5cCm6PQjaaohOYFWfYjVS+kc+zDTyhn98O2GRMv6
xMVLB8Qfk1QlQTgExXz1iYuNgpecQ9KgPCr9QU7qgwnMr77u0rJMNjw/x7wP1GkhxeMqFgrJGiIK
pkB9+SZ1nt8jEyyWex4os3V101IdnQD3emCFya7l1b7VfQWkUXFFUrPMr2+InovNXo+8hTwkxI5f
E5r0gaeFD4rAg1mhmZE3whxfQPYSvNOcCEeV2NANNp7ldYf5EXE/qq67lpMNK1QIrfIaREWzvsD9
Tp/TRUtm9Sc9sqIGupf8y3wVe0RfFdKNPyKEtX2Dkc9YxbxGDgAfmG478qfRilW92Q8kkkd2FttH
Gcyklus+A5R4dzFspG473dpu62np522WZg0XUBIrh7K7Xsy5RuV0Pm+k+c3QjnloUGO+ItiTc6eV
C0CSKYkHQQu3BnSPDo08vSJkhvOXs/XMetO+lkqpntjRseVc5yy42FFg9/xbV9+0UIhErMCE/XY7
wPu1676wefBlQsUV2cMxjTv9160IsuedFlKS/60qBVebHL68sYhk+SJ6U564J/FkyNDKIQI//LVp
Pxx+L3QGgZ0J31faBJDKErUaYeuxzxNLKkBVdksBCs4BDg1Y/r4pqtI3vxfOuOgjvCBa0KHDU8F7
iMnoocUkeMBNHikeSBDNP5e6i+w9kivUhHL1thHyHyWNVINigpHUXShr6dEEJsoCnkur4k4QFzeK
y/DOAdaRE9HACzgeuOORDM5ipqJnzFAOKIflv0Mm2/Ap+awm678UBcPPF56Nvzm0qppkWDj99poa
LEsVKtAl/GgApmwPpX8aFb4kw+r/CvRNmiJkHAKBSo7mhGdqOTZLMaWP6N1cYQ/3hI+XmGO5wSQE
K7jjOBRM6vWShW7roFF5lkmMkGLxlgW/ky/ZKA8Q+G7WzT1T0av9HN/WC3hWmAI1ExliPVonw1NC
/amxboo8EnpUze7Yu8BBxVNEfjB/S7Pk2/m3YvpTUfpVStZQISAybXtg+mlJaHT5zgzOl6gFdC6h
JDYyjGAmERDLPRy1N5EDwrLjfqoIxujJ3hV9JVzmwoaPvqmdlDI8cyRbEm2rbjx8NVpWfRux+tiR
7brBVJ8taizyHZWtdDuTMN9IqCzETG82pP2BYneZvaNdG2oIZtyZMQVRQ47DQNIAEv1Y1i8s01yF
2qQrkVaNdnyFuKqcep7rzxWL92CinodnPPfzljBVuZZnBBPPObMwqNPpl37+3z7GIbbTjw4fTfYY
s3RD+MgQfiiFFbxqtZ5CW3DtneHxx6DRH08ngxtAiu5A/u9nMa/MNmHYTRX6RkAgL+Fh4W3gV8yD
0IR144emvudA/e+6M65VFhmrmYFgyO27zGzvu6GRxixXgBLPRYaf0YuQAYHw0F0bojtbSg94a2Id
gvrDUX7ANvqjUq0wvF08NCJQXN9dX0VcDs/yw5fkoBhhdarNWZHJEYEPe9uTePqjQAWdKlWZ4hdU
uxHE5jLtFoEpkd3sf0t10WcWeA5mDVCdBX+MvTpGMgekRoXhaq4NaFJCO5jKrYbYLrSoDTV9kOkD
boMDK9yW+aGmWsFSXPyLPR5dZTm+YEl1CrN8Wt2vE/hAu6F5jsbPu3cbOCb2UrpTYJzcA6CLRcpI
Ld65bRE6Sf4fz/8L2vtWJtdghk2Z2X/VQhtEjanoq8NAa4keA/msD+Xz9UMbZBLKKkba+m1UIYDl
GeamSEzQ9Xz1T/+9Ts/jpKHCrJCc+b+n9nchbJpaIMLuFXcYKTnUjOGLhC6KsLrm2d40pxtZhj4J
SG/2TWz+QPJm+TQsVJRQwUpYpR/TSZ0Z+l3xp8lDHI5rapFL/cnEPGAcw4f6PIoTaW8QeCw+I/D9
+1mrRWkZ22qMdRZIUtQmGBjAqrc7MqxgV4hLrttqwEGNPRdBNoN2EgW0D5uCPUtHIn1GtANhCtj6
308S2UPQj43Xx2KsKhgrJ54lXI+YtSKUgWn4cQfkfTY/e0WiLRWjKjA667EibpCdkwwK0uVio1bf
/Isy0G4NCpdpxZEExV0si9+nsOxVhI8ve/3J3xqcMLXkxxWuaXysSBSv+4Ova3J1mS64CJoH5A/R
Cdi6mG+83rz+wwesBAKVy7NeEybWvIgE/UxhDmqzAm50KsxHlnrwgHlbmjr97Uz5Wpd6nvFYEsw+
21lp8u6ClA1Y8Lnps6+Wuiupc3gbyRt5zkhIkooiA595J5f7vy1T64VhMnYe28lOj5yyGVFt09bc
hAvzHB/d9/fY2U48/bR54YhARq/JtNGg+NeNoXi/57yKKDd+eKG4h/FvCRqnPLgunPSpMdPQWLvj
/QRyQvdDDBrqIJH1+NIWKmgZy/i1iw7go+ijb1tfARzgC0TGXg5bLU1Tj8/Uei4Zbsmg+ER0ymCT
Wy8lEMjD9EwexNBk84ndZ2iaHxIIUwuN1TenAcylMM3ENV00GfGNiL1gMAJd2ZUqYNcCDYj09KQ3
fHauyBGcCAH7tG0Kr13QXu41c5Cl/GcKZWklldeHzyiz/Ye/VAZHmgbIDEhQNTAn/SkE5h8NL9si
jt2qzsvPsOjc/yRJftp1/VV/yQyCNoZtoJfoscHX+MXARs+g96Ru0vxSyWq+Sz7oZRrR9+sGXR14
6X3qGGK40ZRGrRjr/4VTLne9bWCkNb+TRMjQcCHRN2bp/k9vMMyzfTiBz16xIvzmOAIaWGEnj8EV
uQIyhS9e24sBIx3DfzfXSIIAZRkDh7gKH71lhVaLn4u2bxBqvEZ1GksXZ33XCVwt6P/WWdrlOajA
neHHHs6ZvZQcJ7v6SsO6PdTF2D3kV4KqMuSBMbnPkKspYBjHYAkm3WmUZ7aD8F/msIE9jp1Hk+mH
h4r4Z6n83wF01TDVHoEkF5qFl3oX1jbl4qN3DCy6ttr15fSMO8semQmYPQJog8GakB5tDy2vZkl3
eG52wZjRgQelFmEIuoO9QqnTLIAGTC82GyHT5ZPAeEVyL6pZPeXVKXX6lLiqqG5qBO6fK6Vr8ij6
pjn6nDkj3+xghfCWe7MB+YzmKPN4jypjcCUWGDbMBWKvUmX7AGJjR9kFlA9V2mTRJCjxxrHywZPu
SvR/djWDfdHfJdRxYaG/Rc1aoe8K/laQnJWvwqdgq6IBH2GRPHDouDm5RQjn7DPCP+NfDg9SHEjA
ACkxImGIm6ZAc+cEvxD2eLbpwV+8ApM+PBkiRe1U+FeXLY0HrkE6Fdf/52CXAAw4o1P5AfOIYhpq
tvrgAymwHodSBsVLOkELm9UVHvWxF0TwM3XGsKI+bpF3Jd+qgPCDGFXtveFpXmtYAiv85/5Wb+qb
OJtzUcLPIGglnTLlCdKx/YDE3WdxQNZuHeguQrs6dCeoWUB9DOpH7rkCDX3iItX7j+QbSR6oBkz1
CsjGUmtPGpYphFHyzy2I5OxpE2vbl5loG3IjeIIxIg5OlUakB71gvA20RpNKySn8/bI6f8LhgLZi
buOeiB3XP9ZNANazWxLnlSm+ICc3EEyNMeQbqIljdGjyZw3IMTy8+E2DNTXUJIKNHwrv5VOYBS1o
sYERGjLTl/4EoGPrXi8Awd9SSfGkdjTf3svD+i3+EbSA7m6X9s2InY+76C1eUj8jbTW/koXmENXL
QvKshaYt1ZdWElZShXUqGyp2M+s8hrcLOdTuE5+M+J+FZ0Zb99jxktFb6+YgWFkbuBmps0O6sU2U
JwlsRNtcb+KXzgD2QFfEYB9U0x8obKhIzHITGwkDA0+wSxuhBiSOndxYt7o7VOb+khjEY74ExSwa
Y4sHAQn8NDdE85y4TgzibQ0rLBFzTl7kWx0JhPcdaMGL0RZSKidrZebX/gnw6BrOhwie9sPs99xt
kqFMqH/HyYjyX8jVVSm8MvoLFIGhhxcBj14ZnZ2QPSHIoHyPfYmFrkNf7ANMCnbaFU1wQHBj5rw2
bk35oIb13yg8qGz9YCrbX8UV37PasyueQmt8MbIQm8zwJLHUAgxQ3kEcLg7BRopJT0Pv4cFeoBH4
oExAhn1mJRgP/sMnkfxahgwWFrBsDsBvNJFdtdki+miCOUD5Lfmip6UvHL1Kxc/WvQvmnTEn7c+9
vvfTG1i7mk35VHRBbNhIzLuLN/fgwg3S/mqJqV9dAL+nN0QJuDnXNWr4wJf6tMD9UW17MNJZXH1G
s1AAJb9S+kEH7k2Q0X0KWVirT2VtiwwcWfxSr38ETP3bDDZrPDUk2pmaMkVgd10ppP3xCrTOHZfQ
vZHM/0dgbsKZAQemzztLchF8oWFhEB6p6G8W7ia+uaRfHJGeNgqm71U8RLqPa3Fvu08Jai9cdJx2
t6MCNcyWpBbYZF8smy7VX2uEulgCvSM1QYNPCzlMy5aW/qvHYr5ZcfJQGmtMCnyR5OTC1SOAYmm5
pO4WUXFe3Pm3WyJoewn5UaadW2y1JYuxMfw4axGR1YFvJadO2TDr9uCaiwXk7J6vXAt3I9V95e6o
wSXKdiv3t4ITPkGIQBfOjUt0DpxzwxxOVpHvt41G/x+MMyYFgYu7qUvJOEHPPdc61EZbJrj4Kjbn
Bg1N/0lC+uz9E72CbEB3F1nZiBqxyMEJIBnz9/9/kSOMG18XbwoVf/fRTS7JgXEGkX0zQufaPl64
LxXR1ypXxz1EXIroOpDReBBPvd8MRAWYVmO4c6EkvMqPEH2ch0zIFN/rynJCATbLFlwpcKvPZBZt
4r4E9AbwOZf2Ainp+tVfzHC9lbL7DIGgzo1l/pizqlrwiJyTVMlSfGuQsyCvD+4khcD4+RrbzsU5
kjfiaFCHJ435+9hXoHpybzNFGrRqrQYDPRMPhR56lfh5Cl+Lbb8V1CAiOx59mrYe2JN1FLLbILh4
rWZU2l6qzN6usB0Qe+0PafZ3x6dMA2QCgSrAHttn8bTyYNrLx+Zu/gXFY91uVPSNHLC6SnEAtHpB
VOyxYh2211Yw0NaKcj5bzpo77Zs8LTlLu518T/OvWttwyXCeP36jVHnZEGZVQe1zweI7jwxkcncg
Yp20Hcg3vnQH/YeG1ZQwSo4uOgK6USagcezLXETK4+lHRLiTLeQx3MOyvZ2cdYvJqH7Trogh6b9g
odTk/T0ix1hKD+A5mIkCYq7ISXnKjWMsolkY5vrPvJSk+inMCbqp5wjn0SKrXuMc8MhN4s/qXdTD
Dt2GxJVItqPwQ8OQnmCTW0SCtkjxalr9Mq3p4tXgMg95nS637JNmBaMctaqsP2BjsSE5OrgXRco6
Ptc72GJXZP4Rgc4hgel3Qa75V4WiUTogqopDm1qLVwzTO6q8ZZ4uf2+9zrKLM9NxOND8+bp4ZtPf
IEACdO4FdxkaJQYBcFAA1kdqugZUukNPEydmCH6FaPTODG72D8vC3loJ+SetvKbj1/AJ2XwYXY9h
8JWk+62JOa9cE/v0X1/2gWA6oktc4RB6putgu3meiCryz3ughxYJiVK3r7h9JDDL9GhAjJOFEOsk
9bf9J46geA5KLGcaYWlNeb2+1xLB+KhK8lbMUsWJZmc5J1BGi2I1cY7qKmBviqSrCIpjVnWN2kg+
Y/61P9dhSOeLbHzEOFyxeDv+XnH3T437ow1d/CAz/Kaq4+no1KwzQExUn8R5gGqBJ3DKcdBAW5/D
IaNEDTQhcuXPQX98QCdItTC3zF8x7h02MF6hDzoKLB/NheANMknB2v6o63YQaV/Q0QVW/DtxsKpP
D7gLzKCHa1CLCJTbKC7oVAlg125JtYRLiEySifVChuSYaWgkvXQmF4ex6hq2u1dQHuXO1Fj3qY1x
KxdjayWGcArg+/9esIs1DaEw/8w7VuSCcapZZWFsOi8bgHyLzg6IMxWPxXH9YHgn9rgsAGbG1yKF
wysCLON0oyHMhtVhlxTX2nTEoLdjS9LOtbS6Oo04McdWMRJjf0PkZMNMftFDNKpSRaaxYUsbeYDW
/+Xvnxj+ZxZPtcoLXoEDlX5ozBnZZLSgVV8dhde4GQ7DiA7zvrseBZsFjaFZTqiVfM5L71o2xOan
xNvsR99uYICfQJcxmgLQ0nWwabIlcxaEIn0tx15Xq6UJCen6lpiESvyti2bRv3NyJbUfKoLxFKAT
do1U3mg9tHYm8fpKWiOuTtuxYEkQPx45OtmlxE10hKhg3EqKSL8j4W+e8Y3L7v6uIAzHCVb4vIzi
fwVtw1Wxm3cIZay/UEaARAQFEK43FgdoMeMq4tgmy1SbufigB4yWU9y/z8+MhvZDN64rfzoBWV2k
+HJ9mLM0QP77HSB5HFkc8pIRhx/ams3n1mb4SlhSWYvP+YAv40fbExbXhxIt6JOnkHWYF8NzvtEJ
I4A1quGW7taxOrtBRDGMJ64Gc/wFYt2KWy202dU2S8w616Sm+EEcbjoJSMynBjLIrr5GFJKSvknn
NB8IWzpI5JTCW44Dc1f+mEgVGlVhraeKirzITQPMEYd82HKtUp7Dm78dXqirhLfG1kkXZfKikyzJ
kA910MD/0UOkaDN29jlpAoUlvMl5E7EdUKcdwkGtyWfr6ljXpkiJmuE9+DtuTUm1STiwakT6e3mD
ZCHSuO1gof827GScAAoBlTFjVgKgJVizehK+jPE+k4PJ4Qo2AKfwl2VImCUlIDHxqYxgUGrdVpJn
bbmc4jCdhkhSpQ8RBDNoMi4BcCan30ynVX8gni4cWt+aRlVuU5qh2jRMDkeP4vPs7vLGaFn9pQZ2
YV6ZBcCfz50IwmzXGGAbJoCANBsg34GLoePf1UgHjaRt+glgaMb4O7y3SGOiccpC5DfYEQvJpGjc
rpl+/mEyHS46oveo3CjG5A1MhcQyS+4oaVB1HoiHs4z3+baw3YZ2V2vIsOyrYkr7q96TpLAbYjxs
Apx9M7gTPlLUavoHjhvCNk8QDb5qvR0uJtrcfHr8ntiTRG4XBZiAxEWPN0rg62kGRvv8Ld7Sh8ni
PCcBuBQyyKEhBpKChtLH6CVpDFPBUJkNYW0ZfCiYA9W0McsnDp4Mt40FT/7lKpGqedFY1DGo4Is1
4BnoNgv9DKugR2cul+KFmM4l/8zCRAyorq5GjWa8r88KE927oVEED9WpGKAgmKr0f9t2Q+UtQd3Q
fZiZb5JfVbCl8kHaSVGh2DCQHr3LnMUoHM4SxgvBMIJAYNvGF5p4iGGqP5Hql1aLKyD921F3KM1Z
al7rzRrkhesvao6ejvFmzq+vg3LmHoCmP3Apn33OrFQTzl+5olrUe0jLt+kLevcAsrq7Wv0XpvOk
8KdPzZEAqqCWwNGsl2rQif9KMEgps3OsVx8sgeutzAlThIaWFJg3mBjKVILKs9Abp01oBnnKwyE6
BOMc9yx6sKZwUGeCff2aTY8YcUrPbQO+doLWlOsDyvATYv0Ut5Zz/dOvujqPAIq9BNdxC1ka4D4A
eBuNnO6hO2HUKYn6BHFUBS9R7zOEayrvLe4Fx1YwRwFJe+QyCmy6w2fXUFvnOTh1E9MHY/aLMaeN
zUWxc9FA0QBTVclxU74+ewCJ633+CCOPIksv30DrTbhJihA280CqJaXZpEKRVN544Hb6t5EGlRcv
tzmRYDrBTOwS9TtQka5YDfYTS05w/4EX1v6OLXGy9G8VKKcJcYg2CK3wj3f4PqhRDyfhqQz6Nv0K
pM8mYw6+7htU/ZsgIe00Qk5L/2h4PsVfYqBeMe5nrPqSuyYj7PQE/wzNc+QYbRsAQwb0znE+CRE2
RpgOqk53UCMjTbjm+5tgyjHBsx+WeCCtS/L2nJ9tNeX80Lk/clK0isl1B2l7UO8iO4RYOqT5RIly
pIiGBqtlXUyMKXxHWBQuSD18toCF9jnZxudNj1INT00hyDdSvOlzh+VWijV+5ERfpHoeYTDcPS9I
hM1xlzPqUNM+M9YfU/hg6uj0V2enifp/yA6lHP21In5ydvu+5CVB++Ts2hKsN8SSdoTLzMMkZ7ax
+YwNLzTCGqDd8Xbd66AhuScKkWJ7I7XZ5bsiUIO7uoV4P3Gci7slSYNXdzwFMgmmtgj09rkaPx9A
3K4keiSixJYa+gehCZ6vwziBfy7QC9mgdylq5N0e/MGR1J28COKESGtAklh3sif5NCMZk/axAAxc
iuIAhK/cJSWLe+5cQ+eMve6hx7w1UnpMtp2bCx79EhuatYmIvJ3OXTcDEe0pGCf9otuc59QB1bN2
XKdGVPnPzEIOWUc788aP9o/3iwRTV/DZTpQS25eZn+BkWT4sAmbqvokIrtcx/3sOPDDBF5uQc0Ch
flCRfQPXtFqwJ5Hychd92Gr5Gm1IKwoF63AR0WcOYy6Mgq2nkb63NVtjL0366h1zDAnR9KqQnRHD
V623hfKsbtopR07T+t/fM4cEjahBB0b0EGzeB3aYQBqgeeE5ZEkOmP5JEQtmOaRDJIFrKLOWrogn
8XLWOizQbACuw0XkwBZq3eP7tjd5Mq1XR85cO2NI9AYyeo3yeww+npvmmf87wQDjOIp7R4gzogwp
cklFIeXttJ6H6T6HPZmj81JRY8qilDEDL9QS8/1B3Ap48TltgViA5EoGN7Yepm95gL7fSvemheTI
mQYOYbQ79i3TFLjBKDAgzmbFUAXj4Gft0Iv9YNB4PwFPafrtRz1pk3DrP/SvzR2vcX7EewCS/aUd
HLsLYif8UsKFWDPGswVtepIq9xCPn6gXg21ueR5KEUZJkClIY/79qNrSpIv0HSnTKLkyxTUNpORR
5OM5hdUt7jhC+M8D22aZ0XSw82Rmbb8b1nhtmGzJKWbOCgeAuxEiNZbLHhJy+17h3KmzRL7KHJj+
T40rwBKwBmd47c4eDAlVwlsHzgEAWOKCE69AGXhnqmdVrfjTPw9JX/1QASYp6F/NrU3ObKV65aSG
o7hxqVfYRDfYXDBmWsR9xVKZ0eqCLVxpnN9ZnJzUqVUh1QCKhQlVthX5db6Dr5F7mwccsC2324fj
RQL9KFpC65mGwgrOIufyeRgGzMSgfNjzondkWKCrbUBLZFGrwUe3NUaIFspiQN7DlCWBCJIBiK1+
EudS8SZ8yOfrbTdc+cOTANfJfAN2z8mXx8EDcbSUhnlozQ7M8nFvLFKtXcxvjDQvzBubwIJ2ZVQD
yp+LSdUnOQXn11w41S3Gxj0jHqv3cCjc+SP8CIk2McGH6uMCyYTW8NyEham4spUFg/BPDmxTGExY
2hyHDGfMUaoECYLP3jF4Jf0N4XWGxfWVvqmfxIZqJAATD5TFuUG+ttTwiJJXIp8w+EhZukq7q6mZ
CUMDq1L394t07bCdk9tFHhaZQmubfGLdcg42b4A5nRk0kBAIK5EOG5jiIUhyH8ohV3gXWy+s8yuM
PHkJyrGRNq1zB3yQFfZhQrJsa2DFaXWJvHsbuYBeZgZ9KfNC22U6lX4ztdKTLnVcvR2peLVJOIA6
AxfH0rifP59tLFVa1aGmOy3XUhLZgTBptb+xHqNWJYAZacrh1TTRGrQL3nTxwaPMhSuX9hzNgWD1
ECo4Qd9cAWi2p+vR5DoHNmW4DPctzpYCAxs8bcZn6v94d28EkuwOMuXixeox5Rt3jZPJDlrf9xiJ
Ds07Gdsc4uQj6OMZevIIsSO6RmDzVpdEymoeZMp/j0s2pT0iw2Bvh80BRCJML14sP/ChcpY9JkSH
tQ+RHlSvl3Xn8a5rrlBmvGizkShcwis5+aRWVX/RuJqtNtoxremdq4DfWqMAmQN42/aNzV0Vyal0
Eah9g3Mtg2UJ5NZIl2T8od3F9pLD9ZuUxrZhVGu0tuwrCOxzHhtwBKyXnY70aHLU7adFLMSuRznQ
TEf/HkwqOMeKVeFUfj6ViInJRyXYBLW7XBTPXEsBsScMowwwjTRHMojY1btz4ZCZ6VZx+RsnXZrK
0TCdEixM0Rq5Ts5x+HHYnRM2vhJhCLm10gEEP7ALYoyHCrF39KNNiOu1G3kVutcnawyz0DccxmPr
tyPFjrnY+wZO0NdSxbXY8ruR5Ec0JJqVjY9HTswDZWgAkeqVe1O59OIC9h0sYk4tDmNeLVylc/Y2
gQSeq+dlHUqcpMfokkETfb8jSHo6F+FJT0vR2YevYyLuDPFEO72+iI0yhSAHeQzOWdLNnVItfI//
wQXiAJQYVRHpCerpdAZPQeZy+Zooz1F9fZTqwbET/SSb//wJhrHdM6VSQfCZeHXOOsB51oxeAsH0
E8vuFIYhefBO+wVyi3vQ/9YpXaHvuV3+aOCKxeWSPLWQPQloDOfnKyf7vGM6C+WnvFX/m/cR0PYE
4LoXPfWtGzjOv97wRxgVJ4511+m29Sa4ceAMeowPXk5eKBIYWGMOwiD0IvmC4u4K8LacEgX+4w4c
/te+VQxlkXGtjPZ3ff0RPcPh2saDJQ8K7a98tCODRWweb9jg3cnBxDKJD3fH8xZUhWhYoVSCEl40
MgTi4OKi8oe7ShF1P1EwtHYusAIwjSaNQIuowYl2xthu2Gai5eSXE24Rs6CC1SLYTiAttSTXMcdM
rqHVDjFhZHc1xkGZkxqRnPwkWC2I2CjL5RIlMTVnqc3H4gwi6lQ1n3L7fwKsDkrUgyDCfTYTZ58v
jLFcjt+d+iHs/R0WiFAf9IdBRFBnAp4e3gbQWGhrsWPyOaYanXfnfuuiwRwp2/M2E158fFtGdf9z
kj4FIRRVlUxIZ2lQI+ym7X+KxwY6ZWff8YIbF0wMrQAYJY3Pv/nSatx2RXtp9m8VzMIwB3iMrZY6
UIIU9/8npPQenk0oUzciCmUjHaIuYuErxHxRsRj9jgH+aeZfbHeviOWk+547EwD+4fsZr1YKh4G7
4+ixCfSDhkuAL98zYR0ZZ5VJcwCUfzYna7Jg2TM3NgwM6nrJzcPpL5QOHOq/TrvhW7yJY1Oj/HAT
5wlDYLRWbp/1Y8iiuwMma+5+6xk/vDcBY0Hd5g5u9F+mA0bf9mpISa0kPJHnnQUD9mG8XsRac0aP
9kC8hsUVsR3NjNWo5UHTqce4Y/rG2lI75teM3C3q7JUAaGcDCnEvhowCfFUaisk7MKorUJ8UazRK
gnzqFr5NxVmqW0AOURDBhULQ1LegAh7VS+Eoid3A0X3yPM1a9Xf4nNbAjTwhBTsc4Z+qM+gV6kYT
Jlf6FTUCdvQaCNELPIGaQLz/2lVXglUPEXonZ1kFRDw4WlOU4uqBsGTRV9ZnSsBD1ifJmwC4TP+c
cVIfULqDIZ0YGYOHcCkpOP05CTFHtwPmc6hEjDr7Xg87hH/r2X+mMvhX9guyVWQVQm+6kDwpkq/S
x0ZAzPOgpo2B09ZYdpn4w5wgoXuBno2u4x5Hy5+YMUuXe1OLj9XtDlKh3UQ5z/0zF6ugbMs62tAf
S/hxr8J8Q61NB5p5hC90zHhFzLvZnlWwx6EGYEId0D4UIJTni9EJYVJYeYn1IHHxOSTCZwUbORak
p+nIx9hLW5meahbRxO7wK4jJ3osUOECQfui/aqV+QHW5sr4LDsnwGKRdTe613rJWRrx5EnNWO477
2O1M61uNe2kHFG5vCTS1W+dCcS1kz66VLqlNObT7AQMYSonwcYDH/XxylJt2IxLAg0hhNYA0Ybf+
Vl1WEgPH6vvWLZSlUZvR6kXrc7e1+aDIrbneq+1ZulrP+q2Felh6pGgGJoVrNLyDonTKs+6LzlT4
OmBMZ0aCuUGYUFxkZ5YZaGBqXPzW8iOc4pPjAkGkenIbEDSKHWGAFomWp9ZzVsSnd9XuF1HxpUC3
mXULXY8mcVBT06s6rSJ57F24Bwk9wgJTGjBRm8iXq8AuxOEL/c1r5yJmftJS+fJwejuX5TCkoyj7
8Alf0UKSHsZ5+s/baUn5kbSZUEW/mJ/0rY3CJflAmU8mP618s0Ba3OIGrvaah6rYy9n1I1kF977p
jD4hwNHEtCCtkwiCUEpMmL1pPrr+qZxYN4Zk/Wy+lO7Vl5unZo90e+YrZK4cv/3LimKlZEiBUJiz
YgGj4kvNLR9Es1n47zKCt1rxpKIkQ/LmiSUIJdMr2wUga8h6awIZ1rh0KaOAOD/m+5Lx+c7+Coqn
sHqcAV5PYXgS1UcdrcYms7SKbKd3A09pwyfxbJdZnqXX6XM21eQtktUqQly8Jy5/+25JlEY4B4c4
c2ajG2lMsjPo4A1j9h0a99h/E7rKocFzSHHaYFo6RBS8UKzfGRZCeChOun0WohSCrSG7ehGz9aCZ
wTe8xSQ1ixlTvIMIcsifd4NBxj7V0RaYZCwrJ+NoIhOTMva08hL++87js5ARM2DFLgQtmqW4SNoa
M1DUBPpiWgXAoRkNfYhmkTNJopsooe1GeOPOEuDjANe3x5KRBFJiOk/E7SfLGSQOunMicjjGFu7S
0wEYkeC3Z0tAb1h87jTPhrDLvzpcSL2JEiksbuDIKABVmVdf3ZkS0R+4wzJCbiYqFLKwAA7ZFIzm
2lVITE8tdEl+c44tbnpfMQsNVP356m+gl+mkkT8z+usAHFZu7OI/Oo3NsVBWr1o80iBz8GG7SYO6
vHk2IJphvN6/l7aLb6hipKc2/Ayfoeb8AfXN7ce6gXtrgjWpi5GwE8zUEWXx5p+mccbU5lyayeh4
WN++GvgjlHzIK7snTKug4t85OeWF2bUo3Sps6hhvLe3QEu+dIlzs5K34a6CWtoYfvmBid3MEMMPd
adamKw0Td9xQeiQ3GH5Rungkx0+FEcuddLjR53XRvspAgjUw3SRmSc9DE6vptydG7P7nUtPxkHth
y6x6P/hwHe0fjra3RIoeuQ+tk/ximBTUp7ufIR/ApszOB+ipEgpHLvBE7t0sqHI23VCeJ9dL0iVR
NTMd+iLA9Gm8N/reViuKXqkmsxKi8oYYzS9uvs1CUaoqhR/01QHPzn/YzsJ8gi+dONKSpDKVj4tX
RJ87m+xJIkg6B1F0ksOehva40LlK3FuqzT/BrpX9v1pXe/R/K6zOhr15nO8tgr2shBBiZYh7aYBX
w11jJd/aLkq4OJNMyRS0L8MQLe/h85neHSKwEmK/TWHPUxFxoALzBrdfdF/J9CU7h0xxLTkF3KgY
SvOI3jwmEVOFcuuQV2rNBUXXvqYHQxEVCr/qRcN1gYUNAuVxe1bldWdy9/WFXCl7D5U8kj3I3BoD
ISMGev2YDCXZl49wsFOtJZ71YjKP8dxjKWlteWpl7KTW8NzgNvt/wdDed/XavVBtWTLpSMIIUCY7
Qk3Xpfmz7IXSfNZP3gDa2IVTRrg5PG3yKYHCl06mIXL9WAHWRmmDLfDKAV/A5XBf0ZlxuoAxNRem
AMaITXQM1qaluC1O2Zm7DItfyJbX27bxDL227Ue/+AW0GykldGUlzlOLotzX1WoK+gDfClt28yy0
kEmNnuTtkr5kvTrtT2gL/c30iFfAhkW/KsDPLMCrhonCCUL05hXNZb92r2ETckhNGEGiJI4//2xh
uY5VTzpxyrQHeorhgr8ivAoi7vyhsCsBPrETLVUyEszDEdgTU6J+2fOTekqrC3uJc6FUCaFAm1Wa
sKQ6212EN4WuU+Gao605TWm3fgSjQTMPcFHENzD0KmhFLHXvnTDXmuPxGM8ywvGNOBz/nFqZ3mgW
+guDqzBgIE9T9UfW27Imtwum3p50Fq0FWDhkdcpzK/qi9yGfCxE0BzUtNuHE/w4dmAnUOFSxy5ZL
vkZapjnW+NynJZuU207hgGhkMcVXtXBbdSrxtIcKkYq4FtMv6Ciwg7mjI+ZCj2lpCG+MPSspULwO
xm3y/Ky6Ir0Gdx2rZRg85Sby4aCPsuACYr16dZWaxOaKjw0NUByTnr/tNf8tniE9DH4gujj1Oe/S
bnDLlUk+PIKgBAqvwdySyeD1Y8FuAeFT6zbCh0736VK16KV/6ZjMQ3rDaD6RmDfZXBBsoSbWtu0J
PUAiHF/iVWQ/B5qwiV+1WUUHYk1+gNoMezGd7WvJ0xbzFqcfKpF8PjGSir7ZoXt3hRgjvjuwP6eI
Ca6LdgOXF08is+9ywfBRzu8qGthOWzyasV5i67H+a0vNoihMGThQq+1M1SzyCNSNE5TlJ+CgLEDO
2KKwvKPEFxt3tqIalYRUHOGaPsbaGzrgAQOSVYC8j3H3+awDBY7PJjpJ8/SnBhkyjHPyLtfcZaRq
qDaC2ZYxsK9FfsmKTaPvftc7b0eaZYe1QiuMflkUL4c4tFabUFrtSlV78fHq0u8AWUBtvbcAt4OE
7IrT122vCufHFAjZD4Lr7nrygo1/AdRMJoAoQ4cR0FzQk9bulWJW/mX8n08KYYBvuim48f6cNyul
2fjRkdWAddz+tP+b/6XAwriSnNN2bAliusavI3HAeB8Z+wHfjM0lrniqVaBu2jsOOl9W+fKlw5Lq
3sFl9AcVNS7rWi3dC0nZecvNkfeJsDwMFCbGDbFHFDRDOwHiKPlRsxvd3doqwbxKWLa1Qdv5e29c
4VORzImDmo0hPRKphKKlnGC76s0GIRVYH7EuI8Hq2e64QK4pynKzPUQ5mC+py/7dMlN7QsERc7zE
z97+5VAJIxlGiTb+X55Px21XdUq+mQv4sCdTqE+zwRhApWQvE6qPVhiu6U0hYCa3Ta+rvoEWtyO7
RSrTiQCchjFvkuSS/AgDVFC1GNhaP5smTK6xvJyzS8ajA29y8VrVKaYSGzBXwjtDKuFC7zfxpMlA
GTQX7oIe0VoAcV7GXgtWg7JVtj8cwWh5oMnaKkY7B1bydh0vvesOAhsRsVx0Gk0fApMZShaGSE63
WP4eXT3L7qr12vNZ0VcblCSPG91O7vJS9fjYgfXNTXrsfyLa48vw+31YvFyONBMYbTXV7azZdIF1
foh1IfnghLjDghJKm+OLj00nrbwuu/F0iQ4gxqzl+wfzjT7Rx6wDsv60N406+UydqLCHph+QHhrZ
TXosI0koiirriNbYvMvYnjLPRfWD0nmxiWnoHn5O7IDNRAJNQwub9fdsAEJGjo94GhVNncIxradF
WfSBHKPrhI11Q09Xc1MSiW1VDnb6btUSkJkpGl6leeiG208T3p1n8G7q2Aa7NUIcAe2XEMb94bLy
K/MLidhGFdTsMg4BOQzOFRWREaqxFVZUQrttatrZskImDhmMwaALZmMSjyFZQSYDKRjUorgZk2Ke
uTtUS9l6fecdnrrXshbS2FSyiONPv0927aJNtqwwXFVfsx02j6Ga6qYFJgqz5c6Clk0Jf2d+1Ler
Q57nYwyAwJ1Sb+7i0IMz7i26DC7y9d1RPiv0C/zyDqmnsa7kCgxGo/MzOewl+OsWkj9eP5luL7C3
Cdwq4Z0L2M6vCEVn4fuZ3RlIpe1zksNDiXH2wfz6X0Wb5ACO/LI/DvlOu0Wm2KGy+wOBXWu+Svre
0FQhqSYboRT/wJHCo7beNA/UXsfU9xzo0dNMnVGI+9pz04OwX8G7l3bkmCq30Mc48MFsich+60sY
PrKjLcAK5Pda1i+EWznHTZreOPCwwdiqoXsaar4fYB9F4v9jq0SG9pU0fuBYg765slx6+eXv2uj4
gpAon94NFFSYSFGOpjsCMbFjfjlwSPiR4n4T7B5ffy1AB9+4W67K5QV6s68w1YO4UeL08XDN3NLo
vC7NSxNzurljMPDeEYlZDW8ng0O5u+fH8GjGmjSo6626sj/s7ebtRhjJ5sGyXtJMxBycRa7erp6t
SspKCMiTcmAX4uB8B27ZsSB9GBpQ1v6aolJJhlPF96EkSBCLyqAFTkhcYFnEVHOdMSyPpu1d46wZ
Qzh989ek+9zsVLL2QzmraPIrEwtSQipfNJDJf33tJqZG7NOExwECdeK4BV+mBSP0WVNoQGUZKxAS
i4djCSbB39UFnztV2vYFh6es8BNM5f0PJfqoR7l5k0mhGtM0euxPA6xOCgmirV52ryamHUEzwqWw
W4XiFwtiZCKUzkXjMOaCHLsWgFAZA7/fQjV2m59JRIVMSaIIBXj99KjviJZL4v5/GgrKoxbDRz8A
7u2QRTIPc1YQvTuEUijxRTbcArXLL6tDZ76DUU3mLBIR/2xschzbrTo0IUMiHFBz5rDKOoJJAoax
Ge8jfPMdmTfMx+V34MDRxnPi3Pyz/HahgZQR3kMxKOahAZX59HhPobrtmiU20cTRD/NKV6IgbC4k
/XfiLIuLsn7pDkKkJ24adbj/F/c5apsvURIkCU2zbLLW469wp7Cja0zmxj54t6Cpy0+u1jACASlE
w1q3gde7sAzXGgFFrWQ/5so4iSE1hVp5kVeFM9WTS29FfYAF6xZKPqFAYv/4O6H4GwDu8W6TjNvu
e9XhdOmt877kKaYtLhRDXX4VOJb2YpOH/GM5QqOHLU1nzapEJYVR845cgOeA6751RupgQ3bKyTte
qclb3YjKgGTrGT8MuC86zwzSnPUItr8u0iVrnVvI4UCfNb4wi8AziRr/PuqcrjMXzDpEA1scgpUU
QAF7GMKdshd02WGBS2NljSp5KH3MZcr1CRiZRKc/oEhh5pnTUULsF3jbPQk1XUqZZU8/PaRGZAKr
8FyRdxRS2JqOJbGigxH6tRC4CC1a5u96ZOzu8hs90vwyeUlerIM8ymWsqYMegCzOKdqjClLzilnS
6gJenMA/fiauYXlSq4oAzcxTPDX+h4LN//U3bDoEyv0v1g06EafRyQOIGoSiTGvIQFV0a5+i34Gm
d9OikxFDRiCZKp4uwB60Wm3jd6OGgzu0uvr5EPS4eSbAS69OAvWpDk/2xjQlOWXX2/D5q6MPXa0/
4A/qelHz2rZYOyCMujYo75CB2Ptk5O5cFLKjNbIpkJCSya3NswptL/BCBr3iKFn0V+q8vvlsxyeh
LIZ5o3B3IsoL2N37Sc6O0xjXLVdSUzWsXhiehcx6OOEjUS0Tz1m/HjWRFDHWS+wWBowbdcnp58nd
k6RtnF17jJuUSYVGaHlM9I6Vw84eTUjqNF1M+XBX3/Qsp/rS6N34ZcV9mwHKrB2F5hVBdUNNb7oi
k5eGz0whluhs7TUtMuQysIjzYdmG/zdAunAGZwEz0uDD0X4qtYlm7BknZbHtAyHgF5kvy418Nz7i
A+oRXCITRbWyEell7yONohB45apl4czfZkQRiEAqoPYc6ysoQJaJNbvZTH9rtbR31JlDe7T1jvh2
K681tE76HW3JFvsP0ZKlZI7ZzjA2BEoCZEwSz/4tw2zzgDm6ya2UxXm/ZZLylFq+eWvXKs3NEFn7
Atz5HyB/7/j8lj1HnzeoPB9pixU4TIAXwC0Ge/BAMWulBBB4cYxiaqFyVX8ISDU0hHqJdZn/j3rz
8t5UUAcAX+6f4cu0mi62buZ/1NsRABw3VRJJVi85XIgvRQARnPp/qEl7FBipLPVIQW0jjLLRFgGo
h0o1/qxNYzTusYc5WmOmMiqI8hoj+WwVWWUZpAnjTFmUASBJqFcVttrF6pUMMyoqN+Iv//FztiAt
n2YxK3yvjblpW+1eGxhdA26rT3juiDoBCkKvxT9/uMKExVkMFSU+eFWotmR/cfNjowHXoUllvt6j
9IX62MS4kvG8VchS8ztAGgVrGNWPsOyuWReqzASFB5ywu0wPe5qbkVjVNEUk/opuIs0WXkYBUaEr
jcES5w2AD1iZs8S1v0L+blza1IpxY83SsAylPfh4B5g0Dc3NNuZz7LmnOQGeZ1CYSN/xbcmYiv5g
7yAKD7fP6FpTGDECtvAvCcU0nFRb/G2jUvvi5e7sZW9Ndeq5dBo9TbZAtiN6UavN6PqQ205fbszL
8DYGjbRSaNajIpZCM2Yd6INenoRv0PJn2UkQWEb/VSV1Ro+MzR68zv1uojA2azsJF6LFxVQCDWlZ
tIZlIuYBQ0pO+LeO6PUNtEq/faKmBvKggF7cJAA8/wRSGSBL0jPbcYa0J6xCrFiKlHsd7eqgLXdT
3uiAgq/SFjuOLEbLvbSVLxuIOIrzsGSGYxDNJ5dphrxOCdE6V23ByJw3Xo2mm/aB2MHSPMV3xK76
7/Lv8FgGjispIXunL8GbawvBt2wOHrFD0tfU0MNoTuccM+B5QIr9eL52JpjFipT1nmEpTelVMbPC
I8SaopD/ERVfj4+U7WvTZUElMtkaq99jx9sF4ntyQ+EjxoshDW3OlzqCXnqrgvXfV/jTVG9PrSQ6
jtiAbG+dtbJSXpQ7LZppBCYiC+rwryhkvCp2GbnG1LP8yw6paqWNPmMCVmaqraiSHzHhlcyT7kM2
DRzXYIVcbXZeFvQxajhxpvTDqGEzZkfFKFaNoFti35bO8M4SN8yV9PwgjywHPPnVx7CrQbfTzUrT
HGfhd6oTa/B/sO1/mx1bNPtPKsfF/qLDk1B5zyaRNtq5of/P5Y6/3MxqGrhRDRaT1hFGwqhZxsLL
qWxIf0WtSl3fo+64E/690imTYIwQ5khvJvCRE7xUDmQeOV74Aw9A50KH1zFa2EO/4KDWPv8SWdNV
5CN7ot0Rqvt8zwe4JFQwTWbhUoIXri7lW5iG/Jc5mDdMQqqGtkzHEmaDukHdy/yXS96jjGW5OgUc
D2/vFZvE3pCZ6Kk5PxUj0ujsrfmSCcxBL5rnimSOS0VgJqdekMk/qqo+b0htgXPW2UekbA5qCIT1
8qw/WBZ4g60MD/IHlaFMeXi0w6UYWd6EiwKWdIZ8Q351vtDGAUNiUyiKWE1rrcyIk4fRguaT+61k
nKI6mUxoHW/tCR6qoJSuoCcTQiALvMLZG00kehBaBcH+U8R67fmuP8L4PNoj873QjNlrHlG4RgYe
PFivf7zO+uuF2yMDpSpzuC+yP1rkWa1KcDRCVxpNAD+EPff4ZpQ15xFB1g9FG73ooJaa/TPFiuTr
tHujMOiGA/o0ksAKL0/cAER2CsQku7pX12Tb3b2xrCVFqFbEwHmGRKS6tH3fdkm2sjFHyHA8bgCo
oMRhSiZ0zucH/jyVxzlkBw7lPXpLur7Rj0AOP39sAh6rdyZMwyuR8LUR6nnlUE4giGZmwRjHo0et
tMfGWnwsVBVLNB8YBZAZrcrWULlJITv2X1TYHmMsegQxsG55JZwswwNRXO6PTgfEPfBG15jqtR7O
Ou/fWXnY6qM4bne6O/VBjKhAJmJesC7+DFgB1SpvmSWqXscL+UtldslCZURDupVRbvtUGeVPl/dP
h+uPXpA6xsBEDz2KlRZrLNskXpogeCssMLofdGAyYoaJc+IMIPK5cS6r6YGpjJb5DpqCAau7d2se
fRPeHEapSkKUu/pxoKSzm/WssQL2wh6gCT9MueH0tcDCnsC6sPud4bMT60zGNtT4145bJHhOchbH
MLXrqSCG2di9s0gRncvh5Pru6Ry17yTxt5ar13yDRvD1/XgkFfhQzB4cvENNGxFT369X161rZk5H
a0xKcf61qYg6tIe7V/ULT6mh87HfijYJlf3EA9SpUKV3WyFJao8aj5oetiXYDZPzxR1L3RMTLrmA
5ncWxqzOX8jnh+1ach+hb//7pCnmN+2HxWNPEuTg/cPvtyKWztUI4AnAT7WsbNiIkINqudL4odj3
drkiI1kILO4DRnTfbtAUwrQkzSraY3fN4nyEylJCl3iqM/XVMg6KhDkFZoYSdBwN5dAKUL/U7H5n
ODmGNSMAdPcwkQqudRwbji8r02SaWVnIpjUWU55iA3Oc+lmTd0d2hsyaEhcYbG79RAyQz8gkM4cW
NEG//XEbuAW+w8yzoq3dtvKvAt0pwLP2jNw39La28n6Eu5/BKqFOazA0/NMatx6FXbs6427XFPSU
f1mSbGF2ON9ceryW9fu6cZ3MQFHa4xYU3BYYSWbXgg22DYRY3hj78o0czbGJgdXycx+Lz5Pk5jZI
hvjkxXhUxzQ3y3OESU8GPoIHvXxOO2x1WzAgXIe7F1lttqe7ZDNyKjMuKGs9Jtq34PgnI6x8RHMl
LIuhvmaYyGfRhvAweFcyzRYrDi3Kd/tOyGaOrP7UE02npQvoswQAyI7UpZFaXJxx963cQgFRR9wQ
6eVeeKl0TxPlHpdCunzkIrEfcvtNdVXrBiZTGa4a8eU1wSBLCjUNYJItRunf3L+RX1Zxy7qlgfgg
cCjfQlNj0h+x6NO7Bc0V5QHy+hcqDyEnUcUIzua7bPACxYCaQQ/DPGYZw6I6MSz1LiWrryiq4eaI
H92SVhZX5inDjGQiDrEaOPdL/8ggxvyduACEasFqGnAX1A/JbGohprN9SpdepmFfuhI+nQ1BS2SH
fK9/FF2vxlTZeW7zwclvKP3eF0GfmWobI023awInhmfwyb2cpyyr9ZVDvOAY85Sn9FpjXNbTKJAo
ooGJ70DyapE8akKU/W7ER6c8h1LbcE70ro4A9YSWUvATR6dJB5x8UIePMv5p3R24oz9cafmJb5Lw
0hWxWEpnDnm6M3Fq2FEy31GVhQxmLBZOBdo8OqRt2HvgLvWTHp0Izi2LLQZM34E/ze37pWwTfSFV
QbGUY8cksVWybhl+kmOttAI+NIcRt7KIr6GVNm7Lev+QaJvHGR4Ov+RWlUEZRYF2dujAvPsLQisz
AL/3dO0V80yzIwRc7fh3r2hege0YVBUJMT/D2cTlSwh4Tu7Q6xPO/txpIsGODts7zS1LxNPkR7cU
qSgWbJfzs/d7Fv/fXyyGCN4v5XESb1MQly2+tyPREbS7HGsiywLRxlxQD6mS1j1P+VTauJkTLkm2
0tsJrNYYOV/vvKBKZFuoiaYL6yT1AupFqxCj6dmndLIwVOfnDoSCzWs8z6QjnKewx73oqSdgH5xV
xZ69+18qM0J0RDzSX2v3n1TfB1was+UR4nN3yDIVxoP54HcA5Z9/bshstiCEOmD34qswBDfJE4Cp
KZAXgEkgXiLD2kHufry4yXA/12DR93L9NqC9eL0D+1W6Ft/aDy1NX9eZsWxOnNieqAW3FuLb+d2Q
phWxI24kzqGKG7s7IQLJQvlSLE7yw6ooRnIc4q1ziinbfBjEdsOhJgo8tAJSQQmT9ilGU+m1LXvg
2DM6NM0T8wRmFYTcQrY2Aqv+VNeSGQQedD1FlKh0iwtSMh3cx3psBEz4mKTgE8f9BwwupxhJigi6
mnLSsP31IXeqtO7/zQpgLdnRoJh5IcBbKM/MEVe3LHvf7QiOu5utjweVGwVQYV3lP4SePm8E7cRW
rCHQcs2HSSJ2BualoXeSSe+a7GMldc/SG1zXc+87BO+SjAHzzZUzZ3mfi6unDp9MPAjJ3bb1rjtG
E3gjgRy70P4OMj5aBCjtkVrqDV/OHCNbc1BuB+MApSSCRjL6Lp2pC+MyYIIH/jQxlznwUWxA56BH
ZjTdJulUjtMKI4Ncxg374kqN1g/sMH7tllvbpqzRTF3+pQNMoKq18N4rmGSH+FjK0AuHvkAP5BK1
7ITDgaGngOix8pf8Uf3O+eAWlh9jEx3Ra10enjXT1zfw7cwf5EBQ9hdq0DdHfai0WWiCAyn/EQyB
sSYOvY5DkZsae8G9Pg3xs6bOSZVjhj1xh40PDpVuO9DFxDMQ7OkUpQfp2Nck7vRHH/lElgYJlzcy
U9B+6gxss9AO8vU3o59+OrM65hrqGgUaOZnbL4VGeayKT3Jbw/VfSYKICl4YHPaNqWEm5MIWstpC
vohm8elzuSDMS1Tm9+9MAqOzsAZrpyDtq+FCTw08I87gnZws5Gn0O9UIezHR8zl5xt7uufNHYUe/
y9qf3TpGRCo6mlNRlzW/xgVk2UwvPEJnIwVhQrfF8b3jeJzZ/GawqFP8oKYcgJHVUM0QZU+O7s+G
y6MQm8t36RWprF+cJhhecZUBsUKw7bfZjAaQC6UN1yEY14zQ9FXOZAmj/wHiPAopfrCdQU8Llb61
uBTCFrNjv8BrQ8x36+GL7JK8bnjRBYs1BpZKT1E30/0srnaw3Iq9z5wj2Tq/gAANxaBIzLfttZRa
LjZrQa/GzBbjLsa2eYjeyu28JGnDgQq2MvHGKp6LXCjLfw0aIMiA4BfVwx6NcY6muUX0A7E/xk6r
qmTjlOAboh/oBaWqQvp5pon/EHipcZEUba4GXYDKJHrXHytosM4R/InEyO0KoB5DuMnF/lm4vWFf
hq/e9FcDCGM4KlstNoxSr8zy44l3VpfBT/i4vH/4lar4WEW6baCCpGbDqD0mLJ88/INpw3AOAIve
KH2354gqV2VJzcdRf6X+F/eTM7fQqjZIR0oxkD7SeTtirAQ8jYi4+CX2GVUWBRiWtHF0QnG5wRXe
WkapThq2WiZJUDFtTpxPShVIklwE8e3JsBeZ7GG8T02bN88KrBqdl8uI4caoUNLPjBuDvYENJn+w
ci+u8oRb4glw/Vot/nu5QyILWr44Actg1Jt99ZQEflRBCWBB9N4T9rGDfx23YeRUmYZo6pvNMusC
33tPiiW5GM67I1CVeAJ7kOwxXkDFZlKAeZLXL2bu8Tx4fkZ2ixSxp2vNnLiHzahcG0whXjsxoNrX
WzZOzc+A4CAbZZL0RLuBPCNq2gj21bR1ISphvji5123opRg4YAnFKr9OQcDIs29BrTwUe3Ck8HWX
T2aqipr08P2MiEOhXUlfWBlm2z3jcVrKqIiWmCuxSC67klJnbpX4RDaiO/aBjqiaoOQKY+61UymP
csTBCvi6Iq9GXRvVh9FxDxMw8ADAM9M7+uRWo24nHK56RUzSMPRKVHnEHhmra+QDwt1hAr6sXroe
xzXuhQ+3D0TTaRQcyf5bs0mqGvH61qkO6Rl4MatvP6k6sbIg1Os//sJq5RpnlpxiMgvInbe2++Ca
RHVi0GrbD3hDl3qOYq9KVVFd3cH4I2AcN4WNe4Lrk/tWdtAQKMzfTFYrHlTpcqhXMaFPQaepWk55
n1dqDYq7IXMxsU2M/MQuicoYo+Ti5a88KxDbyKwQ9Lq96AzCoxl/Kws1jDS1TFCSYjIPLZgzWAqN
fMjT1MF4rv6FlW+jF9bhn0F/3V3QgVewOnAiU/r0kZT7UR5ADooSUxsD6j9EKHzc10JgFPSmKDz4
NnTqzFbiOe6vtE+EWCUeOkSv+s3sNJP7pif48L7CoJ58P4mkH2TTzi6lURoZLzM48TeA5L1wTu6r
a56HOTrdN3I+s6Nah57YqUGI585itidHxeVrYlbMs1g7nA85AHEMtXDg0MOoSjB0hQVcXNAGG8uS
SSRLzXLIiTG0axsaApplbn0yojjMtNl25NgjvipRbSyG8BXh4/VR63Op9qJ7xT18hvt1J+89WpKU
T4grXMnSFzyjDg19msy3ydGH0CeZSWJq1fCtBrbfl/ag/9QXa3y26Z+l/B+1n0Jnqj67zTvytHwy
2Dxg5OaizZtouOxO0Y+VJv66/DCUl5zFs4rEX8Ql3EroRCtMq0bbxNgwQy+IYx1zN2/GQNKzFKHL
xJLxeYWiwOUnfGG9FTYML/CvKnYh1l2pwW+L495c3pJXCJo4IZq5wow7pyy4jf8T2TUHZCnyUbiO
8EcLfozT44eV++tc5FQI9tnIEJM6tz/tBLUFpjCZ7fUoQWC0n2IOlu1B1iZLj4M3j55vFfOTW6i+
n/CSMNii7sos4+OW+ytzOf1Y2WlrKL0xKob/7X/8Ie/PPNwTkszr8v1BC64Go+Q7M6SxsZ5VJvJW
9zXYolJTaOZk2/GufQY7XXFZbu3TNRuQHj6IYJ7yRHuOKNBNGDjBS2WvPQEM8Htd0CTAtGTAPXQq
NFAkilchP4OuAHtAdimssaGLm40/jHq4RKwqiKf/molQ2Wgqrf8xDxJyqemvkOdKWDMktmrZqB8H
hKAWB4MvLVQOo4hPRrYNnY+rhscUXdmFfJ0TRT7rail+8/FNHd0XziBE4Y/ppjuIUXNsetaoDtWo
CTycQqCsPwtQfSqU1rurTaSmUf5Wr8ViDMZt4yVHE6PKPHmxVkro+bjADYkIUH7obVe13XbwuwyJ
oatbWTNFJYzRPu4SwVx7S08YD0J4Mvn6j1g7AjCVV4iq+M2Qt3+0oW5Ga7RdeIuQd4+ylbBM4O8m
GDkk65h9J79cV0qvQ4qyj8Qdou+9VTZXLEao06nJkqXBZKxoRFQn7/cbTeIZcapCROEw1DnwvWn3
oN6ZKQH+99/41My/K4B5EpmmMgGFVorfEUqO2rULln66nXdErXWri4f6d5SPDKySPMltNyw7IPE7
72ynkmmmkW/73+paUvII8QoZqcRi8fKkXQEzRVfspXh1yH1RcPA243J2qND+m/O6/wGqeGUbrUJp
w4gv08c2Ktrtd0qBikr5vp6AzS/HIBPY4G/u4IT4C7L/UB6DGKy1QOc8XU6uVG9V6Ro0IJsGaXis
FlwlVDWLo3NSWA03Cly131XfgOT6DlCq94BsorONRv7Nt8Y3qAclcGFg4oufOSaVOByscRdoSMmJ
gIs4bcVBNWK/189MmnLWaglwpXiDkNj2ImuUisQgO2jRihQ/eyDgAvcw8HSX0VkXgTxbeszVQvYn
AthnetlefXmIOCafmlWOw80JUCtuH+jvanZJhIwt+Mv8sv8Fm88T2QlJ5c9fZVtA4h5aofkZH2t7
RtrjGdEYJvzEH2xTrzPYX7lAnCxfbUjZVKH+yir9r/NvkN91am6f1fRTnEUAASJ6M3/xihVY4bqB
98TcP8e2D3TP/ZBbmyq1ASMLQCsl76BORRyvwD+MVWPhXRsQOyb9pbN69voLlmw0KtwaElo6oN62
W6xQXM0vlVC+KfpneAdzLrZUqy58v4+oyb3Ept6STbiL1QpUFZ98EoaiEVaxygsA8Vtfua0B/q9N
OxN7wmUnuhd/czzdGc01qXlUHwhIpLYOjUsFj2sdBLkccWEa5aJZ+5BuUvlsRel7p+64BtqPvE7r
YGX4RmcOciuxpSNjEM6fziCW7R0RbicK2LaoZg7dGJoREMHEfkhPHohmyqZCgnthmRLa5eGXmsca
RAH7wpSpWlhv0Nnzfk6bjXx1a5UDWOkufa3+UxOPwktfTHnncvtyPEs5MwAlsVSIYfhVrOWlqvAP
iFq9z1U71q2Je1Nl+jJACLFPP5hdikoPJbkhgqmQ7tr4TKH/bCN09Gtvqn6AMOC/32l4rZ7XAZQ6
uzmTe+uZqkKzNzz6ziLxHQB9u2ItYuE79G7o1E3IplLroAeSWRC/HgqSCjwE0AsKet+w9+moCwFj
L+09/JvwS6ukJP4O9h2u/hJnhmPTtj12uJ94z4cYrLkIvj56zWKaEkbrtj0VxT8ShM24i3MPMDqj
7FzJWY4Bjn4+hNFa92UcqnPbdyveE7Lz7k7iuW6hfoQ+1aLj8H7TkM6j91v/1vwuosYunt9n4wmo
ItXi7mDjceuQhrV6KLtPzMjSCCkNjTSTgyQFK7WU0ipyInZOS2KQwdo/ra3rGcz8zceEL+72ZUzI
1U/hMs9SoxegHV2oooUHeQWAvjKMS17H9GQ+q9vZrq0E3XtXdYSSdiG275kMhyu1JFP47M9qj1wZ
8petR5zWG7b60rQ9YZRseZcovBWo98HQEd9r73Oc5D/yDZk4BrEJcbpXV1sKBzIEksDi/IzTxjsE
eZC1IcxwRjmdVjqTsSiHj0PWJeQOlMtdoHVlD3aZSMfKStgjBFtEWGgGwiwrnOuRlmgRR0QdvkCc
CkAOCZymHAUclFyOVueFvkTldsrEvbJI6yyEVnByxXpk9khoeWfxSmfo3Rod4CyfOcIbvo9selRP
YFfLGHqJ+X8X55yldfmew2OPJT3X/ckJPLGxuFKQJ1MbVwQFXj4N8Vl9e8FXXVUH3prxsMKCDOM0
YgqIc9BQdqd2rISxuvNbr3zp0uBeYR3JsmoHVCVaFY73TodB4jPWvvzhLVvjyWW4vgqqcp4PfpYy
7wp37ia7STT7F4fL2bkwsX2hugBJ9KuzhdzvQvMNfGEeC7Rmo9O3wTYDV/npN4y9JBfxNg3myS6m
fHeDow21knKnkXzRbpziP0kJLzUJ9gFg9+MHaSrFdZ+c+N3Dck8jo1pbypYiyYIGaIwDJAqV5lCz
46NBwHTAWFJsnlRzO57IiiWwvAwvgGdNkQGgaWCmn3otRdTajNzoO+JISekSiFZBQaU54rXEGY2/
ZI1KclSaK78QRFeJ7tQhv8Zk6uYZIMqqBwg+X1ANwgRPxYUUcrWeW2JpXbVcO39P+MzVVSgrGgLo
HJ4tV+40XOIWuOu14D88jB0jRXhaOxQSYyCUJBaBGGqNbqzjbhg7ja94FtzmiJBrP43i2UcSieUk
NCRNjuFSGYy7Dp4x/Q1K5VPEb0svmdFmXmKWM6gFWvf0oiGV2wAe/Gq9d38rRg2OfKEJ3pE2cUxi
c87OAybEWjwlQjYXoP2JCAXFPgMlJ5Ndi9oy4HSLfvUhX3bnN0ky+pwPPCm8K22yhnpJ9MUYQQMX
0JqoS157tW/3E4jDUoHXav0CMPu2iaPQFXUSE4B/FfXm9XDIka4MF3drTQUcIq1pVY3osPoAKnZt
H4YNtPfZQhFmsFECgcFRMDqU/dlX9vN1RT27EzHaPmkGcs5PMbKxXJKSrjUqYY/BV7XFfBv+ONQP
QaeL2MebnJ8Zcx6e5KDMr2hoVkfRCcknpjdi7C9ilnALcCimALi+K5cG4a7SGyv1GOej2n/bCdz8
8FaHGKGE7WQqkdeiv1h69ubTPRnmXGEJ6A6zqYsuAPlfmc5VhmzpJqq6LdOn7ppi4BGx02qJEdKt
AaVzV+8x0C+1wvCidsFR+idFO+dnpE17M+Bgipxs/0pTBhnC5jQIFPC/OfF50vqStWeGcXwxkdAN
uJUOT/4ZSZy5RYlDvik4h8f96TL6o3lXPWrsbCUVvfL8ZIG36BclGLuRFixwhsaAXdio3zXi0teG
S559o4tOptCqsL7iiyi6i9onIsK0bwP4lT81ig6b/3AULqquWb3DaGbgCxFihgmWL1lfJnN+Dq+1
Iano4bAU8CJFESF+41YDIIjXtoLP06CU54FeHQcC+8drojsXrnNASyhiyHeNxdVNRkQBOowVuxLq
FA7Y4cv8bvgMq0kbENpjIIPj1nTXZ7ppR7cDT9Nf4bTE4IQYKJr4qgw2kD3utQMHf2hrv0O8HDqo
eN3vke99a7PF8/5ySLLMH2zKZ747qOVEjn26mkLfVyfsbS/4WD/YJ/gPiQzqEooYJFmXilGIgCw1
9AOxwOyylvE/6zwbCD4HxZ4hTxkfHm65/Q9NCb6Jb6JZH/+bSojgrGDBn4tg+fD/1TSYBOVKc349
3tfoYqzCBsjNmy57r4A7Av8TpVpYFD/eUcG+KbAU7gwhXjLpFuPY5C91c+U+wdFjKz3AulT5mc7a
O/UkUq95s4Lse7+2Ulj5RvELUR7luiHO+sQdMP0h1Io0plYiNBsRDeq1CTMPxq5IA9qv8Sk8FLht
KzHnwYT2033bgNsq7l4MK5mga4q0aAJsktFOR3s/gRevCSAXGm+gj7waWVBC+IuFSjosJL1w5qV7
vPeEdQug+1doyJ4Lco0dfUQAaC+AnLwP1sfjj2JBb5KPAhvwyihdZ3raJNPfUBnw4BDoqV+LwYGM
v+YOFc3UxIKBCKEYcWXdPIXOI6RNSRiL8FmegebQPR0pdkIzbnSf05T96ROV81wEQu/T/ZuMafOR
V1Uz/EOxJ0OlWECVqVbSXueA/h1IvKBuyOsWGhnQmd81qbpvVw205+yLIp1ucmmZYH6qykADx2b4
VqrQTulT7AvW+ziEAbMt9mi6LaotMyipZihQCLjh+CIfyLBpXLYPLVjYglrb4ZnfYpXZHdDkVB7O
C6Q6mvm6iqsoqqjIz9J5EZuBkbA/SjC+ZiRhsIbnwOv0oNdk26p5vAVsmDT01rudzaA9E5wp3yfW
MfUrQATC39Dzdx0gIwJFcChEk2QIgHRBkPeEKdaUi2Uyv9bkUvyYw/hxqLIyQ/7psXlyQfafyQS0
0yonvBfxXiZtNmRaLHDR1yfA8QoJVIToczGPqGXnFCdIY9/T4Je7OxFXPtO4LOqaXfFrckJNW9/G
aiAAamhy1sxNKTaPG2FMizdyd8LZRT5tXuidROL/ssKpQpQXX+7tOO8GUGr662o/KDC6gYueBd4I
sHErUMZ5x6WWSpPI0d+mOUbxr8NbMBLRzBz7CP7mwlTg8sa+x6+bpqDNXeyV/FvaOmeWHG95qur2
yiSdYR9StKQj+ZUSRpnFri6DEsE0bvKV+VhMehAVaJzb1dwLlCcNcpvXgLPu/fF3g5LXtZ9ILKgj
+QiTwW8D252MrxklKaRWUNqxv6/mz5DH3owW0lw1OwKm3UHiAnouzhC6mgoIXncrvxSyqNy6n34w
G1DdbT9kiV8vDCME29AQ4dUXOU2s3uT6mZ+FVbMjy+yIbxGq0AdF+w8tuyIjKdrnHJOBPss8er6E
3tw+Mv9A9wFJb4xrqebhfGGXQ+jjCaFyDeTxmQ21Nhz+9FiraEp/LuDj+OzJ+J9KxDDcgwA35677
ElaIK132n4H72xUiDNEKuaX/Vb9txJv3eg/TrWKhJw4KzmXvE2fTgD7AQj2PTcoIQfDY3nDB2hcF
f2JlGghdmD7oGVl87cNVo+o00lmzJlWWNlsNb7UHhzAo508geRZQzSCHolW3KDwGiZHbC0EePNmC
SM4ZZcCGbx7hNvMjYnFK2elbC+HUV10VAmG7Jgc5oSc89ofFkS2UfdxVloCXEBqmQ5jcY1pSxHTH
le40PtbbA7TDzS8OeoZ8/MaI1crQnyoZKyNt9FpqfzB3ahscqCqqcGp2zoKXkn754ecNzdNcCRPh
lrlOCtzARQHfaB8vJD+wQAo164qNHri+awC3602DvvPQ3YN0E+7CPtSzfs8KuhhT5upQ+0UTErG1
fFucTgDqgeyuYVgik+MVMbxK2wvtyVL09yZ2AwGsMPEo4iaB+JbKRLCie+KJPyyGSmZssxENYt5i
szv0yI4c4pJOUEl/3s1cVJn3fVgHG7YAlgFcIxWJHIefGku9kUsVXu0JL8fOdDTJYhmShEFSuj0z
cVzBWRQlUQRtNOU2hHzxgraHfCHcjjV5vzmDEpyIRAqmSQdrLvOIiA1E2mbxTubNFwhN/ziMm2cG
0pKqzzwZvDw5iXpcBOwz+cQdIkiyjo6ql7y2u29u1JCMH1MifEGqfY1c7YncI73u4kRX04BVPYcg
jDPKzY53npdsX10YwyBATahkLot96CHjGnLk9p0vQ4fMOM3GCf6GmC29YZK1gdj9AscX7R1KY8ax
pwy3S96Ia/KAwHENylMvAcYnCqyZ39BWvf1kEa6e3f5R0ZtTuUzRtpHe7P0/uCGL4Rky2S1m7zZw
dkj3w3FgjSWMFKKAg83ssqSMwIHstPfR3AuLBNhyYS0aqOYKweiCS2JH3jpfSEv+zj5q61BrakG2
5yjblwB3+PR1tDSFPQXSuO9By8UBO6ZeLxrEFH6Z7SGudd+tfp4kB6uSGX/VSiy8jBptft8atgwk
WIoWRAr7LahQqSgeHsx1R1RHD+29XjJEGCSNJBzNXd2Io6uoznotLItJM7LYCngbizEt9G9KdKoI
LbRZkXYUAdVMLFDK/5wOqAoNvNW2EdOD8D7M4CKg9G7GqCSydRx2JmWNDIHm6aLTygpOKwG4dDAa
fjTL2EXMYQv3X2XzvpcCKzxbdW9Rg5o9c9nxeKNo1riq8S8JM2TsbDdVmiFDvmwK7LQqC/rzAktg
kBt/5bSfCAV4nTGtuIu/n2T0bj3qdPrJ41qCugFstPV4MzH6Yk4c81b16uT9RSerajcsG0Pc0jPU
/OOi7fzhC7qfH+2eovaqFzoyoipNXi3YhzIj8S6jColn579S2KXnIvF7LCkIYVct+5GxetluUrQP
C8dxGOBDHaKv2MYJXsdQZO2CUQITpvsrlLQxoqtDVpmHVKUNUnOo52hH3S/Hl8tnBwL9J4U+Vcqb
DbiBYaT/9bMN2iXRoFIWDh+eIMaIIn4gd291kLDKyB7atexPaiQpAVNh23D85nayecmYEmMM0Bo5
arxIzOYtyPp5LKB4E2YaDsWBe1rGsDrUy4cgdRxYvgeEQHWhTRg1xMkUNFoP+B3avCH+WgMfxmtl
3peC/3Nl7vpYBlgDBb6ce0vghQClZ/G1PW8YuJbm08yxuC331gxOIUU1P+XFJ9Boih9P/Xws3a5l
noO1wnqm6JCHeozjPsp/25bc7vcxkzH8RfsYpFSROzDh0ylZlkdYoWTwc4n0BJMMCf9Dks7R4LxI
CTCJ6KtduH4IwQzj78V+sTZh5tUrHUdGS37lLqHiJ39YqLUueDxDTvPmaVD/FwpRvUxjV/ywMz50
FDhOJvTnoGzO9KIazn4aUTdMa2vNguJ698iwJu4rWXwmFDz0Jyj0fST6OjaW8gBp19GNe/z0kHuw
EBeQwpXRt1LP6FIyFlCrQvAKNIQDj6CssOx4hXztqk/McVUtdicfyH2jyYUxv7b2ZEmHtk+mGXEu
iDHBkpqdKmjZs643BvR/lI81UwuAIV3GBhhQ7RPx2CMT6yZBA4bjckotVBcj+3TuBTFXy4GbjI18
jWrfEdNX4vfA7dGU/9IdZNZaaW98jCKJasUHh1tMdRskf0w/WTxMqwbn22GXijiHQgLi2gOrNbQQ
NKUuzPU4Z9VFKS0Ze4pE/ejeqiTAm3/zp//95W89AfZHjzfHuUMxmFWMYRnnB2ljClijLypbTO+h
QKddQXXqqOj1GYOlnulxvHcAuC+7LCyAqtOBzLuEgVCsaM0GdNoJJc1jhgBtI/R7E1SXqGvfq7ak
wwqbX6chnF3U8OXIOlgOGbPUSjDY6Vgtjye6fOcyBGereK7fmCKktVB8sTEEyYRfVOofsva97cTD
6W1kpDyMEpHGUSGcyDqcgT+oE9KmwdfgseTThgIX1rYhZSVdzEeZgg55W7lb2sdw4OqH+fcCclws
lINYkWvtlCupZUS5MT3FfqaMa+AgcDlmIfxBNVTSOyNTxWsTjMtJq2nLhoVRnaobg79CQcHhlkcf
LEE3ly1afde3SN9kParKyvE7xG5VugsrmuZbEQgQniCINrGyPSWaHN6dReX0TqCvNF69b1A1H+3g
YcM/q4EDU4pfh0Pk5IeCLFSnJYbb445sv6oSZfhc6MAa6eHp7ZE6uv1ODkX5mQifWyJ6xvUpbBCw
AjiPWyfK73c8gmKiTu7lY/w8pm9l9eDXJu3p7whK/FNN6+MQEDQMDveXcqg0bTdJZjxSJIzPyF+Z
pT9I0rXePKsInI/yk/U8nSXVnNzKvfzHP8E9FJ+B9bdokheGWtQyGm54dnCy0oIiE4izw1qNM1Mg
vFs+2NuFdsyoEAGGlfdHrGMpBNSIfGBMVAYqEFp4cS6ObiFOqjC6eUYDJKRh6FUSawCHAQIR7S+C
nxtXrA5NDI56zYyls6n78Tqp1D7MeWSNWyGUBhFzTRnJ9nkTERMVt7/Owbab6kdUYBMAj9Zw4RYl
WNPl+WBUJZLFIPPlfmVYEMZ9QuIi9zphTvUYRgpjxuSim55Ntxtqkwon/Hrt85nZOVK9o15/316A
YQnqHhWN3QMSNXdZMpWTYscHMh2LFB0f/oDXrSsWI+dbSNXO1zPDqW6OFdqwY9Qn4Saf/qeSWyJ5
wNOQ4CQG8QYYdKZzhAKvbk8qD87Kz++zBjTzVD5vnA5nwIWdtHGPb7uJ0TCHvHsUAObrIuh8uODA
n4aeWC9XEOsFQCe8jQxgwetKTCtz+emqitj2sCCwlU7MaGuzSm84kLYvNvw7aluPyaF7S81O7fhv
wTG3GGDiFMFmijTLxb3bSIpgInRBIIsbcSz8uPV6GWPuj6WVdLb4JQjEQqcvIkprlKtuKGSAwCzZ
r+BkgdwpYgpCoFvtDfCbg8tLnljeS2Y+L9O5e96oYnPvBPrbrn+UEXoycpgZ39W9nKQazOkL0EXK
+aInxY1y07PVyjEpVjltJL3nI+Do1yg+FilrLhW57j0XmiaApCahMOOX751uN75ulZ/cZkhkNDpj
xiQ6v1EMZ4Mj3Q1r2UmfEZdMqHH/CzRMSlWT1BwCoFIgsw0IuUFIqiAvUV4Qm4T0KBpa63wAC1Dm
df924FMbnfCreyjn/1SsYewIHAHFXI5cs9jQqzQ2A976qSLrdbfaxwmQJtT0Xg2VPoM75ZK3Vay6
99P2Fqet3qwRq4HEd1ks1EGjCSS4MsZ23p2ZEDu9o5D9hjCt4TWEwjWMEPz0ZrMwXpE39vd9adF9
lvH8yLTjTnBIY/KFxcXQfiEgTo8xK9npDJlQ80hzPEex6iQMqjGf1C6rAOM9OcYelJC4CApZohpF
Aedj0nM1jK0J4YHx9+hGDFj4GXRQ75ZLOgwQxWBhbj15axFMFD7Kx5bGohumEVYQL1eEGlYyEJUr
3Xw5Z2/8LkvRB8rNcqVmCrTn/h8G4eBpEtj0msSKaAOmZkbcaT84Ae4NopLBZ+SA9WZg7xCzRl58
3kLpGEACB3V9I7z70dfkUIPYkB4j5af4GmeamHAX9Zx+Pd2d7VoyPl65/BRXQZQ0+zxJMy7P/oqF
8A/4kd80PSc3JKNcL00Lio63E66Oy3jza61ZVZCBlgaeFQnj+cOb45d0imbzQ/KlFeq0DLIquVjq
0n41+Wo4P9WHh8wmoUEGIL5UyNw8P9rKFGtkhxzapN3fVMXXh4ysQxgZkKGlsNodgfKqp/89HzQR
gwMc4e1qjQ+xXUqoZPs9bdDGA4bZgg8cfhboWMVBjVnQyIn6ttKV4WHx8qeAa0VaNNDmQYqEqAaX
Ft5IMpsJDTcO6n06BCeQuwPeYQnS3k6+UU3fF0cHZUmcmnef2nW9M2Owyt9Re44IyMuuW6y4atuE
7r/ejYcEgdJmRrRBhBUhA/qxDv/0cKjqy9LACXUJtN4Ww73vqtahb8b7CgulBWI0rutlPi2PYsMR
+T+SX/dLlq4/sroeJkIK5B8auPOxyoq+N8EttccwOO20NPgC5hDunWSIFF/2rfXlvjW3JQRtqOlK
ElRX4utw9JgwnaXnaM0Huat05RQVqf2O53zxIBBgOxTzh/ZgX1hUS1DSEkquLh/AVt5XA/AwzTd2
/kbSjP7R60b5U1EWsVltveU5/SdgJ+4Wer5DM8VV7aM0tNU2FgI98HrZ7/DexUAEf32IM/H6Y8/e
L/rwo7NC46I1wl7Kp/v5YcdS5FaqlpQFmhfoa7XSdG78Wdgps2LiEn8HAhAcDySB/3QWpwNyAot+
aB/dFe8mtW4g2KYoCfAHxeLI0cpICP1XBbhTWPrjMOIUY7Izrsuqd9lRNwl62LiyHywcG6MpNQub
9jMipgtb2xsksCidxnw9RJqKADY0JgtbrCFBt9VvyQZciC4L7wiZitiy/HYvz7GWgbM0kJHDqyqx
7JSbiEYO5edjlNo7rzNYctdPkH6AKSWYV/uK1ayQkUNRvhxuvbwQLModbcrvWelNhJOSMtv2RtMp
HLf3pLS6aLMUp+zlObkMfH/xQFdUsii1oT/i7Xbim9WW21Zqypgc5Cvs0w0e20YZ/AjUV4e1Oams
8LE7bf/D7X0goPs6/HbRQurJVlsnMWrP1YeSNzPX/eJcn8QzNVwFcyjMI3/z5SxLnXQnZgn/15du
d2wqpp4Y0HzhYr9cat0DBtemFniGzHpqtl3wPubTkIm68bcZ+U3bFG9xgbaoXEFDVsYQl6R0QOjv
xJaOh2qsJ5V1t2fZJHdh7ZGq5iAi7pyWDANi+2LFe5tiEDTr6M1tOjuygMmSEsrCFNFuMWu1uwt0
esT9tPx/Pbo4ZpGytOrNSMZ70oFy26T1xNN5tq8s3QT6Zmx9OhBuHDyn2pNIYkiRrt30mA0p7LKm
fcvw/ahvkcYTPANPw4gmRtLiuHN5igGpuiF6Ri2NWGaELO76eS4P9ldNHCvQ+/cPcVTkv1UkdKRy
2EPSOVd9YNBeA7gKLgHIeujpoTwRm+ts6cR+AmB1frKGY3Qht4X/vYAQ3L6vPbllWicT66oCPA81
uBblRL2jE8s3OqH6p6GWNWNRHvZahtUJWMWvamM1s5oaHhVo6MqOOo6W6IOqrKYbFhI4Pg1ZKaSn
ABYS/fazThMzF8KLbGI3ZpM66jMCpQKams+Fl6zu+fvecYmjnV33acQZBY8/Wd9R4Mw71W2ZKylH
nlyCc2DDTz4UeS455QNc+8K5/8jlacGiT5IiLxMiPs3BbAh83+nAeTBSJzWtn7X0hNMAjuKJ1iyp
C/eOqKOm1Nbfcpcn/T1mYO3eCAxyRHywGyOKSiHCrdJLqWunRqCn+YollJd43+H7y5GUJ1U1e+Jy
VP7k+TobNFt1fOieWWpt1Jfea9J/ZUXHlGCdA6yahgJ8g8uo66bj6PkVYLxcVBjxiKCp2xSXbBr+
HqRXr2/UIkBwz43FJ5IJtYpZBdf2R4wUahV1cUsB6K4R7h8RwOEjcY9BDan1zmPeEX1JiWiFLPRU
qk+EPDmqJXwcV9t0+rTEg+RmVE1Jcv2X/aZyfNam2VUJuahU5bzC2yPPTXvt+gz00oQ/M50Fl0Qs
xgevMqfHCL/fZmiejuO2O/ttMUrtBJhCHjWY8+hN0YtNMjgpkaRerjACQPZJ0TaAHqRqCBeKYq7T
PVgd6iby0WMqqo7bdF3mSnw5w9FHGrzlhhtCKZyD4misJpWAAy+PaiaKvg+YzpToHhVmcS6aFQpg
2/zq0Q7Kb1Cdgmc/KRvXDvXtOQhC91Zhaw15blc618eWZE8RXqzlvZzgy3BNwH/5zraKGMvN7M4Q
4eizzpv+N8DvKkXE4o58QC/NM+1gJ9JTebrfvm8SVbOtLhnvQEf1c7gQUnv3QNZZV8jmEtGCmn5T
qbkWCxxVlF775cNvv4QA7LU6/2z6smnc3bTu/aw5Hs0hnUTd3k4XfnHKqPLz/G/DWB25gqlmbzLf
WL4f7VopRtFD3NYGfZl5hlj2m5VBMbR2xOQdBTINJGUCMJNORGjlQ7KJg0HhKfuegMIczp8enjvQ
w/xB0lvhQGsWqyH9ImUisR4VSArTmjTen5YQgUIr/ZNwY98NkdHNsd2iI67BpTUXVKZrwhfKGayo
JZfhP5eTGO3ErQphR8Iun82OIB4gr6g3Ntn5O1j09lYIph3zHp9z0Of8/Z5xDFs5CKircgJdadNV
pxPFcL+ckOF3l6y89u8gXTSO1iTuBQZ2N6hwjH7fBMYCMUf1yDunACXZ54ZYpC9v6YmMxaRo3onF
+u7mcgwUuUTjEVM1RsenXksUmCkPJleQARX42vJrRCR0qVvIhQ4WKyR3Sn8J1Yk9UqNXUkLFtW66
DdL2Dhx4bUNktQXKdcQSi6a0mcHoVqxSecZQRovokgTjAe7s1qv8szNequWTQd5WaQzkQEEJ9eXr
t4Y0mBBKzVYLsxukF6ly1Iab5HOwsQeaC1FBMH5PY7GkQY4Ku2ljmVQFjbcg+kT9DMy+vhQM9Hz5
QVWy0AEPhG2i5Fiwf47VrQk6ZBevrsAwB01djzJKptVbobAFElSu/CJnk2ssgm3ZkAS2Xw9BDJVn
KMbJnZ36kisfm+dtrNIVcnpEY2kAs1RuI6sj1jJJCI5iBtODpgl5i90wpq1jWMTmumil1AgcP/R2
WUHDDLw5iKAMCJDy2mKJ0KZwE96iy1Chju4Alrbflle8q+Q69NY2vPKD05e2ec8gSwZoQx3B1o1Y
o7iJuAvry0a6tru/t5QdPKc50/yl/M8KwUQgyg87oa577WyJc0inzHATn6HsG1vXaskS6XMcDbHi
dkPEVyBBQVUlcVCaclw+ULWhQWE5WixqvrHAMW/02un0qzQ2/Rt2BFJDL6cyitI/YSvS9vZSrtuA
8DX5Q5Md2blXpdhAfD2i1GlvRr0BunXx7CA82vDtP854i11Oy/CY5Y6AcUc66nojnp/MIJ/JZ47H
bPYPS5U/OjOggIWNh6zx3QRnvOL8J0fkysCEYG/I4CBr9+7TCwYsUo/grSqYYbgcdnOEuYkB7q3H
pz5XaT7Kyp11/mZyMJz49uXju0trzWbSSp4kjgLOwdzwhL7u0MXFyPfqWWdqbVgbiunbDeRsWzFI
0LiFn1YX4o6L9ynih3vfVm+PmlLdEWxNXHC7mQjqT2au0Z6N3h0qH+zZ3n9yAqfkhsO5CaZLe6sn
hEoo1U73k9xb7XzMpdZMManXt8g8y+TF7mpXl3IxueIUUhem5Nm6zAqWJgfUPkSSzmkGopTp8SQo
ApLCZFlpyYo9WIF0x66/7pZfIT315KO8XYBrxaqqnCxy3LyqQkT9tZQ4S7Qo0ovUey2thkSlKDMS
PjCqyxPhmk1FCMNWiRNYTlBvpvncZwBqK0XlI2fh6mV27E92XZFCvVPMVmmQHh4E/uBnd2g4LSAc
eYbFOs4nHPp/LMKt/TrcStNBOL+cyz3iGEETexjSr7eR/VKx9K6D4dttuOHqibMEXkdjrhAgakMY
ruaPjiXoH0yFhlVXkJGEzvlge8MfhOakW+MpgcN1Lhc3LHkRDvt5BWOwPbn1MnkWg/axyY4QEHdN
NuDEO91m69kVxTKbVv48RjbPXi4Ri1vDVxVk0pYyNjdTN2sGJHBaxZGmZpxQdcvIK1ydxNoIJu7d
Ug/+87mdGnZUZr2mBMhE0AkzCFPpuYlDhhN0KciLzeFkRzRjwp2LvujJvX28XBgam29PkeE2a+VU
yo6ZCehnO7JT6LvEXq2z1dHS6LK0jbXGyIByzOofXC+Y09vCUMCgmGhcs4dROPe5m4NKkb1jywye
oJn8+dojFwuCh5X0QYwVCNCfh/+uoV8fcwwtjqQhMWIxFqdY5soCQyYJGK+ANro/lbw3dUqVtVxb
MudhBDYRFsaIEGW1v7KV0nADbrjidfZN0/mJt4SjwfBCO7Fur7xx8DyEK+UI+gL178ezqyaEFo9K
g+Eso5x/FCHtXwg9Vv4a/8HlzyWP8xcGsmbmJ5WnQIJ+6yV960oPRtiSpN72LjIuKBQFdDwBLP5r
kYr48VEymb2Z4RM8ZVOGPW2hPAFU9+RxS+HRfo+8hqicZzlAvva51F65BLTntxNl2gzhuw330hs5
eIeodA/mvK71zzMgJ6gHk6jlX0rqRRZtGujaIWu78mDRuwZa1J+kyXmOy4Wr5s6i85T1c0SgSqWx
JyX3+DQeSjbZpVumP0wbYaY10cqW31ZW1V9luXLlY9IMPHqK6jPOWZ2VK3JIRF0jRRzqbmnA2r9S
pf9R2YbwjVAM76ZztSrWFDRpR6dySAIGegHKuWnilPs40X799la6vJECE+N6tlSPDDG7Xi+5ojmZ
PfDUBbJHdV6qfeTHWpswJWMLRn7/cQK7BtXRbfLcztzIr3gJRLMfrPQtBugXpDzScmcESC2D5Fn0
FSN0Y2FRYK1hXNc/fpvGL7k/kdzU0XFFA+Ko0/x9PwvmLgZP6wGpBoZuN8asJXmJ/m8XiC2+4Kwg
Er95Qn8SRAHAKzcaLhSTQ5ssJB9hg+ydnghWklvxUXWxHafAHseZH2nLD86e7lTAfqk+AxVvhqu5
b5H1IMOeGQUwiPOnv0kr6AXZbfz01xmwl0nnRREXGL/l3FE9d8XaIZmxPqVW1eRMj6nRqGQiujRi
PGGTw6vwrcbEYFB62amy9Yuj9cjqUbckQ50VNucCmXN+YuBfCnNQV0mTUw0w/4m2uvY3B+AYeHg4
MmA3t/tjq+yAgadnDQv0TThuJ/xCnfWLIFCoUDm3InpYlmR+X8ByXFubQYUfhrIboRMTNi7pqsjJ
oMBcumJ6J5pUpMmCcpJjqcfku1FP6eoADOL1xc3SkLFVjrbWQJGRmCXvx6cvXlJbwPHggXEBAqCn
DnP8DflTzoW9fqszPOLinDUIiDYcyUvHwj4Lh57IAS559G5CNfVYy9BT5yb/iXtYITCbql80JF8U
1tdkXIXyCygL8933po66WhzTBWUBASNgzzLDUwZEn3wyVmPkzY4rrlCsi+3G8gKcd4+vKX3s51Zv
9Ys4w8GHqZ0kf7zTIohm2v+kWQjzmj+H3ziPda9AU9C86HqGyLv6gl2HH20tL7daksg1Kaf8r1qv
xtsalV43WOxTYaV1P3MNWayLaF0CtZkQIhRUrCkqicut85tkUDT+OR44vFBX2V4EMtOSrWLKq0Nx
qCpkMrjXUs1Fn0xRRtJVo1Hh9260C1ilO6TT5+99jtbNq1dfkoYQTBwC9/DWb2qGgH2VssSl+Vn6
8LUte7VuBFtHnIviHSVmp+6IEZpitFdOhGY6yMqEcUrvL9WSNbr/pMV6YZI0lHRx0aU4uCuTkj5G
coCxkaDsRNLcyk6LYtQSAa7zBSD4kL/aiTSZJWHDeRzGahpT1BrFANEkr5EMkEKBajVYPq8ttO9q
Hd4czOjjvs1u0zwG/nN8rgN4TINWCZJYuxix8lAQb8l5udnuoXlUCKyXKpcI3V90tQRhuSREHEBC
rMfbRgRACtaEdVF8KZjEEvLk173y5ZMG0cfFqeucyibQUN+Qv4/8ThP/iBAgmcby1S9b0Tu5U+VZ
WfcsfJ1Hh38r0sZNToDfa0j0BlR0zDmq5QghkJHbBp5FajvyovTjWToIX79fqf2ZQ2RxZG+nj3Eg
eDa43btW7hCO9+d0RNq0W9qfEMUJX9KiSbV/3fwvlZJmjbaMIQJxbTL0rnnlqo0GE/Rhy1/Sr3sL
MhGSNTXACcKyV+Zgr0JzoN1oR4THqoDZ93XukI1G2+upz0U3oOG9zoAT0WZkQ24OstZYsMshFu1h
Ut42pnd6OdUqDsLQHCh7iH+kGBjGSxPbgFbIpqHSejzj4eA361kRgDDxIOZXqBv65VVZxSj2kN53
ijBemYm25nQokYIsfdFyGBo1Pv+CvG7SIBPp42IstoIht797Hk5iziX7G/ULS5DKO+pa9XaEbkr6
eBYlEVa6QMb3bAz3J8RN+08pXL7l8c3i/dpfJus4EdtF/Y9M53iEFc5WAtAYkPd3GiTGkD3UxjK0
ELiU5Fo7UvOv1AKh4M9OUkR8Zl6j2jF1G6QWiuU+lh2T565IJ2d3cOXXjsU4GAibWHnJePh7w0s+
naItwlq5yBCWcGt+EvGSSd2ewNZB3l3AcgPNsY0Zm+QfmDfSUqQW/PmD2lFagqPT6cxGKpaNj5uY
iiSPqjpaHBU9WH12E9jjjPrPGv5xuwh/TW9C8fh9VwGoq0JsEiR9F9DkGaV89Ssm9z3IDloRkZbg
N/s1MVy6PMOT2kyqrBqva363tBOYVNhMZNGJuXERdKEF445qo4VBpxwQY1Zhw6OpZfPbjp74/CYE
zQoj8MOmAYpNQ/rhRXVFQ4Yzfg/tuOCMzChvr1HfS/3IRiUZl+euJxMqsSF9lwV/v7g3DeqDCotI
JNOeDrpa6w7RMKX8TeeAgc7vxPyj1RUsJhbAJKtb5savhsrY6/WtPhyCKX6bCP3Q5VsrwPIQTnz8
87FZ87bfaixu2QvchDrbYxaW3GLVOlGDcrQSrqYade1z2oyYfgFdqFoiuqF67Gal+YmgYFQLf9Xe
J8GQxL80U8hHR66lYUi7Kmwv9O5f00177NzEouDs+xk8Qd5trnHD8v+fEVB0+HpsR63wzjlAark8
IqQfyQhnGeSENZ44Ln42yU7Y+Nv4UFrprN+ng5yrwlLHEBLLqpZ8CJBfZ3jwd49RgoCNBXF+hoVD
Xg7nEkvpneVZqxuzKW4MshPlkpaxE4yVdWO3XoIQSryuFw6WdUlFejtFfF+AmcnJPLupsk8EbLsg
YMPjxvFaMJE8keadqJapqyYD1w6IuNnQVm5PgAqlFIAU3YhD9Y1vpplY4WSTJUZQU0eiUWUjpg0X
GU9/SV9Moow11WVlyDpo4Y+Fhc+usJoSEpaxfdFFdRanXXW/IapQGjvaC04VTsEYTfk9qURY3jbm
HHuOo2cCoKols9Ml0DRIQ+wG7B/U10zY3jMiYvpRSLnpvrx3V7vzRrUEt6skWL/ukby1mgKuc3nF
6s/MHgwqL1wnpI17ECMjkPv09Rhh7tNF3xgpctZMUaAmudihG3Ras05Ky6Ct5RxYE0KMIK7A9gyY
O9pvXOV4Vs40E5DMLMs/bHHVE6I3QUWJhTKiF2FLq/D8k+IlJ4Fk8VkTvCqFjAMQhQVaQB357ASv
rJPE+ttt0yy3UH93QQrUEiRiX7PCdU2gqgxOXwF7kik+J6Vt1q9KyxUPg5HG9RY7skixrqw+BbWq
t5xKqbFKeeFAHdv4B63xeCO5Whe7u/2eE1JF1ufLGdndwE3ViX3EmyMZkvOKD2nxKpVuFrtu1lVi
nSIP2IlvbAFTZ4mluRC6UvbVFeLLPTZsNmm/4DO1QhYWAICy/lclPNXP4Expq+csYasxJ68KiPfz
w8QKEpgEPaYOl+hmIgapmnh09bITNP9TA1PcCmUxTe6FCRCSR9BoLOECb2eY3B9wzI0gO4uZczx9
vPKdMJ2CRj7cn/+esalSpC8PnohBFnK6XglOaLTUjyPYxYxnfLpAoRbihXTkkdQ+bAZziW1HhiOR
kta2y0n+NDjnaGfZIglmnM4iEKmyjxuujnEfVDWyIquJYEFFVt/vBEdzNw839ftGeSxZOGtsqYYF
LxYyB4qfwudzSjH2lWg1HRaWwevBy5lJ0FETA6E8G367gjLpFG2oZPzXLnZDoztD50i0YCPaDNRK
3PBJ+TLEdS32U6M+l0vOGxIXHgCeg1yigWni+ROGd3nU4tGEFUUhAz3cA6KroTQitjWgkbyI4qM8
oTQcvQIc9GquvAbfMdqzAlhQ4t6c4E1BTB613SqqVXk2NIdgWoxcw38kiC1D5m452Zx3+FwiB9F+
S9GNejb2Rq28Y+pGt42ygpPIugQJkBcgSEfLM5/yuz8abCYqFtFsaOnbhUthcoLTW6jx0nfV3tcO
tVwg5a38YG/hiEheWuhxCtuaQrRJ/IhbNp9Zkdqg8agQdpVGpNwkDctHHGA4NiUE6XMSA9rI4Z0n
dfX0XxW2wc1+jkD5bwJ8VoYRPYJTggT+kon1/aC7V7DCO0a81jnV6/2yAaMHkkUh6keeBY+c5WMS
SSi1x6r6FzRW3ZlJX66Htl9uUUXO7UT/RWZLUtOwWowDPJcXW3Kr9eP8cw2CwFTvQJnZegst4FDH
zsDyPCiYoqQ0tUc76PEpyUD6osw9Wf+m5X8NhGDpQvLmO64VbhQuEdp+X/AutwJuf/0qIgaV01So
YLt92Ivm7M2k0nMblf+aw8/Hnuz/Nc6TP/hUTG5gtVh6cc7WW24BBItamTfbHQNWydYaUfGGIh3c
v0iPsqkDjjkRxVplbdKoh/I0MMkhTEIEm7gzgFxaGLwlf1ItgcIeD0koeFJVNbHGuDBOfYv3CxD4
2j9izyxz+gBNvgQmHXWsiU355QRvbu6tdUc0fgCpcVfozbW1PgrFLrR7pS577gpeO7uRnGFBzeJS
fu1PFhZjkm0Cs4FtqFK7oo9AI45D8KvQo7TRP82z1abgtAj5fYmnrmJsj5ttRxzcRzflCkeuMxAl
m9KGd1ICgqPPqPq2kE7aSs00mZqJFpMdzIxp3XDpEUKoPrSIlapt+t07+EHoLKz64zpQFtagKSLj
sfXstpDVZoa3e09gO225UHa8acW8haOu0VwSJTlO3KO41ociT2OTbxlQR8u37ryZlzUqrFsJLNtU
ec/F64QRdILoXltr/0LV9k2cSnYUIjG1aqz8jmclyz9kiXV/3kEI2+Pz22Noieg0liZjWBHF7X6q
u4L6nJq8xn2k+1ihxA/sEs6sHB0Nfq9ED2g0ABvKjA8zMApTeLRcCnfv5UYTXW0x84yO0AlqFyVo
t4PjL1CJIrK5IUgGcIO70rzbKEyhVGnmqFPqLdicsS9ojREVDLRCAPMG6gQD87PSj0VcFs4V9/Ij
+/Bl9CnxTmgQvQV+RAuN3Gh/Gd3dEb9eWooxq78PAl1E0URs7lSKa544vxOjLEi2I/e4ySiRWh4k
jzbvLC3SPUa5Qx/9Brr/TW4lKf4SWjonkN/ENHDOjr6fhfXLKge9pvuhgKcfO5ZyS+uYQ+MePVt7
5T43g1XCYSu20kq2Pcy+p+zHATjGqnw8xGC323abKTEOflrubaF+V8q/IPAVG1ZEazfyFG8aWFPA
SfWKb8BJq0LRwobhmd4yiCAqdzvOz5LqtJ60sWLyjPbHdRzMMpb8jP0l0dy7vdkTdLqV0us6eV4r
kmxSU6xcArkzv1pVLxg1EOR62dhSbiNxGjXurKrcVK9hTnv2RU5+AVkUa91darjb4nvxAglDcPv0
TvRPUeTR6v3hEAl7RpXmi7S1mxfUGfyAs2K06BTrpcc27328X4crnf04qWwX55zC/TJfrN5l+G5o
nFCPcUlqrrKG9jcGehN+c59nM5i+GXN182ZsIFokCVdvO4klgT351PrfM9/kQXtqKdDyIRRr/c6s
NIw7ZtNzwlFaNd5RsWxZOJGVuiQSYbtwEM1cjNY5SjJYQIotUQMUgpkMV9MigL3rP5JHmfDHUPQy
YpxjgJ0QEOrjiRSxCgJMSbz7K2hCSd2bic5U5e+0xACGnE0d62t0BAQJ6a1LexkaYs4/PSGhQgZS
iTSgHT1fJJ3Zr5CIZP5+Vz5BftFyIdhq7LYk7q2YrAE9iugrgcMj9j9H8cqO/iXFpASHjoPkHKUv
C2n8XS1UZWb4qck6tZLS7GdeyTZizyUrZk5sSvrwjP7qjeKtS6CEiDqyGw7L3eDQN8tJsI/4xGYf
s5L/JwZrnbsRFF5N++5nBXAMivZ5UktndTsl/+EMdvODfYk0qJX0fkvMsjaRMhSWAYVBQzhPJh9S
qhypQc3Rc49fLhPi8U2DEBMN9lFPUJ4EiKDjEihaEtgK2byEflRdMSI0z38lAq5/M1WgG1ix67NL
smM9u2JmAGxnZAEawIDiLZigIuopA8FHU9L/4btqhsb/c+rY9lFJpl/YLIVdWctgRvqNWIc8dB9b
OliVfiXsiQ/lCwof20ksxo9Em//Q2rtUlWs36vmw5pzyEK/NPmYGvL6ZUhcy8eZFJ4BvzrWSbk1K
FmebO2tHDh30ZRrrkGGzet3K7+lyREJuYk8U21Ic4TTODkd+0hiNXD2EfTaISRhl6oSrtwF5Sh8e
dt1gBQrkn4ggKZ0infS5gUO76EUlQE8E8JLHzfRN/WRoLGt4nR5NcaP6ur2PdUTAKaWYcx35iief
jgRsqEL8mn4C6/dcfnCNAFGXbHDdKaCsaDLpJ5GyZwdQXC679ago+/RfrMg8Fhw4s/eyrGt+471H
qBGQFe93kzB/rEbF8mx8ybN9LqZDjkUuHkRAyqWMyhu3H3O9DubcHFf5XEd2dQx2QCwAnLeWvO4Z
gEXju42b1hJeiXuQHhSeiRZkJ4+khKmhi+WZq8td+g/sfTd7l3RHg6wwoXmx57GGb8ElO6uZkGCw
ifEvWpgD9gleFsNEvKy70fZqi2/CLsQyhgA6FeLTjG4z+n3oL7NaZ2RptbpPfP3YuPGdPgjB0rm6
ECso5HDs+/mf7Wv0QrKvQw5JRfhD8SJIWHzEWpOAeu4byX61YbMR4xn1PdsNqq3PHtVMwwpYinQd
7Xo/azTtoktvtLnweVOns7lxDBWR6e8UNnfNYaFm+l+E4CCorqOoeAh4XXUnIOeepsFMHSN3WZjc
7bDEEQpn+PNRWPRc0hSGkL1Kwjj0ct7mqlpBPI4UhPhyF0mWubiiKu8zWXAsZL3NUxMoVqP14D+m
r8k4KepWE0ltYK0YHhAYldU/7207xiJ/5hPNbyNyTxMPx3ubV0XeLmoxagkooungGSli4C/MLukA
QXQosUfqit80myFaww7oDJzjniUeybSvzRZcBhIRsN7VBFDEb5EC7AEpeVNkzeVL/sBlg+pdkbJ9
EvJqYx0pqtDZgFgPV+4hc0LzI5PukoaY1mXSKGPXnH8r4vjUNN3dzaA7nBdbD3jHt+2yAIwMYQ4n
32FdJb87U3rKSmfBkv773Kh8DnzB+rPYpldnA4dbelApqZ5mOlPtluPTiSxoxtLwUmJI1EIXFzrj
5+JDpVMpk+arAlhUZZ1XMFxKgUHRYDr3fB+GOwBHdf7gpSJaa1qTFbIdPqwQ2Zhx6VsEh3NsdLZr
uUOLydyELoGr+SBql0VSpYimM8HHN1aFnp15DhpUFZvox23kEszFglMkNnv/O3ojmOcK4DIi4/xb
Vrq1qVjgWIiZFvsoKdtBgoVJO7yqwDS7rCF8szkbbnnCZIr2ufkcUGvnGIbhijfK6oid3vTE6amR
S1i8jyUsq0WoCd+0lUqYB3ftfY5TCGauDqrwFbl0ngkWEBNEesyf5ovpeJuYs4sy1mkLQ6jOtsB1
ztKOJNqkqajkoFcNRAVWAaXQ0bAARFsCxxTSEISBhaflED48MwerXJ3wzIqj1zWCfQ+aIS4YSbgH
CThvfx82CP1HF3ONUvpJAMgu6Ri9vI9tegRV1swL14tNXcH4hD6Qd55RyiskoP/fudzeX5D7uinL
QBNnWRvVoAQT/a5k8ceVznYfaLEgLHYGsOjongH352/5l1tADW3AOZVXMGmUQmrMsV7nNqD8G6XF
U9nEFok96chLfp06/1tJAwEkCUWSU7ILCtvuV5polLebj5W55h65AjoN91afHAdW/87z1vz6CxPR
jcrtF18EsQSUutFuo9DqGDycFSXnlFWr1QbFzANujkgb6pse3sGwwYJNVEhsXZEOqjYThx9ANKQO
HuCRT2yqr71TUJ8trmWxlOSQ4CNS4DScTA6SP+w5rd/60FzHAXCtmgT6oCLMGtNtmqKwSWdVmg8G
2xfmZMxIzZhnnQtFxZxq2RNDLeeHm5lGbipqZLvUnFDJC4VqE02ATxaN6iYgGLmUNugbzswhAGh0
ftip5aZ85QsPelOXrVxNYBh8Of67XC70OtOxQIjwGereB4ImN4cHf6B8z/7/XrXnfXf/zWQdtMmo
d78XulPCVKF9/KZreWHD5Xik6/dPI/dukd7U0sIs0P8OHARRx6g9cR15wo8sdEWDPhsz5h+uFAB+
UIQrnPTvTNrEH5Hg9/eTpo67JArEXpc2Z3vMGNuKNrOSsZxk2DdGw5M8dVt7w/nH60mlaAFZZYnr
VwbdUbL29N8yD+R/AoqCe8HSdhZoLlPg1yVFIQRXWAjzmWnjrotY4ZiKrR/HPnxbY+OHzHwpkcKW
ZBqg1OuQdp7VvUv4266Fiz+Ph2CvLdBgPjR8B5v07a4AoxjYqg2HPdPdKdOeuuOUFe5dLSGKADqa
b/E0tdi/yP8fOBFUdf6hT+xJBeX8hMqJKF8u0xPpaTJt+BA00J2elAhgcONdvNs1okM/+kf5bwBi
XcpRzh5hibmBxvPpKbBDuMvgNVYZxI+Yq3lFjeHVFWcsLV5IE+KnqWBowCyWXivDWXKtPygn29fA
b+SvP7AwRYjN1J4dLBoYf+etPYdr+5jMTp8Z7GI6IaxkDqr1G/RdYLjcTODFDVL190fWsZlfvn1I
6NU5OupDG9iJt0pKmBYDnZrrNeJ+HOPRgyKf4Fn9P7CJOa2znaVGYEkK+Qjw4nmiyYiQoTvKWWk0
oOZge/fcfz2JLahnNioXicJELph0L6PVuFtH2zPUAwIwLbFra5R7Aiy6q/5aQ0Dpqh1woKsCtcRa
bynlxy4ICmxbfj4vVzxo6uF4RYZtvGpWR+D5YRRNKKmZtzndAuFUJOYZmuNdOkAYioA+qIhqxuO7
qsFJ/gOqyyRyPVBl33r84JwgbBnz7btHoQOhMKC/cJWkFp0ybN44IckXx2XHflis5dmh7Him/VNn
Fsfz+0n4f1UXmMOPbqtUkSeQa7ghy16plmYTCnieQbf0LgYAjm8CfHZk1Ujqbe95QRsXFz4D3FgO
ke3cd7D6wHA/Kf5ul/m7XZBDwlH5TvDO3VNbtiC1In0T1Yz0d/1bXeOt3Kb3RYOcsAKS3Z3Ev1kf
fxhQtFaw6z4VsIn+/pwGW3zLRpN09ahcLvYJu+jybI4UEYqNGDCcl+cGX70+CZOtIMSwYl1ChL00
+m2N8L1aDBb6LzvOBfXIFJsigROMPeoAOvUivJD8HZCH+zpe1ww4lCmSN5Ro2xhZ00EMfqglsTcI
2ZbgQIQZN/UiOY9UFgkCjqvbriSFoz0o3Mnyw1nGRt85Yfh0xn4hQCElI81BH1IQdVRW/z8CsSvD
k3M3eadOd5WU5LHpvAHh5PNF3HuuLQFVzGto6HtIjZSGPP/q2bo8SzCxTL+2eeEuETWLX6bEQUX+
drrdj8kY+oIH15o8jET6AMxrez8KZiNI+IVdrBQkK1wYnIgyODbQ+a1K5NFYdTKVD7TGsMzjhY5k
GzBBEosRySjiKuzR09u7Ast6ltzoF5bTfimZqEOTD1ph5x0FQqBET/MrDfPN91XLskrmdhiWhMbG
431AN0m8aBychoVZbZ1ppKCTbmI1kI39NV3flxo/eqCuCuOzd+JOCV7emNdTdvdiJgO8kaKcCUgp
Na++Xf2W3AAzUzlznXO9ccMWefNz8JJBeWyvZIi9201qYmPYpOlK6B2BPefoYRBRsJfOkUsBq2ad
CCmTSHr/KhyIdvASiS4CAVT2zngP5gYOifTlf6bPLblC8/Iw9Pi4dNV3a12+P5QzqVHle/c/REQg
JUkpC5/8vOsxCw0ceacJ3N7JJWr1NsnjbM4wwBu/TY3+L/MFhdumVBIG/Cbj7HvJ0oaG6zUvQ3Kn
oz7JqVdBJYhMmUo17yIoFWSjjE7ppEnlR8vH8Enlb3eGjgG4WXguLIX6uPbK4APP4FJiAsd+9ux2
og+IkktHiEYJA/XMe7K78wb0O9CM7LEeMjIAHRzvRNt4rfDQp6awCBC2mROUgVeJ8ycP5Zm9W4oe
ZnzlWk+ydWMHLblTXKlQ1Mt+ahEcm/aXb9XlMEdHLFTb2ST7/ln0yQitO5QfhoAMaTwiaqvuVRG9
RXYDbO0GKQUxwcSpb6w8Y9hr9Ky6CrMqSprRknkL8iGPPUkZoHCclJQ9vOIyoGOQH4gDGiZyE1Gb
u4B0eefvZoN3UfdHspFWy8v6N0EtlWq7mdKa6RyXchXMtJjA1/2LjrhPvIYZSn6EUrgdrmLYk4t4
soILA6vrKZs/49UxuxbqeAD47HLx4ClQyVLqgN0ZCC/KaF0qkBzRRDZm8bXT6qoLjjvSNwVTOIpu
Axw7oRXX4T/5rt/le6IdyzeDVIfOXUT7JU4rpAXh8oGug0mGWkNLmfnyoWIkpInsDzdIde1JSD0l
dPNAbUzWAJp6OeqSq/jWJ/6gElWl7t9r38j6NYm9Oxvs46Ng+9lbxD8V/4AgWnqf9O6SQrxdl5zr
kaDsSiavIBkdBfgQKjAMONHoYRD567khtNXsUMHGGj0GFoDHqbCpYmvXRTKQEFST4zsa0WE7bBzD
lRlxNwAHIiIurJ8/vI5en8IXVrcmBzgMpKyuYWZ5Z9D3AzbNmK+DquROyoJ99i/wbvEtL9Yaq4FH
hHfHbmCIwacUf6HZIflT5HvSA7TJm1vOx+M1V11ZhXcRrz8hwVIEbz3tGz4hmwtXnbxlw325Duob
NgnUgQ9PfhSzk7p0a8YlAXVKFiB3mfSeNDWqZop30/b3O8x/QqeN9xtS78KN/WoD499wwluAeLbb
LN8Xs0g3cMgqHSHyHMXb5fZ+1vWJ7WD0HC34PU70zb4ASRyZhHLVhmpLCtQzbrMsr5irXxtwTXZ4
WaHKvwprM+WKeYBRDGQTnE2TXJp74Ck6IO0xFqeOWbmZKGRQ/mFGWe7fiKr5pab6mD/O+u8SEaRJ
SM+EtHSvOEy0HXPitn9IdYK7X69YxdnD2smRiRkxHRRFOMVTsPQQcg8X21cx6InayzFt8ahWmSzC
QUlkPcRCi7zjkrkj7DA4/1PTaCCV/5TXHDWiCfNthqtrkle6C4OWONMk2IUFRHMXBWkIgFiTbDzK
hxewGwWGso2WK8WGthyvdKfbCl0nbANoQNCrWcufjRMxw4T6/J0FT1W53z/LLJcs3RLiLZTJSY9x
gxen/QzHiFWJwiuy3RO9ZPtvVL7mSSCPO/lQyUR7BJgLEjNbTI73G/nritmFXirGO/rSs2esuvV0
xQbA1WnNp21NieuGqOo8ZpFpxfzpSdN08y1O5d5oqGA4eQUNmBbIQ6mtX0vGkE8Tb7sGHFgu2J3A
/c8NoslghFIQrrnWwiwKY9RzoubTKTcbyDh95oBTPl5dxmufJxWN9yhEq3bVGgDfmemGxWmjooDh
Z+1/hFBV5AcRC2iged1NlJqMk1ADY/ERSts2dZcIolN3MLTpucKc0oAn+X+YYPHN7ibYgfIITu5A
5x2/CgWlkdJsXYI0h997PSOJTECBQWlU0i1j3BMRwQsvlc5G2RQGX/DA4G73pfuqF3dI7TclLxiU
pAZc4UX/w8mURnIvjMrX2s9qwqoV3gIRwE9oeiEkmEtDPPl3EIvFZgYYZ+d08pCzeZehOGJPZsJr
iasPBOi8Ord/RQPv4Dju1p+2gnDuJy/FdiktYm/bMLVI2lDydmK/Gr1+W4XWP3N+zKpoZSupOE0l
J4DjXDAJb9nTODlV5pUVbT5Lg8n8r1OrzzMfze3jR0JAPV766hIC5SbbOe1zPcPMV02YPkaT09zp
54yHPaFKUk/paMnzmUoVuCazcIfk4sqF8VO2VDqzJdHhOACw0TX9WArcubCF8HYxt5+9cIcoodwK
UvXt/y4IjGgk41z/Kmpwt0Eal4/HkVbAX0Q6GHcmzCfIZ2Pq3Fhfhn1dBCONCcmGhjZuyqLRTuqv
8ZJbtpfpGCvOgAr92fXi644hGlQrTYVfrKxVh/QrDJu2ewcoaEpLy+L5NC+yiyX6MNYyVb4bWvlE
6PeCqJQHfwJvt89oNOnFq847UHp8y63Pz0lFmLdZj52HUKpBGtr4yhimewSclyKJwk1eqFThvC7w
Ejbb39UCN/hhLPg1F3YP4dcVIvpGYDQY9/IVhaG3OizgXMHuX57AqC9OsUl6H2QYZmyFxhFZhUZq
/4amrpDN2HvEFsq1BW/OxfNuJtvBB82+Oq02X8O1unLDN6Hkb9D9njsAxH5GN/fr2UQUmDjzTXNN
1awfS03xgxNQhby/p3qrz67YY6+IV238839q8QAfYb+q/paaTjxN0ERdnNkYw2ANvkwYw7uMqc7f
QV7mKFacSBxLSqWsQOqVNZfMumS+J0/f/2naQTRU16LbJOJc24ECsGKKZtzjPMFSLqOYiwDejZoT
3PrkqKU/8KNzoqHhTltNCFdmv4e6PlKxzYu9/lLsP+ZZd0Mqq41xxNbCIpt1AgqQ9xdlVLJiCWbY
6DInijz/UAJyHr1xWpcdppLJxnIOYPeFCVuDZwHNM66bowIykzW6n8QwUKptvFQLlbYwp4/h+OJX
aJOxNOZaArY89qxFb1n0v100ozOnsuCb062/clXjug9p/O5pM942YIxehDzWt7xT2Ny5wNhupRJy
mBdWytVNc1y9gRBVGQdTcNb2eC8m6trHAwUlmiINdcQfwtrjjTT+mCUEc0zIfniLpyzyYYvjrGsK
696Y4NoaGmrksUNRv0tU3RlPsAE129/RXdBCqQh+kAmNU35kiFWhBUZ5CR4FYpGzcrISBcF4rnFy
LMlyw4v3NmEgIU7NtjITJFOI7ilY8GxzWtRmOkBVAZ+YVq14dRbWJOkHt1k8B3TRcb2nxGxNYezx
4Ko7z3Cmox82d+ftMffHugLD0QVqw/d2JareI2wX8Fexbrn3o8iAzprsEFVrBZKy6Y8R9SdenZ29
3vFVae8ZIn5CK9bWWewAnabzPJPu8BKJEXeV7zmgKUbameAg8m19S5kH+L/3HOt4q1yM87MpcP3T
L+jt089bCpMsv8eIO+o+jYQj5UL8+X0EPLCCq/9KKIXicifqe/zRBw59eG3pJxcyjSc6TZ+T76nL
GLp0INh3ic2tDGn+UOg9V5hjUNDxf2EkTvaBBYmc+WOS9Divy+wvAT19yuhYeYb4onOQtdw6aBx2
ZcxzwuleOrfYhnDJFXJbWcy6HuL+3WZoVpEjKK22Am3+ceark9Hu4kKfACpnDfUSgHAt1wrqXNnM
GiqXDQ6N0EecwV2dI+4ybcT1aX1y2alf5pDpxenJpnnSwu3xnhQgJvMinF6qgW82YFAH89ITw5LK
U2J2hmtfAkb+Zu1xVkQPhXgJhF6oOOQ8Yz628BJ2k3R10loWIVIZ1P1Uz2uIwuYO+W0eOK9jsl08
X23tt1Ow4fi6WlPy95eqya5DOakARTJBtw6cma3l4P3EGwg12zFseN5BPXUTZTbLoKxfbI+RxiGH
s5POOCLZUqFXlw6i8Tswg0vkxmrwI22+LjzD8HF8vw/Or8ZqUlQR7F1KsU+9V+36ZQ1OpwCNuD6p
Fg6jSJdZFd93dE0onqCuIhs1SybStwPBL7TvYTLut+dAoKysMWKe1wB8ErKrUq9DjIYK9xj2nBIL
hBqCopxLeXsT67OvEr33N5PppBSDXs2W+MQwq3SVYhib2dKnShHJcUXzZ3rDUWMt9i3HyoRtjHsQ
6YwTu32vMkOL/+Mjq8c6nlov1IN6YcBUBgQbghssaGp9ZTXkQbJ2rZnsTelwnSeb72Tl93a0WCx0
dSHtFt3wZKySSx18pVvU5Fex3b0SpN7OVdB/vpWupBzQAS/pK6p5cIcwER7XbuomlBiK1IHNaXop
HhfmJcQMlAAPWpQo+mg/OutyWGWbqodjIGPOM5BdVoYXMPDRFWwrwGfYimG4OvYC4MgBR1nBsiyu
F5XK3neVcjKqyY20/ra6bpGrqK+Sla4u+modgMtcNG0xY+lZQiK4occnHx8VvsEC1pr3IOpqAq3K
BXEMLLSQN7EDOf6axLMLnczy4TPmuP6zIMTgNzNbWSlE8cxcYtOsAHR4ThKM+F4vxu+M+7c0TsIZ
cj3fG1nw6nVkTT52oIPxMsqCam0RIvNgOKfZY6g7DtQk5GZTTxE3OLYUcwQxa9huaA/suikXa951
tc7udfTI+ljKTGRJRkBAxl9PS/qbUTwnj4q8BTkVYVQDBps9Z6pgwCiaDYbzhGCbvVp/EppYsK73
8OZ8wh+Du7jmFy3EotGi3ZTvdjlpbTAlbdz7hl4O0mFhp84RnrdMYaeb/p0il47FOUQpcHc3zMtJ
6XvCMfo2lr4ykLAePW1VnYg9pRHGJ5Jjo9posDuwim1lmulRYWKM8LpoedcqXtxL7vgAbMcA9AJj
tKpFf3jogKjEZubAhafVmxmhEmxx4Lt76ormvpZGPQagnOylvL8Cq8Zk4XvNudu9XbHv8FONPi6b
UpOm83zRE1SVT5ORO7dRmkGNPs0984HKqxyD+NbTOCAoS1a3OR26MsZa88SMkhNEduArWz/n8hMW
auEFEbiA30TMULi7OjY/3CVsizrixmVFAoRUtArk7iz2ZYqb3wBzXiwYWEzr/qyLL2lZnej6WXgj
+6IM+halXvoIfhs0hS+krQgfcl0hQ7uhpfW/MthhbnmaQFmZNVy+A8CHm06j/mPy6YeiPeClFYtu
0WAiKu1b0NgS/DjnXdTCDwBk/6RfCQGEHgA4R15CDZ11V7h6tGpA3SSg4ixvuwAsCiXsNmIfQwEW
+2iTcxY6EDOmFQOcLzXwuXwmCVZUxIGZMJ1Ul+DCB3mzJ8LfHZMjqnvzFfOucirWrPfU0kcSijj1
qGETBF2FP1v9T1SQOt5/aXwaNWR7LQ2M+P3HkpqKf4w5iT4nfOuFoLGWCwx34VlOIZgcx45bC2zx
HzGO+vcmVFCl5CCeD2kQM9apGRcF6nnM8MqF1UtScvMf3iqeOqUWIVvIYSNkGTNHssqD+Ev1lI0I
KWHMHiTvTgWAziWcKdYVCUSVPl8nxw+jhfGUfXz0xzgzMK2+7UnGUM+TmeiNwaeiF2k0WSzLh4bT
tx7MTiZ4/C9dvkhisz2ZL3NpPdY94xKOCka+/WIJrBTJTRphLzAW+jyKGOeHvCzidlPh+CYJ7ckb
hXwkIgZ5/W6WuwWqwDhngm4nynl3k1tX0X0Pk0HfWMlOIIMBv6TOQzDLV2e4IQVFokbH9lgsedJu
iIWEhcZXOeJUpWSyAaJglC6/ArWWlqMIP4+YfWobV6d1OIia+i5TX3uO59phlbpZD9p8i/hge3ps
H3ognOc0TssAjGe0FSXle4CJNpe9sPYRC2O21cZgFvMciiVqQAMh8FjdgjTz/g/gFuag4+Lvzsq6
Wezcq1qeN3PI6wd7nDXAvbcYsbze8XH4xCy5Re4TC2bYPEj5OCohTcK22ZDQCGjIclnqLUznbo2b
waAFkxOqI6TtwG+oLCfRR+U/JG8DzjbFLyS6Ts+nUZRcDC/N8nLAT4BmbQqdWViUPuZrG5aQVi0Q
0zPqswvGef8l17d/vCAPFrHIJlMehr8zm4iYm7TX2UpcuQJ/do7f+gK8G4Vj/XpXP8a5/BdwYG7u
0sSpF4hEwlvynj4cexXOOUAE3KKN7kmL6KQsj5d6svKhq6pdSnzYOWy+qgWCniyJ1jeF71g2RwJA
dIgX7WO+LFDqCf5+4q2XiXTNQGJ9kxueRqJNHjB7CUdpxg7N8loOo2W/DfiSd+JThtzRBJ3iE1yR
J2w1ulKZcJndcBLxR8XB4V5E1OhAryLHUPlw1jgAQyjzw2c/Tr1ck/G2bGDGhxvP7LLnIELVqhaz
kpu0C4fcHVEgzo2PF8Eb/DueWmPcowVRvO0/KZ7xPHchEIeDIevL7L0nd+SkxKnTnEJ2sBLorM6h
XXDTkHj+1fD1hxNuOy9rp5CUDPbVjfeFpGrn+LWocwEJlLdH15UqnPrhHjDuUNJS3t5mWa+bXtYq
DB/iOtIqEq2Ye7q3sQVtrCcV5PKJWwIfA9pKiEFGIuV4AgZEaTnX4PD4PfPZiZCAhxQUZB8rCKwj
5oTLe96BVolSxB2gKvw4AJlYYaT4FW4wkbARE1IfLR68smIWx9aRJlMqtkOCTKOPwhS788i6LUPs
2Ga2FyvjSrZnqLq0+/nr/5PnqNB72kLLfVxXRmmXAp+60q5Fe8Axw5dEf/Xpl8hRMIo+stHi+cm2
OXCec6C4/dftYu3TZPOBMqjzMTMya1rxtVyypYVRmGpZf2RldVlwIKmKRZFspS6l1o4yRpKDYnzw
uH2DQs/5i24GubObM47SkVT6lVaiZ+1o2DT14ALs5S8WAcaOa6EaXC9Pw3DWsQiaSqpagbF9eejW
3RyQLHPxbOz2oSpkIw8A3Z2pjL+imDkK2Tipbv0ti7XLykchiYtnelG4OtZ60vQgic5gmI3DuiZF
vsEx0tRN7EdEOWwi1UGJ4galFemfyDScDz9KVgS/mYfLGbyNvip3NGb73FR7y0U7QusmTArfHf31
5g6J/oPAYv42O2lt3NPoDUHPnwUZOSJdrsN3DaxTKlYagYmD/HgvQwh2mB1l/JjKYhN8GMnFIQ7L
9hNFLdVcMB+eDvRSfJfv8yfH+ZvxvDA4IwclpGzH0wW9tk1rqJIra8s3+GaFxwFy5i8tPAQues6I
6cKR5DAQ6r1nEhVfc02bXyEGIHSgE7k4oz8RwyIsr0tT0THt0Oivjn78TQUtok1I3MZMkP5wWW8w
KBl53kNf8dpiookq/wRQp+tCvO5dmhUqXo/76UoWqzztI1gXqb1dgee1YBZLlxThaHTUbj8d1TgZ
Fm05UuAPCQOikj5WjlKo8aQI4QeRZYeXTN3g4vzUfIWEIBODxw7ISkNudY63iRtE2iRYJD7LU0LW
ENFJddaYhfKHmGakcEN1ju+ED2HT0bCHhtoQV7xfGSke7LEWCjotDFoxanQkHwVLFZHjOAB+iNmN
dpmDpegD/LcN4DMAoASRDanB3unDr8KZzCfNKij9Y9uS9ZJzCj6VjGO4QEnVYreEh7wMdjwf4wTB
8xiBn0ZyRTK5AUjo8HIjtR/u5Av81BhES+OL7YLBM4cXXR/T29gRmijgmFB+m4lBF+C8FnGnB6Ey
vJkQd3mIeK9yt2UXLqqQOLWRl6e+eZtx2HJIs6kv2+TulBDLhH7hIJ5gyS/2ymyrax0i91ZzHKpm
JMLgcacdzPQZi60p58xO7mZRqM4e7jTi0b3kvZwMhHusloh8HdhnpeY5vD/l74g4KnoDzY/gAgTL
08VEKFsWaGRhbapUAGCkM9AdQpsScmp+YRaiCIA/23v1dIA4A6m6pByMOV8WBsejZfECCG1JdGKi
0B1cdjoQobqfBoOyBfimxOn5/7qc+wOSY6IM80GXdgyVBT/OONQYUlKcu0Brx4lDNcte+aJg6AYp
ebo3bQdZ/pChlSbA16bOx2NlQTsINZ3HKf4ykJ2HTvnN/sIIlyuUMWCuVWC4cfMJiaywyShTKMCI
o50jWLEkvOulqQR1Vf5AX8hq0TDtULFWs4xqQ/wfd/8Tg4iEltckf76HyM4qOuEGJl6pYBlW0wT1
YlucfC7H7OWAgfWvh4A6+FQ8w/UAkP5ISefO+e80LKrGZ1U1PrVWoCaqBuwg5zfYMxXkI3VTdd8J
MgudC3fJkUuWdOStiVB0wlJZZ+AlltYDb2WBln9BPjT1Qe5qDTZLDSDgLiZg3C4XVyCJ+MDYKLXw
ZeeV9XPCCI/jU3zrsxAG4xA4ziILVM4ItOE5L2UdOIwIiF9GEAlb70YT8vyfR1yQx6RxA1FKTwKX
rVBheROuSwxga/Vq6WBjBCfHldlN0NG3BteBcsTiF6FYl1NJVvksKKDo6HJ2wri9CIcJNz4OqksB
MZ2u+DPXGyNYNkGYmj8zHSiXCc2sVXoRAIz+TSP3yF7IIuQfFpSBKlYmI0tAJg7CWyXix7bmugZQ
arEIAkVdcLRP2nNTyXJdZk+u3JDsBazEhAuDtMqKGZ+ouxGRdrqRzVeSNYoPCnZzmGfqYFQNaZas
Ij5cQSpz9it1maAlmZB8yLRZfmwX/5CCV/CZ3RxX8K+sV6Yi/35Qlpj8asOENHyBUexP/4fRphhe
RG5oiPMLpz5qHy4kK+gZsoc1mzWTiMudRcWI92hPJmELTENR3+DdkRBteh31NeNNqvPy8mbTH/BZ
dawVt7uD7nz5WVLe0r13v94uDFlkJtCCGU74tDKzeA4vdsGpaZOMPdXuRhRnTp1ohAWXdWce+PkQ
WoY/GSn6ZBqsct3D90v1Wyl/BgsWg8MkhZgI4/mYc9VcjV+IAic4852M8wuzbDb8qULBlvZA1R9k
ilo84BAJl4uTL5v76uya82kmc719S0SSVPjU6vZCeaze7oVafSPLHqp5HNEziqz6S/ycDR71jhau
s8z7XEcVBnl4JtfTIaqzoNBw6CCDbJ7Lfr1i1HOIP0Ek/BDTTtY4mrNS5RN3d59pVSoq3WDVfR+C
IdJYUhNBmOJyXR3ZS4gXo53H84KuFb2pzEJEiEf8gnbXymn8SGvHrR7iXENLSJ3irfMaVWiOhAPr
xjhc/2gptabqTzqAy1BxQO7XiW0X4nyGX21ma0JyViMod5vGMJ6EAUbwkR0Q1U/eJJLXGi6WNG1D
j2L9vJ/LJlAZ3vFpBSVOKBdZfjCe+8iVMi0g8b4gzpO1WBMcynSrA3AsVg0U4+hXl1GW3fM/xuyv
xfKYGzIeveXvKRjDNwrzcw1FJ7GEQEIcOlWJVvJvbiG76C0GYp1KjWq+eCBDXASPbJjNpKaDlh8S
cW2cPw9pzlkw45J+Yr/jS3ayaFLy+BenFC2dmn9rYzv2Wy7WsKS4PCLn12EpBjUiESH8d9JV0W6b
4rHjTL4crvftIQ3gESLZwFbpEOGwSBM0kcz3HevDJP1Dc/nzrHZxtQ8YII+yNepy/UsdAqrP6XnW
C7o/YCafH22YzbULQb7901ya/5baXkQD0QnPrSnE383JkkqXh83fqIni1RGahP7OK5n4lZakoypL
Zm5qskYdonkLcxwk1SfftObcWzbIX0IXymkfN4STblIhIGh7rU4PrSFLRlHmBS97SoXsN1LDaLeq
WDp6/x98TV+1tuASMRjYIgLtpiwwZp9Db3gpWAfZbscOaXe2iUOPz18qlcrzLDlCn2iL2ehZhIfc
TPfQ9GUFaAy5FzJbRg+YEZc+SkehN6NSU9B1WT6Bqq4p051omJk2lPzDNwe3fhYKMJz9jO6CRjFv
D9IM+CfCVbVeEr0X3b0m6zcYItQj4W5/YKyJZNBilHqwsB7+rCy08Hgz/9sAgZl53jAbcyQuK+8H
X5fYEvOHV2No1CI1i9KV2Z8hO9IIUcyZtjEXALu4/4BfObMW5W5yLcPlFBVmQ2ybpdrttfkzrPvI
E3y9Cn/jrfn+qMK+qFJi1JavHaLkMrCtkoIXTDDBKBN3EeOp7YMjK7ExRdGiYt4tQCVhhDZptmQZ
boIWAYK9RFfx4M9Gt12hvAamxJWiQ6GJ9z0X0cF3HnIhmnraAeBCh3zhXFg69qJoQhCUkEPusmBM
WnQQQT1oLF37Yq2e0C7SFpPW/TdJPCHVm3vqyLtmpG3LJQkCWtIk8OGU94KOjZ3jaMtMJtU2WXlq
2oVF/BKD9xFUSXqzSoFr43lvxlGOiMb/6hNnOI9jhbCR1113qNRJGNybxx0EWMgGqwdsaPBtw7pz
LSUeor/YvGhq9spXcbs88NETMg1Rwbp6NIRWGVgAs7zhmPqPRa5FuiawEZ5ukd/zPQUSC6VqnFPs
7/95+hcEJH56dx6jYz8q4ERo5qHcDZ0W+IwQLc10i/ldAgQra9BZXQKnASS886xlu74x79A4iILa
UI62Lp77wR22oWdWmTrJjPNIqKaySnl9vBOV4x1R/4KBVMXZ3zdatE2SXs7YQYf5LE8TbHVat0u5
el44R41ESZvJtVb9D+s2g/KPqo5KVruZOSpJqpr2LI6KFVtQRhYb4vEdwb8MokpZPR3z0DA83KKt
6Kx/jPpl9cMUBZcQ8bWo8iLf2GiIJcEJlilLJbVU7LkIiQFwZJs7/q//pBEwHum1Oo8iUyqZx0aL
1PeBJtordibQ03UsB1k7j00gEDJShTW0++a7sz0ssNbO19pAyK12lnSLqKBKYbDg6Xd5vMNlo+5m
5M0uktcTf36N+4uFV0aSIlVm/LfSY6dvrZcjmPT25lTuzi3lerrbHAvyjCeq0+pATNMspmKQM872
+4Y1JuO5IdXn/HUUZt0Kqde84TsR9hoZviu6Zup953CBV+7P46TGkKSo3oH3gZ7v2pCAhCaS+fQ8
yb0qP+M53Rbu8XdohmH2/UyVGzlgvSknzfcFCcW6AdkigICQpEq0MxPxR9pxm8oPeKH1TIJ8UyN/
0t6Bi1dqhceZ4US+LnAQPZNmlhsmkwl/caMIegeHwHW/yVzsM9BFlp2+0m8OaMF9nLwQg9FPXLBN
KGBgZ4EGLzNoxi8glTrwAzL8N+4EzABzSxgWGJutV2wc9scCnUMm55mg43la95mBKtr0xMDvSmxL
gmVOh1xAfjDzG4uW1fH/vkpRRXI9b5PGfqZTIAo1sLXN4huLLoYoqlD5WTm6hK+huiPND055P6yz
ODDm+t5fmlXMfkIUx67bbc/O/OvUEgfnFIldaIVv0DboUr3QQAXPDNF283nur3tqALKEYDXcyNTe
Li1wWcPCYsWMcpuMCK52L0oqejPr2Lg1LomX5ebdOh4Qzzosm0Z4V26nRhLJLnOmwA1cfLrjQXz6
yiJKTR0W2vL4gJ1xGcoGTbBTYSQnRwWpKnGkDWpRCz3+LwFra79QTdJV92udJ3MFUNk6LHknYVI8
9pMNOyjlycldvJWtHgn2tkK+5D7LJ7n8i+SraEDbUCuE4HcTuLD6EYV7ZRcTMLd5BLfzGhQ+Az+H
F89mOdDKwm6ckIZhkKp2jjhIrN9jsdWrlv80GnJiHrI4EAzudZw2fTZuySDi6jzNvn7czErhLZlB
38JsrMR3dpwPhqT6zBZSUPjSGw2hYH9huSBl0EFBs70jCVazcea8noxcB+rxSCluIK+VltuHju0O
g87yENOPryuFg4+7tg+MxlEyWTof7a2ly0bP+tcCcxGwAb0Pd20EW0ysbLbRDSjjAELvjFzT4YzQ
PU8hLNO8Ad2pLhSbB1FlvRfGpmLNc6xJHlSQxjABKK3HMmN1zHuf1MsQe42IC16b8oFVOa6EdYee
ROil8zvmTZfzXxDp7YGxF56XsDHD7xfVQxjbL3nD8YsTGAyq1BSaoEQoa4KCXow/yrTQRbbkpmpf
G7KAVeaadfQZyozy3ES1UwGdR8NmzicFR74lPXwgx6mm/BC40EdAHnjnPhmbsNWZhvEhH33GxavM
WdTCH3UqIxxslgU7zkxvY6TzmhESHcTYR/cQgkZsE3MK4yqqE738cjeb3C5JzQBAZsvUSoHzD36X
1ZdDqwQXqmF2uJnReJW1GK408zm8kBP9DAagN92zFcWh3ZS4QsvU6tuKNQchEchPpTWPWZFExouR
VEBKkatwp4llGS9AtnqqwFzhz4hChZpw9Rm7IHADkmRHKoHmsA2/j+mKVApxGkovEo9oRsvat7CM
HzRkXFpglpOAhrVbYdq+KHMjJQqc4WdGisL5iVefz6b1Z4S518Sbxn0vIgAYw0Su//K1IaUe+8YD
v4XNkdTSbMg/RwbXl3hnK38zPII4mXeMJdpnSOan08s9GKwAR9CyHo5BozduvmnMeHcNkzhSS0m4
5pL2ic3gIQxYj0G8hyxKMIqrTFXlCuTgAKdvCemX/tXDOgo4gDn4mdoKMCNWLTxGXYjhL/IGkSPI
9PYtb6GblZK2/txuuMyy7tCCGiCZP57zxfoD+InRhz3zzRCuG4kT5zSdI9jIEE7AICHGB+p0kNpD
EPZdVRmBY6iGAhEV1mA26kie4VkpizooLlH8kGoADZdnTySGC6uZ/kBpmBcUcHiZssLMfo/mp0OX
lostVgU13nM4nZyZcW9CUK6qzNo3mkgal7J6D5zY7VCMYwFRSM778V1F1J/aZeqWyHaGr/hK3q1c
GDbanrGrn801uDaDfX2PSIAOVgn+0HQoF7JUJkKIrfhv8gGa3ZPhNvRzYlndpATexryroCcvSzIa
QdR85WNWEoKYCNEDFI7taPPBixk1rJr0DY5d04riUiF5MD5YiU6zh29pOt+vPxHp2A/Gzdo0cD07
Xa2Ey0y0mrs7oh46+Idj7zVZtxoTFvbKsKQ/FENe9dP5qblQPppWvWARSAczTK2kZo7CjcaItz9B
hNoZ/nwhoJZ3tbLxy5a9zSzyK5DEjfQIOQX/uhzFw/H53o1jAlm/kEEn7wMGUOBuM+3gYEjjEqQv
R7YVH82/Ux3JxUJc8xzSmZmHH3fw3rLO7WE/cvgQa3rHW8twvYQArq79bLIAWZ/RHB5sHl9mUWk4
kDBeHkX045hTYVRGtSkYVF5ELooW1q6SVGq/qILQxycIfQzTrSUzsLq5JRpQZ2UCqWJCUF3G4QPd
gqAwDtTQJu9Q3Ks4wZpU2GLgz0u/82UX5Z1H/dhJKm+89kL+D/ii0NAk+Icu9YGA3TjAsud8zcqC
btUPKCbQ/ZcQIBtYBTlPWnB2pzf0hqIEaw8jRgMTtUZEoM67+6bLbSZenfd8Zmxp4iVRdH+35bKa
hhCJ7RjGNd0B3heKy1N4YJXRtxYCdJwkUTwSQbcF7slIKDYcT33uje8HmcfRzEhXJsCJSR3lw/55
9fyuw0dIJHeZj2YOdS97NHZpZ8O9Ldc72dSEouX5a2bNYRPp9i/Lzty0CLb/BpCV0rhNPr5O0lvz
f85F/ZznaicZ0PtzwDiSUw5tBtHMYEBefuI+pXqSok2CH2UIL/s9elx2zlLvAXUucTAXizTOgCga
WxbGj8sAIoWYZ8MeJDY/NiOAJm3WTxdr7ap7MSNAbc8YGfCKZxAr8PsYdjOo5abiMrvnRhrew39r
6EDKVSpKjtbUMm6gBUonvxznx8Qi7VEBx1US9z0rBgfC7i+hzPZHh8m6WsXoIXypJfOoRsPBrc97
ogyFFQ4liIkEk5SMAMFAO8gzGTe7JFC3NY9u+RLGNN+7s/OkqI1MngOHcRjpZAdEqq2EUAmV3gZd
r3bLJ14R9ocNpf57SwRmFM5wsBmWaez0MXRz2o7C2/vNcJkuy01J3mf81D5VQERRGyCVBse/fROx
9FoPU+iehM0rpn4dFjY0Wd7DjycpgD+G8DZ5+ONZxIA2nZe6ItBlcuSJWAxVFlPl1k3RoQlcr3Vl
nvujPF4U8yZbTIqIHoc0xuxMhB8wKUlPp/fID9kmORhw9azckUdUdw+lvSlHim6AhLcuGvd+/URB
4eVbsS+1P+7vM90bFjkip2Y4pM/3lwj4c6ejCe/L0FlelPjjwCzVwKU4zlbljASUxxMKLfab9mgb
kLBge6ihEcT0QgpFvx+FCrZjGMxzATpPVOeDdyqa7mKeEIPLoQFyCyZI1iBzMVkQ2HvaBb2S7e9V
AP2y8j/XFY7l3nUNp3HbdhJGbo3R+WF6wCt6Hz0gQVJ97T8qMjiWXfUnHDbqZDjoYzm7tPdRRwcq
4of68t9OI3RdszySccPWnzPBn0Ib2uKHE2PEGEQ6lO+z132r5jIPqQzTT9hfWGu57zbBuNPabXop
kIRViKyQ0RNba9Od0p617g82ZNT+VnHPUpgcIecfeWd0gTGq0Eyujphr32Rxxnu66/5xTHdbohvX
I2ToBzqwEZwSm0n1LnIuwS497s490sbkQC8IzpJg9z2ay7eldwZfjmdzlQPa3EF2dT4FFIT2GySA
Z4oLgvnQAWnu/vYXl2zHJld6QrQwpzfabjlz3GnI/CkQbqpgMIZqvdGAjFFW9kNQP8y715azk2f7
pgy5As2fcQBaa/Epj56hJo8/y4obRmiqK3KScbdYvdYgjWC/PNUBkqSa7Zpy1NKNgSQstcp0y4zJ
FDF6D728y8jiOLCiFJrhWV+I9ZJlsMsjrvLLwRE1T+yFhxq81hts/4yvWrwUzDHgS2vrFwBV4pJD
2b5ilc/qi7q7Mse10Y2NmuQuBbSGRmF1fpvqrglza9f+T28Al9X6N5XXshe9Iv8LOOIUps/inEiu
TKManhlNDFSw7pKG5iNH+NVIU5xgzCC2o+hOEMuuPlWxnMyAPohr1eN8GdgNNuBkdDa7nDSWGm7y
qN1K6YKbS3TMkqtDjKwvHfGxgAdMY6ODOXb82YF8Bty9gAMSzoLD79JJwiqqYlvHVatxAmd05l23
jayKFQ1X/wIzG9L5flMGl/GXZvJs/cOHc89HPQK5kqRv+HestqEu4Mx7FhJ/kYUCKK6teoHMlH6g
EMLqcm1lWvxWNpryZxfoGWIAtm1uxEwaOBuZugYymCKHES3+w0cmstLfilAaGfYVmSS9otyCHff9
jRGMaYV20uCOHqTkm7fO5rYi3KXAlQkR9kN5Y52eGWzawS3pX6r+VVcIqX7G+rLtL24PU5OFxgec
t/mVCC68ZW4X8V5ELnkkgLEHpZY1Yd6JqwhExg54fToKq7/jqywm+nqsffoYABHBAohfRKmiutaV
JBZoBvuja8I1zikIou6UltN4OFbTB/7FVNcgFCyZHSGPW9rirXDVBKm0McN5LEpBtq4H7BajH8VN
7N6nTyy61drVRpJ4lY0Oy/ZWQxicVLsVOvi4djsiO1ZZ8DxGRMSsTA4hJ2j+UQo50S5OyLyA2Q3h
URv7tZ293Z94GDtZ+ct3uGHByN5/e67RU9xUqMcn3AGYVj6HoubvPEWkMvwLj5W462l1d3d7rkv/
b2uZboo5xiBxQeig03sNhju1tjY3Tj+ELXwXYZM7/H2LjT1ufD2TZSEggyPx/Ctjl2mEicLkq9KU
ZKYKCgouQAwBobzfYV4/SbKZYMyZMOZqFXhD1eT6qDq7Eme+HecyTQilKZ8CtF12NMVK68N5yemb
UqBOLQwzdSMoAFiP9jsWEyr0cBvVIWK5Diegc3rbSqpkjbmUM2pEPi606PJXN9EhX7kVpunuEn7N
S45dsrXXDklnyTt6MdXOxiODA95MCmkabvAfdMUa6HWiO6S8PTi+6fAKnlu64Ck6JnprRQSx+Rzj
u6MMLDlwozGngLjHn07h8TbdK/iVV/nDivIh7S6nGFxM0Zh5dJbx0yyxAK7tlGZ6Mvs3DPdDaoE0
g/TQFMV3GZi48M1IgwZ6mzh9gOXXwOLkTms5P4CIHcm71h2unj4j1hriypQaODCC6BHV7oUMYvcS
IjXJtoYDYdGV3Z1+jKmdis1xC/GzWDCx+P+Rkvqyz/+zCN6iq3ttUQjnNV7lrKncfRC0uInSa6+6
e/fEurSuoZP920378TuX+S7T7u/C7LwbHBhEWibcK1LAGaSaRLOOgYvBdeN+0Mjp1oJDmDfQL7me
QbPnAdJBK6z4t49TVLDW1/Yf5uMvcSjWT0RwlU3MykpSIIFiDNqg0P89QgQFiSjB5Hf1idFiHHc5
iUsP1feKeERoS9NpiEMp5Tv5WYGWddG+tZwXlaf5oufDQ15/ivl4przOgvwIpUzRpWkb2NKJalsw
gK20SGB+v9Go9fyqenph0tkW1+462WgH9HJwuy5cQoSAF7YbrRHdC+yDrC45EY8QjJ79c9JH4dwl
c9NATxIxkqBbCeo1D80DjcgUGq1wP7ZA/rtLC/YVfzmzVaTtTINU1Ykn/wV/+JSB4D60XdrIwJ44
Il4EcQtcrcrSoiAIOk5FvhORpc6538HdjKGTdviQdTBHIU+joqoLUBxVEWSh0VCxGZzlBFg/xAks
MH1fXQyGk1aZ5JOY8P3qoiGaJf1GRDWII0EQx4amB6zR5ouq8Uim4nGNeiPXnYklDtCGh9gIGVJD
cYN8uo74YdM9HYRCz2TOS0V4rh+q65NgiZe9DpvaPiMYKfsHQelEzHwI/hpUQ1dU+3vd9cdyhoB1
qD1VqtEWG/bSJk087Os8ZDqAGj4lak9M0YLDZw6ds+WLpmiN5qfvBFtOPAbppVp+dv52ceWtjhZ9
6AvCviCj92T8Vd0Tz7aML3FSsQutmlrPfxkKx5c2zM1U/9hy676ahCMa7MkX0Bdawsl64KfnjcOU
9EZ7WG6a51+kvLckoH81TXgxJxripROyI+Qk7eBOdlQEyuf1iir9uGJFW0bFSuktAjmA1JD6RtWS
pzSeRa6AHKfjrsZClJjYL1T1b9L0YS5h4VKl625FT5IuFy3NBdjg9bzSN6ywcP3/lFKAYHNDztB0
etAFc1wtNB3zvyEiaxpnng7kB7pn/G5zxXa748mevY7RLWqIJD9sl/vC3AyuexK06xt2Ku4Vgped
XmmxpkGrOcFrkQLG5knNjyqVohIFxHVPAYxvB34ZDqxVVkH80zmvOcQ04rW7yAZK5w0zwhIYcBli
ApvTsaGUsqRJX8zLkWh+16ccDWKvZv3DZqbM1g/q+Sx/A81HwINhuQNffIECVa7pEw5TZpMtvAwO
XP7rR89J0uEOptR9k7fyZ2zcVgasHSyDqcNRenKFAtobgD/m+PJA876PCPnAMqrgkKlRx8GTsbjK
awT/JTDRJd26I2Fahks+4+PJQT2Da8sHMTs2hASqKhDL8gnImglZJDT+tB+kixsSS7qPwhi2kBGJ
oxDPNrmOcCvChcDvcl7uuXAknfblHFro0rLyEsB8Sb4HCpdQkFNmbu/MkcZ2JI3KkyqHwELN/n2O
rt0k7gDIFuZgg4o+jVJ/RDq+1WSqmlgOUbBWDQDWT7NKwi3ASnyW3vp3ndYx3Nh/o+LH8ktJD5gQ
6aGVWMBAw1qM1FTDT8MIsapEP+gFCdeBz3Y8ie8m57fdtQ7EOW5FX6mUcT9oK4wQelJtz/M/DBzv
PP7oMDR2BYZCIJDXiCuKT1BZH4ozYqSQmlFR3CuDbcQfk4bx16Ndb5Vs6L84YEWog5QRotUkR9in
Y94wvT3K4f8+6wpoPOuFFaJXaW57BScuZSI4/3VGXmEVL8Xs4isQlxDGtFrjLk3qRrk5Ywep0Gl+
e3f2qCI/4n1jJC2bDUTd1WZnRqlOxb1ZBc2rokA4rVLpDtVbyzokrTmAFNpHvvfoy8bA2VNifzwa
0nptorIHpGA9MDdQFjJMdBMuYJrsWwFAha1xvPvpQf7kOjr+RXAQElWXQpUU93Q3ZKceXJplfRff
POO3FRwQdp5ixQTyE1cUP6gGeYVEoIFKzfVhSJvwez5VJQnYcbS+uy+1N9Rs1u8ZpssMWtPV1JqA
eXqDOjq/kQWEy4t6sUrwJEatBW13yPTyGvmLYY6FaUHufuxUZTaszFp3wG41KHfRrD8aW3i5PNzq
m8oNfLq3G/q9zBoZPyLj7WNka/LR+ISeSfMiOf5BpjGglfyfPwDO9a4ynvicG0TzE5/c6uKOsGG4
IseojPTp60fVaKmwWyFLAVc4Qqn0i0HBJ7GOSdu3JaIQGFlcUbr1NMYOH5jx+jJXMl1JWI5db7Nx
H2WeVdyI6mpMkAxsBYFWzM1ivNwAVH5Oz+7V/ySFsZ6jd1uMGamix12QUHrQtjxvCNMdr5RA4Kjs
6uKbzHNfnW7JSZvCV9aVxy3D0nBob+ZBBTFji4MrQiIA+E8PwXsdCYYuFFpTD5MkB23GkYXYctjn
ZJtvpB1RYgJRZgjSgfIXpXWC/SfymtXWGpTz8tqLIKqnfCxzTt74MULMFcSoa0UdMAm4nSYbOcvN
Bxq0+cyzR3wugwRjWVITh23S3O5D64HixtPAZWcSQshQ1RFNCgBJdKM1B4VRPDciGrMLceylnpp3
uBxifCcWiRpRxUREFDbLiYlKiFP96BqgOUrwclgo7pPfdxZVZ3KHDPJbgOpZrmBCdrXoQS8OD1zj
DRFQ+I6GsfVheCKidG9oUAflK1n7Xy6HL86Vn6hebHsHBzA4p/xwukLUkTuLt86uHnmK0K6mFdBT
xevUB7myaecSZDPr9wVyi/sRfuS9fDr/SBCBj/M4hyvODF/PEqE8K4uK/0q+HQTJjJd//4FQyVWY
E7uU/wBBK8JkxJ9bI8VVe5+32q8VyRsyehL31k0hkW7E53bFLHI6TImk1RkmC42UCuSa0Ju0oqQC
IvtB/LvrdJjta2s/WWO7dfQ+CuTTHOkqQlFT89+zs6017SohSjDCts8m0dwI13bL+WwW7Vocc1vB
glnMbiIZxmsZgiXQXpCA06QyqP6KB3/BZH4MDX8Vjfau3XL60p25BBrvyYmlzRMQOxnka1fpHDGA
8PayaT0nTB868K9HcZ5vGHYqlt7rEmHNCKIqN9FTv7kdzaInfZ62VQjAt0x6M3Hd8QpHPg4Nyi7T
Kvq1qjoYH+niUypPZOEm8clORFziqXLioOozwi/DK+hyd5sX91C5cTNGzR64Qy4YfoKGAIRs2Hh9
J134kB3gUp+CeuwSyuSSRDnUq7evBIxp5zvlEyQpxBwNuKhZyjGXhvd2Z684r7Iz8QoYu5IW2yJH
ZOpGdfHsoHrRIrd66PIkizm6PdUe4FzvYkTnxdLp9LDuZ2iamr+PxKoH0k5H9MAPpQhRmvBqm3Lw
U1bB68bS0dNPoQxQbEz7ZsdEx7kw9fvvUWjw8RznlUkZVL1U2sXUxcqTW1J2oaDFabacP+3bDrvg
1u22K0x8LOkt15tq1InlHwyo2DD5c7mtSuBmVgKfK/sAe4h1i4mdYCxJKVZk1IpGO40imeQM9FH3
3mi0Q6Bm6K1/gNK5PNHrARy1Gigub8sg+aioBqeE5vKSflyGTESE+Dt1Y0FOTxTUROr1T7V6nLAK
v2gKSjWPkJYmmjitd+9yafV7JwIQWLmdvbcyrg5mM1m6rUV9p2hg7xJp6k14QTgCK4fgUjYtolEl
G0X3JaKNf5RGwhlgZNJWIAX6PBry6PrBzYTpG0NHQkmJIibGCdfJv6eo+V2qrMQG9o8xiEzCk5ap
lPxH0MfdQPD3N79a70Mjmj7447rODeo6BBj7KdUcimt4D4TnS4e0l7nyd66dyeiXAjHot2qrkUuP
vfxLFDOdhpcDMl9vJHJVUAHp1E7djGdY3giWacwDmgVewaGKqulWfXyNkctdz6eTeXx40aOhbWpg
JYr6SHttycYAjupwOnu5VKr04Pdt568wtKsAhfub1RWqXvbd2o+yk+6egb5DHzvEMi2QiBB3Xh41
TnmHxIZdTbf95tt4LtY5WhSlsbLXYDXEP4hv4PQz4zkO4z+B8s7Qzu8F/+hMkPyS2jJpEAa/x5sP
rpPmrRp84kBTlHs4mJah6YTcn0RlD224h03XmCP4Ky41yFEKTuPdy4oZ/erG5YgTFS91+wLDzDlv
zVl9Af7iEDJ0AyaRIc11ywGMIGq0453ySNK3RsnRkgGyXYOQ7FJuurDm2EkfpwYsnZrwUaW/GT7n
HVUeDYDOG/0aGhgj1xP4XQQoNyyUSMR65ibqEOcxtOdWSII8MDvxi//Ad7dEI61xUPuBm3R5ToOq
LLaaBRk4PBSXqUSvbjOzKHHTBJRz3+j6ybXFt9z0FCirNhYOBTvF0f00XfUAfI8wMdnxL5E5jcqu
Me6SMWiijLUaD/yBz4LbG7nuR1YnokcNA5sF6Kblp/PiYV1hKxm2ef1OD1WnM1O+exYqykb/syoL
/MTYbnyWaOC//WE4aBZumsIzhMaL2OswNDiDsKD2H4Lz9M5GfL1qdhppEtdv6TntfCdpjEL0bFU8
SV6SyAXCVkbv3GpTh0sPa5piqQM0/8L0V//5Expwpwc84swGcBgqRN0gQrDdFhv3v4elrHWAD0M8
99muKetAnFzLV0U/BHdi+iw7t65WHlDR0kni0EUujG9BYoaGc/gwX54MSKkcJKg0r9h79B6I/k2T
n+7iovpbQsjiWTaIdoCJmmZogUAWDzc0EiEf+zAQOeyQzVN+yM1mdfo/YTZSVctPPaj1PZP/ajso
M5PZB+WdlEjtrtad4p2Xm+wuAsj4UOLqqnO1Md8A8fSiBKSyT1gcUGyNgpu10n9Hrlghn70F9GM+
JpLHE7vm+ChoNNlrX9imzsntrzn2MLYsZLJxMubxQ3tlLkE96v2T0avSOMGxHBZ47FRVl3EuukX1
4nrt6H2FXI9gBGQG+BYQH6yjp4MnVRYyg4AnmJJSR5nYiu3BnWx49WsAxg8uhyjFd4/LKH6lH76l
nn4MdhDCQjN4Sgn08a3BPmmkshqlCMuz5HYFRVUxQ6PLxFK/cgRnN48MzqDXy2EGiqI8CXn7u/lq
Sxo6VZIEgTC7RtdcH8bvKG2mAwlZ9gpJTOgKe0rvdZIfT7//z0SCKioNwHyl3+wSrYew8Pk486ZC
qWLilnU5xUPJSZyTDhXGWz3EH70LLtkoxQnJazxwplS48RoF2cpQ3luhiEEA06ukGytr1EskSyAS
oPR9HDG8ALKPhYEn+UZ0KQ2wX2M25ZgeK7Y6+ITy/pYVWMZfoYsC9AnHQdNNMO/Df1rn3t1Lhm8O
IGqEkZvmNllDNOC9fvoDjvf08DGNQSRvNLr6SE9QcAyfC9wpFkZTdYjXuzO0tWQnWqD1zJLOMf80
TW95AiMnf9SsrRewIO8eiJtlFdSPRIh5RgVNxc11dQ38VsT/1wvFRGlP7XP6Qhpxpdm+EoabwHp6
52+rLjZuy7GbOJJxNvGWZIYbT51FHekApJ1HJn4oNVFLskaYEivF5+5q3Z5ow5i/Cn/XY+PTGtBl
1yopLcuXL/1Wrp2arBMOKuL2ZIfOYvhJZXmDgEGj9F2QecKPhEhucdx3pZ3d1QuwSpzqVxAPFhWI
Auq2TDoHtuW+WNIbr2Qj2fjwoBm1tQKTIP/fpBs+K+8uJYsqjZ84oTHXLBuxVsRloIIXE7YOwfO+
wfiEpxBFVTIObeiCTBHskVZ5c3ThvC0ERddj5vRdDVs3NTnx4dRSACUzsVO/psK/4P0m1aAGEpSD
7PsZ02dNu5KP+RAHZ6ATQ5u55GtrurOC9PJNeyPQBuid74kTxlLv4L+tV7lBkt8W4nbDNpGzBSkN
KeNOOuBRZwperoFaLrm9e2TZDAzlT3Xir9CnSzdDgyPFuDtsAqT2wPkOY4pssubIinEAfvtxnDOg
2t3PwvPZWpNRqxmIW2K3ovANPlItwp1QLwJ+AzwZusZWXZKRGpceiK4cbMmpBVE1zAaPVoHQAC6o
ODST/OPl98nesHmB8FHWIhVnWnVvFYX4kxBVBaAcZWGmP2Z96sjX1EBW73eswcNkmYZjiT2DWg7l
Nmjirx5KxX8c2+u2cmEM70JGZW8ViQxSEk2VfaqW5UvOZKeP/BLAXP/zivvPaAEtTBMkQWhZbsja
LEkx1Fj0VuRBhEeiDydFB+OHk9M12XKz7XDA0NRw+p76aU9O+1BT9rQbhtHLcKzrPMpub/a1iuVU
jtQRAwnLCFPhuako3Ld3Nv7G+0LS9VEHJiNyVDufeYU1kkVyxR0OPdxBJS/YQb3IDrMvWyuKSNlb
jQdGX9njIJdz0s7W4BVG5HgQPE0Yz02QFK2BN3SRWBKyv7U6KSBgk85SqqHI3nj4tRsByZVd1iPE
PPypAaL2syFOOVU48DNQjewyieHntL3yD4koSoY/+3mofH15JBhs0j11ImotgBh/SGEA/bI4QfpB
Vs2TrDfQ790AvvXFZ0pqNrFOMDjbva9uc1s+Ln97Ru8v6eyc6d06F9JcU7NAR1xV16DgWg26NKRS
cQM2LdBgLzdiMNk99loL/eaMnk2HqXdDn3ztWC6fRPCUS0rFGmeMI1f6mfKTEp1Zik54XPYyLNQ5
yG35jDvyAymsSvIioHvzq3h8Qu3MECMIGlKT/JhYK6rcLy5w4ZtIJvARndTpZehXFiagQOONzQPJ
+dmLucG7bgG5AXIl5jchc8u7D5m/i5OMAM4nvy5fwT6BfHc1r8pztSR4XSWJMnX+K0cft0OM/ytf
7k0YIzgslZz+8EIxzeFxRN4e8sd6s4+4IUyabhfsTRSBVd01LnQeMvRtwbsY+TSatU63TDTJc9eR
si0OvHTnpYXrLp7lL5SvOfJv405zJKCLeLsiw1f3Re7IU60m0JcrRNL/bdxfGiKtmoyc4KKH0spk
HjPWsvlwN8Ybr3SJZJDTyEKDvMsFwQv5D9FeCZEc+bRgVUgp9pel6jGhpp+n+k1jauJSrFnHy1YM
jBQjX5NHWcGnDsOyp3zZWndp2675I1rM7Xu1AbC1Kk++VQHaQqjenSlMDKrCumvzI6MewSnGRZc0
Q1BcjVsA6fbfmlQWs0ddf+prehF7oFk5qimFKTiBG6lSXzWCVngpdE9WgykF3DBiNU6KsdCtaTec
QN1r1DHTPHPVc/1a4jme3r17aVM0pw1AtabLRCvmVdzpTPUwI7JUxeO1oCZd9+KVXLwVTyJ+3H2L
EvWpQhrenBFkews8KzwbsMRRXnlAt1nAnTGlPHTf2GDvMdXZlOVm6WdCQumC1i8s/omxc3dELq/Y
1FH7KP4WwUoSPP6aXPrRjq5qiWaA+aemGD8qAK3zNhIs3Sk/mePdrMQRvycwOzegmthr0f2QywL+
zbXroNPIO5F/pcTg2eni0xD6tzl1lOKzErJVqQ++0yX+GPr3fOfaCMBu5/ggw4Ni0jurKRtO9Mgh
Kc3MVpSAFYhOtUDQQsB/81ybGZobTDSiLRH6YdVdEo4TmNmRAx0UJB7mGJ372Rsfvuluh/Ng6e3t
JfAXayRNb35E2JS6u+/el9gXOqHtUJ/PP5gQZeeFXu9m8KMWzZ8XlbjIKT0i7o2x8OyZBGyiRXaM
ZUc3Ua5dJ1crGsACbyhkBjOnO2xTIjRCcMZcyaaHogYPY8NzdbJ8eq+y7DDeiS166qn7zjVjyzfS
jL7Fjz5jeCceybI4/45wpriNvLrqV9cF0DIvfE7vzBePVibMQE9Ge2f3DuD+YI4715eT86BqWwNZ
8bDtD9pTryTBLRdwnHudvfat9rvluDqoYkPzkISi0CLn4WoE4TtLRxjE0WDEPdsF18+ytUCa6y7Q
HoOBSAm8731bukzZrsXtxmUFXvEsCtxh998nmdwlCD1VOG47u+A/GXE65FEob0gPA4ISNkrO8klR
GfA32Qa6n2rFwJW1yhQO31xKkjFXh82Y0EvvspyRCxAQEWB1gQMrad7PIMHMUlm3w8CTDfe6rkr0
xR014TbG8wCV6GqqvpHQFh1Hf4kQ19cI9FqTVKI815x8JMYxuJAqMzsDvhFUwuUBAlvQmTefK/En
iJinRFm4UwN1Gl6VSoCT201eLNf/EPBt405hweO0tJ1V/xrZliUVM9jOzj23WB2Gtk5aqCV8IhXD
6jj3nvB1UltpnKwIKB//EuaKz9nmofUrh0s85OeU5vmC9Hl/Gf7+WIiDFTm5Im9fIUqgAOKrSKZ5
gTFEIHELZ7ARLyMfgb9iWNR9dNDChrO8hCR1NDqJHccw+VeW0oM4w58REYzIuMxVc0vEwb/PscJg
ddY9k8Pxj5OIMjhJZAidlG/rHaNgNwUcYHIH2Tb5WqAEzq3eFy/lL1wiy8aga5s2sQWCAByeUsE9
ctUoUz/yBJ96HBrgRh42GzCEfiqDfWMKkUfUgkQa0Rru7ac+0kj7UNQZpBDfLdYfWMvoiiR+TOge
5hQGmdDSSgSMdSGdNI7lXKT+AXRGg0Ee7zHKOrNWq7O42MBEKA56kV5/cIpZmYbN3/buzgBkMzro
nUrJHk3nrIqzUOruhNu/WWV0jSVMU3gvNey0yV3UNZQqzwluuyZa+kREcdoDdky0dEucOs3dMWNt
EkvEaeQCmzRNUdjy0GHUeYWHQPAomj+MPD8/MCikrZNfOg18g8RKBvv2Q/8/UlDijksvTrUmtrwj
Ru2ICZOdFHx4/+9WrqcoVE4ir6mmGCJXykk1zlJtZ4hX9JZYVqE95Yooc87RC/o8Evkkm+Tba2oF
2IuHiUSf3OEWDSxvbPyl/BT+7ZFtJJozJcl0Ysu+3D1JrXdAOd9uVTa0j/XsmBw7BUjfrykc5x8I
LafiRoNT0CKtgJigtuxsLx29NiyRCg6CmAE1UloMVHltl3eBjiReb2BsNMrd+PVwp4ZlJgaG2pdy
bDwWUyoNzYfPJkEugV1IVOM68nj08DoJwsFUc9DMvb29Lcf1gtF3MAFutahbXk0sgWtutgNC4v8p
qcZnCNGVLUdjlpEeYL75+zazP4xXJOYXfvT7SiA3PqVVa86NG40MPZfJ/R5+/B80wPnqlgIQyeqw
K5TqbLhRygmx4eiY3meQItRD7N9r82BpaPlPb01wcUnqPe7Xtf7+Yln7GSPyBoxojHiWTW3yFWVV
ImiegYLbF8yicCIirOX2Sb6GT9tIYSswqjKuhpVES9E2ZHIumc0nYiHDnF1vJST9NUei/2M+WO0n
s6EIvYFBjH64BP2EzM3SR5L+upzVAs/LD1qeJdRejZpHYz/gi1R+7OPVR3rfQIp2iYv2OaOXJHhY
clb41+ODDUjZeofDUmRPj3zir9hC62f9kplX0PmzfFB6h2TvhfoTWNwfxCqp1IPYDt4wL8MPI8Hv
+2FwcHMjPW//UFVtN0+H0lx4JQaT2MkhU1W7aHWfZeW3ZifrDxCCYZxnRMJfRDyhDOVmgIscpxsQ
vXNzhLdY7/QlY8/EzLl+Y7YyeZNcyBxDAUR49HROMVJJaA31TOEeUOf12XrD3iMqf4HsYnYJpDU9
x2cKXu2wIHx3X2Vjt3EXe0XF+eu7nZDwGLkv4+DOLJtyGEsYTtht6Mf2ks6BBqA1+qll74dpLVHO
jkvwt4V0aWrwzUO/qo1g3KcEXfIoSxnJg9o3lJT4ynmuDwB/TOSJSNz07H7Xj9t6/lKWwCIgpcL/
sHGQIiLzUa74Kx+z8Uq7CZOopVuwKsOmu/mudPwTc8nZnP22/K12z9myrYiQUcqldVgWjcrdLQuX
t5X41DIptNKQKwDT/LjxAl6IERPzNowAetyJC8CAskF1Flycjb5E9WK++f6Lb1XHPV/vR7hOAk/9
DKeWCi6TJsdLAJ0NgN0R2PURcPLsESkWg5TIOBGAdkSYxoFeOL9720xa5I/hBVKmDSHaYDUDUi6B
BFFW8RW2K+up4HuhIxxeTsmq2lyWzujYmmrUWHfR8VD1UaPiEfcpf6DJbGtMzKFbiTp83UzEuoH0
7josrsw8asvqcS4dGue0UAgROOLUsoCFSSDl1UWCarI7M+iV1o726PUuv08vhottNyM9aPr2owPw
vvMqe+mWVh65dCs4O+fTFcHtRvXLBNcg2IDw67cyXPyI6XeEEylKSITnluViSLE7aKm7pJawGWUZ
BYWMjllmSouyl0YUacvKdA6/NC/40N7bs2FOT70346WXJzrliRuioLhN2H7JeN9yI4kRYY86P3cU
0oMYDRj01s+VXQCLC0EHzB5twEH9vZpS6ti1BDiRylkHufM3imYWCQhz1i6zagc6mWPGJAaGTS6u
TTNfL8ECfAVUb7yse9xp/KoCkCjnInpD+9eXMYcgFT1DXT2wtN9gUvhKN7R607tUhemqu8axEfrP
vwk4eOhlGasO6KzTTv4guthqEXBDAHwe8LrQ0bieGQGoe7pdBIb+Vx7rbfTdqwXVp9koGRmNxXMu
WtAW8iWvdp5u3OgUSHGUPmSukQ7LOyEQUmWwQYmtKK6SZq05J4wdUx2H90fZQvg09CCKE7fZJJXU
ePmaky/+STgCOfLkrM8W0KbyISDYIATTT2zXZhMgS3gBbq6iUzln+8dKFrxEUewAA6XnF25jtUDx
ddnBtDef4JUrtEUc4ky8xnfgU7ni4K0sW46kjq/CnLQB9TszhAlNboIbAVzCKnd8TLIwwF2USgYO
XRRiSmYRN0bySYx6EhcoqbLlJQjw+M62A8enPUkzJnZqbve0QFDi5oXSedVCkPiUIclgxsRVkR5+
G0freBGeoTiAvDB18F+oozqlRb0huRhJbD+jPyY5mkbguKwPOYiRiR0aeiGRIrI5vLkqAVRN/3He
5J0mwaaB+lwAC5tTQAqBPeMUvoIxQ3Xf5ei//dykAKTGCg+ysGxQONbljuMVvHTh68biy240elQW
H3Sn+M3APrvNbUaBpOHuqJGP/t4MRu0DFuPczPuRGSPC46GL6W1P2UhIJ3dVoCiaEUNKzCd4flOo
8geyExvjhEqkkXNgl41MP1uY1fAth4jdFzRqQ8a+0K1gwat7hBVNLTXKb2JNtxXegalh0qj7ppIb
1prEkWnP800wRyAs1grfhp+FQ6S3QTGgM5v1/hctdo1iFTMxtym68sPposDnyvKRzY5ilvvcZHgt
Cj+Zy5HXVwwZUdYD66A6AUa2tBcTvgSFMXSZY3sJQ9JM2QbgHVTBXpJGzfksUu7qoLyji/M77syM
fHVnFGTm2FE4EdXstkxpFX9bn4VBzpRxsEW5X+mdY8rcalvnB1qIPs6YxlFYC0x4UDd5wT9li7Ks
OoQfqYAnFGrNO10F8U0PfkMbVlGoxjsm5Fqx/sl13ra5EhfGN1v3aJGTr3Yj6dAh8NZEOjFaqybG
btjV+8EEr2iYQFScvP11UdfxMuqV8bcjT80ZiG4WLVKph9Obj/4hUrQk6Cgk0XdNg3RzSzamGlhU
r/GMTOVBxpvAyYEzzI0apLeU3mQOY9R+64IwPF7pXHdwJP1tEyGN3LCDLJxYpdufNwQaZaxiw07V
ZLwEAisrhX3PzijfOXcvD37+z0uA3bu5fmyKhfY6kNRPPh3gJA4YKYnDfDXubb4ogROKFql7H5sO
UrUAaOWZ7xxvMomw2Bgl/c9aPofsIEPe2WauxnJLxW/b/YnbWCSmdkc90RXRNDzl+F1D7jq5mbWM
/xZeu6CbRA71BaX3p1XWJQ5h85GobRoUgxmIMouTfYDp0Vel02bGzpr4TwoKl8GeOvsOUcMDGXSu
+tXZI9381xkzFhhuFsCq+LycLTpHNKUIfDx07HWJv8+BBTSlkcqVJokqtuxKtwxsBnoG+3dfwig+
+X9XtxceWuYupTen2JX7Pl7Zfs13dvd4K85XnNT4jXUQ4drfiJjfD/iSORWaa+ZPoT1JTzdvCFyp
5ImB9eY6XAUr8y34XUsZ0VyUJ8NCYHNYdjWfE3VWoWwaVFk1cgqa5q2M/3oIxcmxcXZstrjr6rYZ
2I/wwgf4TL5GspIldsSQBqGIk8PVYn/vi3xEFPAY1DSj1y020xHnhzLldfW9nWiN6j5pZ7Uznipj
NqnOvNVw85Kp3SjVlaWiWCqDKmKygdo2xNKpLSJ4lCB5phOwYy93S7VhvCZXCt4V04eZ9lN84520
Gy0BOd+SapnI6C9fYUIHAkQVEdbkZdUfwO7+WJkdqHJoAmYFBKx/geJ5U5GTTucATMBQmMWCSPGl
XBFIfMi4mPiMBfkMBPQ2vSxLUqByJcrYcwHJRBiyU2o1M0XoFIeTG5QSWEnVU7isXDCwGA18e7ud
FDCvzCCAv058zH/MoDS0xrPTkELLTdchbEv6LXfhzgzdz82ZjSWo6QXNnMBJUAsntb0F/hFPWA9k
JEHTIe5dajtK8h7g3N+99akt7Drpdx5s69quqM658Z91H/5HEuBCwou8P7NKYS7D/LIyGr/iuPYR
xK6x6jlASjiVtCqlGTjW0cNC/2XYcVIVVCVhTN3qD8XIOZkLRszO4Q9/V75AXXDv1nBBILxQLSyD
We6qr0uMWqQeNd04alXZFK7uZdb/Z2OhoMybPc3y5+5FNsoDnB4AbgzwkTaB436AZXqXYl1hTxnB
U/ZUoZstL8HlgK/1keyLbw4Z82P8snqm48sBJHm4WSE6Aj6yfC/8zPcyTFLF9D7T6SISPIAMzNo8
hB59eZ0+8B/eAJGdUpTLsDwGYzWK7svxDNInMci4jmN9kLs8rLag3uEwJSaimO8i/3qozdXEZR61
I5dzpAKpOA5gZjLWdK5GPq4yk3eL5IBoYgf8CYHnSs3ohnP9d/4/0GqhXnt2qN29oeyGi+BhfFgb
3qC6/7xwhZa6bBQTD2PJY68WKVIrsvWMZizU1uxH7M99BVvyBfRlE3wDFxY6p9abL6eIFEOPSu/w
1nwCm4+x+6cmX7b3Z37da7sKpvyVYTbJWTNwwIAvQmFYulAftRYiNvmC+Mh6HIWfi+JThD2LNl92
XA/PpJIGyXVmAHvmUZFOztf8+Q2QesbEPnNaWNRl7rRVPvvC9JEPYIrjjj1gaaQ1G/0BykNPNYqd
XF9ZZRVrP/iJkJ//LWQnEhD3J9xcMLBj+17cHDxTjkgcJSaRAdkdy+6Ho6qdhW4qFZrsu99joJPn
oL1IRxuyvGfwIoKKD177BDrg5uRgiHl3mZ0l/7dy4uMxisoHm/ms0bVHx5sDyGWo48YOqKgkWmC4
pGsmY97mpGK9h6IEoZ0szDTlhROJ5d2I4K+JHQZKpfbsLEkGpMm2YYRQzWXIgl7NJwVGec5jEywE
4Nmi+CTmQ52RRTVkglxNmw3y+1hTYXGzRlblaYpKkhq96V912FOZ3254tu/GrC0as2lYYcfClmR3
qET+af1dwqaDn13s+Jm9Ukl2buhB7TzpVIVutVjgbIntFJ0A5NWcE2GHqo4O5qWLu/dQ9NrUk732
1kegt6V8uD+go4HHLJVp5oPfSclm3XzuJJEHz/+JHUeFU3nnVFoA0hImwRtVGiapHOOhFICYbhX/
W/C1n9UhatsjHadLb2pbrMLNRsWA6oB1URHoD0H4nW4tUyPdE2O6qxHB5GRVa/BxoZdSgirYhOM2
wh3AwvWsAh9TxSzZLHIhG8zKnZL3VQvuIceoZAJw+RF34L9Ersfq+5UM6VUiGkQPM+WS2LEacwyP
Elqt5GqdofB6UTc/S++FoXuoSlkz20LAQS/zy/x4kuljyF5WQ/Qd83/w3uMx/AqllrvEfjiMMgF1
j9Eg37poLVMS6lXHyQn9sjNtyAN/JQI9WO42/rIId6jhQ+fpobE5iIhsYgVljH1m2ruAcFCzwJA9
PuI9uVgPdWDs/xDixCCSJjtjeUdIeuf2NGd+gucAYPIc4BO978/PbT4G+rsPAv0sBXETFAIiSGWT
WgK+uqb3L6Ge+i4j5k1LsXtv1SnnI85olN6BeWBw5Fdt/E/vPxbPOdL80gJazKHUXPAkVgRYZ0co
dV3s11iNg0r30wkgrRNMGRVacG3E+JVGIfJdg+a7wpdcIVzZqKfFwlyFEJTEs7HVH1jp5g38LTRU
0vVVra1b5j+ZQBnD8Xb+74Oey5Hz37uzgE+5REpoMjS72/RWCU2Jz2awRIIfLQxArKWrg6GtfOWX
wuG9jlLCBC09C0XCZrNTV0WSpPaenqFZKdk+J/d7cgR6tWuCYTpRDmtBH1vUAXRzqnydDlIxm1yp
nwYwLa1IOHUkVACY6PJ6HHADdn0Grj0ffG+wrPmP964L87EXE3DF8A8MNDJHpkDcONkwv4BCZ4Sh
waqCrvigOFsS9rHHmyby8irE1kjgHFNpY/ZIHhcqJ+pTCuGKSaywvSrl8stKJpZxtZqln4cLbDu1
Y4M93TgXC1VG0Asfj5QBQW2uZIrcetPCFnyjytlmHWf0qEwhZereIi7e2m4WzbWzHed3qetFQIMP
eZxrhWbXyK2mqxYImHfHjdj7dicba32OQgjsN0RTw5GV8r3rxL+gSK+S09yPayj37UKm32NQATPh
SKC/JjW17FBbBzYf/2bewgWldCFS+T02/pCfM58qKJeHLTC8biOlDlWEB32FE96+iGA0cMQZITmL
KJdqInRsDMnMmn2VzJiMrT1WNMH4tBKVO2tPQUYodOpOUns0y9zwEPgj1NLRjAyTGCk74ZB4oWD6
ljSTjzM6Bf3k0vqfTr1dQPuXRJsmAbgZrDNOQ57y5h4qWAqCvmA6qYRoUq9txQDLL/VxMg7TLoK7
/AdKLlbQb77i9AoYGPglRfgnQkNLoHIWp8KPN4HxEcdZ+i921lurm5N7MgaG/m2LriDwfvLq0B9q
cCP+3xhnLL4Wys39bbAMJnXDUYBNJFHUwC1dqBn/1oRHI2Gfn9fLLuGi5Ak/Y+MatF5vVfkLKNSf
fptvoxX06AIaCw0pKQCl/RoPXkh31Zq6kgBAzD6H2mjgkm6B7WBje42d4Nm3ZgMsRognAqQWX7aq
TDINtRcWfcvZb3lL7ddIyCK2BQ9gYfluFnZd3cUnH6eibi91XRB17JAozvuCcIDBonVKFvZ9iJ0f
d2u1IDoGFl1kSz01i2fKE+sB0rNHZtaPEOh3aZfkEL8+ijJ+dimjfNJvRlWDttu8S60Adhj4e1m3
sU48E2YxWA+IJLJ+kTAI3GbWlUhA3k4my0z27hJhYXMik0qGdeolrb+6kOZmtKjBsKkRQ/qxfFkk
89V+7UAgDaAL3gw9TwCL86DYyeLyNh0rAvxIbhZp2nLg25Cyg78MwlMqzO5cQ2CfGOWwdoAQyVPX
DXkebD2iVYh9DU+jaPLfy8iNYnBSC04NS6ZIcO4FaqRxNygTOORuiQE9hY/mXJIz/xUcN6ojOS5d
D5lIfY6+EXY7FklkrlfKLFZ1M2jHSK47VOWhxNyjmJ1yZufF7YKpCI9XGV1r+GLDhTjehtV991kA
G8J7eaSXJ1m7dLklKCrCz2LUQUaCsGIjNGs8MKaUSIrUswKg0nfQNH1PGhh88CERjas/TqAz74Nc
tv1tk/H/F/uzmcK43ipBGOes6hURzkdWUtMhumWyH67DFYelkrZgtgxdIjL1ec6u6VrSdpQT49IK
xEFPVBroCtq0teJuZVDhWKrMOF3VaSBNpS+L/zaMTX0URl0GHjOw/QNSKy4nvRoUDnlVOkPI4cFG
hlusTvnvnmyXYfb2CO0/kx1iGVSny/s69omV8cC7DaoO/vczHSsSU+wKXq7Xveu/UlGSSjjEofmT
/G+Nl6akfanrQ3mYFBrsAziXR69gNeoDosCl6QYvp4HpoBlsfBiOxfw6J1JAzgmhALE/Nu/vQSBN
79850zPN96YJNlbPftRXc2WqlOWnJ4gSEGxO0cEQ2bZyiDkNr3c36GdVKLBM02UlRTPuxpSeWLXd
NfJBv+ST9xQgM5oCC9HDdlyef64+BgRxookhfO4hf7U3x2fCcRnoMD3VziTtGZnNq9+K1UR3uNr2
rU+mxC4Y+e+upvosU1XmpFhRC70F2MUDtwM/uP96TWAfuzzJxRpsm3HuMuMzEh/c6hhZOK5yX6X4
WeNgRio+h3JzbG3fyc6tg9wqiKX3qKnghNpnOjFdj3NKl2eiPD40QIWOmDLKDCQjhdUOzgRc//eI
zN2++wISDnfMtBOO08xO7pg5KpOOdn6gUHLvmohYenxjUVjv5skWpiAzWALNd8Rr3DWyhMzonilh
RCq/c1f+f3KGhymAsrR1Iqy8PvcyLhPDPSU1cmcXrfJfUfxshT5zTMo3f0BoSs/QZL2IviANgcBd
2WC2mbyAH0F+3Mzbvjw6388QLXQVq/5hQtFv70RKcma1no5VRreBWdg6XJM7NG9ah0W5/nF8FXFU
qVq60j+Ynnz2YCAZvzopu/tL+1AGRc59o+C4Eg3v7VdbM8NarcomUXgkUFuqaLSYwGEDEpKIuh97
CQDhrrzmYyhMGXZoplvjaiw/qa53XIelw/kpk9o8S0+Gx01XkxbZMcqaZIUkZu87/5SerRtyPu+s
JpctzBQI7GyyTPP8ohIRKvpXU2cb3V9YUI0qs89Kwi1BJXPbSyf1X4KIrJ4A4N1yCkPxgIZoIgqH
2bxl0WvL9p+3grXBykmvwy5C4IkGIl3CCHm+u6nPzIWxFoFrU6Cfc6mVJ8E5HZwYrNKq2SXf8i6e
ck40EUvjfZ3UpjkGJPMYCQdARHbHWToOc2w/nf66Ckwo70zVY8pUXyIy7uLhc15SVI85M5tOmGgQ
z/jaLwRZuzCJ7WTRLIDQnYJ1cwjZeZoSochABlvbGSaSPs/OXYEROHf5dOaDiH4571beFKFXGNA+
UuPTjf9CWLlmb1HH+queMbZ2oMI+oRA7/gJkVOsiM9BrygJiKUPOevxpCuTpDI8i5N6ep6/X24+8
zw79UfSLPxEgXjCwUYZ7bZYycfOSWBetLgJbqQ0O+2aAKyfamlYik8bVksx59LLyLij/zqZorpaS
CUmSr/OcL/SMmvylh4QuCqq2/W6ZBfQSBaS0Odl/ldrGVXHP3MhrTQeKpTOgk1+eg/vLaRi5/Lq6
I2d91ODoeK2INi0Eapf/RPnyGW3kFAWUzqsIbExZ16Qd4vlfjxohWycotdvHN+yQjqbgFRRgYFH3
fClf4Z9yli4QcheFN8L8sVH6/hggGlrhh4RB+J8loakLiCdmwgG5OL0xPWEOgTCaVuWnTPjRlQcD
XCPWY+zSxU6U17dWPdWVnlFztxJRD8CRE2ZiW0JdqA0yMnavwxbfdhL3peulUPnDsJNVxk6mrMeo
Jekn/isXqzYadAR3vPjx8eqybWL2iltLAy9usbtd8qX5YzrPOFTzpbRf9dMvGONH35hj/lilAqiT
SjAn7sLbFxjyx341/NvC/yW7vyGt3IGQ7nXpXtBWFlWWDdXYXjDPdhlS7+N7TKW+mM8lFO4ySiun
aVR4k8RixtVK6s2JF7kqPixWubmrcrWtXVaX5oDHthRq73wdZIkAR3dDYX+2Z0eYyNR29U2pRO5u
5yXEyDSFZ9Pdotb6JxVjNHI0C4MrlZYqy2HK8yX0A+mTMEWsKc4m4waEkP9LDiqKM0MCpEU8ybkc
oBTlttNTs4iCiiBUutEOJLguCeM3MwxeZagCVDfxF0FFD8vWN011QfXGKdeWG0J/cZpzDN5i8ChG
XQ0i8orWxJM8+BEwgGFSmTpM5ZzuIZWlXAnP7B9aj4iEO+JcCukeXm1RN3PGrq0mxelf8YMRt2HT
lDwz/ZRMoBWsb/q8nCD40aD1BrqwlL0NDFGQle17L7X/Aed4Boc5mi/pJ2VJGZ9GIvI6Q9Xxl/6j
GcRH/KVtEUBG29pjqaJEo8mKaUAT1r+/yyN/TG7TotwRjN3BxJUHwhScZRd35mcAlQ/VIvxpkFdL
bzwyeL9dJEUI7Jl4Td0win+nwfhItbnrVxzpx+4LDlUo+94pgtTteyxjlJP/btC08QRtLcqKzJb3
gleMsxwFwAE+I/etOVoxGXEjh7Xi3PBCV8BXTnR9UPSdjMqzWMVJm0M6oIIgbfJFzCHYCoUUxd/Y
SuIAP78AR8N1O9/snS4yZxSRHTXN1KhuZXp6Jw0UGI37TjBc7q9GMgmeiAnQvLMht+ub7kVjHtaX
zihSqn7A+nzk3MRJC8lOS2ZXnVjaNkACBtsnpUsRrk+K0PpVtdZCm20VuE66pfzNtt6pPh0MJjH1
23vQJ6yDkSUM7CiglJBSVUQhYyQxysSamMQFzcTCleZNFveYJP6CyQ6ppuJ90Q3YEClA1w365FCe
1+nZ7FDajdyh78qut5DKZDwnZoP9U0kRO1t+Dco1zMJ8ZXUUI1nHDxe7K8urqWOllRo3Yl9V6NdW
AH3UMs/6EzsYcnVmb0AU9CkFWDOYTMV6Ve8tJ6Gq1Yjs2ujRsjScTLWOzPsuhJldcea/Xk4dK6eq
8g/tzfOEsRR/TbrVHMetaSo3ysT0AElcsFeONjGRFeEsUbJB321cflRERbu4vwIb7sRhgukj4SlR
3MXqqYpKwfry0rE6yHrRyi3n2qKDH54KhV0zFgXW1D2gvWMrguN1gA+Yio9uEPrPrZmxTo1c2i+W
h8X3BK93XXAYi3WvGnuh7WccZsfQXQ9wFaxzquycgm7XGCJPgy4dmzgBLvIEU+IM1raxBrs+Veqj
w3t6YAw8q99E5yMxWsGfZRz+j/7fAE8Dd7HxoKU+GAMPnymWcB73tqKPyr7fxW0YbxBpM9onsATN
4UzsOJSoXfGIAMyBzOSMhqGZGbVhEVyCoB+pPu1XjfctwWV5MWL1PI2EdfWvkoyN5wr5I0Zh1raH
05f56IIw7QM6EZc1ZTeMnCo38YMBQQwfP0SzNCFTgrjq096/dp/gPR5IHsIaodgqLnWT9uPmdH82
pkEGkePfQ1+PYe+2XonaYmV/IYNf9z4CPS/+wMH6zyObLp73HxFv/vme/ryc1Od1wtCbrkFbJCr0
viRwbd5OW0lpu0pc/n7WTxCINLvk7nUIbnNlQ4FbZLBSS0XYhFwH1XOdghHN5pj2KlU61PQBeeCi
V6UOuRbzedqc2Cf0J92QjpuHzxO7l4HBCiaUP5hu4nDIz2gHD1vI+PtDeKz5p1bTy7DWOYmguW1y
kC1iS/SLFHUUpSOG/AZ1MsqKLyXoovGPseHxCyfhIHwYdqGToOVWqYQbypQQHX4Hfv/mwh+4YvMB
70PHzahzOT0eRob6vjcg48wdeML+rAHtsuOWE0gwqR8BLKmxBuV3tXaRkkrfAVO/dMjO6p4FdHQa
qnJAmNSAXLE6HF9XX+OYcnDHwtR7h+pUKPSZpOM417PcX9sWL6XrU7v8HhEw4eR4bwXcNNIjvVJ0
i8eG73sWTk9BawhuolL0UQAKAxJwiS5JWLvEvAb4U1MqjBIAPFv9ighoan9lA/2U18FbSpmpEacY
eMvrkDOACBj3bWfpQedQCVHqP61XZG0j0zfVNvf0p1NCdlJyjDmAVLn4Q9VNo/jaIxc/RxTo0QRA
1jq0Kgc2n0Mllct/wC1dpurOEIglr02bUHjZ5HkUdCelnmWf3EOzTS4Otmv2wv3FEaQte1Csj3io
cyY9ytKY2iNvv95D4f3WYaBNmql7d+8A61mInJO+q+uJi+Cm2GdZ5X/6VXqo34kDcMVUEjR9w83Y
Be07Bd7Vu7GhWmmdmD7L5pGRDPOohECu/uCRmdHEusdp4rrkgnWougpBKs7BNjqxprPgazjv5sK3
jW3qhdQjGIX49HTRREKDybOntQgRHa/RhmccvgQVyiUZo22aC2ndtfz0+KnsaInHhk/J0lLBaEc4
O2RI2hlkTau6vMmssSuL7PutIk2/MZV488xvtvuKQUHojSTZR5Io9fisB0nIyIL6vmSE5fynjotA
KEX2nXdCAg9mce27g8WTmS1l3jO9oo5P9uJzeW1QFPRAZ1Cg/mqoBTIWwK8xqDxfd2fYK/IABjv5
O5KMEJEbZ1NqR6T9d4jXoKHM/js9sSecJ91Iq8MtlmGQ7fmKsfxKUD2L6q0JMf+JeKTyQD1OeL53
9Q46CDgOxJE8vAjW4q95hVWxe0v4e1pYI9Uvtz0ohaMPeWSzJvCznP+J4J5OCxWGusdkLwVWHI5y
+tdgXjFd/SdUWhJv7KVu65axroT306TiLds4gBO1ydGGN1WmSihQE9tgjVk/aBH4oUH/GCUEnLC1
I5G9eNFZjy6A9fHPFp2Kk6002jI1icQ3UDTOYw2WefTuFJfTcLCpwup+fqItIyJRbC0r9oZxfwE5
9+ww4qNLV5KpVfaB8+FOxPEqDEG4Sc1MfLBnMzhST15rpuWhyyTApRXdeOoZ6UjNpuoXrLqgtC2a
pwv5TBZlK7HNQvL546xnovyww9qgTCr6yB5ajk/71BVzDUkwWxwtHiVrcbbW2R3Jj4fzYREoXVtM
SjIMa5rH/4WkI5bACN22McjcBb/SXdQ1Sr3O+aZlw48ur3wJULe1QBWiFVSd4qgxoiJbaCzEOjvo
1Ri37a1+TJNtzcfnkI0r6+icKJkX1CKnLv7Uqm0mGpDFBKnijfMYVpxwSqIRiaAfxHs0ypPJa6hm
44mwZxcnf9kLR0zdN4d9k2lXx60bV40La/lrkrMiQLThU63EsATIjiIJxgxkqUBMykeHEFLxXaHe
sXibMj3Dg1g+F1AoVInF/EEJoVJpkNfE8pj2/rMw/dIupQ8GpIqQoH749BAgM2hQkUVUjCsCbw9Z
GU/rLdIORXWbH2rfN1pxXiTTPYsv41pFigH5NdDBwIwch1urK/11IyfdWnPzHcN+gD00Q8KEFodH
unv/2rFcLSTMDAyS7NQ/Q6gfoTkakMVrOicew0/QSOLiDaHMoH3hOBYhrFrzMibhO2SnsSaRt/ua
2t1Q5TGgAR2MysySwO3ZZAZ1lZjMFXLvvo//p/PGdLu/YI5rC9et+rr28ZICvZM0c6O+m/yXhwHw
f7i0kGi2K1oKFfFj1KuBG6OA/znfSLwWWxsThoFR2OM/Y5kOkHfkMUsQJi6HfrlPP7z/tr8C06qp
Cx9wIHJAqmbJdd/ELjaEXQAKrmV7yCv5w93dN2PgIPK9sX6878LVd3qlJldZw2mHrVYcTVzybHJr
58XSxCwtGhi7Kw4ohlGM47Gt2lmzvJvueixREp4v/5TVLWTy09oNdCoRJs7dCV2POlqUOpys9nZw
I3fQqrwMhxl6RQeJePbWycv4e7ebTedS+abJMbaKSFhbu81vxMrLkZQZTvmC2me6G25RnHZ/iRcW
0PKkmEktuxn8y5UDHOYcFxg+bT4RL9n+bROmNpKanA/+UijfDSOq16ARwMUUzTwG9npTdaWGANGy
rRNpJjleeQgtR7907kj/IWRzE1tTEkXjUkCC6zZH+3d6d3uRD2hGsPv63sZhG2i6wpvnqaIm0/+D
q0KoFo4v5NZ9XE283o5ETA8OCl8BCOSP3tJCwkvWZ0wD65+4nRhNPqrYKUpzqSXyGyflQednpVyp
FmZKBOXKI/jQnzmc9vJE9vCFS8hWc9tESYBcLHQyhGfxRce/ZPczbfA8X5UUFiOZExBKGI4jgxJc
ty2IA9qbMCPNPdXaQ6lx/c5Sqh7v/t2z0yekoHRSKufRmKDcHWgnv4KWCUFVItG2QU9hNZs5Ln7e
B1VuJ9+f7BEiVQyuXuDQ9cWE2AqW8NO2jLnjqhh+ww3BbRK4oEeRZ1Syb0SuEK/yc61Z8UzxLOVj
dC+4oV7KsYQsBHuo7ixPJejSZB2Bwdjl2XdLzMkMe0c/Ga1ICZzhdayrGaJN/8ZhJXPo5NJKif/x
B8beMy3gjAaS65hEWbs1idW0QO+83tOa+dah1Cyj2V1u7JfINKiwJ53UVrJoWtfBuMCskBYDufkP
/qrlRxtyq46Y3kRR2PC2ant/6H4+YNTYKxbGlYfYvYdiHDALbaY8U0yzIN8gFA/bDG+1V4Ck1/tv
mZN/AgSl3dXH7HtmmE3GR0UzkA0pjjai+K7uhGWdtMFC9wHTGX4I2Zv4zUmgKcH9XMbXz2IWrWb7
Hun561TEPNH8xhzo5Pjvz8zj9ECVsSjNC9hPW861fyy8+P0Urb/gsi257b6Ey6ruI0K4glvREuI6
yhyketKpzoPLu9WpA2zsQtG78+9hBOiHqZNBh85e5G5rWGaxRMEOlE42QeEWlXUOm4npxJ7LAuX4
17C9QENjbUlLTMFjQkNscEF1lYf+PdYtmcr1OZQ/BlhaKocRVN5Vz0lIkQaJ5zXpVVOcUNMyifsz
8fh66fIQ92dq7TBFD9ixTXO/YBN+VoLZms5kXY3PEhX5Kb8KC157YdgeayUbbo6iz5f/5mrh6O4O
STUwqwnEXFh1+yxAcEJFw3pu4qLtqPH3E45t+B2/aI3d6PXSMRFEV7ZUqRkCiz3sj2qFUlVCFzD/
wWqP0lb2b3sJIyw5NhMroc9xbMDloohU/k0QEumQMn7kr4dGlV8LpyD9WWke+IbttG2wdtqIRmTF
NNuLvBMdU1qMG4WdqwqNiszAVCdibxdYaglXDy0rtnN0KFshu/B+fjQ7bkzgRMEw82Ol2LdCeSpF
UpuIHbdLlsBSCIj59+4X+y7axvhoQ+i4GrYfW3IW6EVdkbP0ToNCxqVokQTUA8glDV4BHcuCIo0z
G1FzJYWGoThlgQURfKi6J9ipcm50iGkzPbVilTnycKtszDTpA7Ehdh3kD3+BkqnSTVSDxSeOOcfJ
THvhL7ZNFmvvNNRgxn5xxWIJ9yTra7KZleR0pBvDLNknZ2Lj2uAgIYbY2VcKMD86QQl9K0RiKlln
l9qJtC+OcDCYWnhARVgJHwlz8mLFKecAldMX6h1QHbyz6rem8wh5sC0xwUw05npvwGhc3neKYR5L
3NQ38fr450jHxZLsiKOoOwQZSQa5eGxf5QywqbF2ARnjnopbr/hzrytEFw5cxVTdmbN/4S8bFbqm
uufwi2o6HPgLOGgAUkfuCM9D2YBa6HAf9sY/9FpRvYq8Jy98OYdMazdcnfPnmLxDEB4W0QfBCMmH
Idy4iYs6HJWrv2gCUu33WtiCBJUvLf0FV8+qQ0rQdq4VeAZIBk0DEQ08f8i7IqlN9tmc5vpe95iF
egs5jzRqv6/k6boCOKAvYATITVtb1wKxRpDkkq/bzE5qq1B6cjZZdcqgoJd3POU7UWxvPgIFyWsR
zU1BCIO0iWSSj86BnPXDvlNmtrtcCMPNuya5f7L6Sn6ansLqFg2zlYJH0a1hfCNhGmiPwdqn4KX4
W/9DO0vcoC/fNV2RWuexPOq/ZkLbR1wjsIZ414KrQ4cRMihLQFr2PaDlSCCapk0U9oHJuTitotu6
tqOsZWWGvAmrtUfKHLFj7zaljj1kGFb2u7eCHLI0WSmjeyZG2RSG7pm6+i2/PYAQaiK1YeYHq4u+
I2tZ5P+rk48q0pPgE/3kcuTbNb/iOmgRDoYkOoOq8HLcFa8EXYB4xEF2kEVvj8XUb7XW3LGahGW9
BWnfLPMgtqjknvtbc+pXmVFcY5FD64YWkK+fioT4ll9+UxBHWvkVN+xZI1ry/LIrtX0qMXEB6Dzi
roSNTBeHdeYxENLw0+AF7uNfDID/eROzp8g7Zfhk6pZ2IzJbUI9hjCN03bl/tWI/diR9/PcGKRA4
bmvlhwL5UU/dITstoSThXzZ2Db7TUZPWxT7yBlr9mSsOuhv9dzaK8Kat+6iBpjRMatYv+MIwhkTR
O1H6OHVr7VESsvqKxChI3fDzNTXIydSKuqnauV4UV/uWnSc3bOaVIvl3L/VX+wlY4mS2ayloxdHW
p9B6p+eBU7dgez/Kkgu01e3rm6b3+u6Q3vtYbU7ylgK3i/vxZmnouYb8BBk6muhP3vMQ+fm2Se8e
13rDON0zfTBdt9vjcGydVIPBHh3drioZFniUH9o15tmE40qkjfRF+7ZepAxBxdKhA5njtH1l50yH
PODK5pCiEtRK1t8hk2U/UyvjTIgiojWwlgxgWx9Yi34YY7UQ/bgpFaGm047zvuqxchxyGvlFOyTT
7Wmh7no5iYWV4kfuRWAy1QAo4akgjSX8O5Rt01YAbQOdoj65yXhlg6i9g7yXXTawAcPwSQcXpaYG
mZukazQod58A8An3/mHlkqI0oacnDNrAhuL+VzqSdHcpWbkQa3lO/NuY0WXbNaA+N6Bf9aPsZVRA
hOxnoQ2X8VwVVLhVnbBFYsCfEZJY2Hrui6gnsSgAM669Daj860XsdSEPMNVdFBjUgi6rm0WX4tkO
xoCoHzlqOFD6XnhUjHJoQpkj35LZYT7W6G12xULpVAba8LslJLfMoqz4mPD89IWpoCNCIdEThk0I
LbWLASWAaKFB2gZ7dQIDMJ7yEd6/RQKT223hwpraJphABcZEl9hoxiHnMWbwMjiX0E4hhTugdqVV
mvu+vgR2mrIrh1rpcRJXvPuN1ynYk0LWjShcY7Cr0yzKhi+SE4TzaDFkts1LwlLaKIu4O8HDgSIi
ZfmA4a63e6diZediw7oflY7OEnJKFS+Kzsdc4GqiXQmHfMAW0WjPgPQOK29En0udm49ZluyWBH2k
FSIVjT75XYkKTU5UJudCkJ5w0EtQx50tZvDtxkNkqr9N1jpAGXZIQS9BPovJQ4XfVVWxFATdNxyY
AgVwStBN/jYT+G5im1ciuzyoGurtgsIemnfbdnX8BpXwxqrdtduIsOUIhx/BN0fzAr1yslPHFHyI
OwCV5ycHPzWTWYnfXjKOOB+69RhcdWSUKgJFtwcCh356lLDob0kcDH1KgBxw9kTbO/dJXKpXq2En
vfZWhRpkNFJTkl6Ik5wdxCP/JadIXPc0lpX6buTSWPgxvYxNe/YmgBrpD1zswGaw8NpHh1Su0IF5
WJMh5b4jzpu89dFEcSU/JfGpQd2KBup557QS9aNeh/L0hHKmU2cDEOKQdPfhppAzeAAnSbejpsxB
ZIGs2v1EHiSQNUggJdPbI32OSxnDxJs3Cwzhysa/zZZzxIjyWVOtIJdHK5PZpPrhfR9/xq4ah6IJ
yCb91TqsFmihhz6KUuPmbaQNDgStWWOwGKT4KaQ9JiiViUjagg11IcL65BFZsn6COa8kd8qEBx/G
k2Jm0rGGiB/3GHbB2nSZGH9kp89uIMjdrtovAAtrKBZUbaDGCnV+sgb6fSwDy2uTASw5n/S18VlW
PfGvaNVu/b8H0oTMQG8flvRA+uc2Jy8/HsTiXfHO5+xRnT95a6oiq2lAAMg5ZgVfTyLCz9dskffs
DpQu+spMhOQyokeeede0El6RjuiRQG2GiY21sEJfkk0fPzMFqWiGB4pqXRBUWz9jMENj28jvFj4j
LkZiL5qsy7W4Y/S6GTKOotpltESApB8tr2yiHOnI6whORFezkU+3TF/YjUaQm0MgYojxPkxBGk3A
13V80VPD6TgvESdRPGLYEbfbfGSOca55cDrHjBuuZyQbZKfIlbremnjohODfSX4t6kGIEgAPOozu
5Gn+dUy74ypuJlA8WfsmKXRSQpZ52D1zFmFdf45u9RkcTxoZeB+U8P13OYyDOX1+2zAHbm0VJKDJ
j2CHz/xX35wvQbMBn+O5vszsPx2PtVwrRmsuUr47IGrvLkj7AZrHQhw2n1xg8tbIWtIETLh8LlH9
WjuT8dVhs+iHio/qC6BzIcgTjb9r9BmiNJVPF8YCgNOqPhkEdEeRl7F48RO7kpLpngycdV66XP+f
nPSeCw1Dd9o7oCNT05eES5lnGquwVLSUjTfxQBUmMk1rcqLSjlkc8+96aXMOSTWNaD739YzNyV5Y
iETWxYycm/oXuT1wMJMeoxh66NHEM9fwqdzrhkF3blSZNVNrnu8ZvhI5Rgagey/o3IJODmKTqs6B
M4TgS3gNht5sc5Nyfd5hmpxiWYlSRtebpr6WW7OxUFsC8CzTJzSJfW/8EgXkx50PLBlrfcn17c2X
hkc+6IvyQdyogRz1qM4K28Og8QydL6xYZAC5Z7YEdRzIFLVBVeSRDnEeZSSkyInnDjNpyzdrA6Lc
rHIwbrGf17wEiW/9/EKmJqZtg9/raa8Dho9QQQA2zrc7FHKLbtUP3JrjK5S5duhqfIOiSt+koEsW
UPlDx7rQ8Rk4CvjJv/QmIrQ7v3pnwsDGOlyY19C+6f1ow+KAFSlnq3C3+gG9fHja6SHqUbRlWqKo
KbM2ucn+rW8TSC8UvXZ9DQQzd5HmlreKc5iaXAD10DKUHCiyYLPDKMPdkDqMerRZlcqNYi01WrCd
Xg21sLeh3JNQGaNyLTdUAMUqR1StH519CJs8ERFT3kQuBLMxO9lRuPhQVSeAuul+nvHG9IEtMlVq
tElQXW5Cueeg3Q2hZYfYRyWWZVIYYCvjhYzSJd0Yxgl90tTa65pbwJy+U4kq8BJugcXrBlw07xKq
kgoJHg5E4yW9akklds7gLXYXKkLxP1RGvamDeqN/U0hrRHixvX5bmyCdZESyz9c94gKVw2Ghp2E/
rb+mD94428qbSyy7dTaSyIj3f7qLpzq1lFAPECdGvL5zRaUZe/1eI89OwqtDPz1VWxeP842KSWWm
YQQzb7pErU1zcctIOqQz+XVchgAeHhkqodSkNX63lVhh4o4sml01a1FVpaIn+P56GoKRgFv6ZIZV
50sQ03IBd/6fvxPFBw0WulgwRgFTm0qgJBxJZflbfn3g7yAmBPSl0YrNW3ZmoPz0DvMgfeyuoC/j
9DsEIIW3HnBfxcKWKsMLMesP1YZKNZLZZwfrbagp1psQehAHm2ZPbxieg+SIaksy2/s8vu62dMaM
i0LAKp+YEVaRCD8htRtgkYfVHVKo1AkhlWqdBrQkSSTRJxTLOyx4/mZHO/G/qj9SQ4hOBhGGfZgq
+ka1JP9he6X3SC9VYYi1nqFgE85nITCfDo1+9qLn3DCofkRsBJt3wxJ+mb/snMeQa+wG4WHlTnWH
naWvsguFYQ+loXbrOswfZFe1JGkN7h9lqr3EZpKhhQV3ORQg90FJ9E4/ZOAQouEivwjHl0WOIiKT
OfOrm5kTYYhzzWsJQ943U7h2swDsh6sKa5/HQgPEXmkMs39kLG4oLtJPSoivWZzCuBNOjSXyaP28
7h6gbNswFBFQECzd+Fr1M+oI10cyhUKj4/XJNw+98MX8D+V2XGM+mU35zS1XlYTyNq3pC4T+EtAx
Jx9o07pz+CfxFUcsmBisgjnBdlu11Y+KdUZ62XoT5NB1Heyz2ZxmE7+jLXCgyro+PuJHsSHIHST3
hWsrJrovc2Aprdom0Bynmir3Cnzt+MkJOztPnGHnNpcPcFcoDWApDxvwm1K0jLXbA2gL8PSf2cSx
NcRaIKt64lA/rM/T9m252b5UPMuqgRk8aa88E2DG4eaN5LI4R2n1OsQJM9g0toWaxP3tuhPtSWrf
fVdJPppLAft1n0YRhlupbXTSZfm9vzmm5oVbpz9aQM0Jb3Q5rTLAGHi/mJksKEZpgKRyACNoIHUA
jZDljrJGZIuiR1QOxJEyurInbnnCzA7E4yuqQZ+LgKwJBcJNfkP7fdsxr+6oYx/hu5kMZ8QKmN2n
GlPs1BGLWX7lJc3yrn8UpXuWyqJ2pSgGuW1c2d3Q2oP7vDS0eRyxsQXep51yCIm41BOd/LD4rK41
TGe+uoHWEzEOQK6mb3yotjD54gRO6OPcb30d+AVbkJJQ7KqnWy2otP4nOBXFKoX3oxSKS7nFSYHW
tlTScdAjgLv/GY33Q48ipd/QCmYllcUakxt/Z3tzhW+CK6uAKPbRWtPV0gLHHp0lh8alOsqtxG5D
O1yB1eqGVJiVdAwG/yObRMDwU8jTYfVTUopBOYyQE9T70YgYzeRzst3YnST6UqUuu2LNOSmdXtTo
WZ1TdNtuH0LWWypVb+dNmN5xKC48z7UWfCrl5aojy8ayVOCQ0Hbl3ofB3iSOytHjSCi6kYlIlCQL
EEO8DfNHX0QAbB+W6jNgVspXM1Bldn/fKmqi/Hpkzt0dON2StDpfM8XY2q0RFwgodpmd9t+2oEdZ
b9/jC9hRFLy+gy585I3XuSCxtO0erPL/xyl8qSGO0ziumc2FrNy7+GW5YkLVhE4s5i5W88HXmqmK
mS/wY100xuU7Gv++UZHAS84LJgfu2UoHDXjfNW3xFttY0LFjKkB+iEsNfOsSsebzwGmn2XZHizIt
S4H95YKQ4u/0JU8ej3l6sUL2FzfpI8Dc/ybiQPHNy0/gWJuHXUL84GZeflEKJt8WpflEvpmI0S+c
gvAE1dlZnIE+gCI30gQj1Hb77EUrIkxP8CEp3aCugqPIFnQNa/sEa4RslF5yeMO1vSiwDawXUvLL
0KBQPU6/9hdl9uMy51HEkKyyYgnhrlH0W8guS6Pb1Aot+bjH8n36oxy2HOvEmniheT4gmloV3unK
E47zMX3vXSAIA7LbFVjlBl4fzBLS9V7G/8iLNup5mf2ChYB8kT4VvvD0GERgyAqIloZ3rHTwxoBW
lVAdwfMVeWwI1sWxLxucNQJ6aQBUUx3neY1Iqnpoos9+aFxY4ZZwobpzi16G8c8/+HrL8UNmTK8t
L+I5I9cvoE+N1M7ik1SYSFyDTGSxSQLr/u1h0Y/HN3UWj/AQTWzFasvZ+aOC+3uCMDzkPfoNvRmv
0fQgUjnhz4jR7Ru70pyBPnncKsPU83Jy94JGejvB/5t3zH2wG9AH5EQMPfyY5sDQ8Jyp9p2LDYfU
d8Krwb2icA8kJHeggOvqO42BQa7f+B2j5Zs77Pow2JUWb8ZR8yp5dv6XXKi7NSb9NFwkDpkQyr4G
CdiUz7Q241dChfCBpoOxIt3GuI7AomKq+c4s3PYa/N9RegvV+1wThrdhg8YvROKLEKdy3sFYJki/
hV7JJCZPI9SCbr+RPtKIMLrd4LD3SH0NWJXNX/h9IlDwuCTCDvV9wCFoBE6wAIwNG94jbpQa7ofP
1aO3ygwmG2VnwWZAX6qNmVOqfzQg9p0ooFBqdNuvt00W/xbckG1wQfiphjPO2i8ifC+1N7hVoL0S
Utx3M4Baj1wVvbaUcCWALCCMD/rOD1SMkfJrIuGQzHZOfVLnxWek+kyTfc/3XUIvqdtwIvN/f9ut
yk865YkGAK/jdMP+LzDJmKdv8JBeqYPzy4/vyVCgXVCow+O5956t1YLSS0WRo5ifnn71C9SXn827
WKsFj1/jKlyG3+9K4MNJbTxS4sWnaCXeIUrlZKhUnDwg1HqfIgfUje1OQxKxD6SqEft9zhyz3RpW
AwoBJD/s08gIFRdFxx6xIdDgkPB33e+ZyrZHns3FpTuNXydNz8/+mo1YejtIbIu6p1639dVYLrnC
NiwuoAHut3xpSQlBy/QKUiL4EkgjeImPodBKG4RK3eapRho/Njyyvlpb62lKYlvS8/8kDMJ3/ugC
+wgHLK1fyRpEkJBXV8wDBYoxFYqfl78sqXbsgxHZivHqCUiIRHLqh69d+A4XGBvO5XGZuh7ShEon
FDmOzsx0pvbuCD50Nl1/RJeDtymuGhM+5HofAlekGEdVnJ9MDz2iK1BbmnFcHk9EZza8YuPTi5D8
AfPiKVRk1eG4/B9CwUtLugO0N7EHsqt6/aqgDQj8B8jrjhklsd1iBefPLozciX/23Qtgd1FFw7W9
sl9VO4yXZ+OpQ/wL+RT4xKz/sBuvGbCBlI+louhK2oa6IaMJED60qwuuBv+LwBfu7DLNJPauKMGO
2XssADmU1YrbcYw/9osEyBh8br5nunzSw+8b65jK3vULfOWkXxbUz7INkdqxV3riJOFcngFKPhCp
rksokCb8UiiNmJoIV7oTCFLSP3tWxCLKDC7+PdASnB1rfEzIEaFRNMDyA9gOh4smK2UPSlguJEoZ
5Wrp+zX2zUsjOJ0Uge6RXwxgkDfIYtgBFeWykpq8E+huI5LIr8cgtpiCUs5yNTKykpe7zZvokVC7
0vWc62GUWmeIEtU6Upqxc8F2MHqyVzrWwPdQGBZHVVRecRaNsQAlM4OD/xzKdsEl/YsnMVVEH1fo
ruskRvYrZjerhY77DcUJGCY+i3glQ4jN0+pBq5VGJuZ37Ba0sx4MFNvMGDLFLBiqU7yVd8F5ghWn
x3ZLKvKkc+x5QZjyxV+bsMSV5v+aMOq9HNcbKrniecmp3vGzLaJrK/k8xv2FW6K+xNpVxOit6a/3
m3JlFHDif/PcMo0ZMz6nvK9YlXWpU/2+gCcuMLulgKqhmHAVppJVXEukuU0cvXtIZ/M1ZTyZtOGR
/r/qcuQLqIafUI3xQs8v8W9xOyK37V4aIDCF6LH5dgwxgjOMVlvPs3CMFeQ51fRE2iL9bXgBfQ98
Ftm5v75wtTJdi6SXQi2aFNI23bGl0beg6EMTSm6I+EGF/w7RCA6Jf/DKls2cEe3gIhiyxxgpyWLE
LAk9fveqgxxsE0PPo6tZkjwPfXHTJqIp3bn+OtwiGYns8t02KenR47KSpyUVLIcMvrTL/LK1sN2Y
G9YWGrg882wWB43OWkSIuk2Nl6Icsx2nJRjUWiHskZIcc3o+PVrK80ihYMkMZYUZFXyMlk4FIfV6
ykEI01JipbV2ysPDHOtHNE7RSY8fxJMdNtkv+LrTXXxtoBCOHG6Ea8ISh3a5XviE9WYnjkWrjKEM
uIQFIEDjzriUmgSPisxJ25xjBHlHw/K+ZcM67I2wNWrOWu5VAOQubTzs26GYYFBNHAkEyTckalzL
RBVHVCQHRuiLo1os0BXrHKPF3qLgURScAWTmEMlWY9VmqF3dU1vgqT1gZXAxSpUz8rqlRWXc1VBN
Ioy+284dnbaL+fwOq7YwDv5+o3oogj7zUmJEwG+04LONQK7gpLmeAiOfIhvHVGh0aAgSM642nhn3
W6cc2xMYZbU50DGSCzK99DntYrtOC9LDdRckJNby7yqbtvE3XV1nr6PhNrqw3IZSbZq5hkCOvVUr
awpmrfnVGxMw7R3vM0ihrG/VJfL9fTUnSkTswIwo8ZhyYDEF6ak72u5Y5FDZPo9snMdlf2DRsm//
yilZuvvTPJ/7ISzCmzk4QWMChBzChOocB+rm/DdqMBQFtZ8rJRGvDDyl5T1zObKAuuvF/pNKSbEv
5qc2M8qZicdJrvo+qHMbB8ooFA8ePUSpQZna52PawGvFLohe98nkzI2vZcZf6Qutf5TcRhe55QLZ
W40PcNxIP6Nbflg6366Msbpi7Bc8KBlj8RVW1l4kLnvDZPjJk4+FvguRx+HAagIOlpLJDTOZRJNe
do2gJGs3uYZcu00/c8ckfuEmdH/jAgQ9WQuQrWUUa+TtWleNzlinBHcDYy/Gi4qSq3gTC3uq/GTZ
oKEBdSeBkPnzY38gDgh+DNrJJ0/uBRmAjt+aw3MOyGTXIzpvlRGF491pUwNAUOaQir0MwmvgT2QQ
GtCa8Jl/onqwMW2e7Wyhek8AVeQI88ANpr3Cwxtdin4fdF6GbxP5JJvsjD5C+PMPgpVMoCaS5cQs
mU7gCZGPPnE5HkVPD+kxWgpyZh/toSZNy8zAJTV6sg4cPPBrgmhxOhW9TZK7aBiV5jQ+MC3AZwA7
kALwUdyPc+BzBDT0/bQdKOKQi9qIFsTnbyoGiYD84Zm/EE0cviYBFa0tKUu7PswHYwW+jLrFSE0x
IOHK2AjwUH7IFeCVSR6AJhG4+Yn+Pgnni9TZGhC5bio+MFiRoz6fJ1i2wtcqQVtJTQba7LgMNe7D
nb4kubGYg0Lz/2BVUo6HaTvc5WZkHmtI9L8q8Y82mAvkjauNF9MKx3ySZ7fFoif2o6XPMVYefGOZ
qxIyD+chDchY1/knPHYUcIHRxFGQEgHYeawnYeIAPcRbBapJ1cS2+VmgpJ1z8vZpG1I+Iy9KoGkv
F26B+y9fR5gTaR+xAbo+BCcn/2yNnVia1garai0D2hbd+Q5EzhV9eTX2gXGysIAR0qwGbpF/mwWN
f5dciz+paiPEC7Awh7jgJMm/L28CQwPNztAl5Y1al6xZmdxtGGgriHNe4KUlAyKHnkJVtXptE0A8
PGiagWVSVN7eLOKyWii+qXa0/i/VtrOUeQQP0wH9u88sOv1C2rOPESNbaHzkMYlnZfIQ7swMhuh+
jFLgEPICRPpQRLPQCkCY8TF/dEbCo9d9N9yFwYgqBLWV2ki6fv2rDmcJ0C1tiyeABWrvCsjmkL28
ZbOX2oNBlkLMU4j/bnKBiwysqh/q54uqaOg06YXbbcWc0fwvWiCSVVEVw6x/d1BrYQfl/7psYSol
jVzjtpzKIfGHfPrVrsQknAf7BaIHOHT+uKAL5VywzuRr0dgPkTH6h2WdW92Ahi7huZ2qhJqH7FLk
+2zP4KxyAmdHLC5ctxQZ4a9XaFUQSBbeYppglkEoJw3RUR/s0PzO03brUMt/TfOIWHwFjOgydYjy
cceCkyow16hzuASXdEi7ynx9ltwhxS03NfoeAUZNCE6BfBaBFbYu2/oXqCEx8hQwYVUywxbeaKH8
5P0muH0+nK9kluy9tuY4HNrawrXdg1T72hB/eJwFb1bD6HHC22WlLWM/a9r9QJDkM2CfJI+IiQKq
Egr8SZE66u9C3+HuPgZgubHchr9uTeTta1nYYl19Ycp69MCg+68HxI59NEcDZnEMxxw2npKy2ZUl
d5tSUXj7z0kQ4WUwBOXsS4+Rxg2iJloY4YFU7Ae3GgDFiCAHPnzC5qEHaifEf98ntoEDkLi3VjD8
TMRrZDRX1csQo+8jCBzyQskFMKHcTmrYRusBGXTy81WuldfmZpUaIolqV7XPdMqFU2qWUD4dhtpa
IWLLm99axtAl0bFKu9/o1i48LWQLj2RQ19zCBKbtrI9giEKvL2lW17knqvADfEf8i1WXrHrReUt6
vYYWx07Co6PQno61bzzx95eHo6Li/qudwWouIvcFv4a6B9XSQpovEaUnYOC+Novz3zj9mjLILsbD
ICmRUf3XZnUMCVEv2nVCsArs1mEMVkMkK9pddcyru4IoQn9lZx7+eIrNCCYr/ul5tTDsIKuTzDi3
uO3+mPVNObvhAnu1D3hkBU1tIxc5s5WrGexGJUl5B8pYz0npObyyFoLVa86cvYi+NaEDg+gDfQMS
kRCoaT2I0PzbjX7Ilt/fj+DYWGz2mgiK3nn8clRZzQJty2agutbjRvBv7hBbW0u4K4UrPyoZdRtl
B/a18JvJrAn1c9+WJjS0fvc7N25sZu8BqOtsdZftttvwlAInHypKxrWLgkKiWPlkmTPgMNlVyA2Z
EjMyQou2ZJ7OjAAOZLege+c/s9MwGtGbtlJhGFlFOxbRxNo/vYA1ISxWKqaVoQTPyyr8Lc+9zKzJ
HNe2hzrSiG13NjUsT53YZkJ7BP0g+jHJPzLyCVYKbvetUkAb7ftPpD7gO/iK4KWp+1qQU9T25i/Z
erkwGk1AuMhkaax52G4PT/F3x4dLdEpJy/9i8FHFPZovn4SJ/oxPdTxMFBnr0STSHnyBRa/Pq6Sc
IEL/7fyO2edvGpTWZklA7qF/AF+L4SrEXQhjc3mQ0QfqI6OioviY++Al686f1+N30GZATNUO/Hpm
h/FPkQd3yHQrJZ5NlBR+2XVTUZBy54+2h8gqxX90Wa31g4jCZ6n7fIFYNyAxHxfNIkh5sD4qYhd8
dIH4jrMjBTANaSj2JXYyFAUoFT2xNT7k1Spw2HzO2g4W2RaGcXgm6706TLGFo2N0t6bTYeoWclD2
EO0GSITBRs4q2+vaMUNisxxo+WPfJ/mgvsOKZZyk83DpL1in05EFWUdhTOrqqpvJYE7+a3z5nRAY
JQ5b5bN1X/HHPI6MkWO2G60BM8wAFgfnlA02JbnpZDtZPUUgwuhtlcUyqsrWZxSy+3DK7lM6GfSI
BXdBIF7mC2RJXKxxr7qvicD6EKU9VCAz9k9cgwnLHHcGs5dzopC/DSBglRNnE2WrD89GmQ3k8PR/
zLo0YUCrP/rvZuuBkJMfzFsXDfR+sq/RnfBlbwWNFUijqquowS24NhttzRADJhnu8X2QY1hGxPQR
h8yMB4BTAXtgNgXnN/9oL0MDOpzxtKCzavGD8luqoNgIDmg1dAmkqUyFj9C5tzfXNw7Em7DS/5Gi
By3cj2oinsMnWsnslJxcfFBDiECqBqtEloimzcpbox3FRffOtpZGH/ssRQfO7aVrcwhYPeGwgnUw
8KzoMRcwMOlKt7mWmdvn5mh2t2q0genQzZfLLDxfLm74936M8N04Frrdt0yDWr1qv46bYMqhtpeA
HDUnh6kJ7tsrQ+J+l+WiFyH+wLtCAPgsXZvnHzOJC9C6bKWhpVcadnACWt8K+G0UZSMwGoaHTuob
iX1hU4T3n9PHU/V0QNmKF31YlEBpkWaVtgpxSYi5khxfBDB8+K67GpTC0ko7wsqF5Nv/RqlVcodX
mKzPUpHGbc3KZdJRSHjvu5Htx8A8bKhnW8ZlQhDusnEEY/qP8/dbel2kDMqVe3wyp6pYFaX0BVMa
wNm0rMUdsD2aBKF8Z4irnajuS3587LheZ6hzmWCM0Dfi1/5qPGPSV5LC5Kzz0TyiYYTI+Zrne2Ew
Fcl/R7/pXyb6n7Kb5psPlmzkI1Uumv9dWzfj55tIwSlAIUZpBjnmm2ovjWzrkXkaVqVav7DumcWW
9Y+rjuEh547jaJoxT0k08s5tK40SJSpSsArvSZO60sRVRJxG0Ar+UXrBAPCxNs/YFHxbeuXI+Q2f
mO5ZC0zKKqj79dH1/lplsNK+kfl5yfDKYhrrOdToGRBMhQO9UN9vMKwd3O0wAiJgtgVuAQjxwcmX
d/YEHz4uxtydTfvjp8T503scIey/FLgog5LxB+ru1fqqUkV16Zb0JtpVr/9dupF7GEQ8wYw2ZOk7
kQAarQG7C61HwRhSuU7mKy21dlwXhiR/e0fZ+hjH++YyT8Kbn87XGSAC3NklBhvI4K4kJvkNycye
bdRdt5CS6JJjBJ0FnPP3xt9nJj478ebk9vNfX179zO16aQnW6pJu7hK6kh7DetK370+wjrUHjX1+
lbkYqlAp3R3nOqx1d1xuAxQ1GMbmV78IqValabFGAwa33XCetQONdT1od+YUCTwmLNwhF+FTzxSa
4LSv13zlNwvs8Ii+DI+R1EZ+FepTIS2s6WUHTGUSKz8/yyfcv/qpOZag0QHpXLzxdTHh9vOxOtAn
1t7Xw4hqIt/c7zBf/088S0FFYX/94eRuh3sWlZZNS/vlzqNrK4Zg4CkzCnckgRnqEFtEtyWkQsnE
U0rW5lmYuddLdGJeGoORYaS/eECUUlxkld2MqmO5EhitbTCk9hFVhon5d623qibklCy/9MSYrELk
H/STQIE8LDTzFMV4qkKsXwFLmI1J9Dc7lcQLzI1Y4IOuXAEE8AVo2fG8Q6WFQ5uQErW053L1zmXo
Gwn0T2n8jIMHB15ZkgO8YChdRDMvyFtDwL/32FoRM+UsqNNll8Tff4xk5Ejl17ZWt4SDDNdRDIql
cNryPKuUXOd9FPusx7V8oVPyuLtnVmbQW0yhK29I/hPJQKGsQOt3PU6aWwUkDGg/POwg8fTGT+iy
vryLgYnDlb0Bu71ScaT6NnMA0ABT1W3htyoDXcKWvW9GEAuxNmuy4oAyxTdMijKf/C5NPqJkoNQq
Kc8d+eKtiiICmDRbMHGEdzgmoNp8qPZL91UAmL9EaXo382+ZarQILmTfuCm13CXjMJn9OOxFMNOX
2etIWd21OTCTfx7GUVYaHKqTDOF4U/6QERXGDWusRf/XfFRmGpJLgSXfaUczhzyGR0T4InvjAhsW
QrQA6HSeX5B8hRnWUncEporYJ8uBgL9nOjjmr642i+4lnNFoVzeTYk22NIHD6bqFFm/RFPSASdMN
tf3zzmqoemn5cYlbhmPyvzSt6NlVBOK1AbGUSMZ9flISkG4yceQmmXAlSJ8dOj1/CauxuLFjVe2c
AU8Pni2RwXGwES2T10VKLc3Xow+9JvtobefemiUVUDQDhqMJKcKRXuPprZgmKgG0R24mBxyOUDnJ
eO4DQsBZ/OXzpvwSGRH1Mi5kmmpPrBjQLR7/6lOe8tpflyL7pQ2RRfzxfcSpjYzoQtGpJRtwatyv
UJ1MyBNT6rQH3gq2jZ+yp4+dvzegXwDj0YUYd/KTj7RgFr9AK42Zv6hdsM5jPnrI1UE7OCDrUTHz
5G9PVqu4/7xbqMms5rNoRS7daQEVwuFu3YD8dbEwtwp7B8Vfpq2F0VXYEWfzY/fWXefQrDXhEhnk
9/9m6pc0sSU1LHpx/QueN0ggG9omgCSghLTo++Nj07sQSldZ0/Dng2mDCekKWmOAhX07qAvwhTh6
yxifkU3Wg0ITqmY+ry1OuoZfhww+otTzsSJFY+dhUgW4m1tCzhmR8XQWupLp82bLRM12iovtPHKA
trmh1bVQIis5CRgpdEt/mGdPn9cktgmCjhsZX0EvUzV27+J19q03wQ5bAUI51Qs5Kw0LeCusoP4b
X/noFJcrlZFpEwvfUOS8tpDKM+6gej1fs1FN/SLkTBbHd9Jm559pFVKBAtQ4CljO70IhE8sgemCK
hahbtuGCXlPaIV1o2SetBF2ajmv2hHF1vi6QhE/LZncZhu7dYGS2zGtotQ0lCzuQX4SE+ztIFEao
qxVgtX+xvYbsmT23M8hOzTkYWeF98+i/Wzo8fRBN5ph7R283hEJFAyNMvsfbQwsZj7110FmYysRe
LuM+52gmC4tFoY/c+P3zvpbD6WgLG/4m74DRActTqrDz90n1uA2iN7qQK1I3BfOMsDAn0ic47Aa+
wTjBbDgFWFcCaln+jb1MyAEOkC2Gr8eKIArt6qO4DbUuzwERQrL1ZT8s08yEc7yzyRNRI8kEXCNc
qZ1vFMJg0lxq8RFQJr85ipkFHTwYjxyfenjIHqLfrX4Jg5VMhfsoiYW1cPGkKU7yZSGQWuEQtSpM
oUOrBid0Pr7JU3q5tnmMUohFqrAnSTquvPvVj/TSJyYl/jtkPBELoAQf+Hgm8AZep9pQyMvHxKMK
qK1o7Gm6NiTQJUbn6iMd28Syhnuq8UWwG6opceZYNS9qxWisr5gw0Ec1uspp8HMRuqZAgQTvAZHV
QkdQzlo9Ihh6ElBjhKBf7tX904HFFM4xgTW9NmPMiQELF8ME9Yu8xOuFxd+qZqGjR48TSYoPim6/
5fzsNqN7TSxZLS5tWF+Ju4JhlsD4oLO1hVkrfDaWxJWGcJxon9beAOu3+pPDJo7CJ5NPVTaCEXAu
3yzTVe88ZAcE8K0gAL7HETzpfOQjHDwoqBEtUX9X77ymEzYZ8xcoBpmpkF9HkV2bcc+yKJusRpW/
+15m3P679F8d+ie+eEXFV/vDOUmfmYuoIfbtLPd/XAru+DWEEY6uqSJlEStxf9QDknMWdVieCo5+
UAVu4jNO/6vEvGKPss+gbMSbr2kd7scsT2TLQeUF9zXcl6ClzxlQxbaDJ35ql1pD077ovcCNOBa5
JedGkjvD+UOFxtnq2z4WTF04posOLQTCwNNPZ5QogIqwGxh5ZjlegLBowtyOBL44Zlpxlpl52v9h
E9vIb5rEffMlX+Lh26iFaEzSGk0A3AYupWKCiQshyhYdnXeqxwDbFfFgVeSxTi8NbJlsaf6lZpzN
2z2EOyzCtv/r+yLIaMvWwWl5U5L1uKEO+yxShxtQ/TPpRXZ01ppkljgRGXE0pMyMQDZa2U9FnPr4
JbqfGAiYHcsU6BDmJ59AzWDhT+a3GVNbt6ysEZY1KYrj9vzZG8hOjIXL94WUiaxGEX7G4qghcQ/O
kVQ5fzRUBvMMP+AKaIYNkXK2Ml5QAKYDK+KqCJ8lll4T9t+gv6sHbk9465d5cUVNk92RtscQz+eQ
dnRQTUjzJf9DyHOIbEJmBuA1rlTD6bhXavXNzIxr0NZV7l7KpxqghBXtT3QLrdD7bW0o+mvY9WDe
5hrl6qLBiXbvPt5e3scwRJsgfUlAnvsLFPh3rzgBEGkHNhY3ZgB/MHzc5026TdLY8xz0+4CLpVjK
RGTqaTXjz2QIYiSVMxkzF56PG9cR/MxEKvHrXrrWm0WQFx8t1w7b4hP2jCNrT1yNvBq1eVu2oWKc
4/3itewMJmCqbb4x0qg02ykBYMQhN5b6K7fGIfqckp5b9UkUgcCV2Und/mweU+0loOUhMyYOxUxe
baBL+W0j/WvNqoyhog1KZ6EvZUl/L9eap24SMZoeQx29R8BxNHg5F5I76n0JYehybfpKejXyB46N
gMQZ+jPafVTVTRU7YlVfBV09GqI5FUG8P4euZyFNW5uqVAztJpcXnrcqUKeNFC9US013LSg9kI+7
vS/Cu928drDEaV/KU4/e78QLVAUFF3PIi08O9AzfnwPPf6qajAxqbbhBHKzVunYsdb85jMnCKf8o
We6T4Ux2k0WgMCo6B2rUW2qz8CdBlZq+1niNj6wTeQXVOohoVG5DCjagjqlVSJknvcoUs5WKQJi5
M6QxQ6l/B+gpCSx2ugzeshcpsVFJ6YzsdUGwCfpKUi9sOCK4XRjg0WK7Du+HtZqjHZhetq9tkLXN
4wLUaHQ4RVLlL2YShmd0e9kgHFAass7qqaHpo23F/SEaaiFZ91CkHloElgqahrwfBl/peMWLK+37
zNQvESZfUBKqI3nWVPzAQeWF8NRQSO9wtgCWQvJvqR/haM+ja1Zf8AIrjerDWK9Tqi9tg4JZPw78
LwO6G/K8QhVlsuGQoPFfI8FqO/adic8tYofbgSkYj//B67aubjxrQEyg4X2f1XhC7/Sh3pd2VWMw
Bo+2LxvFrzBxkwesvBePL8InJMXh8cC7uEfBE/fvLf4KMxFp0qWpkvnlBOEVCWlCchkV9rRttBu5
CMUCzYZGfxOy9XbTcMryML4Qch5UbtYCEsErC6OjY/uIBWHr3XbL09DsaxbTUcINEEgVr//ujWKk
nX5ynqbGRZHFqN7FwaZqJQz/5aIC28QrTMSFFRRsKfDDo3/480n12QjWb3wX7P1yoAq0mz9IJ6+8
OcjEfb3V7Dt0PBwGeqn/LR0rk77/c/sSDvA+xR7peTi36Uym6eifq2W8Mb3ieM4DTwfj9EGUKMNz
tVYtiB7fvaXdvrcBOWlYUqdYmEdT7UFO6CUKeCU+J1WdZfrkYFqJ2jkdqpaWgOLiVOFamCIaZUFQ
jiJo6HVBmrFnGS+Q2rR1g0E/Up9o/beArHTyXLb0xuUI22OnBgrCKzg/jDU90OFciiXJ2EbwkPqD
IBDwqMzClvpgwgWHWUBydf7eTZAdK30Q/12E+zZ+lOCo0h2Pxpz3EvfK63khX7lUt1WfigFLhdFf
dqmMQVdpmggBLmH/LQJJW/FvTXuGOfSaYs9GrUW2jwNKID6n14/S/vDMEOs6bsjTYEeH7fLX9+n0
dH6srZr1a+ADA4cAMe6wWoMWiciIc0qJceIBIZs8p1YYCfNqRGqRZL2WBLSr04/XlZWNmR9arD9Y
p9YnC3BQP5s1kaXaAjdO0aL02ePsY6SG5E8VC/I5NKBoeKDaVLzEDK4gEJb29OkC7ZzsOvpj6ODm
Dtdox2XcRC1w3ya5kh0GlLKZAFMzbTKfoofBd/E53DRkwCesMJxeoNE1kiy6uUwJWP7Sn4IGYIy5
3etk9+y+NNLfw4YbP6XEsk1pA4bAhJ6lxkBhQi7Wq+f57ynGatv0DEx1O03PsNsyQXLk0uEOO5AL
/CB/DJYwp7kfJMaP9ficzwTFjOtwDh0M1Wh5G9eBQkskoCzohrVPokf219pUwpzxD/5QAblK7gPO
5bsubH+wrwOXJg49T6uqynDLgCxo5zZHsYh4YUTJKwoo3S6OR9ZWY27UtebUBufm91JBfviAWGRc
qZne7ac8WdTdcoRLUWKM0+xdzc7uxY/p3BvBQ866yp/t+je94qatg1qvBHS8JQ1aDflkQ4tEJkt9
XkCWfggFBfXx8C3QSgqL1ERWedAACc/7Kp/NHILTaD0Du0HKJlQcJNAJaNT6j3p5wxvHnTDTM2j1
+RyXif568ZEeInT3RBscypMRAWP6MuWU4vi1wNA/07gjeLXs9OW+ZOElhCnWA2ZZEDrV3brXraaz
8yJ/6L1vo6OF/eXLZ0y7OxGYYuxOREvaQVXlPeMImRyT9AWHmt5O7d0bzAfZbL4AQBpEkI7e5sJr
s8J20AfXii2uQhbh0qcVprnzZOjKP4/32VrmeIhCEZmqvTFLNQiWpNqkVOR11KGpfS8IEQfcTfFb
nWZDMWpdckmQ75rphTktSQq8tccbPpkkZzbB+cAd42cp7di3JChlPTia+wT2aT+0WPMYSUSV670M
tMXmgWqyTGu8y2lJVYDRc73SbWWiWDPH1wbLoRZajpnc6w1F6R2KPNOWn5toG1YLzOBzpkpJGG8E
Flja7YYeqN3P4iJaZUEBjWdB9YpQbPYWBWIoz2oQQ86UM7k8rBNUFSM9FpqIF7IQYqsRzh7ok39u
BGVKga4RzZHEJ9mYeTAhorQ+8znboGhetRDZ8Vo+PNXDMgGcpoEpUJBS2eNpIfyfgVwSTGvReiLd
ox+chDDBte6I6aLGBlRkiDUn0V8LXehHK8sNwSfsIUoFC+803Zxsa+F70UybYcNUd9GYEYuXrxSG
QhH/lg+caRyDEMsA9aCs1jhq5FRp9XmkvQUBnj0EeSMtsUssIjPfWyoIbl03sqQ5n0+MeMrhk7j8
Ai6Tc2QjxZnde144VDc9xq9z4YA52MOZGlpvYUkSLnGm6JE6REhA8AbvXVXLm4eFE+q3VshsIR+y
pjurBEFL/WjS/kbuOfiG2gQMxX4prmWHzyUmKfgVbwzuwViJnXLj1zOLFbDxB1o3vJiD5O8Pk/oL
kMIspZHBpE2YFe/jUUEXI1Dh1trnOFq5C9bB6VdX81htjJ7rAA+Yhhbg46ebZ9l1n/6lReJ/ujMX
ADegzOdLJr1yIjMb53dR+87PSwann1YLF/P/VgdgxMnybI3t/YxKEhYpcRRJQYk4dHyT9uyOMpIg
H6j9KBHDO1bLLdYEtzqJolg9NpzdRhOjeb1hBO0JJHufho7u6Eg1OmgZPb7Ox+732NsloaRPkvXX
jwjsRPpwa8I+I6oy4ydHM41xOxqAD3i2zJRZw0fX1VLoVFMMEm65YDoSP+Z7VoR7f/Tw8UKat1ja
2Scvnr6ypdLDLYG46Gz3FthbseROs9jL/mttAPbQiF1eJQvaEzb60zTvYjghUf/SX5F/PdkFEmW8
+c2OHDbH16HCOwr3mxacdy5huf8hX7JFinLhcLGXod5abudkaA+uHEVRNxuIvZ/71SQpuRJujCcU
IVXFLlPDZAGDZEBErJTZWNar/AhDAqI+HSb4ReA286eFWsxB16vfiHkqqaHG3QxLnjRSo/WFXogE
aWHCuCxYF7D+7Mj62Vwj46guVeqkinsckF99zlX3tdsgYqZgHV/K7LBoZMQcoLIUElMExi0V66Fk
lvuCxvJk5VrfX7DGSXp4CuuBHGYFOqBvXeBBerNDx+ReHS4lfDaQKYYcjROpe9CNxb8wCRS57Lrx
NxtMlrobz9M4Un1Kv71XNPH0iZFwGxIk1/18epITjuXTW6AV/a/sYIZOdaVIMgf8X/Yt5jVZimHu
qKZGD1F6mKRiZsv2hbJWMz2+gDc/stqUOGgztInCeCmcYsZ6l72XMVqsiQMTVzu8rPfoLcx/4rZf
OnQZn54V960tIvFKCFtvIyYNHVIu5FB+w5NAlFa6tRq6bZ+pmGJ0yX1ozRH6ofGoUZMTUOEmjyCv
KmhRjUWqwD4v2NY9Ovp9ZkXkW8oPSOy9mljp9VuQajlCQhwtXvG2z9TeQAiCxfoN9gR6IfoDoWuj
4d/wcakmVLikO8SOss/VQMk/1KJnudWV65JzqhqEUNKSSgLIFY1tq4n63Ah1h+4AfRHFuaqqNqTK
t8WfUhEz4NJQUTeSIpR2M5NpxulJcJHGu1aduh7/pHiaVVQMFEcT4jtTeA4G21fm1acbNnEDPIlJ
Tmi8eq+Qpacbd6nJ9dUaJmQTAOeFmEkneVTDmNBqAVuL4Q9rHPlPLZDbj8rHrXLIGBW703hzdBQO
+YuWOCGJqNY645tmqd3OrPLrDu2dgaz+pD7dvzGANT41ORaoOuaAaJy2RQHofh3NdgrP2fj5gV7k
Neqw1Cq1OrMZm2yHeCQQb2ECAfjLsuNFr+srpRu6mDoJJuMIHxyESd3CteT8MZKMiSmDv7frw2u4
ULkG86X+JhdWpbLyRJiHiozib0Y/1E7hrw1o7ggJswfBd/yFO1v3ggPGquP8eeIDuTJF7ur/f17l
w4+p2JdJIVBfHcGrz6Eq9nEtAa/PruK6SQat7OkCs725/2aLdgBqR0d9aCfxBk0CR7hKKn9u8CPA
kNVZrA2ln33ubfsvP86v9NQNufT9afFzPaZS7yKE8Wa1CW++jrjCPE+C8rfNJirHvJ7B5rzB3VuG
IYtp1xLZV4LF3ceipUsqnoIsBM+Ql1SS6MlOF0mzbJj+9xHJnW7ZAkAIzn0+jOkwMcFFXbm9256b
YCA7vIerk9Rt4ofJbf7NgV1XebKunVL82aR/CJbd0kEl8dhYfgl4yYZNSWElhmE63InwH2MaUzRJ
L7sGOUEl3+ggFBTszvFeBlJVO2WhrlSBIiKCPzfyr24UZMfLXyAu/3PLV/tnMrlVxuDWOny2yvxw
ABK6JBEqGB/RFwL5JC+cXt4nVZZQQ3ng2Upl9D1kumdzSxH9rkFFkshWoDWbMz1aOhMbMCb6vBwk
4d0qgtEqOhfqO6TfEMTymSFWq6GyGobKTO8dhJMVjcqSC+flMx77afsZVIkLL+vrzF4GHKybazS1
ZQW1hZZZN/ZdYs57bD12eeBNz2o6bTs0ecHkYxmr/eEXiB6/6SuYMpbpnLF955kTotXKXoeskkZN
dZkyZpSlhaimWclIlBYy9+PUhgCqRfv09V4CbdSPo1untAaRcayofv2Yto8nZ+Mg+IB0v8+jN/OJ
7Mbtd85UIzflDSkDgQ1VaRsaA4ObBguh3c/vB1R6/oZjzNxDFxsTBdfM2bDqxSqFDWhIe6QiFWxI
xwlbhQPdQH8Rb0E+DVqFTWOPW62y89ezfY0LlllapFj5UqSYceiNAJuMbAc0x1aWZfuuuURckVpp
rNZP1YgT9d12JBmBfdqi+Umlk12TvWjQWDdbaYdpN7EAyVO5e1iOektZuxNTgKfR+qqDTG5Sl4pc
vcqp6FHmcrSpYLeCzghpn+A+BJKPYiYOCIcs1p4w/Upn4Jyz037Yps++7nB4fiFqI12549fEFg4Y
186qRTZAHLC6o7lCcJ3rgoAo+TOChIVRA3BuUF3rUp8gEtBHkqjIrlgfDHOcW2SiSATswD9r/41H
medZC9qd0hSoT4ZNSus9fO5/amYHckCxBz1j0/Du+T0lX6D2y2zK7xNMxKrK05slzHSdzD4l3KfT
cluOD6nIRcQ9eq3bfgHL4PSc3EePP5Ap7GD2HYfiq1CuyomaDEV+zCx7lM2slTIbLbo5gjOkKTN3
AKgJAlirlOa6DBhihNwUuo+U2kQRdRSw6hWpmRlSDCObdu8+IMK/7V2XrPu/ev5mjYF9OJEkLOOD
nk6XfaXEXiNuVM06k65yCkAsSSDDQhFeadg0lL7rY1QqywV6gHzfiGVxf7XTVaHZdGWEMDYTAzC0
cQLt8nz4HXVCpIZRigQNjjX6vaTQ8RhDwbXEUNo7ynuERQvxRuUYqBWLp6oUWhmgKoSuB9nllTh6
/70T2YhNQngASZrOxqhxPeNr9ErMI5QI8GbEs3MdkeJoFDUIEtFAbHqLufLp1Irxbb6ubRjuUYsP
IVLuFSsd5O+VWU2dJAwvLkT1j+FpXRDkOST3t1kUJH/8EKjjhWrP1LVlYtlfypLtKQZyTNkWxysL
xgnWyBrbCdJnjFXSM3OlVZBkevfeVyTM8H+pqCvsbrws7RhAM3Ey2Gph8E6gd9T/PjrgCsZwdMNi
xNTLmekYMAayqpGO2Bn6fijGAf3dqPZyfD+CSbvebeDlfpyLdGxbrSQ1khiHBMRJed1L80WOde5H
aMJNz1LQt9r6H3E3BdiqsnglYP9RItpQLjfusBeLTsyxhdFi0NW030oeNOAyPwWT+A9mL1BmtuT/
z53QUTmtVapuEyYA1fokQPwBM7eqFS0txUm89nNW9aZCp/+UKPpqnrVPhS7ncWo5tAPw81rW4qIH
gYxZiaI0lw09oVDZ32LRQbFRSqRO4OW6sQVhE8tX5/gHVg3WjKQaO5iEMWVDoMxkuVbkOEKc7F8H
vjtXUI2qQ6FVhrtqhtj7NIBw/B5QTkoFLu43Bb7B25M3msJWglxOmfeD8FCsCE9C4PGeGy3Dbahm
5YGnDE4TkqsdXk0vK+snvnS2gKTqzIR3FDgltHqDaK1l50Y+L4YRam+Aj7i18/OSqtiFZMeg0lws
COpI/xRwC6z/CGvAQ9G1N1vnJ6Vyt858qdJiZMzDsrAgmzj5Am0C4OVZkbbIp1a67MVUKj/cllDo
5cBn9VSWmQiMiolFKdtiGty/b2uDJ9DhXJwZ+8wDlbscgjQVC9DBcK6/V5S0VoWJtx35r6D8J1Ut
AFKDz3XBdjlrkuziOhRSZc5ffDSF8t0MR3H8eobnD7i2P6oPla/brR6HuvzLWabs8wmv7gwqkL5E
pyKJvZ0gg0GZPLP5aBVdwL3WKhHox9y5DjS8NXWFtktHIvQUv6XhBrIBohp6PHT4BatyGqVPwt9V
lM05tW4BGag+atHlB9+GByeVdf4N4XmLJ5qTLA/gVSqlE9XMKl39g/49mci86bvK8qpQxXM4cJ8d
qH4pitRhZ3O8sQhfteZ+6pfyoZkmIIlTlfJ8xxMurp3UA7VIWcqfysfJh355t6wML8cSBkd4TPf2
9mEmee+VEJKIJi5Cl5egaTwdQhfIM/yzgSFrIuMZuWWq96Q3KHx8XJiNsYtM1oJVcgtIittTYQEz
8iqbAZOzvKRlZp0fNsQ9/jcY1hLbQHNK1Tfu9TP/5QifJwCc1wXPMsRCV4r4vYqdYWNBfMb2//iD
DAxnywbSSwL9dFO9b91QiRyqf5L/YlwB/2jhoGWna3iJI4peRo/wQfVe5KzZo811gZLeJD5SlfBc
dXPhw5TpNomgJkgnU/o5qLd/+3nOe9JPPONBXTyF+jxkfP84lUTI3VcQS9ACo6b2nAhg71wpJDpl
IagnCWjagB4qRKzRglOYURW+4wrTfgnSCwi/UUYuU4Zo5/ERloVVloMblpc/QzbNCW/gyjfjQUqP
d2SfKvSp6zcPevXnIo20RVWQoB/WH8D/vOy1lNDu6dqe3Wu2FeJy4eiXpwiXsqyUau5tojNnuKJq
aQtd9mWzoj5zpwZldd80LlcWDK9WmIfMWJ5hmlqVYLrhzTY67A7+wJk0dYFBTPxY77XJ1tEz2mYA
Oqj9mEV7jEM2QIi0a9u9HZZFb2bVJ0gfXtNl2OF19PMwWaY5EBgkZxbS41zKxcfq5PPY7JJ+OfX9
BhN4ezrIxOtOuaREqr9XUUxwT+Uepv19srt/L3AJ+BS0YGIhQnU/F1VmDIe2lfd4X0GlwABb4HKz
h4zYZrCrRAo6d69/a4qgkBYGTZlmKsX3TvFKcxnIWTOUDPMpkIYxODwvXuceNBNQ6gIw82W6v1bm
4kd/rffCdli5KWNPLPOgQ7p7txQAP7BOwbP1i7y0rgdhXVbjg9+twOpv41PBpxKHuES55yYvT9Qi
CZaITwIPOB0C+XLrDnVekDJXLJo8G1l/HToeggnOldT0O42kyu5+mq1xWp3TQzo/Exgd2waX+PZn
XxYyCEYN6/daiQLWp0xWYa14p6On0FKFN6UhGlhfx7d5Q67FDQPA+tE/wHPwJXcmgL667Ytn/NXa
V7+O0gd+jIRKuLfq1yt5LFC32IfpDoWXmJ+Y8nEHdyabG+Jd4hO+2RoHEXdBi6QwtanHfbtbQbwS
yNOoQVnLpPtG54GzMvZm45NWRWeWHq/esFLLfoZa8o8gRaz541ZN+ewjUIXMAQoo7x6748ES8i+D
r6Xm/ZMe4jQ9dhlFaVsum6u3FlJ+xexlkwwm1I/uPGeaROdD7YCmsckiNr5s/9OnfyxfZ92Z8GrH
e7h/mj9juen2dNhze8X6crtWwV45cWaz4Wh0fD4/go4/CgR48rlJXlthruY3I6ekPHVids6SYvC6
5f5x8hewMdgz+QMhcW29l2bL6tVrkuzfAxDQBRPMAnCQAeknwvoqZ89k7J06rWNJcjVWBeeSk7YU
vEwXu1mio+o33iWKB7zrua9FPNm/dv5uJ55eGnbsuMdHXf76BpZEiXGpgH2FdYC0HhwJILdcYBOs
GpDXbCGzN8OS7zfM9VspdnbYrioFp3aW1afxWW9o7ToQ0MX3JeRGUnlDcEuBJwe6SAlBrruIGasU
a0Yl7yTtkHaW2C9cKTa/AXrAtyHjPWdJTc50aolO8SBWW/GsQxA2sjmBQRoUlwC7SBtWC1w/fImc
lUWS4aTJJU9Pp05aWzhrpu0v9fZq/c+DHSbvzY19117MIB6T5L0EJyJqd5ICHMi6R4cu+F5CM4Sb
krR2YOfWILmX8bzhM9d2MmJvFtGB8seNaxb9g6BxW8y6F8FYqy0ArJEcTkdF/tTVgi/9IeH4LoRU
yE0quo3w3CsnzaJbdrMWbwTeq8U+E8rOKjNcu49GMTI1nztBLLdGBNo2adoEABXrEpHDNdll8t5v
7/XDpJOXtWtkWsCxsNMlbAE5fTPayCDXmMS+A0bTB4Fpx/aDp88ZerODZzwPkwA6rJxmwyMdnTIL
JrO55u8Zhqzn2xIKJ2fUJEQ27mLR6D8czDfHSd/gpL6hqn5CWVa8lTBlxp3VmkgG5hq7YIKfGS7c
O+tEQq6VWiNwUkO88FWtwzsm0QNtGMRY2iIWnompKF2w9AQu/KdQgtVnqFd4M/jj0gW9KkefQigK
nIQcrDdYCaykb1zqfK9knL1XyF8XE8F3ZN5xUNEKFP2cGd9iZ0lazslcVP8uEafLs7z0FUw9aemV
+yFKnmhkYKl/OPcqwqEzjqb5Pk/yee8Ne+K4xji2oNA6KekmNqz6jdjneE1sgySzVVBngmGgW2Ea
eyVw6nmEutOFb8ZnKD3SVcH5mLq45LMFsdJcDlSSxZMV0IjWtTFbJD8W5Ky+fF4RGf/FtlObZCJ5
AQrhFmjuaZlhTffOY1btYygTHsNHABAiptxUeba2PQg936EIk35+ueHhDSmk69TtYy+ErJVNuqQd
s8o80R4Pu9iRo/HAYdldEQKIcruGdH+cXbKlMKAvj2SvponP9v519hFQ/R5/ZDVNOdoc+jC5CYEL
4l0dbA+UzdMscWyZ+BAfditTrkOLkkCWv+v0y/DYcNFwvfcFYv8tLm8UnwhJU9awk+U9h3VEWvat
ZgzpZfZV0xE8Ad4EwNfhQdRc9EmAHBe5l825ZdcNfOpt4n2oLIbzWxhL3rmeW0EzDWKMBAAd55/Y
ONTs6AEGT8sESVW2NxtP3oF5qvc1EU3mhDIpCEQpPxTQmG8hYhC56k2umwnppUHYBM5P0QBi/VLY
iHX8h9c+lQrNDUTgGYpdLyqz4wyrCu9mCcVBBii6ESvrpWynYEdCa24tqwYDBmxQHUEjM8PCfGS5
V/kch+26EhmDyFtgdgTjyBAtYLm9XOoOz3hU+yaw3/INfeV+EvE/zq3sZGtT8scMVr7F/Ho6LFgt
w2eRoTPdL/iLw54SFXs/BPjy6cjLkABuLOIJUQvFc0mL+yK3iUbuDc5Ikp13wa/xLMrnU+3p6S/q
3cUK/rGKydngGWuLVsgCVH0WI7OWHqospCzUycBrjKQK5oZu1xZ3/dvUeHcuNuXpG81IE73Gsu5k
g9rPwU4RYePKM7yBIm+gNO2ueuwW86rhev2uj0+BT8la5mfVhYSUzeGiIsJQFUounDN43wj613ot
nKc4RawbQW9dIHl4M6bO/YuJBeURIgSOZDlJoA18jV1I+Asa74O3GLe5FeueZFoTnKmZ5CEqyARY
ISVeXPd7MpuJchVJefjtpeeozgXQVU+zL2NfRXTUyHNYtrqiqsaRPxIn23LwW0Dzawn7CD6Ft0od
dsy7SkwLuv7h1Arh2iPZmVh8G7i6TY4u2PqeNZi0tpPZsec35n9b+Xhwtu6NBVkY+fdelVXOi0Lk
4EOqlzlSca1N4vmevDTtOh1HGAsPqxh6fF3A8IVyShrarqRCT2JJkb5C4D2CC2sArW5P+JGtnpZ2
C4e4gKuKzx47+RnCcPtyZm7GhrUBs/wUEKtxGSQy9Fh7XubeuayBK/r1By+8VmrXLfIPSMbL8Vwi
lGWDfFvcWvk8RB/4/PANirfKBl4I1iDA+2c718QbLw4BFMlBlXtH/RKsXOc98mN9VzwK84yiyKJF
4x76xniv9nrvSUg3nDUl1neD0tmqCqvk5lSnNiGSTX8WN965z+7dlgQWoNn+cHO4P0irJH07Friq
Ue6bUfuKRSWPIvN4TCZz+9JbxejHNId1zilEo5MhGUpsQ9CpvHyE7XuHMenheWHc/mzk1ZwDpEB5
d7gTjZvemfeD5WFSOLq8zWyNcQ4P29bGI0msuEET7OJMfk3HgoCsEuUUbUweKM/YMByV+KMjCM3z
S9wTai4BPrqT+7WGbjNwMn0b4w4Mf7/KgMLiCKtiMAcA2MsfF/51lFfyQAHqOw6510BK0n+204/9
GjfyLehZT89ays5laLf49Dy7oXvLWJIN7Fvo2vrunQGh+eeHVG2EAtUYjZvFLaUuHvDyDNCPGt85
L/tIlVb2gEop96yVPb6+TSOkM16ywevMgQkP6CkbltbvioDXwRtqyE+/KhBb2hAiJz/wWLmM6jSj
HRKxzC1bD/4EHmchZqLWduhYBtoI8bQdy1EYLGD8zlxfWIxGlqkkuqjVr7Din8OGzBlAUTZtxZKi
X0sFIL8SKRER0bwiE5otZzhS5QnkiB7PqsGMi8mD6bNDaK1UAQiqmt6dUmkCba5SIxIVRUfW/UIJ
E7dXdeM8OTSXO+zOrNLhlaNFnrbxxvN/MtJmuiTDSAouvhCyvbQLWpI/2dU/ZQiS28J/mZinjSe5
EmsrKKM9FzQJZYlv5b8x2sH5daqwDR1vVBNeSoLgv6qpMPQ41ZWaU4LlX6GUrY++atdQ2JLXfQBz
4ySqkLT3JEYBDrgrxEfL+7wfKk5YydxM27F3p3ebIIM71J3OUR22x40CRdXi6k9YBqlohVlNIziQ
tyRBceT9aBLk3Ty2ZpgGXNX5XUWsc8bfLpZSMg+NYT9xKMRORJZIeIMYc/uaCHEnT8UvxvKi8J3d
q6Q7T99UcUAh1kgMfePLtbvKjz5/wtVWwbL87bRkRStuY3SsbxoZuiXB1OGCftE0WyOKfWuZS1JI
p6Q1/1dSWgRibnVmTcNu2N3vsgQAcbMrbuetd8JUkhy4LAUp006qCaN42NL16V1ZvuXRteLh+W6m
ZvAsQCg61QoB+7AkW1i2bQvrlMSNnEMKyLivTD2NxLdLNexFe7ILzC8GmhTv5sHagck1xkimlN+x
DLzxn1xmgS7/vGjUdfpVSSC3KfKA5Hpp6GGqpJAU4Y06uINCFBKOJTwqMC44241JPBnVUg/ojPWS
djFSYZMJJRdGl/7hxVrcyHfD0bLu49pHH/Ti026i2Y/oA/yt4jojl0R+t7fblKv0NiGUd/hc1axD
Kd3tqkad4wCCwBKTbJdPAeghJ4AD1HL9GnEGWAXGdGnSL6E3tw05VS/IAWnk81gpi0qJ7KbBl0e3
GHV8ySZsfZ4Za1wGDiM++0g6QOQY5ZA2dQEuDY2Mu2hXSOAYt8FP+D03fm0rwDMWsFzXtpib0zKt
F+fVBqlp8BymmnHzovAJB8Nq3/i9BMZrzvUfG3yG03Y4F+xH77vzPYoMtreNRJRpz21RaIF0/sUa
osDewLSAkFyf2nvzL6zRiV92pzdk3+ePMWl/3C0/KjmfnSFN7cP7CsyZFOx6Tq7ibY/glJdpXVaZ
sAfPwD4KYNvHIRWaJbgyrEVAsxF45Sh9jEaGAbZl53dbqTXmZWN5aAeyyG2YOhZuZgWwB8rXIqa1
RfXxehgdMbxh1hrlteI9oomTXAeJog3o7sRRIs0xYCrWzG6KAV+f+rc2ePFJsgJaZy2wa7Io/qz/
R0O/CnV7QQIn/LwZCfjltfRQNzVBbIgLXN0e5cozWWLXxua5bSxqFlpdL+0K+dxbBCq6+YU+T6rs
LHnCZY7LHqeWXB0v/rRzhRlDqKeT2yJjcp51hwjvoafj4ur8Tqs8aHNrJMAgLEEgOtzsVx4oVXsN
j2K+QCUIDMG2VGif1yf+AOLQaM6lwkIAP9uzDe3xfKNn5mOrTAZCsMyHrx9LyJ04qY8j581PeU1z
S77S5FNKqR7Tfo2jK7ml6iQk3b4rkeEeL6bWwjugszH0D82Ah6Vk7ouPOURRE4TYmNoSFPvr3HuS
ZJXUxhY25NYDWVlIrjuwK0Y/R6orRL6duLfzDtKrcEo0jzvTBAkPPvJZ3WJWv/PAbQH7Bh619ZAv
i8Y/qXz+85tSwcVLZkV2phsJLKwbBJWQWjkYbZqNSIojTeQksDMT1a5/R5V00AKd6lqXQGxy//WT
D4WzxoZl4azf2iCwkrfZoHqmHQphiczRddpkVdjpJSEIpt0R4WN2yqB+AeeSKSxGYucosyvZeH6P
mKOGAjyXpz7NMl22BFccPwpMi9y5E0Y7DG+4KqizNnAPZpZ4zx+MJQJ1O56Jq+3O+cfynkbkwzLx
oISNn8ujfvMdAE1483rS9SchGL/9AR4ncfpKRZ5j7TN1cgSlUyRFftzIR0J/VjC4MjKGYTqp85EO
8WJyRAL1+krP1Mz5nKzSBZAkDA30GewYe44Rsfa+ERZ+RM1UaRpVI5E/rsaMgXmJSwHRM/riQUAF
xgRoyO1VCOE3O72Pdj8VIf/CGhqwQni7S9hXOKcggXdj6A6S2llcz6JLnV7308i9cJLzvF+2YVLt
mmRIcrquvdo/Z4C2KsEi0uFgj/Z2E/1HIAclQrZbbeLJEQ5g92WQLPkkCIfdBBQkbxTVYRTIxGS7
XMVXTlwQSn8vdddkdwugJ9WHg9zZImlCn7eXgBFrpubSH5HH5L9gHiiHR3l4eEKyA9/dL8ShbMzg
skpa+F1Z4grr5rYH1T/Ja8QfwJZkQVmg9wMiElFOxbTaMW40wXt5788iOaSIkV57L9vnN45ZHtfz
YEiD54bXLEdH/KTd5glwr3jT6ciHpnTWIHjvey5j8qvnbeeEYUU4ZV1mUA0Mx+UFjVJ8XVbNZCk8
/GLXIv/+GBKbYKBeaBZWrquvbTqeA6K7sqScAJPCBApDwRaBarQD/Z7BfBXzqT0jjv9lZ1oyYJAg
BB4AGwjR/+5M9zFhJGF2UjZtKaw7yv0EjsTjclaVilBHdZAiLGAPXUZl6ZSm5+I/iRmTfxDQjsgH
JRW7/bdz99INcsrJ2akAWBJDMgkdUauUF6DRIZWxtrNrrEytXN9SImoAzjaWpl5OShh5D2NS5jIr
W1MxJ+WUVLjnruSBLk2GkoW4h2h5e1NBTjWeDbSZFOL4w813+jyZQSD2cF+A7umajOeeYHj9Euzd
JpMQTN/zjjK8q4SLYdaQ9+2M9aSbEsIZfPMYsggDM70Px4hYtUUvVBK/lq07pFToDEhgBHqVn792
q1lqC+XvTMOHvV1wbDEYJbRqkyVOHFZS9iynt4m8m+Ah72xP6ocBg7wzYuiCOzm7miPEzQcXcaVD
SaIu7auw1ZAmaaQK/A4cQEafYyYheOGrFQXdv6krqwgrYfSxvp5B3yMgBjaSlbwhpMv27dCvuugO
ON0ZDTChHTaYfMlQKtSeczkwqxynQQs5jlG5pV9XaxLa8K2I/AxmE7YxqGuFfRXPhHPptKv9YlXd
TlF7OaotxuCniuwRGc4Yd9iUOdZJJHAoi5YtJRCg0g3lHpvYWEJwj5qdKMZBQLbpOb3SRc/AN7hK
pFnByOnj1kTC6Gcc8Mfp/AYW7mMUm3pWFuc+tDGhyYwMUjzR4SqgLXYfS33j9rQc61jtWIVCFEo5
zYIMu0CD5deDlQHc4qIinm7+CqNljpNTNRLRRFw0sCOt6k4xyyDQpJOpbBKUINOHfgbntJw2uAgG
3vJKPgewM+i/LO0QYfqr85ZiXD0u/z3Sq5IelSGAwxQi4WOmVvKqCUebj6GxP0MxoGTAn5quK2Pk
qVnn4bGfrARRioEdmSjCfKdlgUmo5NC7cZcPxslPMi2upwyrpATDOXO7NRglD1Fzu/3umCUqBXFm
OxtxrZ3Qt09XcHx0rRQ12QMAdAM0Lw/moohwng7DM+NEhWD15CDeDjZJAWx7F5Mkqg+Plre6VcRA
ijloPb+HqP//11f3xOGTrBZZRqsTxH7BhGqfvbd2lQYhu11OIhXf/c9iPHOc69/wRWOD517o3YuC
VM079WrYGrIdpSHeE7TIk60opE5Vrbn82PEVBCQ5PpgcpYYD5MJK9+P/j1VZNC89PVODkyPbiqra
/WFGJx+DJAqlpGRO2ixyYjV+VlS8LdYprQRLyCNdcowpYQc3g44WKSp1Z7tO73GfMpQzD7KsQQIz
s7oXYYlfakGnoQ4AY+5vxJjHl6gWkWTdNOkSiH51kuQFG615kpzLTuLa4I98tpoHpTPIgAmQdqD2
/TMat0qqT+UwLYw9E1URabvGk6yCyJHGcl3/AiV5xDJvxDd3J0oQEombvq9evXfzrfONuukrtJX8
yqnmW/fWyD0+Lka7KZyO1jY0olnwppY4FjRSfYKjDLiN4xF4psso+T+4XDpsJyJ+hVq5/MDmcpaH
PPqTpVLyBhSgsQ7mQ54Nb8giOfckBeoPraOGeuOJgDVTtFX0SHcdRRtZdWPSCSoGLZ9ayDDUKXRm
TcsVe6YL7bEpuFc8+9L9yd9ehLKTBmplgw5/hSsNcmhjaFKcOZyyuncD/JgeLCqX9rSHTLPA873R
nnZowXIUvkNeT3rgeWZrKyLRTEhQl+Hki5nI7TDUyxR3dixqoKAMt9eyZxnlxUqt+zYZaE1wOaEY
/nf60zC7zyO2/c63kDXifSwzBcbhGXy5vwb5VRjWhKfFK4o7rx624dCtfs/5uBLVwXzpcZAY2SII
hwMEeApNktbWUB/ckUkLYp+4FWg34L9OQGq3p2Hq2ugbEzKkMTVjDRB2JpcmP4zm2jqTmxZKn0GP
ll0cbRfbizcL0X5Ddk1wUjBufM4NT7xwHFWR/+pxVwDJk0nU4UaNAMi/JyDd7sq7utDX2lnV0bIK
Z8wtjY3UdzdR2+Jl5wg0igauX5taQGMelC95fNsss9pqulrcS02oCOuCJLzYBw7I8aZpYARkyche
QHl/FoTz6sm5jgyt2Brd/n9aYW47vuQr586lk15FoTFAWE/6AiSubr7ikUjwOEf8FjV5wK7fbNJF
zgN2LkeKNEJta6xxQOPNeVePaMI/EVfkskTuKcgA7OWRuWHWECbsECOjsi8kyClcm7mhWybbvOj0
kmlhIrHyvnzXuMcCbQUSydJ3UlpPodXQwa4gTsk0bsh9Q1JNZ7n/yR5BVX44MoJ4V+eNrb4Pt3DD
aJBJo3T43vDGraZdKInGv7fvNSlIFKYy1iM7gxp0tU9IbjaVMh8ehbmnzSLn57kVQunJ3b3HtbKc
9D+yHCZ/4QHeW2kLLHtUBz9ILRS5lcZ7HtCsPhxaPMRb17s9gFO+kP+AknYZlMS6tBAXRzJjiS/1
k6tFgKhbNQOqSL15rbVxSeyPAM2u5ztPgzR7ftMwqJrwaVVab00QSYVo6hzit7Q+6lSLscfysYI7
5E1aubWFlMavN3Iasegm6l8GSZVH2CthfhTDCEcMAl8INWndnjqZy5Y2705iTc8futExIfwKH023
9Fwskbrq5xIwVljk7U7d4dp38baVyelviiLsxLFoiY80Ld8/aC4dPo2xpO3kSq3bkwfCpP+FnIdL
FIb64jS/LuHW1oA1Lz6l8ggnH0FKxmmhpNSfhBNrWntzKvckZSagwcBrL4t75l5XWP4jlp+7U66+
KqMK6d9dEZy9h+rjTvPJZSXI8aBh1c1Qnq11E7cqeZHOb5j+a+i9PvFshmmNRaJbQSdvvGWPiLl6
MeS92r0wUemaQ8CSCMGQan3qrDDtU317swq5nHXpMZT+LGkLSgPVlAC7BU1HTvxnyVK2Cg1dNzIx
esCPfbRnginKbxETYwU+dc2tL8XQA3+xmM+9tXMXjLBH8BlU6P57f2+GmvPJxJitav4D8EC5F7mN
duijFEotv7oIXHUX36iChL0Kh0CuwdHYN1H3C7hksKnzhH14hjvG40lwmNnESFMDeRSw+Y8+McrX
9awJude3mtFPJKtd//8KZNKQMC4eX7w0gNaFpRswkfo3tR9AM7skz8Z1l0STMry/cX5aDuqk5oz0
RdRs+PuJO7eCixJKsUA7QZHC9SNl/rjZzOqBvNC2JcFd/zoJaXpITQfjMYMfzJZQgX1PTRQL0IWm
cUZV63QKvk3D42wSjk3e2w3zlk4IIHBypSddRacm3f9y5Q1Y4uTl8faPqnVCmQi9RB+06aTyjpD9
Hkt1Zv2VgWtiAA6wLhEiVt072LqV3h4igocim8K5l+jbuMYWde5i6t6JfPl15wUvkwpB0Yqlk2VR
oobDZneDvMOvjPl/bWv/FxtwO/YwMdhEC/77jjnoEE3Kj5WMFoCINthX4bTjdaySZaDReYZzggao
Wf8dIwKdjyCddjYEspHUUJHjUWWHKEhQqcw8YS07TLowkrr3YKzlc/FE21DO9MHdKHdBK53nvE/5
y50UqIbSo10wA89+5FcCyCCMxlTlPVcl6a9A4X9seSee3KgWLBhSS3sw6R0BYKpkEeuTYEJ1i5H+
AWuww7m1V+9QlEeCMXYi8Vq6+Zcnso3JfNoRCpvzl7zIqOoTChhB0llLG21VM8ro+QK32erfnFks
9NXq7snIuVfPajaYgUtP1QmEx/BYbkXIrDYfray6ysdFXvY26/0rCoSJOBbhaS2bmFhZCeWt4WOi
J4Wrs4WAS+Aff39yGzvHxe9uvi4j/D3GB+3O57dFbXMfgepIhzZDiwm8TxBGqeDIj4QPHbj2hyCZ
htka53yqqjxim+hr9Tl1q3+NYpVAvJflt6r2tjPP/eHf7Z3LjGeCahZZNhAz6m85Zrbl8arsBxXd
inQQIgIwbu1buWjRds+rDO6S9Vc1hsDx8zLlRivxNX+ZkWDWsYwcHtoOfSggv1andchOaHFNPVzq
CVk2t8IEP+NnGIKXJAEmd8ch2bW2SawgguRCTo5pyc64wSXGPJwr4yzazUEK471L+0JiKNdu/0ud
1waIF5Es0LLNLVrEHEQDQLUMN6H4LdFd9DxULaHAb8N4OimNDdMnOgHR9GgjlKHQLtR3IjZqw2S6
sFyZCTo0BZmIycl2jRQP40oe/8zhVOJVwDC40l5LmM+C0hRHrTKejTzS0WMrq09alPBKRblzvAXs
ajZCRoAdWX/Ghs1URX5WhU2r0pDhZ7KpZ8wMCduhfdG5cJ+2X3ap9ukGNmgLL1bKQl2hagoZGQDT
YD3md3AklCpDtUjP33LFKSy/ztZzCraFDJEEhEc+B89747EY0gji0+xvFy8bDU0F3OLF77dA6tW3
nZ85YPcCRhA5XxTwkv8PXWH+UR/ax7adOrMyzSmwR00iplg/oVPN9/N5WENASUIFGz7AvKmcH9iX
XYdNODX9w30tO6x/E3wnkJr3FtYg82pIqe+ehrjsNPNyi/VTaUMXtZWINWPzByPG8z2oJ1dVEvCp
8IVUMXdvxlxhcIux/2mROymgDdwmBR+UZ9VZ8iXR5OtTsUOvgKuAmR+C57N9bJhMBOi5btxdGY2Z
B8E1GoFCoLUrOsj+iMLjLIzS8kEZnXI1xSvXTFYbVFGrO5/esj3EZ0NK3PuceSCHRxEfqF2p12YQ
KJM0G7lEIo5636ud/7yTElzzDVVjSkqZyDTnR5v31ZF0XhlRg4Z/j3j/7Vrn4S2egdmk90jekVZT
qmU6m1BEc80WOwhmT0b+QTZwip/4dZ7PVcNL+f0N6xiBks1fTmZZ/H3PWJEQGC43b0zBXRzJM2VG
/l3owKla5lQxricTCj2AhvJeoEYu5PhxsyCRmD93xkH5xt0mXwxJoYSTTjUl6kHTsHqq0Jkt80xk
h/22ThqY8POhq9GGE9IJK9We644iYoyM+Q5UK/0wMaR1WV7U41Lssp32d+p3ydN94LKzxezuyVOG
DAoC5jyCKQxDhCFM9S+jQL0beu7vOvrF8c9zziy89glkIcanqjOdnBUZHhVK7KK4sQPMD/WCU0D0
U+o+dHQIIAZNxwlPYVXoYsv7gJNo2nQPOgj63ilMvUtIh8SxJ1SOLfj/L1NGzIMDE8oDA121dddr
pC5u0yY0eTeZLUA9J7eCe8otNeNTwrMSjNXne2fzYOJetGVOpJkeRjRV5Uno7+brEwvTfjohXHoC
G2YzAxyrwa+xW3ocMSUmVrUFW75/DJEYRiNYf7f1O1QkTrOLRKmcjbpbYvezBBMPuOqK1I2FjIHx
lFQBC/2Hij/CgmG53lk2cqT2f5EXX+kH9saWJe5cu9QhAuR6Lvg7+OojXeFHGHYFHCDjEnexinMS
V12PoqmtcKJMHEidXvOJUtCNBXJyOaeCwV0R5zq7TEX7SxK7vqATS69w5ULwr0+2dpq2tnvjXzWz
EhhmqINsrd6ezOactURh5uUTpbnV6a65SO08wR9F/N1eWhkn096jXMrplxZwUQ00LXOM0guVuzMu
/3WE8ibf2HKCHxAmTeDDMxknty3o219oKloBNpQQnkeGpR1uzFWVJ1Twg8taf+bQC/IEdlktY986
A9kNnsZMczM3jL5jKYmb62EvAb51BMF75cuoE6mzx0jFeTJ7sEnNfDU6o42FeOdIj1CZP8X2sAZ+
DoxL/1j4eNgs5dKBD6QEoQfjHgtyesllVzMHZy97Cd9dgZBQ1dCHfdu0yr1QI34kq9EItyf7l7Z8
Uhy/u4zmOGk+FWDKsGd2r8wi6mly/GUxl1VZpVZAAAfIo0UBNt0Jhx6l3WgfLCZeaXbsoQjs298X
6iRGRBUPJrWbPHsOByaSuic5Zst/OdCh5/+x6w6GhxREvhsQc+L9ybt+VBwb8fDjKqLh4HhG/K3p
rXfdraLqza/5oUiKyIjZYrUY55jQCBUQOuZJ5m8HxBC7kQzSL4tH5yi78vTn2Zjhmaj8Xx6Pi3gA
dToqGZORZ/wAmWqSm7wvFhiEuD8/irIfMVnfyWI5ndU0b2spTsnt63JCn4a2/bcd9+XpvU+yYCs0
PbuyqUhudikuOX6Y6BsTcO52A9FzDoaCj/GwCOhdC5JUArDMFMSUnCMuoyl2/QxZepbYwnKsqoLR
GTsRxQqqIMjfBiipOOTZTIO8cNm/4WZ8WccMhQnfi1dPBzxiiL+AKkEgoab6iwF549gA0yTgZXbV
GCkjViPKvDKVJ7BRv/z/WNugGGUJq5il8qz/bL/ZGJ63nBDSV8GLn8VUvsuE2+Vuyk21oBla0mee
Dz9l4fsxE3FX9sbwkoZ5RNIPWUkh6WbedN43ZLgMr10zItQU5LacS2ZQy4IfWjloLKIOjCMo6+mE
zDho8xT6LbwvyYZ4LCNzdY9K+nWGovjS1Es/6MrUkv2XE9qhNWZ+5eDv4CKvYYAeg0px11KhJf5b
KAtqIha4KOpgBW2uZRuqAIhKdABwseUxzzX4KOXI6YX1se9t+W4Zhb9U/8EGwCJwoqHzIGmQy1Nn
5u5ypgAYoquqUTZ3VhpN4ZZcJ3uu4QQGWQ8xxH3ceqjA2S3g4iVze2HVWWEY5M9J1vAYxgsCD08h
42ClbCk7MZgkrbb2ZrLBj/LZFULN0U7ttQ6WBQNW/+2Pg7mES8uTytOnjGbTIyt/YhLajlblZmvo
30yN8Q98zD86eZ+1CkKB93joc5z3YYhl3fu8rRSBm5hPO0ecZbSUGxW/FREHJUBUINMiyfAVYfmg
TvY3HVXcuI3OKeTNJIIMB0w0vVvLLKVnfoWZXs7wyvcOhFCSk/acq08j6qs+CKlrrRBSd+WOyMHa
U9FoWsguG56I1jTO/jpx8xgfjW/IU34XizVIGCJZlz8JpyXCRj1S4gfoWyXN8hBJQZZhi7QoNL7b
7ZlgePVHaOQW2ozxZDZ+2EIjA7wxRUih0+YY3eVJPg+rTNnqZXzNj29pjZcb3MPEUkg9tDun3uQL
YUuHdNnEiACETSlUQymZl/q3xhB+o/bJgP3dgaMWpfNw3foUQ+pnFbg0Mguusjmczr+zDmkRKpFs
48fpBLdcsLaIDnSTNqbdtr//a/RlslXO0i0J0/R/vTzYoYDVSPqFmpUDBpU2Bq/dLzXQkB2oNll8
GFDOkFt65ExdNEHviGpihX1vd1RrTWZ8j2tDgsZJO2NJbQqfSFoynx/w2HHI+xln9qxwZZW6loTh
YIzJ2noH9N+83ubTqMleoh39n6LmA89aPKEDxKdDvjTg4oaJUXTJiiXSQ3eSltJyOxTsHqCuCJrp
ywv5OrQds8fHB3cof8IMS+WLXdPNfBU0Oa6xKxuPzoBGlsTtVGaAYrZtkpSLfgSdNXxrul9HZ0LO
I34Rhbw7oNrC9nqSQJybi0IXmOmTnJjFRrKOBcsg2+zp3r02JU8Kdh2V8M0VHFIghfzcQYLI21cs
AyIvtIaDcg5s1keJOHDs6moovIp/oXGj5YfIjpDZtZ/Jm1NxQMZZ4FjEzs/z4J7ywEQYHe8voPwR
Gjc+CYMAzcwlY1SIHNVMu4EB+HkwAEzArNrUXLtaRLL/LKoy8zkIbDCyqMRYK6oVfGecPK6f10oF
sy5kvKWZJnt3CVitwKlCUEy2hZnvy/obJF8AmWGzi+mQhL7DZBFbOgBp5txFKsCFTrzWJMADVPMC
hlC6MM4X6bg6esdlrg0ax+SVM4s4j9XR9+KzK4riW7VKRbTSxCMrwOMpHFS23wy9wFWsmOxF/dFB
RpCSLusvdA5TdLm/D61yOCQAXD63HrTsYemPC9d9ybXjbV7/ojLfvqxUSGsotWwaKQ5tyvzhVBq7
eAIhe2QvBDWJMVcpIoj+sRpZzG9dJBSd0ZfLIlpi1UZaSqj3LO9siZBlfgIxG7RnUEeuy4HdzEWN
QlhWyaawsWnmq81zglrYxHHkUbMS1kULm/FSX84xW6tF+ORssqBLNhAvcGOk050CwydolRKCt4Ow
caxtdHptDlrIxXJlc+OmJpCupiugxnBOf7WcMQR4r54nBzJHK6JzDIh2pdWUFzsJsdMuD113eJkC
YNVzS/zuYHIzDpXW6V1ITq9bWqs57O7HNnLPqNGvkOCT4U1wfI3MS8RdynKBMpHAPLl1RWQUiF5K
OOiUsmOHwJ8V4fA9BBS2BK9TK16c8rgloIfMEjrJMaYc0W+xDF1r67svs78fm9SWtL7agCDiGdN1
pBeysiyt4cSOv20cYfqcsluqxViQgou78gWjzCTj+myRn/UK9lJr1GFzvyc7K1QWnCXPgdjWL6xE
dOw4h3jPK4xuPdLV4zvJTwZdQX8DUOo/SXbA/gyMRMrbD9EFzRaHodSs+Jphemfx36Di+uRBr5KH
2jgbpt0JtlMOZBnZqJ6M/29v+kCik+KRQ5jI2foTe7uvYQeRsxgv75/LD5k+7AwccJzfX/yh0olY
QxM3n+8i8t4ugQYFtSMR9W3UYDUeYzU6oYr1AHCP8B1EuGPcRs9y2w3Pruzn4o0hUXK870JcJ7pZ
BhDLv5qTZswMxWlCRrD/6dBJePvyW6rwR4w9vDrglDWuiq7PVyFd3UcagALNRCdNQATv+BgyX/ga
1iFsYIEes33llAa7dPn04OkqSYSG5p92zg029Wpn2O9FzmVY7OWLCRtPswH7MdF9TSqOUKNVvn5Y
i8Z0db0Z0JAGMxjCA8/7+LT/ozyfcSHvpUPIoG6ZpK2yRdVRT1/lV6dGyXQHlitO744AVBUV2Z09
NpkosUHtv1N9KwRS1s6Gm3NgF8oynGaeO1he/zfR3f8SagpcmyMTZ//xDJ5brATNsKGElwwYSa1R
UrFcFtg1h1f6PK2o/wAYUT0aHJQ8I7lPfhfxILLmApTxom4M+Ia0d7h76R3NN4ZWKc2YbOXbgwFG
slY6Z20vitlJLuKjoMO46+gYzWz61DCn/71rAo4x3dC7bCgU/NqQaRFjwup7WyBa9S83Gjqc4UmZ
AR3cFWGDOP9ZzwrPu1+WhZ5QtUNwkO4fYbqxIVcpxaDLVmz2NGIj91Mi9xAoYl7XGYl3vuSu8mwy
s8lY81tY19QnLOZ1iKmPaXs6ObzcxhLJibLhnlwj/OswFN7sKNNQoEcnbYDZRz6zNixOTVe9Vm4N
wfIBpNxSorKHg9gF2ms0ZxHxXUmbaAReG7DLfgQQNJBanO0UHY3wZAn8daXx03XM7Judedyv2OBJ
/I5sJJKkkpHv6raxFry4EwyVoIIrJwDjK+hV8ROrG1jnz6XwutEdabXdvS7Fd/OwL2GrndH1KbG+
RQDzMwRbA4MBPdUs2Uy07kQRfv/MSxCfYvFnRP2yzkmFcJtbhJuH0qj8c84ppUpR/wQHItXOVmuz
RVqkyaVpOU9lL83qLfIXlY47OUNPmSl0DX4l+VvBe5F1+l6Cj7eJZLyrrPT5duY5zkGu8Pi5JJix
YETja+ff6LeF0Q9nfzJu97cL7tMtc/x4wd7p3leuh9Scvp8XsorkRjUe0vKhVUFY/CZkXpmmDhZY
XGM1ulgkfOF58j/6KlGFH7wHEdlCf7CRehgsCe6hZt2v48aspuld5n+iakT3pDGZtmiwkYGVD9Mb
LuXbcPUgPYBd6SEGPtFr98jcG1gPE7gJjqCaEYSobzV5Go/VoFw5WEPkOpyCQKPOI3oPPRV1VdyS
QKD9xUq3jnQA8LC0VdI7Cd42OGJ8Axzk+jWuR0fNw/oWDFBukgQArkpLsWyyRpVll3gTe1jnV1fh
C+H7TC2HluzAyafyEbJCfPclr5utD/E2xiJDsYuRiY3gsdNcMEG9PiFmHt/z4AR/lzhncx0W2i/i
Zi9u5I4Cjo/WDFVLyuixg5ZcSyTtkLXePYXs+OhAmoFMHOOQBkfzaz4R6HjKuBYElT38OECF8iPe
8P8YS/9lHZhO1ppgmVpqwoh833UeRbZwGj2TNHUXl+GhhQAoi6FjR6z6WkVMAwlTGtL6m25MbLnD
cFvDDtYfsH4xBMdyAZ8JnCa1Tb0bCZwyd3DHdJI7SaB2tiOVirz2UQgpSMJhlMBBGJKq+jqgTe5R
96Bg6aJ3+/7CAxEK5+AOpuXaK67U9gjWxNWBXgd21RelPwpeaDcSdMu05jb5Q2KCKuptRWSxIjBx
Fudlb5WSuE0WcibhdFRwIrWuncLV8V15TvMGXu7KLp9Z/dOYDIkJGtBg30Wajl4HKeb2exuqNYZy
q/tForLUpRwcUv3VkGt2Hy5LYK7yp8Ch4xGtKMG9U/nJkRdGeGwXkSn2pdu/fPXuaB3X8AdZbl5V
ABUtJ05HVosKBnIoPGK90H6yJk2hG+k3ojYtoKEBYxRqPAaZZyY4qmNcQga39UA+LVFlnsQ6sUlm
fOfFbvI/LdjUwAPmaNHWpTmmqEfzFtUSVMPpDLA3KW01P+iutYmcglxbOwPR/LWQZ/ilpFbvLdL5
zJujWeHIKJVJoQsPKYBPny0vEEXHIXZBkWvtQZ4oNug/P6WlVMQ+SS5buw4vqkHRk2mVC5exxIr1
WE7RaPm7lk1dNY9lSs3ydm/81AWh8at1DiyRit6EJ7O6i94KzPz5te0OxAuR4na1wOltO7KGb71m
33JFy4GWs6MUh5pHpRWFooCOxeWU8vG+BVsgFKJF7/f1eKL3aq3cTihl5Jiel51E5tLJMnXAl/Sg
0bbdM1VjFzH/CB5zg6jZT9Wu8ChXU0TPtgye3h9864jv8BUEEUgiQIym0M5vZeCJ9FWLUBr7Vx1Y
p4aoY62PbhF1zWwmBV6e6RE/7a0PbHwaNuHmelEix5Fmblne4U5XaBrnuIGpqCRSr3uswCcH7THv
dVZuAgGzzh+GK2WBCdZ3r7D4g0nI9mxDF6cMb0etd/oBwwS3p+DivL04rbCuKQBzCccpJcUKUObO
CfXNiEppHo3TPrS5dncwGgQyeRdsOVJYDYGHToS74jWiUnxlPs2zmp0+0OGIJF9KaUlwKuZnSPrS
cqb52ihwIq0Kfnj2cFOAPPxM/YFrsk0ztSxNClUUT3nXmqwp8GAC4yjCDFvVJYQTn+nd4/sBjo+A
pEIyAUM3DPBRepXqFRN/MUCld9nqopWBxXaefwGYlJl6UctKUBPMLRfrDdiHEOm1zeoFf2wgjAuv
QMU3/c/lnYqFbsq8PzsJ133J4sUYCUdxXfczqIMs87fACeQggAiIP7HzixBFRlU6JGFWv8xGp0AS
RDa0N0GtegZPE+PMhUAiRMmAur89B1Lwf5A/vbIRfB37WRSI6QHGZrnlvAU3b4K9ebYyei+535Uo
ZM5X8wUMiG2Ee+Vu+OXlZd2S7jJjM0MyYOFvcDXNb2XwFporkmqZwB9cUgwV13nfgPj2i6pF/OvR
PRcnLk4gRWlQ0LuOw6S6z9/if/EasxsP9OwHLeI+Ty2ptY26ZQ1wkY3zfjtRqW2BUxj8YBPJHZgl
gdj18ICLByvCTNSos6wWBCim3TBcFooBbKNm/8sPZ3+DpcY8dwhpoZicLNWlUIGnpIR6RfXLmLUM
dyRHqIvMi72+PmPFUdj9S0fN5nKwbNfValDq1WYOXHlzeqJnC3JSPqwBzfIBEYBt+27yslbk3WcF
lCRiNeidIOfz6hO8GUp04K/mRwXLZ4kGWVBVj+12AiV4iHX+kxE6smpUyjAhGiKMmfY2fWfvYoNd
Ez+arLQopSto3XpHuUlClZvrNTFsUIB+mvv0MSr9uX1HJX3Apryd+wqDWPL2EhhyF34aRqErTyQk
TOszLmlEAVGY6LGGkKrPiO6KBDsNlQ/OcDQrXyK+mhFVqpqn66IEQqypSBThe+mkZwBWkmPoSpvf
l0t8GEov35dBZDR4t6MniRBGlquiAIdvwPNbUWxJTxpKxcTXzZDA/rhtYmqeSzEe2SRq8rdgZ628
JhmPHK0nBGIwlkfb31HmA/s9mXyxNPIjFz9qdhjv6MKEpRhkIEhRKencHgE+7fKv83eRIYi/Qbvp
rZAcEXuFR3TdqwjG3atyhjIzzmPQkJLfHGyEvCZZorHJU4tL4vOYWWFtbVtSdHAKKSY0PluWqBpu
nI0LPqx+T/tle/uqr425FTqjaZhlMTvvSvgnS9jiicDVgX4QERkxaNWwJRAXo5rJLOtQejk28Qk3
vwf81THvDgwcd1dxD4Le6fESB951xJtRa70k2p/Lxr0R6YkmoLtHTLBUVdUDyUjgZtFGmORCD+Sy
sKbQa+0kW7bE0cgHEcd6Kn5u9XZ6N7p9AlvTxlRXU3DrPVVPk8e7Ppnm9FvoG8wNv6d8VkRQoBZh
TPS4vbFlnW9vNgAET6apBISFycqBNY0B134B9FoQcb8IFIIUXKupav4EEzGEujWXJvI4Z9rJdXQb
VhULeGq6K/zMcypuUL6ypOI5HwrLhENfduoHUiRHb+VbqfAVQfToi/tM6Vk06NSE0TmxGFJJE7he
NtWI0+bRnwYdRjRNqOP2jtMdS65xvtylIZ4kLpwMO0TCnnOpKWwNqAjWt6J6i/A0YkBotduJJL4p
S6Tpa9Le+4yCwjM5W5mWOHuzs2L6ElHIek6NFBsp7DbnEc/Q99hZhjgNTVeiBp6QBlDpfkiEiWd5
DppTOQ4vYApJnLGc/fIxunEm76AmgswNxF/Us+FnBIVpXY2k/8684+B/A4NaoxnAzIWtXbALQesV
z1/ZJXdYSnMIWJRJLPUTyAJ0ILZa+ElUjOy+S4nZTB12OnrS7d8F/zaoioTyGHoJxzeq0zZ2V9lN
rERbQUsYnL4pJxRX1WQ/qQ9ThYVCkXOSSPOdc099XZp42lE6DRraAgkMb3ZaCCWBJDNWHOe7ABso
5F0Nvz/6HxdwsEZ8Ncrm8+SBzx6DySJiNMI52SB4CnocjpaQHGFWaTWrz/76VcX5pl2o+F6FhvRC
FoYtIE7lNjWwOpLJgFURN8+f1z6ZdbCEaOVFo6pZh/jt3Vr409RJVIFAwh7SNcf+DnmpEGx+RwL/
1oeMRasYXSrnuV4+uW+bzs5wXMlorozUSThyxr/QU2W0o1Ej/YC7dQYpGjoWgIVutJTK3d1Hb+/S
I8dq2nYAVhTpUTwuMrNlgi1k0MMNv9NiELn4txG/eoJJsSLe5tlINKCgKLX+Zm+Hjd9dscYeGdFh
XLAVpyd3havRErdpY6eJPgt7b58gJ1BC4ZP5Wg4lrF7JtGpvMtnCfO5d5n84uG3b5JCWc0KZfdQL
PDyt5dPi5I5pIYO4oqSr8Mw+QkzXUd0yZQFo6IaygXmsm249//m/CeQN7OPfuM5SlyQIfUA3Y141
9Nv3sxToLQL50poPyHSqowIVZD9d86oLA2tyqUzF6thsK4sJrtXb0xachQ1DQk3qPbGI6XMvgsNQ
9IF5HCRV7dKqYmlP5iaWcdtMQdXurKTLAc/5vErV/OahJl3Sbu2BAH/GbXxzt9cljr1Gv3Dt0SDc
RsVr2mda3UumRjoWe5ykUNXZ9PMMo0Q3vkk2HKUtBoBhBAgcpWGP5F7Os2yJgqlkLYlzTNg2IhpI
CUNyFHU5jRZMe/oy6uAv/nDo3ocmqkRz9+L/Y9WKasYCvlAT0+2wFm45Sg2m1qrV5XV3+vAjuL+4
nAfYtN9kIolMTKeLazWRjBAxINVpBhXLTWFqbwHsorRmvB6J++NYb6GQnCXRW50L4s3cg0KPeVNo
VVspEEUg4HMr3tiD66isnjYOAYrdM154h9Sxc0jrI9y+OHFSbk9hN+HjWzAeL4hcSunkbeRRytdP
JjjbnPz+T/SqrWHiE6s1gHD9w2Tn89ogF+7NzalRDqC55Q/Lu6Sj86Ut3BFUchaLypcc9j6IIfIg
ppuEYkHrpSgJbfYOLyL24mQ0LAQrnuLcTmhBqwQO9AljNebpQ4xXw+pVo5Qga4SO2dZNMQN3OTGM
ZpofhCKpnVVMvezGO+7RLKWdhvtScA/cW+U8lgvCZamSSiCjfiix8l1HbbIoHqdn+Kfh2eKa6Xgz
9ucfqB510S8DEKHYGkMdyq01eL6z71O9D+A/9kQcPsG5d4Zjj2UqjVrJ/IddlyyYKP50RCvPyw8N
+2MDdPyZ3vCXZ6esuQvOfIsn40luj8Yoc1CiZAQUWf1dgjaVMrZbjY3c2D9GgA02hZqk3ib5ZUq+
BAoDzYbzkmxNW5sY0jhgN5M2iGICg+efXD3LNe2gQsgy3WlfZz99MH78NO9W4BNqs0Ti6bKMZ2aa
d+BvhnnIcQ51kD0QzRjjLSeXZwgqG9K1msYY723Fu796F8KCcnoMjjyqDszk+oTcER+QCA2jdOU9
7CY3KeGdIjj5BE4vaHDp+vrlzgv5BL8nk40I0/T+ecKWaNI6dd4aPkYPB3GtISRZYPakYNqMwz47
7VMZe416n4a4nB1xwjYbecVpw1nAbji6WL0kKR1f6CjFw+IPgH6qfikwgy207jKF4CIq52aCwFN0
MkkGS4HWaGVLPy7WPNd0hPrlR7us5x5sIbX8U2FjjJGwF9P8HeA0dSkFVf0hgnivC2nTuqbUdsmM
ik+lZjKSU0urS7h6bUrg9rT6rKqFZPvfYjQhqmhdqc8Khb3+uiZxmp3EUXDx1fCFg81OySwCqy68
WQUDviFR5nezvKCMmp85XJRsqnwkgz4HSraD1sJ3ixZ5dXUB2MQ2TYIl/sxWJzSrF2spvBUDYZPP
489nyZLGg3jfMSn7U9E5Vuiq+w0+paNtiHyCG9bVI1NrryJncNcuMOjSpzJ9Kv2mBlFhID1SJPvl
X1JOvJ8wjSKB1gfTqY+YPfysq6LiXVcQo7+4NbSiWB1JQ5bgqq3AhRoFqugKTjG/RhczrqVffDnh
W/zQ/zIEo2lpJE+ppyOpl7UagrFoJqQTD906fGF3ewSYp8BN1IC0wAeDXMAWUW00q05J2Z1e4PRd
5J5g4QVeoNbdmGgprmO+HQwm/6uPYWOD0obbtnP9JJdLgEB7yV55fSLr8i38lnCXyPNENvD6/S6x
S8toJ8XB75To6Wp0EwjEN2VNxzjeQ1wCtBUz0n2RfpcdJwOiSvZsuSBMM+qMHCzwtHvjoHmCV7nd
DmL9wk6SCx16bCPm2/1MASqJcqOC/1PoIlCEf/qtewZVGsQU/6BzqOGP0K3RaOPZCG8ZRyPGlAi1
XB74iTznXn4ih+OoozjscR5pqMaByN7ZHEkTRwcn7le/gdOUAfk5Y2gfstSG80ytEE+UwHTn4NRp
KVs1QG1pIjKx2EIp2aQMfqa9tT5NIwQm1gPkSoR/GXKljZGxmVMMG+i6MRwEs6m9wcosPD0O5pD/
HsHfyrjwZoULzl3oqB3L/BQxrRhhkik7Ut15oa+Zr1ci1TAXRhWoazgR8i1W0PSLtsyGLs4JstRi
yVC/c5JkJkuUYOeEMsAYVaiqk6h67SsHGSpiAQKJ+BcmShRIinp+1y8yrXpL/dbAk2+5SztU5s4S
B/zS7/rYzFHoqXYqUbmgjvOj9XGxH7FpOLRWw2rWqhjRAp/x17f31H7v2vSP6kX3U41HxIW4gGH1
0XSRw/85VmJjItEkAdaf47gCsgyiUse5gv+H0WeZdqoBBfpVVCxQUaxDELzWe/w7uOCmnNOKV3kt
gBzsQs8VovvsYQjLMyxDsODhp6mwvG706ZCXEd+jcXhz7CKnoCsuKqZ3rsDumqPNxWH5UR/GyYVB
CPr2qZIklY9AEd11tPuA8Q0W+qb3YvQ2BZxG+YBX7HRs9Pywjfe3c/Gxcqc6AVpNR/QyHsbZxhkn
RL1fMz/9v5wkzQl+qfsTwMxnC5qG+OfplhqkCiHOSQ5TZuY7PbTBz45wc0Ykv+kGFs/+BjSFK+X8
lIHVS5YKWqoYa0h3PPPFpFVxP3sKi7QWUiyri5VUKRmxD00kOSHBBDa+OxSpC+nxDKy0R2EkMAc2
HunnMgq+X6KbGQAsFlhKgjInmYkuuDhPB8FbGjC3zYcLm48NlfIb/addoMBXzupL0Gjdhqmn4RkC
v1h6lfMsM46IH6mMmj/ujZj2GgUO27VXIlZ7s/t8VBknXnNuq5h1VuROb6dASV5qchVUsyRDQKie
G7D93nzaTOZJBimENPayBm9hV8laflG22jGUWyzM1k9mJTTF4e3Yl/fRjusvxBvYtgGqwIzEQX7+
Q9lotUx7HRhn38OXTPRNOtWhgQz3SU8yzebIu8SBNswDXjedHaM5smd0Z7zUJFLouGsSKKHp0k/a
6sR42kqFeSekOtDdJK8omi5XOwwdhrTg9ibluK/zl61o82t2z/Z0/A6KPQofTVVdoF/sPNcSLcob
t0mnhuYUjHRt1ofgtdoZgaJhtnnTaAqbPB+s8/+2ZcpA2rqqGm2/ASk+7go1I95voyFeBztbQ2gB
Vuy6pdM7yggYmUcVMfJ0kN8rlPrcEJ9eHRoRTWv0Q5An4PfTzSSjUiS9R4uAoCDpykFA5Fhipviz
ntH8T7x+cA8G1aR3Wa9copUGtVtRH32fhzTXHURkqhvolpiJoT5CV3HK+QFa+u17Bd8O54zRAxYz
BeZT/ubJYWXomSxLREzY4qVE4INkzr9kaEdYbZZ+LLIh/Q3nbA1UtLhkJsU43mezLoAIGDZIAMYR
C+QDH0zP4z+4O0cs59ECDgidRMZwxp6VpfzEZeOkVTtF3cttFK5hFHJI3gZMmd4wjnP7MZEqX9VZ
fspYOG1jZHj917kEzkC8bPTJ8acToBUAP9TuedWXrpuYfPnX1QvtdRsHvY6ujiATTc8+mxiDlA5S
ZyhFeAX4jenf7CYCypby6gVJjree0WhSQ7WzMUbu0U46Gg8HeaSTzPO29uvSaf9sKOBugbJmy2DG
AZVJT62oOtZl8D42L2v6voA/Q87DhH+W+rp4RcO5HNyJKfLkzGa0KqSB72URbYs4TEEhdHOm9TlG
uGFgo79DFQNgRd/IlWyUFtRRQOduUPOSELB+xO6PRdox39dXB59oZABd5H5aCZ1G4BU/KBdo7D41
KrLVj7wWg/Lb7dpaBAvL9hg34MjoxT3E/+JNPUWT3b9djSt2mCb3WxCGu1OhKaHCHXJl7mTheT0q
8d0Gk0RlzfLfbe36hBnQacB0yidc5z6r7mlMLjSPR7PACWBr+xAqLKCFll7NvGkYhGWUHLZgxoic
8smP3f/ppWZs5ZkxXWTUPsEDAkdOF4cjvyvLHJfy8dVGi9FjVmHjvFFq1Hbqmh4dCO6101eBJra+
focqU0RG5BVSAnunbk9uEGHlB6nYse7MDYnz6W/BDRi6PoRwOQWnrasbh2sUaOvgW2aND4XM3hcP
MlNf+4U3nBS37KaYjRJ6d6LeMrOWG5mxKSzyi2+MK5gAV1RWM7hCMFtS+GllE1P0G9Idp2uNVeN4
KxSwuU5VHF0lZ2gDi2TJOtA/mBns5xbqhgze52D8ptVEB/Y+sPV97JlR0ovgMQTSf/HEljwi44FG
VfizsfhQ1o7CGVO6tkBBLyRD7LckTd9zB2C4Aztt3iZswd3/6YSnPGuvDhPyl+P4QRp2Pyt+NZyL
04V41Ko14yWEu3LTx6u+Uj+Gqw0iO0NwCvQn88u5olkTbo3eVqv4aq3kpmBwU7KR+hC0G7jMAuxf
VmMDkTBNYd3xkdzaXr9VapTue92uYy1Q03p9UuAVsm1LPF0lD6KHssN23CC12AoHfOS9QI+856Vy
A2ledTtaT295XmdROIK8+1tq/wRzuU96A0gDYmTWLrKkNVTzliFsZ1hD+mqBudJL3YkvNbkj2Kkq
x4jY2ktTK3LlOXYNFNfnn2boEo6CTefcmLkpOv7IuBytG+X8GLkLSnm8RPuGlTvLB5ksbcgeZozN
EzcgWgBliPw7AT/7hT/2bvfIa5PPypz7XjU4LANkL3EES26//HldTw6zj/2fmhwyJy06lWiww6Jy
c1X1VNDN4qhQk3p2eANrA/Ck1UrHxxDJDGUQ66wKZyRKet3O4d0niP0crl2cjOSnJm5tvo6fnXT1
1pgFk1nY6QRp3wrLkztmX1B62g3Rc9+8nnhzI8gV8Wyg1I1XGl7oXdqOnMc57grPNyZT+fW5ry+O
8sNRruSem79R3sY1/AXojxXbkJtl3CebUsAE7KhYGUM6TMCZ3LmquIKBDYYkXLkJPjjweepC4vVd
1HA5rUYxR9xUVFx1/CpWjY5XrlGM8r1uUuTvQiUrcetYFR3MeUTB4l4lWE+OWyDMAsId5mJSXFRb
tjBgqukgd8gsR4S7pqR97jN/8jUeVcMGCHNovC15T4nJ4Xw5hi+jZ4GXRT3BVYxFhKT/6SqSgs27
X31/4hLCekFIv7TfxxVEWFhpGcaaFDUpW8ZGuIbP5iicMx6wDsAzX5CMkSjee/Jo9WnmF5E6hawn
pxSRkcDX/zKOzJs9Zp5hv/h2/9d7wYKPVH/XgGOFUBkAUityW+K77geoASTu49n73YIv473wlPxr
Mv9HRIRIN2YVhbK+5MpH730S2ZoHTssmm672TAdGxPDggGIyuhni2jgzszQYhxeo4Rp4/5N7z2Or
NUhaAwW5efOkuAu4D+QT9Nph1M3nkj03SsOjEoat5ncvJ3wtgL5SWOtq5cnk9J4n4p1hh17ihICy
0mV7vvya9n7lo22B0Nwrfle3lontoUFxB5xc3Rb/KyoRGWrIl/KDp/Egm7ookcfUyX6nf+i0LEQL
+8MoAacEN3VkvyaoZPZJAoD2NVMQrTEvaPgEnpJrkS0ZB2HDCERgg/+ShOFT6jepb0UAcnTxWsYS
E8q+X7czov3Q0R7qBGXBnQDMF+eTBpwSVeDfU3gweIvyljXslV2FKIn5oZUMwDK9nTdruK6HoScQ
XV11Bc3xCVi6ha6332egSJChq7T5RX1P0lNOvsqWjnU3zG5Ri2mZ0Nf92JiTp53DD3l0MkjRaWtG
M4GX3Lv6A+sTNoROmAr1/vQMV9juZLixkimll7Zt5VFag2rrczxPMmtx5dUb1CtE2cScopJmz8yT
ipJDa9I7ItVngVT//dai5hT00BM3aW2BnG6lu5kI7EsmLjkkSGx0ZjiaVwwjUyhZHSNVb3GyBprP
GXM5gld9j81lu4A8/iiQUpFJ/OZRBoV4ztsaqcXi2EoALTCy3fTBIC6CVpr/QW2EdZbwf3Eg+cjT
IONclglvIr1ERelbI+KDFjxp4tlnPzx1KaRJXbEvSyBpYIL46Sy+jkM6UJvGhpUnRbyLuu0FMzt3
vvFKxPFD/6VWpfq1SVoX6flVbPeyQB2eEgfYevDJC6N23vF0214xJWY/8xHohq0R+nxUz3CogP39
fhgF86aX7jrpb4tKlzUC5nItXXzx/pqdDHwD8zVFiF1PVXAyP2GcW/imepBI2E5uMNq9Copjy3Hm
PP5K/gqZZlHUPmHJCViHQRjB2AF1ir5rIOP3LDUBOwcz4DlGZK3DkmVF7JqYjxs3uHTRLBSZeO7A
ul7FBx+tCbZAZ8Mqs2+0ncXdfBtlJhXwxVG6PguhSD3AhsE5brtTKDBBfSdg4iCRYKYCRra2TPqy
M+bWkdQ174X5ejyOQx1FjD1BmpRWPxnzW2S7hz1Z1csGbOaTeUi1C1wxOS97SSaBk2SujPmlrHXc
TyuoEgb09AvO2Tm5QmrztTfFmnjRS31VD738jx8Qq5Z/TqK5lzxKhlLHlSo4MINJJAzkT5fqjyxk
nhtx1cs0BGE9yXEzc9fc0ATIGkJWw9yBVEbVUsyutFP5zPxjgcRHt1697REUYBMFOELVCwTZMkRx
AtU2W4/LCAtMusDTTqEeMWyoHoVgAP54nkKnZ6PfaSNoRUCO8TRxYfd2ml1D1MEtHYWfYfFdKsO9
OvampoWuiyaAwY0bfqwwJ7csOHh+UbHVyY0qctfgWbOtyCg8j4QpBunhX0emEQFfnNvNVw9yFtnf
4aBRV0wZVVy+zVaSffvYJ4z1bh79R3AeTw8bZqASyCo/fTWeyRiKVz9iVjHowb1ZReUV4WfI1Ssg
IYfuzN9+GV/D5htvU8Eo5F/F2hTQ9JfoPYSxaOqxnYl2tb2SuaCTFjxNeTUTDpoGie4c33cn3V70
cNAue8l/9heCy+Di/p6AEJa2zHsieEja74Q77j1IN9qhY/bIz27jPP1thSoCFFb+Uhrz6l/XtA72
6XTtFvHA3w9Q/mTnQY772e+NKC7yXYaebr+FFJ40yCJxhPflU3IP321Zt4x5JRoAOj3/RZkz8t97
rLnuNmsCIsizRAANX1zfcjQBDBy07nkYOXiFviczgBIDwxM25T6ncvDRwKpkpXYVuS+LAJ1vkE+U
yuvzXBQxL9gpBQZXuurlaONDWiP+dl1mPTWeOOsygh4SKr6uPKsICdXPgX9QdCoUEOo8e4zzTC4r
R73vxbeUsN2/WFe89620kAeaNDOm946y7K35NSsJFDyS6qFH0rXRO1+K/v82jpXkH1IrO3td/ywC
KYSqWVEtUod73W4PG5IAw0/SA7SygmItBiDDxIF92af5IUg37KYHPmqjJvsRYY4SKgzZIcAqkU56
xPVZDI5/rRmRO/+ETdh7nbf00SSP5xhR/jpmr85fNDgayjPrTUDLxDA1u3HdTQMMWiObuGFkA3+Q
9V8QmqV1kVC5/tIJMXB9UKZbHkujSjD0NuB6fGYbv0tJwFDAmnVanvwfnmKkgKYUV8+uboYXJiTk
UTprRyWvJ1K+95WPm9qFFo3Cei0+HodkZH1glzD7EeOvvvq19iYQm9RSZqEYbE+QDcLLON1POmV2
c2JKhg4xO/TtzMbe6Fo6o9wrwPPMtgK+FbLsixzMGTaYCmWTmhDSAMV+5GPXaKzqXYVz68vTzetY
AHXduXsQ6Om2eSJOY8pvaKzV1mN2nUsBXrUNPPuB6voUPC8X35Ay6h37w+aNPb+tbHUT4OGRKOxV
zktdBghtlx8iQ0OqVWtMYCey33eX/KXf0mPTnJAG1Zk4kdx3poj4H4jN1+uWtGQFeVQJYz0EmvMh
+7ifz9zpzZWrMSXV/28MQ/LlCCJke1V8B4DSmeKqyKRVvQDYG6hU1slbhuiLe4KFt2CbUSyaxcTd
BhxiHcN+KOVaav43QnrbZ5ObyvVoz2wlefqGQjwhiZDwYa2bmYalxKAdLOAb8yKggX9ZOUJk82eq
35cuvdNWTf6HQB3/HHRoppKdJoBuqX7Yw89mIRPVpdwuNFoKJL0ISlcBsleUfMGHxMDPFVBlgr/r
uh85cUulMMLRB0y7CYqGJk+NhE9KmU1Ipgtei8zT8A3qfJrslm416SfqIup+JIAMYO4O0Z0NJXII
uOp+Ies6JktPAPz2aC/oxmtnSR+wmWbdlkCRBxdq1fbqASV8Ldr2g4ixW+wnWNU0imhA2qG8oNV6
oXO8KHubaq6iGIqToFUEBp+z/Uzp22s7ylpra+f3B2llyRS1bGnu8UqYR3X/Bk4gvkGKaSXYfuN8
FUri+RaYaTa7xgHJ/oax09z1PwHmxfBnCzUwfo9SVRTHH7EvU7HrF+KiU2xANIvW9hDb62sv310x
VO6e39/n3bp7RG/3lwSam9W7G8XqbBQKzvIk5Y1suJ1I+ya0vkE/WSdnk91iBMfHh1A7uITgNzey
Y0q03I2ADy93nwEvDGppaeve8qEAlicnaaUnClUdl/m7CeDd0WoGmFe7CWVt96fT2Zz8eh8qJ8CH
3FaeM4L+AelaimM6P9If+dYWsuFEMof4TxbAC46NHU7RG3sryPQ7Bse1Cs//EexS4vLjk1JmavNx
pLxGdFf/aDCKimqeJ9hV6axnLa7vU8VPm5+jgR5eOIFm/ioLrCVX7cu1riI5BDcCbwAib7D+Hdk5
rrBDrrK5s85yn0LDjlfFzjcroeJgiVJgtpLHhEvB/67EZzrbFE1jXro8oT5dzWco6fv/DeJGSScc
lofDKXy4J5eH2kAvo+Ob0HsqQ2lInS0SB28v0AkXHwfhdh+e9WTMRgY5orLBT9bCQVkrtusBbkGk
6KvKTYpzmNiW4q4LI6yPZYAcFkQ/IruEJcWQr1LaFDnQZ3VFTgacTNur8SaT+8mVjxyJKHcbW/Aq
B098MJyiwa0F7higaP1kuafvdr0jV+Vc5YqJcTcWeggJexAiOLR30fMn/cplAEwuVQhKZi1f3VW9
oJwWcXw1PfcCRnXEP1/KDxMV0fFOjd++YIQuHSSyRsk43GvxC6wLwA0ClkA4ydKHU9fh8CwKa4AN
pp8QhrIkhIB7H2htbhP74frPc9yW5mUxOVfo+rv9KrELvR6oAlMD2kScIEqc8WU3VJO0VGpU0NZ+
F39DmlHeIKI6IOpCFO4+I2M/QBhZe3EX7azklnCfcymMcIAQJE7bYF3rK6NssJhf2ft7BVtsnO+E
tA8GA1Ae0ksJwtwc6dhrU6aZazMvwjjFFlIPQMCiJExxo01reRSJ+/bNzPlwVgBcZf13jgzs/pnN
Jw2CvETJ+xdOokohjP4mvy8S6HKDDA/8qkoUw4oP1bFDwXzV3TLOZxYmQzp+oYsYZWa7T2/Wpw9s
5rqOfEBCQB8D3gELK0FD62gzda7VIVWotcRtIYC9MKnN8utEu+2fOpxSbGMe+Xb3JpPWrDj9IKNb
DWT3mT7WcplHL6+Su5Y9LlCmAd5ufNlvkks+sPa0UsvwbMqz+UY948RmEMa4zcM1LgtSIUVdTAXw
XmC6dpUdJxR8NdlV1Y5uuEGbJfylSZNbi62bkW8M4eFdUaZ8q2fkNDsdqCq68Z7p4s5CJpu7FJsu
JVPC68bqzeDZdb6D9QgkCx8Fq6OUgN56en8vpB7RCF/6l119gi5QvHC2ADRB6WZAId5orEoINXUG
xI99JMy2LwncBfTDELUIB+zS8h7lcoCA2WP/l3shdbbYQsN29IKOC5ubTT2oU5C8LZIipoEzPx9r
xCwZuOVXDaZk7TT6x52CFKelsiPBcf53ATLgdcRGqwJMLGGrlDtWUlP0IDkWxtk1xgiLTHSz9Ycf
+jF6PhAwqrA2OwgaaqKdwyJzFAsR6PXfH/wJ352dvLv1G3F8F9y+HwZkdKmfQ6/Nz4wKnFig/+p9
6bKuiBohzKzuE0UHo7lvJzDI5tnJDVVmWRY3UGEL+dVMsrTckaNjkXbbbeDmU+pbglCyTR+B1JZW
OVEpVYKkNcroJylsF6JkdCDnLWIC8iQvU3n9JLjupk2Kd6eK1JqYefJ0156Ozxn1+f+VdKMAIGCS
hUUPlBrSS/9cFxGogD4JwKN5wfnhKjS0MBLWB9QrezpcCGlsil2Y9kOImyDMOomyh/zSCK36x/Eq
6FNlFSbkUpY1GCqcwIpPQXVwfkA7jJ6Q7AjDE7UzPu7tp5xFDbIFlHQKvphy5+LdAfkL1zB/Wgh1
StzQvcy1lsysJVVk8Sk1U8wscrkCO6Qk4B4NPQs8vXoKdpLNgdnj6o9XVuYq8fd0fbT9k6grEV+2
lnsEGaHKWuai9TZQ45jLDvnuEtaHmdiAfxG892WS1jWo/tvEw8VuNQpmaI3WXvlXSefw62jX/neR
J3euhDJ0xVBwx07KYCi0QD/fVN427SCvCy7Od1MpKoVgWMa41vXuTQ4lWA3GUk+IGO9jLC1K7nmt
OMcL9zrp2Cc+GnMBOk0IJwy/mC5iK0s4fuO3TfhsU0iLSV6oKoUOjcHX3At78w5i1WA1rGxrVPYT
ceij3/XBHTR+lCEf1mlI2Pn+eQPGpQCDeZwWLl72YnvAn6u1rl4WW7JBvVFQ1XfEXDH2eJZ13fyP
MPquKum1M3TMnYlVrTk56YozUJG3hX9qnzO/b4zfWHvriHOAltJb8uBLIQasCFWD6DY9jOSAuOJo
TMjAG78BHt/SyCY8zDZEtdWTVzyoECZnmqk48ac249E8epRNyROHUIrdbPj1PsEL460H96oMjij4
ILMxrfzxYrRFUJXgw3He5q6hqOysuVtXxqFKJ9C8jvPnxV79X7pa0Q7VJ5mTeD7DjMeOzH3EDKoy
HKhYomHXtcu0zs7P826tkPG7v+DTguVGOQilZ9xFukEkHuXAbXEs06tTdtA74FF1/aOvJ+tIiuGJ
p04+VuFN0chBRH0rFkRFJHPIAGYHgE0vprUB/s4zXeepuoxQYzj8vu/bAvERT/VLXDUhh+IdiR8B
Yohu1BqmODTcH4LlHig6DSi62lqjPzh/R4sfazUTb9Zy1kK0FhxeWlXZeTT7qU7nBTwbaU9T2/MQ
AI7tRTd23PWtjRtGCvH9WYFep2EldhXT/EyPeGZR9ths+fj8Cd51y6FVnWazBHzxlLIltajoZWc5
ak5L7qtbsqFL9UJ5hBH/M9WzQtlqKQTwNwc+tTjaaSFwgKmV5MTaj0JdgMeV0c4WBh2UOlncNB+R
ga0mcOTNtxr1Rb7/I/J4L8F8zBqlM/JSzHahXtPwb+4wwyAeEEN9/OJFd7vWHnBnxBV5BySd2Za8
kjaNYuUjJnlzsR7H1Ae65fhIzQi0r+yJ3QrYhaUM09PiZPxmKaRiCeuM1pnfRrXDDNV6SAQQ1+wS
EFl9kZIOsFvZn2Rkec6cSfAkEEwtVlWZ4JEIPNQJ7ktnwULGsO3IwnsfaYMzj+XPoSU6jtMdCK6Q
Utv7USKozdL+xQkv/odJPP4RzV+dOR5QQe4uCXsnTYsWcen0Gy5jiJRno6vL+ulsrycYgnViuP28
HKSe2IXVYWMnbgUyRobPVy1ATiTcSGD7m5C1WoPZN3dpJkU7pmpod7+aFaGuXfGqroRMnNHj05ca
tbKybTjo4Zv3Jg5z6RuzNkEYmU04zKPVypRYdwZNPGc3oq5GfFVGWZ2XmakdBHnvQwq4vSygpMpB
O62vT18nO5lN/m3YcitebeyKUTyzACLXaNg4G2wqlZkkYfceilH98wHzosvJhovfyJXXIXm4cLtp
b3fDoj1u0BdXEzL/MXUTR6dTVI6kq/1/aQDYjyoF8dYz9MSpUOGGXRYOLp9Ejijjkcyvdjc0RxmZ
jqxGkHn6D6a1eqthv1zHO6zy0nBLG+KuPNRwrnPDxFXhgZSdA05ikUkLDnOvCvZ1LOwZyvWWQa9U
SMrGN7WDWrMvD1QplwVCqdLUQKGQ/uD/TNfYpYq2db4GIzvJ5/keLgEizB+iDaNfw/sC7Fn2pC2L
Kn9GPKtNwqi5Vv2m8n3pKTD6zY+/B7sgeGnbPyl+uWlkTOxq5YrV8qU5BEzAotff0ReA55639/vD
MUdRvadmGAQBVcioyb0RqT/YcGTyKG1p8BN0JImFxq1zBDBVxB0gcLViMFsvi9Gg0gIoz0o3SnT9
6+IiQYF5ecMm1CtZocoA5XTkg4KaTinvaUaYcn5dmtivlIIMbAMFC0lTLeu3TomTV/e0DleeoyVs
8kA0ZhFqTcap+PT1sg/AgoXOC3YM7eQEwL/x2RtKvEKSUb+Jm8vDlFQUjRJJo7AY82qbtst3RY7o
ask/EtpbbdJGxJOjl4iguWIoRoB3xKUEq+l6++PGjnUYDf8t+77uxwHYpZNsKkybnXVrfDTnpF9Z
6ODlGjMZftfFW6GmT7RZ+zBUI5XGHstfjJ+FBBsdWieTrxExbfyZ9qLUw/Wi6BRGkZpNf7Rgcytb
vKzg8rGRJr5zfQ74U+mW/+aKDp0imRtPWlBqU7Tpze0N/ng+LrK+zK2hWMGviLoCSUH6EL99t+IZ
3iaQIabuD6o6hXLNMunLwWfMGNCf1SEKgFxQnNe7CQgTgAcMArIEJACMsEJ51DPCx0re0UpSGc4p
xpUarkRvK9Y20oy31mEaSZ8HUG4ZM8dwDok9thf5U6leeAtD9jFMrNodKyOwpIjs6cNNUeuPgXnA
M5qTwjWLzadNmjFlHSxZ9f8L+UBQkIz6WM0ksPE8/lqqwqsKopePu5czzsgZ+kMf+WHkepBMCiiD
2cTeDDV/fjleSAdYU/8Ow+VmXNbENjWF4ETtI3DoEnhszyD4l7npK2aS+RVEfGEi3QNpEvfiUnci
UV/XZTsBgp+Fcfnlzd6hvtwdw4DlbmbLROzGqWyBbuT5uPalXsHhf3B0zdgLCK0zM02PKNFrlF01
xEAn1nhCTkMWX/cDmOMoCSJEgV996fxkU6X7G4meimRFs03c0qYL+EDf9scRDGBvZ9UUkOHfst79
22KSIxfX4E2aJovYUAOUy2WaDsnxpvVbLTRU/XAbmGm6nFt1n51dJTx0NHVPy/tZ11JD68UecstQ
bbvU2leprIOyDTWOehpnPQSu6UrrlvfZqxIAezJvCKqPetzSg1RGcoMA9AYl0glD+Vlqiu6PeReV
66V9Z+Z1bXlyQwGKChfvGRDfeveKcRB8Qh71QmzJ3L7EoyM2bCu1PUGeRqbRJtgyp10vMiRGdxyO
InkmStI/rtzZysfwIIGmQQiK3l3n1kzra7iALhDnYAWgc6p4xs+PisyW4k20QflZvncwPOxtUN0a
33k2/0CCkgQzuDn9/RwEoUuAHOxqtgxHioP89+uQloaphveEzfInlCybqps9/2fJEaTsccG4P34c
WFT/1uohXfIc+G2Hlp/gA+Ji23lsCW9BQwAjbrvyW7TghAEA6XcUJHMQXCkLfFsE+RJCbIc4s552
qFXlxqQXgiRRkmN0RmGzAWfRAup9wYFXDQLKceGGFxZFtefpOozqbucbXVA7YTm1jiRUKyRF9AuO
CrORVNwqbNckPkIDCNhMvV7ndiPcfpzkicJXwpymOE4LDCPbH5NtQYi04BzoQ6iqf1hKSpvAPFQu
R34kFeQ/Bhw1QUHXtCI7ztqWHobapZ+gcsRfy48jZLq1q/A8LtF9qZofw9GiO1oYQvvzSeN4DKRL
3QbPzdR0yOiYzxeP+T0pYydgB+aaiCNt6W17OJM5aV6BrDuVhjSNl7hz9i+SrhAhdmJRG+dgdnKL
v39rLlsFhTvKj+eG8r1MxKSXZjilk+t1UBvZwuMGpCG9VIYcYpskQ5vTfs5GzkiHLpwdhnjvIM1u
0et0Bxty76Uh7+SofFFMjI3i5wCeAFD/I/JY1Uy87PA9DW4xsFHJVezA1hBJ9I12OzSqgbXay2sc
wzTrZIFKlXC5waOgK0k79D0MRb/fsHBDk2PEaTJgPkr12lLVhJhGqObLKUFT1HW0MEr2FqYc96Hd
xXFC2aQjZ2OnlAGf4IsbkoZBNzr3DGznZp/KTQ/cenIcjhubM6pi1ifXzE0lVsGyHrGXMn1jcA+P
Kc7p8IpXcFN1AF5jI9jxJ3VLDzj3om0KIurFSgBJufGH4VDuRrrsWiTvZ5hqI3J9GuzNNKKVLxk5
HuZlMCfrr25sK5yn7y+VMZbHJvzr7MflFP4mXibi7QQQFexObT5XHw1Q4opC1TRvEhKbhSyApXU0
qTlR6fS4cQe+zxN+uX2K81GZaIAfwD38EHxm+MBqyw1YgWOojqUGwWMTJyAQaZVaqwA3npHXY/xv
WV7DW6X9AJIrkfbBvWkVy3YyZ1sIZsIi2vaKxg0pD+2jEun/WRU6i+8IeXrzHtv37h4EmkQtQuF2
xT4vlokb+hRw3r0y2tS+Mg1f82Q5iTHLvTMUpkgoJi/zTv6gU7siNc3PsSZDvsG//A3FWr+d6007
cnznPEkZX/I3YFOoa36GHibm0LbBPdMKiOVZbXx4uMXX1e8JSFG2ZGnyoXKHzYp5xWS5pLlX2VdJ
eWxNNA0G+5Xfi2GVa9caDT4xxuy6YzfLOfd4Ov/g2JBmofFjWXw1n4AK+PxnOIzpoTpcNkijsW2c
3EWVx49uSaG3qhw5sFmEQwfehbEmGbcU0e5gkWnHQ9QWiGo4y3G6/c1OVhoayiNBrziJ4bIPqzyW
yZ+PKG7ygX+oy9U5omuQ71pY5ycRVXjGtMiZZA0Q/VSL2UPaYIAhx5E5pzaNxV4FcCytlvoFr5Zr
43omBj2MadUJ0PcL982+FG+1BwzsR5fQdT5iFVh97gsuLF7Ds7aMVjKUdrvkdobN2AbdaejBoTqW
L1V3XLf89oeqbiSW7pEkTyrWu0z/+lkgd6ZZDlPL8pV5oY/8XlxOIH3in8wMt8HrkH2cd8CkC7qh
LaEWFh2Y6Ai1TJtNCApqzIDMXfOwi5tP2LkOzmVCfNjEafrRPReI6UaFcAfqNd1HWp/2EpgZyZQm
Q4dAFM8ZjfNG79zg9EVq+Rk92SNRzeBVM5IlJA5SpCX02IJQiNRm8u4V/xulhOMm4vn9RWymfAoj
oqhQXvIhCOBvlTJ4LxsvFgcL6fHMBGmopLI44TfDGYsNBlixoHyG3woTVSKuO+yPJnpYzwpJS9eI
YSjJt8tYcvinJDF1G/sVnmcrQNYJh4oi05blGXBj77ReMI3UIp2D/FZIE2mtdLpsdIrQP2/dioxT
/KTQIdFvar2ms3mjSBptwaULwhOZyaj3YQKVHpeyTOlr1384NuDfv+c6eutebu7kNwJmHZRa93Wb
mTxrEEqAdWOb8KyhUbp/0R/QNYdkp5KAu0voAQtsIOrdssakWhr/XsmZOkDvl+1UtkbXVYhBYL+l
5Bp+lKC5q7CVVjvfjRspExOSL9s/d8ArPwDaO9Di+mdSdI6BKUsGtF+lrmtXKVtJ0IAefSE00/rR
ksa/zEFV0QFTDEmTI9vOjgztdcTclXq1lQOvkVT7sNGOW7A+YbmKsIn1Qa0dBqBXToclfKJdZPYo
a1wyURB6QhW63PxmzP6anOO4WcAa5ELrkqH7OQyU72aVhhlJ+o6n8FB8yDpaBlhNfl5ye3yMBpKV
+Jrdb7qkYE5zIkYa5RLwN8JpwCeQuiksjWIPiMGyvJNIl/yGW8F1/BJ/ARheMNQXYVdZhKn3CO+B
TcDZCMdMJkjQka3yTOYA6G2XBRJPLGD/Izh4KglK6ru9LvjovCNQQ+wEudZyZPqsvsPxVT3zUrmh
MW6AWtubHTzrn+zzlz9sbUCjNnes+V9olCamNgBKRefHZaGBXZKdpwQZJkM/oHOvnM4MxXQsTPiq
S9bg0vYBnVgiudEYTVJoz1bho7/FVf7pPozd8SdV90CB/281/8QQneyg4itmjoOl6oljgn5j1W7B
FoDEbF/LIhVHQj46qV9gVEIZH/BfxR1EaqlhPYUqNCoLqa8ay4kgQ/GytpARwfBySGD+Jtu8l+Xv
xBfXZDiSnkX3wv5UMVWjoIyHMvXn0n7QuddAwd2Q2xrybppZrIxM6IPBOC2wJ2CaHB3aWh9vJ5S2
O2IVFFSU+3uRksPhrzGA5YCbK1CpWUNDqdNXEtLIOqWCW+shJphzXuN9f61ay4lspn84CWM9DEdA
lFmXwXHMTBaSwNNFpUQa9fYAh+Ej2zQAqZ2r4Sxx+8QMkIHAEsRo4CKmcCHRY/QXzOXrBCGgojSH
KcskxXYJHoPj2KEBOxZNX4iXam8nQ//Kj2WNMbudaFWXWpzjxxKOcrxPWnSwK8hNt6J4nJNwc3iS
sp1ntP9QcGmvyHPY0toaUR12Vx93Q+BIoKStrN4ogRBesFBJ4tItxscaVVsISl3u45FBp98KEA/3
nS7fAbKtWb1Fpr90xWyWvpBtlGSV4ZkUvlTjTvliD1sCc2wjay3qNVXIv4FYwoeTXNIFWvxOnUrB
vSt56t5T8n1i97FofmuUVkHIRkgSYkDw71nwovKVxM99OziH4a2UHs4CYZeQgHJu0a0zLgaOLunc
ZdfaxurLCP/PtqXliLxKEnuwwNLysbO63jkD3/qmdeBAWSGCjRafpaQ/Zbom4rtJXvlSNq9AvUyQ
jyJHK0JAxWx0uEbH48Kt0e3umC9FOQKA/oZ03hGijppyqhgC6G10bj2qxfvkjWsXFr/M9+p53ERD
YqCd5V/7+Eh1MNDAyRJKg2lCKWPqElbkXyNgq3GNnvvvcuLct+PxR0hfF7tbjvkUxqK8mYmH0jQG
Ftm27t5+4QI0F3817jwMvaCnGMP5K/I9SWAOqKVE5X8ltUCAgLdzpLOvqxlZAW8dpy81GBFsL6hN
wKwM/SGT3zXDwxIfpjTY8i+NrVPMfJkn1YXg2JHdNc8NHtus2u55pf6Da9Fh+MQ//jGWsg4a8aTD
NqNeUwu2J18Xvewi5KlfF4LJ6jAC7tKerfmU/xRVjou7LF4QVtEKc5Ha8RctWaQ+h9+W/RpRB2Mw
l6aUqQ3WObrmg/CHcvepKeeC0hbsmvbRdoZ56pdn4z57dJ8ya9XrT0/8fd9+7LT/TXHFuNIBC82h
53J0wvqAJHiGsO+DtZqC3T3/Sbg3maKy0dwBHoH/UVGo5AR/HSPeu+xgCSa0oLJT1N2V3zrHhNL5
IXLFIfmFWMevLo0QdHPWqeo/Kx54AavHQumGI8CjVigflNG0ppe9L7T9KaCiVHAU4y38Xl0djqTV
TezitIwIdY/qvK9WuJIWusPthzlz1dEkWPWMidTm+ZZ1iU8zLYnRQt9FGgK2FbbOYkxEEjLH2Nzi
OqkPGiuX5FvpYVyBNKBgorO51DWtwz1+YKTAuzTArVJf6cdGs/KdoAU32PHvvulVq2hiZZ4DyfdG
ClfFV/nYlmMC7eqtCxka3vZcUcvB57YXqih9yHzDN5Mil+uXbrnRC5iLR/z5lnJBNO0iiiKBC5fr
MBRj/Fgt4Y6PGWdH60wDLT+O2iEBTj08ImHrJsS4uDzmtRwx8uyZ6rMdHpNJIBDU+fcl3DTczo4v
JrrDRHpB9BV8B9DdpQvTYXwJ8L1Kn5621yPXNPSEFQ/asapDm6OmbgL2qwiAegjeCl3zRcn9wAKk
yMi0Rfq0bdyXlUO3gzr8NjyGZQut5jkZB9Hk2BvnOchIaZubA48CKthJv558Ej4PxXpWJgvOY+J9
xz46fXrA0UgKo3XWBtD39syzOWcFoxMINE6uHWkNWjQRXm5VNjkdzWViCZCfLFi/vb9sGwGbLtPq
j/dBojdFF5zP69HarQ/syrofLk8F4Itbyc4ym9fIm3y/hAZp8bN4ZPXVw3cSkpWZQ1uswnhFoJ8d
mD9i9l89TcrgPL/GklTm9H1WqAdsq3t6iyRkjJSwYV1RLuUIep9SaaZNAkhCkF4X/MxKaDSpKEtl
wzNWyLhaIPorQ8hoT4PT9iFPonFCqZUuz9qs1wQoWKBV5ETeyivoSBfFj8WAeKMHnWxQVCbF2Eul
3FcHL2oE/uUVkiyuQLBIhDxfW88s7VBBpsYSglhcN5nj42wLNaQDDxy+R304uTLUd4FWSUW6yxoq
4SR364/IKKHuQgkFxkyoGe33Fnlf3XCV5D/gmLrKtN5fkr6sPOW2ZJHtzXo8Xa+mNyXpFuwSa6M9
U7eO1B7fX1PJulRpFKMXousrCxagx0n7ZgNO15g9HdqHlfpSs+ULmb06sqrqTLoUW2aXNBjgelHI
LK7JynAltO3tYngSO1wYaOSkas6FVOpj7xMrGbXIrLIkiTJSekCG3AmELyUgBT84cAw1sn8qBb6/
5zaIj4W2+HR+zTdNYo0I+CQ1nleYh8goxgrv/cw1Bs9JxJAoK4JFGAM4uYRd8Mt3JFNFFNlS4VlY
5vWqOHnlMrY8JWvHQnq5s5C0Kc1rf5rfSY4XCzdyF/GcNP/mJE+0T5yFgv8X2RT/ttbIJeEvb6zU
PE4Rgk+hxErSA/5KRVttOF8rz4O35g0/QlgRhPQE2kDclnAniQPLrWq03H0OioVB1IBrNcIOBUH9
B4YTYerStFgoP6u54TdaNZ1JFlG7fRozaE+c6ogGKNQvpbC3Q4/1wV8Ke457v0ksS4rANE7JHJvY
T/m/bDoW6915kLPgG89H98dnx0/T4hqLZ9g4q2avMC0SgKxcM2by4AXCzla+pfP8cdBcsETGkMsr
1cd1HvOto5QD6lSdOLc7uwUBhaJKSabVmNhkxaexyyGZcESBEiVPwrHCc29Pj66fufQA8o+xpHRw
hQ2VtR0XW+xTIC/TGnwWXsqfISoiwxRbuw3EUn7SYW249ojAZ23tVXgNJKuB6XmXIAK9d7GqFHrR
9XLeJjh2nzlFIJ62YhfPFOGwGQtzG93p+sRNIKNsvUG+na+LYILUpe9e5pA8RzKXO5XmWAEhzdd4
oWddP+iLEEYulSaKpjCJx3NH59XFgwRX/gTY+qLdVBZAUF5sXnIgR1/gAZJp2/32PROEzc9dCa1z
r3yL5Su5++VVD75GlQw13BNx8rCdznyEENL26X36ohAyiYAuJkeKvMxCu7rcJ9Lxy/UlI3qSY4Ks
wClAE0bf6eW4600QWFaHViGP6z9SGFGf6D7BROr6zIKzdNksQ5LvkXKfIVLFWBRdtPwc0vlc2/SX
m9IuykPjgRKkzccKe4EVeM6K202nTOdeoC72g3YdEWQBGYAOClA9GojChUW0m/CWAOkfRHzq9RsM
ATZN+orHRe2uKutNyNO+FbzpCi+B1v4XhzXQn3BzXYTpnsfD/MfKZo90AbL14eRaDvIzEaKlCff9
KepTfntXSZo0wr98YnudA+/xYHVtXLJJAxHWUk2N5DKQ6LyvoEb5uWcVsuOP42ffJxcIwS+YZNoj
tQS9SE5My9Aqq+lD0tdd2tsJQYXaNBYWE6rSsuOkqMgUlrKBhvS1Q6gGiDxXC76dS0bDz0RaobAJ
iGucKP9mUUoKDk3Oh2n6TnAbQ8iELkqDU3ipR5l7MCOASY9iEuxm4T+mrR1h9g9rXdW63W4DLqSZ
p/ADJQzjn8CmQWlRzon9BVVGOQibokJY6poZnNqtHiGm3AvWhquUyMZQxE50EFvoaFpm5JBTRNWM
rhqHby3GMJhUtI1VygORLhWC9CWTnpqhGHNFxof8PT+2zjKIwgJO4oimS2cn8VlgWtY8go6CKEY2
+obZtqrS8CMRJsI7jH+wrcxPgC4IUj7YCUsHimsO+1iDkvzOtoP/9tuXGn9qLcGaTamYJJHoY1L1
eqgs0T+QV8vxyIoAE6tda0t5Kr8HCfV0Q9Hd/FUn5OXW7X1g4HhdCGhxjOKA/DvbHUYedJITNwAd
h0/NlXAKtax0GJ+e1Q6cKhlYuZ8lZo97s0bdHyxWorO6iH83J0rgnvqP0zxJI4s+783leG1AnWxU
rEeqJjMh+G1XfHT54QpAV2lj5teqgRLCl90ZiUTscjvUsppjD6aombJa7ilAHvCVB2s4Jw5YvRJK
gZaLjdOXX0jR8ew2TVpUaXcfD+maJLyv2xiWxZoty9AOng7050PCSK7DMnXrwkvnaCPwGtHyJ+U0
b5CpMdjNx75nBCJtm237QfOYOwY8mxjxNuj4dujrYuWIkK3u9dNkchxUaF3JlxM3oOBGtc6yR/Tk
VrQmC72VcsjHUQDsaJ34HVUMIH3ML5jUB+lK3u33SjAk7Nb/AoiMTLaYEhu8ZbpK7TjDP0C3l+DQ
dHNn1Zrk42tP0cqCAGvH6OVWTWiJlEStrC+5kO14v/1AvOca6kUVmmnEPoib6d076yUJ5AmDcjUZ
8chUSwLjCfqjChni53HOKVlAoQ1P8tQILzbZ8nQA5hMHoE37WyaFpXAwpQiPtoGfdHQ4t6Bd9quK
xU1Yg0akD9Yqh4ED3y7Z3kQw/Ih8Y5sY7X21O2B5ekUeBrcQzQECiN+9QT/rlgHnNxxvFwmj+OS7
qwQ4RF5KFOa3nzmKit4PHEMTsN3aKQ6wMMdTgxuBDEQSMF/eeJM4TsYgOyJqEC5Re4i8UZ4mR9Zy
7lTqZnbnbhbVzz8XyJ5UkbV1IPwaKlKr2i0c5o19jSkj2vslpl3kQ8qUknbwQGvxr0JXIFj4mKbm
A3M67p8OtV71RjboJlcOX54WZ7bWu+eLzIQlNlf3YqwFGjvbRilwmlZIJYcqopd6VDStX8IwefV/
BvfOCJ5vRfx3de1uSkRvFKW+nYJHST6bX9zXRKfm277FQQdratX4QI6xEyNi9ugw00vzm1HDDado
Fp7OG20fyaQS8z1PA9j78ViMGXoBgQIyLLeDDosEWeLMGx9ZzD3gfNdEPcxKqqVKyR4s+04HsQuW
YenvtZHLPb/CDY9RR9vdnaYrRPsn1lXP1irpZtGHhA6LecDrg3ltr+bsr2r+ZnTcBr5njGMpsWyh
wTqq0MaK8ucAor0siPLWbuxUJg/nEApj/5NgJHuCZ4rZHQaxBWLvbWJ5ABVDP6DwfstQ+WBO9kOS
KWeBfL8MQGXQkm+3iSpxqku5Dt4VqbLuvIb5leDMsN6qHf3PlheFnixQKgFFmF8MjtrwfyMZC9Pe
OHodX0dTTAnD0pjN6FZKpS4rDcrRdwBP3UBVKTZSuh1frIB8xbMIGRE7UjZ/Uku3c6EETLgmGb+N
FW0jwJuZ0LZ+PU93ERUxpq5Vtc8uPzf+hMjrJZ1+YzPSPsq8lUu5Zk1iqoQ5ggfxWtWrnWwXbWwD
xcWqA7VB1GfhY7d7TbFHZ7PqMzaCUJJYRwCEaUBIwMQY34ZwaajfiK//W2X/7iow9sOvRojUFVDs
5VLtaObjJwrt5rSBUiOYJBs12ssv0G1IJtP0dHONi93cwuPxVhEoJ1KFI306U0M1zF5YEyP7RCQt
l3RBh1LDg9gtkCHM1ABWiLFV3X9O5tS1ePcvLE6q1dudAgzs4xbxbuebEmESIhfL4N9U5hy7NZu7
3d6syrU7daQYHfmu968jitlu/1FQyj19hbvW1nQ1PIw4ld8pmpH1t7xGL7azmpMXl69V8Yp8DJJV
MlBMBEsOAB9PD8iQn0Bp5wyeR/qVznxaM3SKZb8IxbZ2TWWjguNP5N9V+sNpSbJgeVnizkTGyBnQ
t29akYmAUChhFQK2QSckZkXxjJowtxSEaRfhrSJKtP63NfymUBONCubNkCgfMHGtgWuWM/yJrosg
abXBDCVSmkzsPL34isqsbjH8eI/rIpEOLd5D7rG7zaReCMcPqZMkapD75xNyVMgOndD4EVt1rgfH
4pWjhetUtrWDrnSch3QlJGNi0TkapGUPoizBfjCd+jN7/OeDDOeMgxbW3lvDemNwUoeivw0xhxrK
B/9rdSZHBJolZyqImdBLyA9OfcfGwgj4WUZ3CkV/gJgP4b68vhbOrR33oE0x9vVrJysS3FrtJ1Xl
TGRlZilkUM0Vori84ARiTpzz3bk4bt6XthEtdIllwY1a5lrckW6fnKettPPO/kSgStwwvYMCLd7+
vaCvSSUWMFSs9firTerwjYYZaeLsnjUHpYgrbTiV2IDdt1usOL/gTqmiXuXuAaB+GMzI+ItXFObY
DQjkpGfTyMjyE1EQpPgM1wz4ch20Ukto2DsQ7zk6bdI4AYEnR0vsOcYQlWtpXbuAzCnFh3qBkB9F
RWcGvK3m+PK0ipmvaHNlwTsh4tmORZlr5yTHXvlaTJGvtmGlPwVDKGEBPaCbkSH/i8vfmhLQkD5x
i0eWZKNDu3ATLRw0hi7D9IuCy6ZOCQODrCFUl29nqZi4qapYUp/OvXA1XS3TKN/N6U+gwWK11LHD
3L0xkQtMAIgqsNdcAmdHsTgB2DznRjOrw0a/dCRbP0DPjZvoVIOtGf1OZfh7APTGgb5lOQfTt8Tu
0wpaP1+nWmU1K0n912gJF59s2dbBnF3VqA236AR3bTX5mWKHs26hBtWz2ftuPBrhb2rUTeYATuyx
gaDDCXD+vuWtpgPFAS+vyjW6zr3BQYtlcr4EnrwUwDq3bfh4IU4c7MMFKVGG9HXvFbHRVTmaade3
Pga6yC/ckxaf6loAiqPgSZdLMvOCR/JKffATJRHCST99Qxi8ALs18DPuy2EOp1hLR+bv5HfZ/N23
yEWQo4n08JMBGTmphvDkKHgMvl+fXvuy8l0y8S/9AUDZjVF/0R2Km+qnMfzDtMBODAEbA5pWctK2
n1A73WCIISA34513TYRE3dm1ykB6BC7z2I0vmjxenRYp/9MhPBDC9STF5FSUmjpCwiHq2E2HR4ta
EvpPuSEhyNrRIDAMPy6OGImwJtt/HlTbIlzW5jh6TjwnkUgRGxj7ASiklVf7jpksx8ztk+kfS3pJ
qb0bg+CyVEhidyyw5DZS0Po8oqmkgL10hG79LR+vt5KHrEScMe2+mAhDj8QOdS8wurFFwbNjpu4k
DbTQ9oB6HwTSM2vKDy2yJ8DOvVNmZscbv8pgp3csLRDtjZUF+nxl7EvhEYU93eIFgSGStZbf04t3
D2iKfAn77Omai+CcetseXaTsN5NE6oSASNTuE9OLnH9ocbxZJZWV/LKMwV4odcffKkL4LTK4fCrr
MH0niOl2NwEA+89IcPyQQ/Yal8HqcVpPnDf8YPW+uWnyTLK9W2fgdmQW+Srk+2AwrV4G0zmF/j/2
b+SYQe+NDs01kaDn7HfUe07EYJkK6S3buLBGwG0z6N+s5oVdM26yeIMds8IrGSyvCqWVFRI+Z1nV
nXi/1cC2qje7KCREwoTmpcmAJ52sMTOydo1daV7YH49j1DF5aiduk2XQI1rA0YQdYhiq6E6MiHVU
8jTE5R1pAijW8OFnVOm+0P/NsS3zJzgT+6cHOAsS3p1r4Y2ASh97iTlpn6oknp2f4bQAANWs8K75
xBROazRA7r3meCRntYLF32/E2zMYuI+PtYjHTOq7/zTtBoIYmPA2SeibBV0uwrCq1WXWEspRBRkV
/KPAZoEA33EPS3NZxRaplCqYwa1LqbR9+rrOTM9mpVPz5+6eM6Sr8q7a21BMwu+YXW3VUW2bNC2D
d1QKTFSInyhriIesMhUM+aZpq0NiXGyzJ/k3hhZiuuMlxzbXCZ4cv1hFyurI9u/DHb0K5dB6vrCf
TUCSfy5ZqmRvAhLRlwBgTcmnsZMBdqQDpsbXanJlwefdUhPOBXnT/TsU3gepdh6FdhOnPTrDI3R4
5GouS+lUulw3mdqUUKElx3Qp63sWpzKO0Mlw0UhBjXv5FqaSQiSx0sYSyokSVTfu9f8mbomyOAqQ
027cJxhSqjMJH0dLN5anEb09eufl0PIrVSgKfJWmggVis6im9KHrM2xrzbOz37hs9o2lEG0WD7Xq
n/Wz/6pIV5F9QOtWuwow7hmLFvhvyefbi2b2DNYT1/Guzo33S++CLgYwzHJjOfLQ9VzvdXKr7gWD
FV1o8Z2BlJGgyIy4fmqIoslJNVX6lLgOAT1MZPxioal4OXPlY+15flBkdFZEOgXkBmdP4Lb8bVSk
mqXh4jfoO9QmyD6dt1f4i0WUJTpqdoLIYJSEDqGHYjycqol3F/z00cIDww4AM/OSebIB9X3WkvKF
IbIr0ckvtjqmj6xAobmeTc6LbZ8/satk9MfzKOaiBJxWvy7e7d3/jJOa1X5SiNUTdcs4dWHpeox7
n/62A+nFVcy8vTXNBzJi4CCkJxFPELeZhIoORTa99BsdxU5m4byoyUAh5bVYyeCTrxtq/eB0EGij
xP/Yp4s3FtqDaC6Kxw1DdrqMtsPu4881Qsl4VJKgTkmU3TdCYOzpG5b1xNdySMg2QFxSkmgZiQzc
MRJBJB7YMdF72Fzxq7+lP3i1qXnpz+DhuEv/OG6UrI0Uyvn7jDgwk3TOkRgPuvGiTjh8QQTGvaHw
dS9hyxIugtnSYcBX/cB0lsUoiBIgrm4asUOc148lSykwd7uW4JXZvjE6e8Ex3A49w5pcNNJwKGtR
+3HJFotUmWFln0OzYSIwdZkWAdREifEWxZkxlw+v6MEo+TF3PIruFug+gxbktXBywK/KljYSInep
QLdjS6mTJQU8oC7t7HaK9I9z/FQRum9uCv95YTaeP+enfL8iHmhBjqDLi758xhFN5xx5WzSyTqAh
GWf9FHGABPjPvfmGGSKTGbWgcqVhOtzQCSAtZ7pmkH5lDVNURCbKWhnq7EXXIvorLHcZu2hNQIQX
33X8X2qmsCnccSkPa08+HajJPP1suROz68+Jim26+NmtdoyG0f3CwIarh8sr3kHdQZnhv0SEPEQl
Nbh2M5Tdk0amD+at+U+XtKTcFCzHv7AzdSxI5G/upD0w7cOgeBA7E3LqRiU2xmxUSdnaXrLUdrhe
kn2ZQ8ytMW6M4+CAiMXWgWMtiHIDjPP2glr8PS4ohuEKOpoj30pIlrBihkeO4QrdikY7qRZziDaj
oHUFx4/0qoLJwKd20+stPkKiYDmRzgZp+6bIlgWSVLfYkVs+ZN8fZvFAEHdTgAThIcgU9xjm9s9s
FSZ5WrJmQ55xjsvPG5HEnrXXHIiIb+84yk4TW87uyE4z84fr4c3bzT7k1eszbRCFIMaKdRxltLKL
3YvKjnb4NShWuL11bFdGkrPnTHvJTIQEbVvrDeqGY/649KVaWfo/vt5pbdTDXwKrN/zws/y+0lza
DWvANnva3qUWBT7hUNcskG2dgV/aMGnfRPjLfbr3SJU8fCp1eU/HGfBgjm/NVBzIYHsS5SmSlX+H
7b+FRNkgShqiGTrj+6f0prt8xlxDhBBG8jYSt7i+aQ1Ravvbp+CR7NRehARPmMjh8oUpSBBycZ0/
mlpFyHyd/iCWHMkI5HAHXzuMg27GToqXMm35LeinKvrV5d1qm7mCKGNw/LG+5cFXtrdMjj08Voal
JiQI3crUZRh9ktRIrdZt0JKoC7EVgbcUsSaTuu242cT3laQEPCE9rD8mDlYtvja5LpCiKJFpOxjf
mCi8WH7MoAxcyQyyrFlIWqenkbzQXqVL1OERjUj5Euy1VP56DVwL48sg0bv/ixkFj+VOsx1PT8Ri
/P+Bvr8exK6Wa0ZVTOvEXDUWPAahL7JTEpGopezrBaesS3a0Pnu+vZKqrVi0U8bw3tr2O+m6Z0b5
ufIoqk0YDdm73a88qeEBgsuR/7/1ljPkI9l1U11cBtnqYHcONWV0+5W98i8P6YPq777SbB/txMZ3
lbNIdNLQRARv06r26uwQsEVdgtUErT+NTT7XIWCXL67hmiL0QKbJ1+280O5UCaEDCuXSUqPm4S0v
/Jppaa3pyRzAGif8HTAhNFV31Sqn6ynhdIKL7Tpvjabo1G6zmZvFEdgxm87mYr5xfZvlPAZnV6+t
E5DAqZVzW2UwPa+ugpgFK5siaysLK1i7x3Bxoob26d4Wr6SwEr/s2NQQaufSyxzzSRIVPPnlzbBb
EBZSqJZx0LT3L7HgXLcRfX+XvC6mhpGbKg8+OySOWMZb4mWBFq58g5sLK63JtdEfh1ROFlCtddF7
AmQnFxm92wf2QEAv/WCFvy1lZPkJzgUZmCKltOgZudWF0bjssocUzMO5YZEoQG/MPHiKaLN4lMBD
3VHaBFstqNoP6TjT3xq9uflc2jhxXzmx+s4SSL93Lyu14Td+73Xglt/OiHiR3XAvkNyAmzjBifKX
/1zfZuTMfCtSXunI2gXRHb/TjsI2p4sfsaeH0hbVpD53LxeB4IGoZt7kRm9HkHKN+UfFJUUkZOFc
0ss5ULd297X2FnekPivvLSk8tFvBkHM+MFO14ApzRSYERqDvYSpExtIoA9DipKjcZtXvDyXAJcZe
CdtwYm8zm3tLbaYxy50kT96nb4cwwHh5ux+kcAmZOIai9tuR/d69xzjt39lNy8Qruk8pENU5LK7u
OWRL16/bdNrQ43o7ybgxZtETFlVTKnYh4dIXocvhGxL/ptJg/fXDyPGDIDQAVk/YPlLey9hX2xFZ
7pfZvwukXHZ5mtsAR6SbPAyGiaA04UtK/bvL5VTretnsjYLPvKBkZpQ98TzMX93fWFBRpAmo7bdF
pWMmapq5OYiROI3vRCqOyXxOQToOCRda4+i5fq2Oz5yNA5ny7CdWNr0DTLqJQecXYHMEHC0jamMZ
BMN+3tTos0vrA43269H+LklR7B/TX95Wu9x2/v+KjOpNhRRP080f1OtRP44InEakzG5W2YP5Isju
FrZEY1BO0hnr+NC70HAX0RMfSVNDcLOlzSepyKumwiGSVEpExdL8FxgCdk3NmZfU5LAB/6lZtUhq
VVlw7b8Wv6uZukYk0FaZCAzxXelUWG7GKB8YOgn57kb615PxGfw8VD2v7VSg1mlPDkRI19vPm/J+
fm5q4t2gSB5YtOPm7dS780QcmKx4yUd20z3aCWPXoc9rKvkfacgJQi7Kp9XP38oSaFCxqoIuOnkZ
yUn5cbtBPA3c21Dw/2l2VQkOJp54xlmGJBkg07qgcSEt5Stjl8ZSipmzfO/b9RXDAokxhxoKF2xi
1Tt3uMf8TNFCuESWLrmsXT81Gu8rUaZYCJNZazx9fn+N6BoQdwQHz/DKgng40w0DhGh4PnZnRF60
UF4m/Z3YIBF2ahBTCz0rvfWi/atjtNWcz03L5mCROuQzQ+bArgghnnI8kYYKUz0Ril+5FxyPIscV
KSZjQwq/YcZ2QLvGxmo9rhVUKI6R8jR4MD5n+F9/G1PzQB77b3Z1j09aKrNjMhht/ZT2GjjCasDM
M7k2ETgTwmDwjPPjEydT0ZVGw42Ym8T7NxVzuazZhYn4ugqB5v9aN1/YSbcb/1d3wE63HHJo/2e7
arRZk07S9ZoATiWIv9HDqpOcy2jRoZh0zMSjLxU1M6oLjuaAs4PaSU+0VpOGdOTzz2lvHX6b4QUC
HByQNBPyQEzULiEFFVKhfNjUaJ7lMHuVIFhSHaSPaol4VO9EKTOlOvD6zTnggyLHlUYtblGg4SPA
M33mlzw92VZz9neoQSHM0xurHjXXwvgBD6bpy4Cp6pMl8bLTBxwH+5n6FhJVqraLXAKBHztHF/fW
RiA7iSQpk98S8RYsqztPd6RSc6C2ZGTOTpO7m6AzPp/UuQEDK/WAPnM4jed2j4Xi5MCVs7EF23Aj
jX+uHvnAonJHDjbgjDm3WjAQwUPfzQp6MsAeBG2pEiVcXoNiTuj2V/YZytGkg3wQLBkLjPkWIOS7
hxwlpiCbLtvPmL0ZlW6w953SJUXFZWCPQxS6n76y0FfawsSq2VrrZPKCM0bMa3f1gAOEGtDoC8dq
Vp0Si18S3JLrqHIhTACoduSmvYsjSRh1QIqaXE1wpl81ZSGPNOUcoDtVFSf/x8ZR837inOGYmGxD
M8o/Bz/3h31+jHG38V2PJ0sJJFZAgtCRXe+cjpbA0NgesSsZ45hwtsVxJO8JJ4xmzgaGlGfu37I+
0Sd5X7YM9WBIMwhSlyAwyWl/tUuwbg5L+SNlLIP9DBcGEWWHEsI30jca74hcYaiFgUpUzrSICirl
MfnGlmu/VtGUBj2oDPWkpObvTtnUCtmuY+qo9cL0pk/D0LzRQY4pCSsbqGxCsTREYaWxeTx0PNIB
cZif7TEb1sp7aK9cF3khGVveNLS7FvMiUNNznKhnTJlgAcMkEmK3TZCc4STAKbyjkey/d3FTYAKN
pbHqpwN/rWCOfnzZvQHoI+5fr+z7aQohBfhrWnKMnPuThlIi36B1p9/vc7+c1nBcaG+6m9pPoRJZ
WJzXW+xiO2X7IZLhA8aKRkQIki5j4DnrB5HBVQHRPToV8pNgYkM7X4HUl2UAfRXJAi++If1Cq2Pc
bPWhnlJb6teAEg+eutfkJYpZdLR8LslLpvIrjvJqggfhqFgBl4w/q5kNoODZY6aj6ufMEcrQhGl3
RpjWfMmQQzmRcp+XDsiUbJ6Mk7ekklYQOdFUJmg4o7/M88fcbjaPl3ifA0qNGYoWxwiLFJ1Sa5f9
KTgVP+sA8T+gWAh5AVRkhzYnyMS0mYAyV8kOfhmQlOp/bPSghhll7HspztWnuh06LBXIjpUu7/3O
XdlA7Ho9T5RvqqWiC+2nclYf/An2VKHsVpz7vmWhPHqOviLHaXyZdY9qz9oWnJ0iLijghjFCjbbd
9uOwgHOsui0OXI4DmtNRTOlO+GSMsqEEefUNImNwD5gsWlpP/QCHl3VUiA65B9VslS7OloBscM8f
SPz38DFc6orOhgvVAhYH6xAHYOrHkYitbmeYdHIsc0hvBpetJ4g86zbqi8OWW/GxHswS7eIY4MTU
GxcTTQurVSA0RW5WnrbOA6EFD6ZXH2kR4e4+xsFM5MPIHy4pHiypQ3QB8/uurqPr8NR3Qq1kFpfq
qOYdmynJR7r4tiOJoEWjPlrnILTlQatkEONSmnxJfIY/HB8mCC3EDCB80xXWGq8N/l1w3Utt/B8j
18WKjF6847J/lgSybfrgS31GBezJsA0ZeG4dKk1V4FKq8Cjey8RnVfO1tJj1yjCj4eMvzRrv+9+I
W5kCwhn87eBE910iBDFeGylqSdRxxdm71oAk99UYQvP58dsBce0VdW+CcXUd7xuB+ZlOx6ouhkhd
mjfstfr8OIaUknB3j1c77EeG3rPq0kq1nATR3V7hVhS9tAFuh4q6BUXlAzIxUdvgLg1IR5NPThwN
MxI2kxg5/3GyWGxGgLSxmZ7Ixqro/SV5L0hfTbIjFOdKnAfaYmaMJzeyEp4586BRSCPpSKQbjNV+
E4KUhkQX9mLAUb5JTdCmJSpjW38HeJFGKlLimOBKHRUPMt4heOyxUwwIBR8STF76ECOBAHwAjYWY
kaq0sQuU3ZkbcHY/V8RG8W3rQoaa/qikE8TI3FDs+IRWHGhRYQItKNy/TLqQevD4cLV2ClIzc+kx
hX7Ffrwo3WBYlIIMwBzU+se6XGPaS+RG6Bd599ZudKLk+k4eSt3Zk9d98eNJjQu/I+I3UzDoLey6
H+zxJH0Ym1Mn8JpPmzSdmox5UqI2iNKxvwA48nwBDfwsLxf9UvVpLFg7FVVTCgZqlkwYEv2fO7wk
Pjwx6zD7XGXv5q8v9HoQf29ogWKg97Ie5SNi9fPj5Rb9sOfnA/dfQyZWF48AEPmAWYiDMvFFfOBu
wGNHvU35VsETeAsF9N3VEA74ewpjH+wI08tH6MfVTETmKSJkJXTYw4II4vBSs2r/vWtqkBB9gXyc
BQ6DomVpdOKCW7732MExd/Wizyge6JmHIHSNCcBHmtji0v4BXq+dH9+vXaUzoxx3ZLAvkVy6rD3J
uvS9tUgu/ekDJlsLEBL3sY9Ai1ytjQ3IWccantltRpYBdu3BzrxoyDByALO3JbzLSwtADzmff1z7
KCTRaayVpA2PSrmvDOg63nXOz09jP5qnZJ0Myeis2x93b+JlsE8Vm9Y5CzR1Q/j/xr39r6uvofqY
1b8DKJAQvw2kObzfGb+buXzZSgt+MBAbsI8qIrwNa2W93l4k8yzcENVaSOrFRS1Xd30w5eVACqGW
fAgwa1+e2NOqKmsAQnxbGQgN3m3inosAG8DOUBGJ35qzATfje0d7nIw5JCy9Lojlq7ri0Wy0nsB1
dLqxoKDE8b5dLX2egNbEXKQvUP4MKdAhoyK9wFGpeJTIlMP0XoAyOBIoSlhyTb9BR2jsECXrGONX
gDsvXWmr1mSP5K7bRKQCw5GhKWCrPYp0GXzdizl4nQ9gU+GkG8K9AxO7gABH2DtsGUPrkCc9ZoWx
F/SFy67Pkm0CkxUZ5uey2kVZ2V5WdpS6suWOhiW1pa03G/+2dxGOaUj37GZBKRXIZ05TX9pB2a+C
vRIjym0pCm1ilti0qIfT6pxpT5u2ULf33n+AOtYL1CsAJ69C4zDODT4Q1EhDmht0pgca91Gvvcuf
CW36ltICZu2pwYxofAmmxrA6BJadPjINtdgawal0TfdNTJiEEBkWlygrbYCmhJUH1BDG3Vzlxly3
TNQcb0ttfcnALgKvEhiPtyQ8kJUQ7JaAmJaTj5dhXFKBn8KkRVa9PPURsoPpFftG8X9oiNr2Eq+K
gz/4P75Fc8AkP+dNqOzvxCPUSQL/6P2+sEXrJ+gocxzjedh8Ba0MaYKRXCIIqbJ+Tgn9BLKSpxZ2
3SGreabuiODzI84DnXmF0ZOr14umtc9Ild2ZedPujSZZNYp5bQwoeyEugJoKx35CD2tAUiLmFYHb
BUdvqrVpmZodQFJCvn1SKFYJ5Air7+OCXCjDa7L+b/T3XnK3jUsF8/EDiCSgVl45F6CcXBQUuBX6
8/FI4f32LendeOIUWWgUaUls2ozGsJN9CGjsecCnREtCXTeBAAf7KuoyrKRK9Ep0TrIqGqJ9QhMN
mRtLytzg1GwnMyzFQ1OvD84pvQCwuGzddri6X7M/l5VV8qBvon+Cmsznq9o+f5NKUMrfWUbSCHRL
VRkuJZlU/alIT9q9hvO3aAUhAwho6wJJ16+Wp0X2H9SI7Y7U3lCpnMWvggXhpzERNkqj+M09Dnck
v+UzjNgWyA5UNsb5KVWkimiVBRPZ7ohQMsfGr5LQUeHuZ9cWv8GEzFP2HN3s4sxmDdBspNnzGB9H
jK24aFJSXOyeEU92E8YNA1oVPgJXy6TgWS6zCSqi6AQRnjL8wM/XOrTWl6Ed9jgh1P98tz71vtxv
5LkIzqfRSu7bld6oSf8HXV43bAIYmW4U0knehioKBm3Y8wiFSiZnQ2HlmIifUk2F2jvyKLMcqUmh
Pm2qm/aCNQr1yqTRzhC/3c3lrrVhMxbzbj8VQRX6FXrsb0qPJMEFW2EHB6KzjdQLlthy8ttyG6Da
JAe/mmEHX6OAwLxWLg4nOejzo/T/ZMdBVSmJxFSn/Tf2zf4HLq3rHNVR6WpnmVxDIIMUXa+BACqQ
X/QwNp7USFOFgVjbKVuIU2TgJKvkH11s7wZMSoGtLHje007lq6jQX8OJBETPYW7wu2S1lHFqwYpY
EFcoKQf+37qOGLJTi95/y2cLHrccR0mCSbboIjrecsHWmIRr2bXlyZFsVWN8ltGKuMHDma2BEJtr
bLkfVBlrhdVaYwrm7D9eVPDc4XSH1m1JMQ2IBz+iv4KwTByJKRmncqefJioGRdv5SVrhJZk/qgGp
GhkHYeWRIoZVQkUjDMbLLlsRQXW+7ibyu5P2qCZl+r3vBeCPilpVk25aFpX+95jtB4LEkWJae5d/
CbHYkt3RsOjGQp28YLxq7t4ngx4uIB+vEt2LXsKewSaXE8Hp3r955DYFMFkIui9oRSlqvXq0zYJa
nBuHEZhJw25tDJBjbQj6bSfNgPxe4xKcYRiJ+fh6Vj50ud4dOZuDZeVUsaQJwsdrSROf291q4gIP
4z6/NIxb1lGal6GOiYeALotUN5r/jvE19HZUxXkazUZsOHcNwfZfTgTFWtjzdNXtfTW9JoMWvVBQ
mNr5IxIBFRh9OrlCVz1PPNPNfd8IvWYXGwAnTBXXoIC3FfXwCP+N3wrio0s3wv6fCxSAwE/MU0ng
eBRF1OJmAzcMS8hNAgm5IYh4KYcHnDtKbGv7c5pchUJLGIc6jVsNvCyVeNjogh1AlOZs1yIFWXFx
SQKO439XvxE1TyjG6GM7+dxxxJ9qtys4r57gWz11HHBr7HUOKlLdOFK8Vt5v/B3YqPN7JyrFa0pp
YpRJ1KWkMsz/tFQHNorn5JzYtUX2jPn8ElNVYrviKZB2VDao3tUdS9QKw2jGeY7bHoE8PiSFg9zU
ZFbhySXT7JJkgWgPblqVi/EHMs9nhRwIAp6hXCP8/ZN+U6KtvH4dn5i3EKzpw9wsfY+k65y5BGbc
MMYVhE4x/nintIOnY8Qo5tNaohgaKB/XaOm4nfn7qhRirGLorJbjCZ239p9IVml8RDvOqrLgz1CM
20JnSLvD/mU2eepsbZz8rfYxLd5PJJnzy6zerCVxkh8eLjwvfZo9nyKXoDJZ//rR0M5386zmHvup
gv1t5ed1sfC+Hd8DPvxlzvQPfqwRlWYWIk7JU6cr6LVFOdRsEEnRKiVcUngpqsuif+dSIP/Ps8Gy
/5VVMgA9vracPO02Hbus67O/EQL+pmPuN6Of/hD/iyrjGDIKgNDLf0p9P3V8YijAkSIExsWlInHo
QQbpmMPPv38kLBBfH6IFAMDD9B0cpGF4xXPgcfzeLD8CxHdjWr/RiEs+DVFfHsewXBpt8aAW+Gyt
wdxEcIh0uwMStjMYvua7BnIri/023sNZVAkMDMj3F4FUIfStl7lR4/oj1ye5j9eJ70mAk3aVhVDk
8/Qj5fpcIgZw4AqTmDny6Ex6XfhSyyvb9EE3HJgawpceQRmVna0fQhrfE19nvokHz2wbQQ5ZxTSB
adeeeb7pszSzJUlA7HL4eNVwNTJtTzEZbrDhbOGSUuuOzngQkEdBRoOAM9PAMM67mnVxU6AJrtw/
5Vi6D9F2kSBGlmhJdCqCQxm0uWN8rQ860KI6u9BlbtsAFfKKgnJqIGPoEH+7hM+t+BEhvvSffOea
dAoIeC0tz1mOt4xSPBUeJMdHDcGg1EY5TXGomRY0OE9k9HubYDxJhY6Vf7QCuS5LRh5tXbJaZ60A
WreZzO1ARF51x/bb/56fX3u41l/uc2rFppgn96dh9TLLsEZvXuMd2SpeY7SiStyBlx8ihLE6obpn
CFDD9oW/H7NDkNZ1Gmv6X6Zfw81/mCi4mlxa3Jv/gvRiYrwo/xKfqLTBSNEp63rE5I5/C3Ievmhp
lgueGqDHIJp5f0EHSVPy+rvSVRBJUsaLCrE3zrWF9d9V8AFcA3KkJz7suYJVzg1lj1caraA+FODT
5FnpPf6Bxm3NvijbAuPMF7gsz4v2tjhlyYVJHh0bXSnbDcZ9eq808XGBe2+CalV2XMOXL7yBiDgO
PHzDCYe53pZXkP+l/TN1AGvwArDrCdcGMt1GF/IGvM8CdO6sZxvJXblKsdGrVVMB0eDz6rYd8xwR
qeFUIxVcigRhhzRFXxab46Ll4ZxvoMInqM1iDcuAzD/u3BwEGVWtzlqAiOeuICVepsJwcCzsTcft
BRI1VKItiD/VVcqmG+8ZKt3mIBlTBPj/udF1bMUYihFWxxkOrbCOSxzNkw7UBJn/6BHz+7JUYRce
MF0SrjHDjU4X3ed4Yd4Eu2Rd+aBjzZRufpm9NI4cU8XMP6rRw8JEe/OFTz+AuGZbaAx+YrzSR7pZ
9j7OBiGyRZvSBxSdf25fgseplw8pCSPBV5Zc8l8VtaSD8z0+UHsrQYJo/RtHzVIQ7cf6lPgPWeGe
oAKgS6G4oTUnTUy0SieDOm81IMd3+5hCQuaa3uxxhQYMYhn3rJ8B4R6vftVYEx1vOkBhyLF4782m
GU/NAOBWiGeDTkm50wbxNEsMpOxSWYH0LFakGZlLOJ7ht8pghVr44n+VvgBk+SLMfvh+4vp5seHS
0ejUI3ORFCmCuiTlvLia3hWh9mwGNtu5VM1K3ZNkjS0yo41RgQpvvAJag4P/qStzylopYJkLDlRI
24hgZJW0WRZDv+Zsbh4Ym4Wc1s4zXOdign+nOI/KSiWLIOn3yYZKaXW0dqYHEJYUU8XLJ8ftY4fb
09MaAI91AqiWXB2X/9igT//wgxvSINTrbreX744mS+SocB3YJBPCRjbRIFDjT27rVPGFty1tcr3J
eLqQBKo2iBiK3/5ju7y6e8tDjE2DqxASv0KrcEWDBOcfPev7in9mtjud7FKopbFKvpRXNHv5HK6g
mFjZ/VMzpIslpEVbYva7dgxgouIVRZmFe4KZ8QY0F7qt9+1gnRFwteulwgRP7EpzsYDcrFwe3oXK
2rV2H7CyeQoCVf9O3AlPFWY9qZtH8bFC7BpHiiCRYUHrO92t1znPXM4wwuxmjM39bd3TRTNNUpeC
qGvEQ6MHu//Y2RvK5LZATiZ8vqwtnd99RouW5QSN2pBVRlqTgPNib/QVokaMCNHdn8vm4fzTS/Pl
o+fduvLB+CYI6K+nf8LiwYOgYCUWaBjHX4kE3B8RxaJ0ZKuu1MViTo9NDCAEfLEoUHalL+WqfytP
u/rNddVDdFPbgGDQD347OKv18+a/WamUexalZHfgDkcihRKdCkeRyraS/QGhCiGziMgd0EDEwaSJ
vkpnCt8Ica33GXAkO32aFqKqWESyIM1BHgBLIZc51uKDCCelNnncvoQXZtz7umRUiLt8GJ9plCPa
w56N8PG4Bv2n6NtNpSTKU3y2d8oGzwjIbVhOgCX5l5dv0mKueijbCR6+AcbVHR6LB8zwYytIPUlm
3frjcOxlmEAw0uSpiDwySCYDnC66hqKyqBLimF1biLKZRXiRIYd+A70kFlXhcgVCyaxDxAjFKt2v
Np7W0OUv1CeBAr8PQHXm3uiph/YgrFIDp4j82V8pHrazwZihsKTaeaz5jsfr77PrcQb3K/iZ43mJ
fI8WxDC6Sc04pW7K9SUgk0aiQqXBa/PrNOrDzviUYa7w528d5aZSaMMYNgxfUtE3ChUVLGgntvQs
tMB2/InpkLOkvlbwiPAWMmMqzNvvdFSHfshmakTRrJtCrMI4mDNYlTOJKcYyS2SGtKMzgJxKfWmt
H4uj7jr8piPAmxqYzBaF6vwmHXYnYDvNr7M25Lpg9iDpUBYTOJM2OgvFqd0ebPDP5Qi0TN2OJ80m
LO8LHy1Csjl4+N+f7J/mKEwvKex9TzGOvzHIX8bfgjlMYc/Y5iAiQid7C/s8TQPUHxrPYeDyHVyB
9A3ekEH8YqFaiQfw4EltB8AeFMb7vAt4QFADWJpQ+iQmxL/QVp2Nkcy/vOfkWAJFJdeoptAVdJkv
384GZt71JDKXR1TGEc4wrDt1Ut7KrXS5odx8QvPJFHwyg6k1cxAMqv6003ZUWEw7v/vHidxJra7a
sVZCAlvaiKvmawteHK9p/wzlxD+blq504G2z5TGjgKDRwF/UhQLk/XcQPLe+qiB1XY8l3OOnbwkP
iugO2Yc4kzrmwf4k7S8A700LqD2VQEaEhZfm5PoENG+NsRDvqErMMyXngMTIDIchNGev7d2jUhtj
BD3ICXJLITqSqgnzaoV51gN4g0WzvXl53MrfkpmVvnngTQqfnDgc//G4wL3XZxH948s8P6wPcaQX
Fb6MrS7C7zEVAa5IRjiPUmWlslYbs4xknrjnBBIOXbWa1syf2c8VNRbBQ5o+YNQMPrr/a3P57qf2
DBXSiF7r8Tw3by0MbJBImOm66GUhfKqRV9kPHv/dmYhLao6PUF4+yRxUE5rD2irkN0dRVcFVGFca
hT98j042XnfYY5muqDj+SJFQ8La9RntV++RtK2ghyCagPRo/Ou1mUqe6NTgxOGtun79njAJS0mxV
36J19WIog0kjfKP5+NmrGQyvkTHSS4i4HoBugfW2vivsvYpHjM8fXU+P2T4oGL6cO12oW4ET3Yhw
nvoPrN3UGo71hafWGoz9yyl3UVAeGEdDyMBKkcrWHGVOyb0rLsshO+HD314fUGoowAbE1j1fjGs5
e55B9Km2coZb9Imiu3i+3gjUoDnflfvixYveIRo2SxSMtVJKhB3dMj8oDOUtTUzCFSbyaS2ucf4n
272nrGG0zaRb7Fq9TCWh09lX0OWRQVMjZjqW0LJSicf2eE7gSRB/L9bCvqwbKUGjKsQUyTsv5mT8
GsGDoz2lpgm3iWch0PM7ekfVnwtQrrPjVQK+0XR/HsAJqkxQfMYSbdBAQw5Ja+i3DM08J9iV2zjV
kl82iSs1ja1mxDgd6+t4Ek6Ihzqm2tbajtCYKiTCgG2Xkp5SIKYN9Sl2N1NLV8SDs7VclmM8cqqZ
g2YXNtsTV4Uq0fl6+WKqjUwCqkYIdg0k0kbQUalmtzcyUQ0RNGSW4+tpEWXeC4soJECmo+/PEPre
Ue1gg1QWL+1+elD/UEJQeEtV1hfz1V5gYHl3jsef6ejqjRnSPZXvVB5wMlYwP82uCH5pBkFokt5j
VdDRl72UklFflk0D/tO9j0n0rorLvNnc+ySML8CDaw51NqPF4EqPiyflU3kO/envNsNoqdwT1ui4
yOq395qR1AVdjjLQtqwnhzqhX6UiKHtu9dGC+rwXOhuHzhy5qat1BAFI5VbSnbUIzAjTNtqsMzzh
8e5Q0fkmOHx00CExBPT3s/aDQ2CuX/zJ8aBZlafxZ56SstOqQ0vjaUTT/t4m6C7/4+DZyCvxtMw6
5KrAcs+68hYj5gLk23c/MRSeBldvl6v3iCKEQ7sPlqjYfZmCj8XdnYIorx5V/NL/XiMxdR2d89g1
L1uSkX5XhdJXavVHHbL6WN10BWwei33MQNjykToJRYv6gYgjH0Jnk54HWQUPz6J7IdwBKVg5Nlyo
CgTO2E84rj8dTh/tL2hzv4Ey9OJuTW/RkRJiCaXnHrGinWfgHEuH/c4wNIVIZ6Ts+6Yth8Qaj6ga
GMOxnvvk7rMV6+vRoVj9/Gpu+qTazrLaDg+JPTDuB19oiW/33OzO83a0Bgv3MacH/qX5PK2OPNA+
SxEZ0ULSTz+Pk/VCzzwAkGNQOknVZ8uWKnamRIbUUSf+n7mU1O28QHNAw7SuKi0ZqT4LCN2TINWD
6W7kqnDiY5kqeJsidoIA2Z9Wr+8UUwoI4XhDCyKsUmfqIa7WqiT1Nsgo9sWpTZdST9GAnMuh7Rym
VEdtPFkUogXCYVxw8jjITm9oLc/AX5RNP7hHmollG4KuBjuuPjDMLU1/lbz/qHIEuGjHF7MeUPx4
NKDpECRltXaM5G9oabHFCZfSs6CkNht6g4Xb3uUZBXuoF6dyI/0Pw5qjTRZIf5ZGqzN7E1RpcMaf
orVQGCO/JTs4fQZBIbiFy0mTT0dGnB/Xr+MTGysYgQ2GksIyiyPMXX2aEaBKcGvxE6pwVtD21k3Z
udB1KCZziHUjnZYAK9riSEaifCwGjXLsBNhFlg19TYX1K9NcgEYgURFbVnPGNrCSmISH3I3QoQ8h
5KpITUd4Cl2N+sfkc4w8CVIcSOo1H4Wk+rDP2hvDXPtdmhk8UO3agiIs9ESUBc7t0i4wLBoyhr8Z
RvSSivF0EFfzybs227urNTwl/yMux+cz9nC1XiXm1ls0kPwlt9QK0IrD9b4q03slYqKAxCQtXN75
Sq//UTXGWsUkr2CJL2QlKqDyyHaid0zZif6RLRjFghKmwyHRBPGZKvS28npX1YFAABC3orT4Rkc2
NbOFb0KGEaabZXhKqjwRmD6aF+QqiNs6oe6aZ+SIZd2EVO4xrozuFs2bpgEoz2Ak9O6jZ7IhscZl
bBDmhzJ8YsbWYwjs4Bcj60THirKpoIfiXfNBLqoQ8zzXD1+wA/LHK4CV+fg5M3lpSu0gyYvj0l5V
npSHQrs/CQUeR2822ZYXUq4O9DzahbTPkszMODlK3avzMmpU9EK4PTBFYeGL1geRyLTQ6snwZe7U
LgUULx0lMWeDf1qInW+GS8dWYfKVMBq8O5TlPaZwDKk8GT9c3EM+CWYm6kZWSGRJ9L0ObZIAq4gJ
7GbqUt903/LVVLEFOEkdJg7AnLwO2itwpOdDfUVQlZqEXpbwYz1NJtxx7LsxgUwEIy9GYaH1XT0U
R0/7lS7FhXQuPiApiMV20EJXIm0joIXThSid9+SXXnIydyTKQ1zQoPehG90Od/qnZg9SC+rqc6+C
VYOJLwd47zgczIEnxtWLj2vST/pK1LHe6TmW4RLp3pCkwaSkmdN26Xbe/N1tcbv5ULQmU4nPjy2F
UJiu+QPq6THbMkqS3LAZMek63Xlk1K3R9LH2kKkrxR+7iOBaum9ZpHMoO9YyOLPebQF8RWjqV0LK
MtYx/KfuLBrB7ml3wWMFvqr3SMYaiSGwKeNdVX2VDvgoi+9ngzQV+RTB05IwCR0mGNjd1nQsnuT6
iGyWxOgp2QHlRfNAXQ7zM5G1Wf545VbEzPI1nYH4B7VNPxof/tyhoqgqG9yrXV9IOtw8q4T4pY4y
01zn76/bsS0krgHh+W4ogOzI0/DrCKZBEGAR684VTvYo5D5BnFMDQmERTaTV2EO13hA6eSaEoPVn
48KKBheWjw0imsxwzakpz7X2lZbzF9iTNShvUPNEQJiPfQ28Z1gHGRydaws0PrTZkBM02MQhQdSk
y0D+DF2SulWQkQ/+D0rdsIqcRCqFdy52pLcBYKYszu/kFobc6+QLTZwk+FvFpqFnP0AAnYH7wUww
Occ7MhFsugDRc3F/X/8qJBhrByfYj/UcOr2nnPFTyfrDwPQvB+6rvbpywYLXs7BT491vYgBsiYfJ
l/eilAvq2+nB+t1Fgg2oRxf46E0T/4z5sfM+576/9+Fw8mRTtVR0pHs6jkaQs6JLE5XGm4h81CMp
dzi38aGADOss2VQziIX3B91K9B55hllhVHn/ySaVeq/VUehl/yIgWgIAHrm10Mqkkw8N4MrAgNoP
Yr8m0XvrWMO8HfW2EhuJUi4Nrbfhqca/oMdaIVDyNsv18lC19L7fwiq6OlPYOoVHpwp8GKtIRbB5
srWPD7hJfYpvi9FQ/wwzjzbt/ONJsN+9FCO5J1/KXl/CyTN1LEq8t1VMx50SQV+z41VOgnrb0swi
yTn4Dea03yaf3u8a320/93lIzfvbkuQDCs02BOF1bpyOozSicZLHE/79dJQHx6xnl7JDmuILanEI
FOUfxC1WpuDKlLXc5+/s65eIy0wMwQtInDoQYsWVCGI32Fmwd3MT7+z0EKqkRYyGocupZ4E2sp4N
PT5qpXhkdAFMoX4eDTI6DVN2x9kd5bJ4+Md5HuNVT+kWFWgVpNYlZixZRZ4o9kaCKMMbEK1ZH7+d
fLKX60HxhmlocEXgqlE9jLvV2jWCiu9vpURLPsz6h1B1I7LONHN5qX8zv+gUR8QC7OEtCRiP8bSd
O/sdNG0om5aeEkTTaJclgT0tqB9SEbJ3CdqAUwNvlkIwKIGgdoM8UamtI+EeWIEtj10H7pvdf04o
nR9+kfpVjN1tmHkSIAhsSITpRcXPBoNenjXNEYHCHgl+0aTnL0aqG9959jtxtg5N4JY2L1FwYN4u
NPKWslaxJMRHCIZSelSFLgmhlfLujqMBMqo2diIeAefyYAwRl2M8S35Y9aORP/oHISVreyzkYslE
LZFGCq7vp4XIbcrI+Rh9aktRVsMy9Z6fFTitSsFzo0DRFEx77nqFoNjVArafEcr1/+Ogy2ZqQLfo
zRQAIb3YtSbfw/6PAULL80knnRBQposCvPPU9iPAwcLO2uvBuMmB28izv/lRh2ZyFh7nc2aV5J3W
A5c9rRUvV2JLMJO1rLMuq2X/wfCXY2Yi9zq4KB2NRszGrMzstSgTTGf+q6U6h5btpFCMsSFEROqM
EJHJyOmbdtrIOTOKhiDhKYCsUP63z7lsMsHjpmgBW/3njq05D8bDdbznptXcyVN8h6Ax2EWA8siu
ZbZolRn9SL2kYwtOzXJUna3L+oR8Ei+5UAepKaBNllEQtnoF5ca1D18NAxTiUnA2ZL147R3I4mo5
wfFVmwRtku+J3RKG3m6F7ka/vcmOsURyM2Tg7yAlrmwB9xgFJat4kJ/v33M57wMKVrLZLp7nkPdV
MTCTlH+r1ay5U3bWP/f8nmVvOkIf97WS6hGir/htv0ootnDQ67+JwoAsHeouiOT82OloJjPrXnCa
dqTNpn9ejpTupKEG3z12zy3bE1SpKaP7GkPFuUQPkTpZcX/QCtFbl86UDAuyUAsFAQbVgojVjStN
wq84o4VlSe9tmdleHF2jcFutdyTvIGBvVR1mQ1pHPrw7lVboJtdMGojRX46bkyU00U+Huu4aJJho
gtmgjmBakBhoY7UNS5sbctSF/louDIrduUShOCyoZklkCHznwT1C3s/KPbklDogQ2ipdZKprlb75
rMptptcXL3iHn8Os+uHwbh21wbRmZKfyV1ZO3FdGCqfmxpnyWrvdNoExVCIpu1SsAFY9ipd6l7ZD
3LTBzhVePQ1UVhNeCOF+LhUyJXOLDhi4dh/ZzkjaK/Izi0z9B0VF14ifTiaPpFH4XiXe1M0ZACiB
noaLhgnPBTepmIcIc/nQHqXSXkhv9Wz0oaO7K4BEBjQH3Xs74KQ48Wc1D16JoKRhNn7j3F5LBulh
yVcilqXqRHmE/U4vkquKaVrmNBLCLlJkP4lLjepjA67Wh9qEcSfPGZEY89tqSquggGA3t47ANsyM
rDibvh0vYPH8wapLXBRKApP9kleHDGoL26I67QSfjEIM2D/U/94D21t46bzxbRCGEVoixy8CT2WD
0ZiZwp/ptlViMgxRXU1cI/YAQzvPkRoq4gJiCoNjSC/RFb/zkkqnOPFF6kGSyC8PFZ5EJLfF4CvP
QyKmKO2fkFshQzylvSZ9Y1rEqGjyvjmpyQI5iAVzi59BkOTNdvnElGq7TOD039ooyudz+rhdy6PU
AVwdIHz4R+p8iYZnggZpLW6CnvDzx7WgJY8RX8173cDwD/6KDtVRlnxZoS239y9EIcNIzI2+zXhj
f8f/e1FhME1NhB31eDfd0WfplzXX2Hh0PVv21xTeV49CaxnKzLL3wKj3CSJLjGN7TpdEkafcyTN+
BXqecyxdmWoNivn+VXTP5/+LQfoiSjwWChNlaTAKgKLItr1zcjbn45/hI+1XCT5mfMicxgMtiQdR
IH4Xo3oITq7q0/bx3sOiNkxiK/oiYbjZpMHAKELE9xvo8PixLsSR7UD5HCyrL3l7FUK6KjonRYZJ
W46fKXlzSPnjU2R4awL+/4m7kMtWZAx4a/FCL5EDm5yIEEdpsprMF42mLrWaU4J8pA20hGuUqdUx
9qfhhMsvqRAgdRoHTXNcljKN3FAyYbwXiVC91MyG/iNU4BHI1oc5KpWW2wQNnEMJrdajqhBYvb1a
ke+drItWKXYj7+6xUzkMK1f8biy9viWrvtSAUtB2CfyRwNZsbWzu3+wsTduw3nqw9olHngMfHIQM
fV1VESt1qNHb+1IxgUvrnk2MseE9BTzg/FPLWxmgqjGjkB7QCPtEeZJD4YTzHAL/N0U6CcwjHK2e
Kwkb7pB7UrfVeyjPzGY/1Uqg3gq1Tqk7K76bstEY32GOHanoMw5e5mPkXWtwc+XSNWepLkvlxRUf
9P44l6SQRmBC4M8gCKuRVJqr4HNv5OYyhTW0jUfGQxf6EhHuthTYBx9zXCCDruliYW6BXoJUdOC9
hPNIeFdyrLkJ6hzjlDypHohjqp9ckY+m3EwBD331SQlSzQN1Uh3Vs/0+SF36zeVBTk/rFYRkKYsm
BTAHeRwiQ2RMohMplumvBBON2OFUyipXMbKtY0oj+tVc9FAiWxepB0t8FwsBlfe6f6+1VIbWESrT
dmgVfIKwMy03YFsBGgKxeYUVllTuEqOY9vskzS3mwVDw80iQy43MMQQF5XRTjC00GpQa7CX8ys4R
a6eTyhbpPUK8R+xB6cn0o5hQZTsT+WH2nOWmQ+wYcYi4QBJBN+ZC9fs9PVIoi8/ZljhfzUQ6tyZB
akxqC23AkWE4bvV+VbAbZSTO4GfC+kv8TZe3iVrqeRKDuY4yV40zaKukrQp9z0QSpU02YMhgDNWi
5p4jMFo9lLQpGTQYyS6ZTnz6klBD+pggsyX+tUnQ/l+5g5nQMK3BT77KOgH32H30TKtKDW5i2Sxb
HDiWZjB3aQDhMIksXoAPGWF2d2XUJarAiqgqDc6+6M7aAScId49eaONQ5pI/q52TcyqM16lyov6p
NsiHAakwPE/4W2oCNuBaTu52ht9e2LulPasMvXTVjIUxV1/syxJT0nHYwCbGBmgW5X1KeU0iHQxn
I17fJYGJafh8nmGgL7J3L6wEDNShiEiBPIHInI1E90ZPkXtMni0Nipm+9540+BwnRXXO5ruilYyB
MGS10PLX83RUYBZ7WRjgE2Z9yJNTm6cQKTkLOLG9TR7vcgodO/UY3i/3ZwE6OOPdXrNd2H3hCJtN
xMcuhxS+VF1WyN+V0/6msjjRgldUHWphEJDX3QFMkXfCTpa8QSMwS7oYFFzfEN20yEUIyVxrqKcr
07nMMx4rx5PchXBUexy0CEgKvRfNClutt1y79/7AyWG2+mSdYEL4teouZ7znNBQoScZSLLtDC+Wc
E+iRzMMJuEWOmkAAgLi3KHC15LOsmFvFzcvfWPiytS0QG5WryKu0/Sd7aQczohRaF1IgaUVDYY1O
00UnVRRza2C2hw1WaXQE4hN0E4jUkH/FCagptodvv58tufRsk4x9wz3K+pJENcv6DjZSq2Ihpjdl
yhKHq1JgcqoCajmXUgKUzUytes9iaL3C7vyWZdTmFSnl+LmArHvgVOiJ/4Sue2ZaJEyHjWaCj/DX
h/bNFPrguCFZe9izVEfABaW2YiFIInBmGcIyMGzQ01xnyUuRwtuezDkhj+oohxMX5fIc8TjSX07G
dXsY6Rh/foJvjlqGMl9Qg4RjOeIFAi4nknkWChKjsDUilB0XanqsO3O/RQTsX/uuyBOChUTm4ucz
lJsRtF7yCT7RsrvkXab+mHTKuE7NTGUYtfH+ARjPEpxaAtadYAYnecMviW5Jz4mCUs8X8xzs4syK
Ru6AUcA9ZWjhIqC/oHleeqHxKTb+3pG6SkNRpwW5N+QWvoGGT2vLsnJA3SXlmbORmXrrn0/ncep+
x+qoIab1gKcfOWuHP6OtAWU+rKLS2MlDCb0Nz54iqQwCm0e28uwELxziuI0wsqQZkaI8CqyKyg1I
g1515GU3G4We2r5Nh5QRwkWvG8a2xzV9BbEfuGC7bo+W5PA9Be13irP7jNmm1b9D0HO2727+DLe/
XqBXege3NVkp5GGn6WlHoIvY3alSqsyxJ1WMKP6F+cuQHtwxTMI8OH48l8MyQ4EJR/Vv+Ixlqxf/
0/haGfezPvERHyfuKbwixH1CLU0SiPxIDIRuHPXGFrVFtJ6ndrykdxdbN2rYVNsE0LhEEj2dVcgP
gypn7rQYCakDrJcnlJfDndITW4uiroCB+Jg7B8e/rmD22Jjkh8U3BNCKUw3V3I/dOv6VhSEascqK
rgUDanch8lIPZJJCgZEBXBhF69kmFiiqqmTJUk+KwHzCuMmWHciVZ0rFl+//of5m5lWacRBLMpGc
tlkLT6eumA5531GFAdXNK/R96jA4Q+h90N+s+IvPTMg2Kct0Jo8Z4ERHivz1Cur7CoOTlK9kStzo
4Ou/d697A85X/CkkA1yNSwV1jF2C/LecFGWHFS/8uSTUPb/lqPqUKfJCu13SfUj13ocJlNLR9jHw
Lhz5Bn3QhggcapNTwro3Qi56skH1qM88EwIyvg/HpqN3xwkRVqpMRJxX/jlFph6Pza9DHf159446
q5sVZT/4Cv0/OyWFvxB8wEvq6RLKul+XrcmUkAzTv7OFAU12/yoIr30MwYYhVcl3/lhZcdmraXzj
djFcieCLS7UIOaOj51WNV9QyQjuyZvBlcYk/UV6Ca9ht4ES4a7u293bGw4PsMBnCm6K0nyZi+NJ4
pbkZzIMhcmNWU+sPVaMAcGaBv1FyoOwyuq9fDPqCASQZTv6dNYvXL0KYuszWszsVf3twRYBC5aDs
YmRn0DEhK5zV6PLQAGMWhZmKMlI3LnuB6dQRssiTSq4gTSum6/0zAczhxW/U9lZ6bDFShw+ISDeo
umQB3RfDPFXer4NeA78bld5kyB0r/s0+4MciqSlO5EOzflZPcslDmKHWJI1x6L/ltUrBghvrXJi7
ZzZjm8yefidgZhbcXrjN80OecQ2aRJyzxC+s14y7o8ivrv60OoK+mhE2FoWDkwB2pBA7C948wxnz
U9mbWEnSM6qL7xmUqBbOB1eHDXmenA0jS/kE9mGP+clJVeOmuCH1vsYj/z2i7J/I9qnyZhJgBSBT
teE4dCisvE2KdHbuoaLyQsY3fwtyLBQ7jBZa/wPiF0Qr7wOjr6AqgrAp3i7IaMh2tfK+DcJYeyTb
owunluuKku0WlHG++0sA96dPCHMrI2Hoz7b29hipWzQJDWez24sG61K5MdaeMF2iphrCe97Iax1f
6/4X3wGy9i+9V8X97KsYHfcU74gj8ucIUpE0PZllJbd4sHbAAYAW5t9RQVBFwJZYu/zJHeKXeISY
Q5dqSyH2QLEgR5zyqy/ojXqq1VB0kpPfuhJUT7TjszcPYyJJxSyALv6x7ngr+CAyemIuIR1ZDwIt
MxC12DthgxAt+XDnADDFUR26uQqCuMt6P5D1ul0OHcqV72fj+efYNtk+Krr2W9tVDjqoTqOnhFBv
UUk+LwqksLfA3pYKuyaVwJbygH2pdCyUKHYL75JOb7UvBDWgAu/lxFD7mnsaD+fieb77JQNfDhCd
tfdvkxveTGMYAvCpa56VDrLARYaBhjLG1noNpauJwSUbjDn0hva43HK/RtKenDQlHQCRTQAjFDX2
opHEJ1czP3NBs4E5xdFvrlVml460YDcfybwLKBJK/+usO4DUUGLLj9IX/4mACRdf0NyzWUaZA2li
nL/OmhdtC/VMXeGRDb3DHnbRsW94Owq5wuWs1ASSASUl9Q81eSMHqoFGWuVlgybDXNdYiEJZm+hs
N5bl9katRZ06pWZaQ/6Z+2AQFBRAZ4G+jD1EowOC5WvsPfdpc8vBiqpc8GtEH1gLOUXmAhtmUXyM
6CxHXWprZKiuLw0elsoKlXahuUobW3U4aooR20tEngVwZcntQlCpQxftUNtVNmAVWXgyXkLylX5J
mfcFEDxbyvo6kWxIFGrTo83PbnKc583rQVlOKzM5BiswF5nhPZIRAI/zWyFuJEFreiH4G53sPp19
+n0k5fbIuCOP8BogW0oqwGKrGwh0wGjerFxAISdHPppw73Da+NKdFVNmtFBU6+CrXqKAUU6AAol2
Aqq+UpHK5bZDQHA7Gy4r+ESzBHUNBBSCygpsYQnC6PqMc1IUYEFknmNqvgZwirVyaRh6GEWXNI1H
QYlBw7nLflAJ+p19KtK+8WICWfIIkqDpCK73X9T7SK3kS914lRA7NxSMTgIFYfrmR3aw4FU3pLoF
tuDCpIXvtF6AOT64zg9ELWgk0AILBosV88SIBzAopqxBmHhmoQzoCGDQnQQyW2Kz5vUGWF8znaJc
1moJwZUJrlhe2r5AfvZX/EIuFKFHojk5WZmTRigg75+iHCBAwqtdNLrG1LtrejhWM8gOiKhrTRrY
0nNJZcCKsw+0M83mJAlrAHvxEYKWU46gimZwFV+s+ZdUP7kWSuujnXpTmfnGFFN6PW3WHBRM1KMm
EZEPGWE32KoTdLkdA7lsAZ8yHbnReZcKbSR63XJdeRGYRqIIQRIvRsOqmYAiBH4hX8FqCFbpj3Jb
HdgzBn6mRifg9rs9jIiFXv6V7ezxwhoVz2Leaz+LPQjAzrQG0dN/5oUKiRFTC3VrgsjgTou/38CZ
HDj3Vt40rmL58Z64xQSXeUMrOFwJvo4cQq6PtE/Kl6Wr1ezo+6LMRgy1VjnEwfqNDO3m8r/0cWaG
/t5h4njroB6b3AFOjUIH5bq1crtVAIlW3weVRv3E6A4608zalHJDb46jEV3qFa0bEA/C3CoEJ3xj
0pWNTRiBwdMTdss7jWmdafDubfjrJlbejvw/WmTGYyW3vLzhR6gQ6qL/FMGzExt1cIZZ4LClIYLq
UlvIuynQj4CKt4/7S+pfHim/gS90fgTJEDHDMkGdwN+8+Iymf3SzZXafIuqbRpVp8HvBP023nPId
M1q0irAckkuOJbyflb3lk74RGw5oJncdlSCO/goc9Z6HByOLGHU475tEjDiM3FWyLo5QdwEZELzw
EOjzlgnMdit8SA+cbw+7lV4NjQWxaM87PQ/rMZIcWCM3aXlSDWHjpVLDaPnGUlmKX/WyXfr7ftgP
zOzpfhiK4Z/TMVheNvAh7MloalJlONWiURJkaT22gSYYnK1UZh2MCrB/1hxWVMpTMBV2bJ38os66
umblKOzU5RkaDbAsYhmTG+ovPIl5jSu+0MswUrj297mvXyAWTN3KTON5a94OE3YhDejbis9NGXRU
GQIu5g9FjkKaeqPQ8yUx/PUTMDErIxTR+l1idofJgq0GbXd2yed8IFTu/O5DTOqvUmtJhBz3VxaU
Yc9ov3V6nOvbrusw96MI77Xhxhzr1PpNDCjvOrwV8I5XkrW/r2mo+/eiQHSelqhgVOJTXzyOp+05
pku0cdorf9f8ixspJVInJhSGVZ9vGMIZgalR6fpssHR3O67pkFcHlHsM2ymoRpP0lxNNnh99vtkU
wsqHwpPi/HZlF3LKHW+Rl++C40RNY2nNOk0CWCdtVt7ifNaCbZp0EvyQwhZvGPTDpOh+wAWdcDwu
JlAwvLYb/U78asQn0eYxxH5KnXeVnX8eixWxnTgftYy14misY83Ixk7Yg5jTtiv+igSpclflf897
Ekgte4PUIxj2ZO8UYsYMv17MC9BpuGqdikLEAbRIjAK3LY414SPOF3ltudKObsyTjVNCT3g8GYCs
0f3JRDKsIkvyiMiwEC3XIO8MhQLYwQ2RawxkqmJIXl1LLppYgJ9Hcq+oZGab4qQZy56ToE8b2Pg9
4RAJIUM/Z4eHFkGXebEyxF4DDGC/ypSpQgNX9W/mgeX3AD30aG3HFSyW83EKLc0eqmL8vu8zXfnU
ikGRZpefEORnizMOH0omWBpQ+tkAey0GCZNWT1XS5R8Cw3qHBNbMz/dXaERyS+OXjmOo49yuvgTt
4UOjmQ9yO7NtSepeNJi46nBgCx2vAg5C0E2jFABem6UpX9ho+rIAN6sgiDV7PP0cixFCW+Xsjptm
haKVaLTgcfPz+LNtAFAvb8knZdOQbcucFDxGDoDZaPu0o8wVk2w0PKP2G73jsar1Hpr+wb+HVtb7
qc3nQFsA+u1LBVTjHng7UpPnPdesqoXJuE32Px9VoF1q6XX1X/J9qF5A0uVZ74+8KPYgExgjS0oM
T1+c8reb9u8F4x0EQ83HBfP2ZJGLjYjqjriZXlkdy3NI3uDpByBB13LyOYP/PA4ZikKl1/py6euF
Yi0MeiyaFMthPF83Rg137YmPDXMnXsCWGZAHW76PRKqyvBQkYFaMbsCNV0VZpy6SE8nSvN3P1XLX
ByqpDbVpm5YXQ4YGjK+eAJPcbDwtA67U8kSlESXZrjh710QzWQOWDH1C2Ay7qVFCXQEqcL7fD6N5
zYj2uygzsP6PpIsQeN3ubtuvPDvBk4BpsiscdNz98fpL4/qLy1pvElD+9vumBKI7Olwgxti4lFIt
WGHGLDjZq2r6ZnN9SU7YcLBKeieebhN86hs31PgyrAt4wmZMp/w/CYIcvf458NWahHCIkuy4q9ZN
YTsah/GMv/GzW2jA8rI9GDoua/SSdvZNwTBtHTJAac01ZQw8uMk+P9bnTBYpnMzulVALqlOMsEU0
3Kbvf/0XazMWzize/XACwnT5PdaMH4s2AZH3f5Q4QX2D5x37MU/d1z9ht589HS8l77OnwPpwycQe
Ibpc4r1wQoLzVwB/deHd6GHZEVzZAyje6qpuEiI5IWJLOYou2ArhpY/vCa8a5Ww01ayESvULuHV8
M/EZxK9mPt4nKqAtkSzYQzkYteBB161IV8U3PWyY8cl/jHLh2sfBnYCEZU6m7alH5rSwjkqAmRFc
WgLa3log+Sd0RlRndDBuy296eLDMnQ0MDps/zlRu5fJ24RB9et84QsKPsw+bCFrxOq1J6xejfnM8
PbOuSyvPNfTKE2AyrAPcybYyiVLVpOS2LPFkM3HSlmFa4C7RpEMPBF+qjCjMljKviqjfEQ4d8DpZ
YtsOC/eXnxQM4KDfPhJGH7Te+FLUDJixXhMv9SbvQcru2Kqb5hISzUp+NGKZcan/2Tu6zgpYX+am
lhxgtnEYym2FdbPNV4NUUuqfls6Z+hbFwr/sBSclM8DANddxUCJI4shbcejV1DPvBY17n6+YomxY
9mborOxYBlJ5W6s5ILpOp+AFskFgavPgNTgzUPwSOJmjqa5wIA1fBk+u7gQS19grTwI5j2rGu8jJ
7QFjbdFtMa+CWOamPXPDE4j9gWyyhQRjgQ7C3eeZB4Ie82MGrGybUKbYSSKDCeqV4lcaPZnbzpKO
91rmQoqjBaUokvW+QhgwQK2a+7hPS9pcv3G3Wx4VHHezBHVT10iQf80NhPe/Ou8kHM2gXj7DrX3N
cLv8FpcIArRUps1I+MFOxkQdEMk9srYzROtikpMgUq8nn+YvmdHME9Rb93OShwlMuoZuihJyvR5O
TBF3Ta4jpGPHd1RNX12tp3Y9pUMuGLKj4ODyvzXh0KCaaH6A5khrHEQAx0UO+UAR7jfvOvK5uvtk
Y74R1FkQqHKu072wznolz9xynIFSgbZxbUrNDIUjh36xxVoyIPEQL0In1Sw0gbQwhpBNNwt3sLvD
mbKB9UZoGaDx16COaHxm+f2DWPS9ndabJPBRKINv7/Fl4O66pbHPAmLM/Aorbl5a2u+EYq4co5eo
H+r/NOk+mjDTbz7ESiDAnhLanEnniQhkpLp4av0Gzdw8OoMi9bLpg9ibVMDAT56cx0i6MTEQlniZ
WgLPqN03NSscmj9w7qo3U1uY51xl+JhjkYZ2H/dh6ZQtr8A5eRA8y3u/LOo5gXy/kK9/u1ogWkTP
GgEZaVw1wDGadW9MkOfwgYrYs0T+LiNktIwEnoL/We5bxWEnm8u7WpMEVD5x8I6S9FnQKFCqYSWh
stXrY0g4kAuoag+ybQFkZP9LJZj7B59LVN5Qk4uYKSPednAdePDjkLVGIgrk3vSFsg8aNfeDiNDI
laEjftWC7I3I0UMJmVjBBj8fski1AG2hy1zDtglsCpVmdJ03lTTUrBUyXeIDdyI7b6a+KNpIhP7/
GhDX6rbg3NFV4f4h4qXbWCOFsrI866r9PXDNaKaticTvcrY1Tarc9J4hoapxuY0O2n8fVW3Kn044
A14c8lNkK63jfXRW/fsb3RaQD8DbUCVjhCpYkuAFg0JLGVMf2Ie2kj38xE0JDAtKkU+UoafKJWrY
tzywAGpgTg8s/5rr06MqjOVm+pCbg7Sl+u2rA/hUQCOS5gCR7/FKCcvbnws8tNg7pJy3du76u6bu
JZMrS2k9rNXoctEOFlS/FKzo8kGtQp+GU6/pL1fPf3/C5zDLE/qKUvk4y6oxTFbSeSo4QUwUo8xS
eVgJoi4SRAqF0pbaDWoH2rQ9coSaZgXy7icAnxTsZ1UlYoFfo/G0xEu2KWnPkpI4DaPA640Iv/8q
zmOVTjHdwXF6Z7RtoaJV5yxEr7G3SvMZh79VVR+NCUBkIQIg3NfT2e2aCGT+aMaVvXEf22XbXiU5
mCaKQoNO+ZWG1LVJ9K2YadJoskKdipMNisINh8T5nTCPz0xn2HO3n9T4E+uJNFPLnRCcNYNOCHnc
eNp2ZYdNTOXtlx6z27hK5jJC/DROCO7WenSIel2SpY0j8wLT1YuXFi9Gqi63QlWtYpaEfdrEuqwX
kPdQ/HrUQAH+gJcimzTqe9hvvxm20av/zLW4se5Df3E92CtrXtDX0yQqdtGmkmJx2bz080WXsS1o
nrTokvPS/pPqSlhoO3xDh74QBh+8G32FnziROyU0ysJV5iQmiozmjGK4Y+Axms2gs0AWjY+zFYAD
l34557RivNasTfvIRhCRIcbY7RTrA8k98tL9YFXP9mF/C/biZHkGNQ9UR1sTJG10AdhSXOwDOT5l
RWW07eehiYGh6/pIisOwW2FB96cl880jvq7abLGnsjgDZPOcnIyd3GGpeFZ1ztwvKJxocRK9TkNW
iEhfsGqfdlDY10oX3SZ6rat33mkw/qaDtq9R4OZklBkhgVn7ttCDV+T9CmF+PRVkTKlK3vleqcuK
Z1NSy7UrpK6hzwEEzrhrvf11nPeWtM+F96qqLzBTFkkkbXBJzv+TwGGosouv27ABmBPskyNdaZZr
y9BaBBH49jcnW+hfPv6sFjMI0TU2rEMCZ/9xYD+I1R8p3fgXbjutF2fUPONyKtcBCE3HcagMDnng
LKYP+4lTpmHjAgiw720qeLNma4z0PeuhQ/LEg7L7u+1lYpfXanIibXcBBlGQJJdKzeY/9oqeE5EN
8Rdnr4OmFH4BxuobA/07o8HfrygL3y0RSONrUhWPju+bEEIfK9KKOzDEs9vDGwE4cpq7/IZjZbWL
2yKtnw/7CahSuZNEuPpHGDMZV8FQb5ZRLLo3IRZFWGyJvbV+kL3BLhGsyOsSo81frHL4kF4l9c1E
LAVGDwVOJk80ETbYuuPVmMNPDoopiayIeCzsmYbv4HGe94PmzBVjLaWBe3uhdtWJGnMKVleypJDF
x9Z/SDYE39zMM9wQlNDqxrNmh7LSIu4HqnKY31k+Bu/wNTqcIXPhoED50sdstV3S44Y0TZg/8Ydc
cS6Au8CMgGUbOwYH6R20y6wDieq4i+m5NHsnvy/vGiPez0+3iGNvbQ2jXxe1iz4SXl+lRb5iQ5PL
Z1+TX7T5IeYr8nYevJZgZNpnfYnC9lDRYTs2QhYr1SuN+oAId+jOlM4K0/GgujvHC1my7ehCpsJW
rI8XT3ppFfKFRKtbKunn/Lqvv7QFG0wTIp2jaMlkfvWkXjvyFAwITIJgSrxj426AFQp95daOhUL3
cX26szxObSDxNjQoL8gtBBRejHv9kN3IAfjJdIL/mKCBFR6QtrvzTg28GD6sjT1os65PsI5DO5ub
zrMTw2VOjR+ksh2vz8UnQdDrkvnIe53db/Me6Cl3Gq31Tb0EyATGgE0wSDg3YuLjbhi2V0IByrJM
975/AHMGC7s8NtZdhL+KMyQUTH5y8N01Pu3frTsE7+YquqrbTejateQ/TyQsB/6MycgwHvr2UNX2
MGoRhz98QN2O76LaZHvmbbv0+a0uxV24C7Q8Fn8TJgdwYwrRKgOOVBY8C1n/blzkP359/GaRf1Si
E/izb4yz5vITS4R6ByIpMDpo6kjhbJL14LeDIKES9XLVlQnQuM+9Rh74WpR8gh32L9nukhCoYRG+
00a2we8uG18qx5orsM+RPddD6EqCDRRPgKLxdwfu+fKQaKpwibCvDE2jd0ISEWO3QMtNETgcWU5b
DIsFZ3D8mhX+yakBid/00gcx/r8DZU+bmmJAnyURSiRXXmaOrFSOFtjVrGm0u+rGVu/pv1P1UkVi
UEEaF6r9ofxgHUer28DKboDIomotDGyDnlFy0jLC4AJEJFgUQsN/vOqEp8fUwJYQufspQ2KwMCkO
LnZ8/ng/g7g3LL5O4U6ffrnsaVRZX+cL6Hn5+3QGeFOn3Z+BI2tLKLUKc8goxUEgZOvCzugUoG0R
BjQena3tnSveD04ise4PIIo8XCu5UcbVUfuwUbDTTyUzNdogBPGaERrcvbAIcAQgfLHaezWA+arK
GaFsL//ejKgSvC9AfjzJ/yYpIbs2XypFeeQaalDOZFJ0Uf0KKj9IUwrZVzcRjDd0cfbmcnocb6h8
+GyQ4L3s1L4GcK4i4zLdn1l1+sLznW1BE1Sv09H5ayLRuEYGrWicdC/J/Qz1xLGMEm1wcKTdHrTX
89Sl9YzL3KVbtU0qf88dkopCEmCzPZaC3Hm0t0yDhON6Wl/uOF51QI//lQeACREQOYljOfQJgjyC
Idl12W4+Sq1Puz1mYhXvAfYA7Qf8MnQAwtGKN/Cpx3yPHl1fjkFeqVC5n361qY8r6pZdHwDldFA3
GK20UWWLywFvBuXJXCRXmyUcOBc1jBGuu0uqgk5hMPtSYwEPVmr++0f1m81e8aQV+XNXnkTKl5nO
KoJlWaOUDK5V7xgH6LQYlnnMh32ZU3mLqm0kXjaUm1EzQxsMxlO/bHLmg/VwRlyAWgQoZH0811bH
FdADG+nmRCVOP74HTRE2S6QVUKoaa+o2kHQ1w6w6UuIIxBXRp1YJWiXD0aZ5N5NZ5o1rx1lATsAR
SLuRk1Q2RE8SOAEhb9TpBxlHxkjaGaHgN724E5RVWxuaUJSlcw+ECgax2Xcmm4Mpgf20Qwuwb+ew
3qItAUko0K3rCSeI++BeckBXy/PA9UK323AnIcLC4qG2Nh3Huae80b5ltpA7l3F71wO40EJMEfvx
lJFhqrG6ue3AiGnooFiJ/zBkxrEnYdLBQRQEXM0wKB2hA+YAs/s3bHZbAQF3GSKQTX5uawR0+CDR
TPp568scnnO62TKp3naZPBbdCJO5zN7fVx7rREKmRjbHmBGsW0t3iV91WP+eG8CXxPPgF6Z+RtPT
wNbHooo8NptUfPcGpJNuA+IxjaUFrX9mP+4ku0bIYVgfl/QHNMHw2vbI0Oj+r1dALk1nD8CFjPA3
wg9tD+KlLLlslSNhUUSWKqt8yH0snHdSthQw4wq8fauIFsZFAcxwCFUSP6ssY7Y6A9tTxLvKYlSO
Zy0BSC38Hl72F4JUrpnJHLNEdocMs3j7fGLF16a89YINF26coe0n9cL3ttmz0yvhjL5DjgF4PvH0
bRPhIv6FDC8C+IO5/11h8jyWXK5H5PQVq6MdfWthyD4oQ+Vr9oUomIUqsULV5I1ZAEdrhhl9U8rB
wZkI3ZU4CM4FQC614Cqm316UvlGiQPUAW9tcYHjqmVL9w+GZs/Pg5K+45+t8njk27k7whBcY0R0m
QyxYbLpqXANm33n4USgH1Q4H/OVapxCiImdJVWosRTTXVQGmnaQMHG1uBgoTCElJgApwlNWOlt7+
J337nq6p6dqjh5QSkN4Jy+M6yU+MQE0e0GjsEFiVDDCa5oAjjZWP5Xc4BKONN0FkzrBElLbwasHP
PzHASJOmMGMXcc8pC64pLcj5hQuDlQMLMTtqqkKHef2+WWZkRiNccL/u+orQFbv/aEGisNww1IhQ
YuZubilA8TqKFGi+Xm6O2Oj7brPkY15eChhSe1BtGAWCPN+AxLN69eRxwKGNaVckw+7Y/7rzUZMd
lLpSIBCcX8pntTwJ1jGXNutt6+5u46uMrQF9fhpFPbOyt6I6XN/UySOmpB1Qi3GM3Ml4tb32tL5s
R1H5JfW2n0b8N4NJfXHXxKWfmpp9ZujJl+VY0jRCi90T1TeC1cUXMSA/92K1koBLj+u827LP9F8l
Cy+H9HQyKpquSsw6BJs2VI+Z9H/52I4GN2zPw7Lk5VaNdZENymov+HpRIWTri/kzAnFA9kCr/39a
4ZSYzTEuH2n1wdJkWgrswswEQ0IEoeGSna4S3fh1MYMSRSPuBjDgiQ94NMw2b5kxaJ5GlPAR+9ER
zJRQ9aAHOhWcC+Z3KrVZG+h2sBvtfwCZRnHJA/7hzHWK6yHspEiCGRy4dCghDAr2CXfgx5XVso7N
SAlSwjFnNppTTZxtq02QYjPsF9ec9r5nf/zycaKKaRREgJBwSNV0zeFGF0x7PfzKy/LNDh9afb5Z
OHjAckosbyS9yvq4/4E5fLmguUELjh6bQugygTkWPy0l6dyq92bnlP7PGogzNZOt3ivGXPY4LqO0
NaIrDZ/eYnYaGTNc9GyIkeRekenziM4fWr8KIV/J3c8bOv2KNMc0B6b/BCIPuX5HEsBBnReyGFDM
lyTF31MgcWt0wsDtHHynm0wOsYpQLkzrMrmg6k1Hb3b8/67b389xhc/4+ccCpL+r0f1XF4iy4+iJ
X2gVaWcfSmUww2Zb5gI3a2gex2hzfoAhoJ7QJyDzzZFm82U3/k4WINOs/y5xu5Q43Q/PZxjQCmmm
CKGz089VI/muzyNSz+0ootee+m8j/Zi164jwyxaOJ3tByY88bgThJMf5/rnTEtyYsL5S9LRlsPMT
BQbTWthgsmUTtnV5a2R9135k53ch24Kk1dAP7zC6KGNH1cXQRo/UwhanHCA+CqyTF+13PQT7FP0O
MuK+0C0HbicAKEkVBlT5T9Bn8ISnhvSU0PeSWaFrbbgfoWJsrDxajCSR/ZG+3/m5AsftUcZeZh4Z
ZT/8H1RgHLQskPJQfHDwYIrNgqSGUeW/veFcEo9/65iA2MtdX/IpiyfBUNR5g8mNzP4G5k2uAWZh
FlvBBbrnaHYPJfxB0rx5+asNc+vA51rdZe6DYa9WoZwZu6yC/UQ/OO8enExmYiVfNJrJCZxWFax6
Jxq7/3PEdY3z12+UDZPMJhAUwjJ2M3NJte+ZR+P4bEUt2YUtmgqvb2RQw9RjUP58V3ndeKtO3v3s
azKQYefbtfn0bkgCzuu92X4NFUqz3tTJYeNtdir4ALmXueE2Y+Q9jpuNcIAB6I816st4PrqEE7Na
9JgjPbfaZV/NVZaZdxY5Wb5Pl65sgdC+qxeCDe2zXdqDFe9zpszYq6a5UWGsDa3u4D2WaKeJ/BXJ
CvWH20rrBA2TCOmlczcSLz4raWxvEcllTvJ+Xh3HWrVVbSyfHJHHXuLjXmjNxiN/A+bwsjccf7KE
MitFf+Y8ckRdt37Wdj0sUfOk+MSY79L1bV76ZQu1NkIUmq062zBr0LWGYlhsvykIKrbfLxudFL+O
YYL+xEmQLTzc9eNlI4m5VzvPzuRIIUUmbhR6guiU3b3cJ02ob6jHB9aGpKQz/w85tRp9P6GmJwzq
5ZmHqSIpQD1HgpNwXsBqW2b6TX/KwO9/M/y2Q5DoL3K57HeuPnnD6TppjD/43TVOvT4Y+FODnJnk
EZss54r4NoAGdoDl0KhsH0Bafa1nW3m0enXns9I3jrip9iHyyNt0rHVHw/j2eZ+vnGRKo4ZB7bjO
0FifG/QcwlB9bfZ7urL2QWDkrCsEpHTErCMO+bLGI/C+FHDf06Db222ZU5kcDPJw43Dpe343CSYd
EcaZ7CPbrl1Paj7ZtjpvCdKOOnpj7t1j81hxxdx8WepirFDlx79NDlkj5nCqxMde1XpxNFto9hzr
DJqKkUTcTvRgVK3wAUmtcvWpAztqw76LdeyD8jn3vc/Mep4jW/Ur5PDdhexRxUu5IWrvMj4VUsZi
0437sSH8fizxayrpyaKqpuvx7rzQ/n7sQjWjHXht33EutOZsbBUQ3sngj/XiMK5HTFR//LtOPigp
SLO53axQVsHWhcnBTE3HLfqdi8xV0UTrfT1KdCH0/wRWjB0IsHksLdiAzCbpz70zKO/tGTBkNLVM
bcidD0OoqDnvU1TQ/igPJMPHbsfeTcEde+on/JqodF5a838vLJKHFBbzM7wcpB0emiQeEP3b7wzs
D/ZhprAkbAHU+2+fub7zeS0lvz+nJHwCTqOTAANMWtPqJfDtexiJ9sEYkGCainlSR/+tY0MHLRmE
GFaeRed+JwVf0j0WGT4uZLiipt5ALOlXbaIngjeFQJ/ByydgvWAbVshIT2u8DoTR/pUq8rLwPC2F
tah31zrWrblEyvq++u7CZPEFomdF0wbUYv4hPtjODBhhiDLcDVYxC8a/9pYE9omEsBA88I6k/l2I
d0nHBVIiox2xlb9x3UuUPC4EPOwEb/Ds/JVXARts3OpQxsNIcPFFLOZhLZwAWgHTnh60GY4T78RG
fOkRgzEL6ziaM0SvgR2tVDBUKQaC65I0m++lClXe/ZPdJ9p4ZBXJCFYXuknwEka8sErhCOAHKy13
T8WZ5ONz99LhYioRdnlr3OmYyVjBh8V7e0BYxlxylALN+Cq4QTvGrkbPPL3sLD/7ZWxythZdm5eU
5eR0YprW3Ls9JnQXpbaDnCkprit5bwfylCrhQbLnC5pbeWdmFdFAlz7pEdyHYacSJB2dRMXGTGAl
JfWApV1nON389aV35up9jHi6l6/DqC08uRb9tkH2ywu1UPZZCqsRxGDA+/f2t393s2bfP1KrTPWn
LZ6L7BS408f2JE8JCN6ppcusP6X/vbyMlyMEFiukagmBYIF9f7mkQN9UFDzAQD2xucZ4vHzKGZfU
wzdTSb2s0n/wFH6BgOasZPFeSLls2hngMbivaYkbpq26+H7GI7kk+ZbNKkP97UQlCwimy89aDbJp
JEwhBGGH82pWS4/HPKbdcw/12KVm/nZqqBHyYYs67Ntx7m+p2GLS9DccEWSECAvxFAfvm22TbpKX
LznzU70sm77/8Jn2OkSctFl/lKXZ5IP2BvqBE0wdfg6aATn+l+/T0lE9Ub5Bjd1nWMcoh3N19bMc
1238b8J5ieaDoUT3RG1LvucXW5amWJOTPst9+YUCkImHSya7EeXzDptJraML/XQg7ovI36uj1fpz
nU0kKs2ns5YxzIHWS8gFnQFN/pia6lDsFQ4+2/18DoN+JTqZjr2o0GUiqbajZz+MyCrNJwAiMP7D
ms2J3B57rP1zpTBRehu2YTMtG2kipoxoJ5FcqriN2LU8Z8Gu/BwhdxIoJFCYcvj/qP5Elx2uzngE
hWjHphn0s8uqxO2z58ark4wQn+/53befGXXZ6l8FLWueX8Zun29BzpKyz1QFJraPIzs9PG9yUeSA
jGfAJ7MCdolP3Qcc8Fj+UPCNznBi7KCdsl8YCwyZVhkelbAF/Va4B4fTdi1uOqzkVTCW27DcoH8i
SfQsI+PvRG57Ef6USzcO/eIz48LTD+YWzOPcmCA279aHwo8bVqOz5bQwqFWNYv9rWDxQdMes71IR
VFZ3Xjcg/OAQWbNJG4k7i6zkmPGuIJwvGem1JiQOhBmQHO2T1jh+TIoowQOIzS6NZ1afKkzNc/xH
euUEu06cplCfAo8mrV9l5mB7REp7HVTSSyC+N64CQFSA9T0+7fVwUOSltVMnVlwzvKFXntKWiFxB
OT4rBd2m58qw2sAT9I9VyuKKi33/xQ87Kqk6njBOICJTBMH+MWQ1aDXDNgvBcw+HGxbLVQt6nofq
7mH6nTEyhYecYMv6wnGFe3DUqmtn521c2KRzZfpDZNpSPt6FM5+4zCN7TeHqf4d+wa3iCga7H/nV
4pNeaq3yiOagA35d0wrqpqL+ejOCcsz2AMpo+apuCWAkzoBHMEYLVeng3PSIC7MVW2rdrU5MbcoF
jhYIToh7dNWWUM/D3g8WejscybIre6rXM4gQZ3y24yHtVpoAHbe0mP7OHuH/D2/kcnpt+18/IC+d
PlY6IiiA/AyhGVNoLYq51ElwvBMl/gpzac+QYqXpNz1dVS8t4FGAhsxTc+FnQt9HfjURUjPUWAuz
IZPluK21wZIuC2ToHJCa86oskRP2KVx+8hXijWoYxxT8INH59Pu17LXUxe+RsS2/bULuRaTt4R6r
YiMxg8RkglsfkKpMTyJuT8Sl6MaesbzyHHiRUiMAgM5VNOWGgG6puFAPXYH+BQZsvhvX7Cpil/ly
3WDau7jLogfKRUykyuMCVDSvYnq8ZsqdjH0qNGvyZeLt/hxr04pSfkBvIlUNuaz62XPyFM+sZqyN
ybydXboctcCXLosOaABNkqNbs4X/iCg6CWKOfdXEV1i4LXvwhK3+66BsZdw0wA2fUWDRVUqTAerS
24QHzLtAwXSXVEnOxTgGhplwlHHXJPGov7cM+WznKufl7rV25DCzlOWyZftHxmqW30a+nl1XhqOQ
a+EL44jWbnBSssri3HUm6FF0akOt6Lg4zH8PKEvtTsXOFNGPahPuLJOgB1CihcczR5rWd1CpDrLd
lISUrKXeXsVC/WZ61Z1FiAm0xIWGSh/+BZvlUiPuFlvdv9+BfM/LjZGsiR9bvXhlatz7swb8K3OD
ULFVnh2bN53EEsh5FKJKKtJ7+T8mM14ESafFVPwyiPJ/ofaVSp0vlygRZr+QiZ2aJMDBig0QCOjw
t9dWo8fpjhKGplfCrUz3ZBspw/9hfTJm1g2cdKcXqh8bxeJChDhCYTKzm5FK/1R0s4hMIXpvA1Zk
36IBflI9CVJp5N3QzKuc/0inBhKPSs20Eb9iqvKKFgdGcvwWJ0ylvFLBbXfTZzb8P2A8GZ/V2a5N
pQO2l6SusL/Y64u+zStpVswwLt4MEamof1ZbWblpdqFHVs7ISmGNZ6YvYyH/q3T8l1wlEBWWtc6B
rfMZZYx7dKTMV3nxnyGYUKsbI6CNRYKotea8RBk9iCV4C3iMpwGKn2MF6zKEOT7HMpDA0DQe7uKx
IhoyUP3fLp2fdJbUxlK2Drbo76BUUUCpsCvHhKZZIX+qNrlGKJw/kLwHEWpSXEh4RQ0rXbNuuAKI
Y2BWHV9Xg0onYTNyTgs0/D/wmgrywiMmiafADZYQvvXTgQA8LoJGhaZlYA66JUO5MEIOlNHO1a7u
cDai7MkIPmnYQkLydbRyZA1jwrDrY5tzLpuaQ/Bi3d+vwAjmlkvcpfdUDNbuhz7x/eM1UqgoB7kG
m0IsMB3dEfUZm6X+7cyRsF5h8vdwaesJkadSy4HYIYCmZulFXyubgN0Tlqu4j1K0/M1sR8LStZlK
esDyvwYU5kJ40dBntZhidhWJCiHtFYyDJjfS2V6dhMB/UiXbzWA2ooFh/285h3qpzRnkfhcZcPAO
YE3wHzpxz2LRCDlJ9dmH9NNNdsMTBYlgtkIwHjkWr/f59Izf1H0VO2rMk7z/7Rnb5ddivGyyHxxQ
1KVpcJnZiqIrfjSFzxxdcP+ZLD1jfUS3YxtKAs5yySqTlaSKFXlPKg2jOcZVOcSh6/ogZP1CISLD
VCBDCImMZH42gPdYbcGt4cSDGpIKpdnIj663vccgwBAqYRyVDKAVvT+hejNM5rRsq1JmOeCSQMHW
g28yt/29SWZId0Mt0bK/W+vU+rb3kbVTHsHyomRkj+LMuI3ihjdfMpfrYlGURnWu2SDaAM6ai6eF
/SMcGU6E1Ke5XFwEExwgcsBUlI1DdoW3T5tKzLTVrO7CfnsD/vzDfWovHZ8Uqu1HttbIc3aDB2rd
DtzEbOuW8bCdXNFca3+8jLop6dCWSEw7uHwto9pdugKtjXO4GbPFpsDKYOIRZ/8wGymBpLZEu/Sl
tQ50VR/libTr0MFbRzPHr2gQsj3kd4RXhbQLMpfezrcmmhIyYIKTrkHB6tPwXOSmDVBWN16IwYkq
R+lNxvApi53JRnygwpl6kNW66bUuNdzDc4mhHcLwipc5t02hL5sJUIrYbRFl66H+eCHpkp0FG2vA
hQnzzM9b12xQew3McAWMeBOZXklelEoWFemgA+J8URW6ASmetzazDUBuBbBybEvJQVd84hcBM21U
1PZSWq1xHMSWgNkoolQxXjFfmwCB+bKcGiKwMadMY9K0j2A/o3GEzmlA2e+LGr+AtTh81I0fzRHd
BkInTnrhTgFARg4EiWLccH5k2nvGDCGWJfBBrZujO207dFkViX3TksxBll3UNrTfbD/ReRs5qt/C
e7mV9gQ3Mv3F95jrOgowSUlJ5k5m9NbTMxerMBRbJlOnqP9TP3qrbNkjf1AxIAKUBeuB7N8uey+B
2Qs0dGoIsUv+852uakfOmtzzIHJ1Fzal8KGWjcM6KBOMxO4CPwdE+GORxvzQRC70FokUkceLh3j/
iSvxdUKbMxLKMoQB9+lvgSMjVqtCyz5w7/1NJIQp6ykae7lWUC16wARrV17SZrikUPFuFmH66fP4
GT9VeL/mCedUhPvl/eqC+DyVnjgV+X2TZNrVbL6/YZohZ4z3HiytV2AEePLbtPN62VM3RP/N2wwo
7K/oX0yA9zLy0EmG/jEvLSf3jJwKtLfF60H1ynQM1PItV127n+GDSBp9HrLRoh5yaJ+FpOdAA2od
/7deQvqLgySJ8lVc42FrjRGR1stVKObP802ZBYdHUTJkDUZYeIq5lU02aqNB7Pc58jfvtfSw/d72
3f7JRTffIWhxVtt1/KXkKPL5zH4/m3BBdGzw5Kqw7tf0H/uziyNM7SmcElX2GAFQLIemPcefNtfd
O6L57Vm09ZZ3qj8AAw/Ye7D9dpy4pMJ14Hh78CbD95z0O21UDRtocktwTB8yCeuzCnY6ftkYvOU+
RPft57RZMJ+4UQ0XKY7hY9o7DNj5uis3Wokgxlos8w7YWervnpUhP7QIrFfkP3dnvMEB/XndLaTn
9V2YoyLS+fxIUFo9ZP5nOclYjyby+BR/xxiDn4NRt970r2GYGsdacVammfaEyMTLTdltqidI/oF6
MntoVsKX6dSlglxCVqNyxWhU8ESJcp/0MMbzKfDIOA8Ff3Wj5ZixtKizPcAsVH9z9LUQ3oBvluTP
ucMAdOia4nFQ0bf8PZo3p2/moP1Rqx6mkdAQ9dhcFGi4a1MVWMDv47gzL3MjHRj8UjBp0xnow3h3
s6tBzaxhVubxtN5AR2dzgim/i4nYIOBjGbf1uOq1fTB1cbc9qw2YfnMRHsNHpfMeXCQwtcnqQpBc
FKhRc2t+Hf6CTThizyEDc9oUkfjvy4m07VSOhNFgnLmKKgy0c7OIUfBn33NbosZK2SCVFuarN3nb
vDjc+4zflwmC6U8Lfvg0H3/OWrzpDIV14nBvZ89cRhtskz64uXq/DM/4ZyBour1lo7WgOoEUm2Ce
c90OS6TO1zOyxQ0q5O+9Wox21YwK25NWiK05h2jHdHNuMmq7FjtoY3/quxob4E4Ln6UreZto3Dab
uXnQLg8r2k8akNc6drLv7OxbskWR2KabTts5iV1akoRLVC7Mv9wrkkoEOPeKs4HcY5Mial//QevT
dM+fl1y3IBxh/TZPwRwzvlzij2HfEaNoxvY8zKdpmX+mehP0FNH6DmOqHu4iM6EGiHEhPu3usS61
oB91UPVWvrkk3Rm8fz4NP5ZM8VZPNX+zdt9wIDg3RxgOPKTvGnefdtuVp/SAKGLqA5r9rz401afz
N0AluxfD7I8UCV2mDzAVoAUokhSYgucAJQoIL1cgpHcg4EQ9aG/VpsWmXupqOs+on2ezdO9gNDVr
bZdB8eokh3fcPAxI0woQIccSkPKVBVPgVK2cQCzzDSU4W/Olvm3Z7zedZTjOHT501GhLmYXaVUNO
0COvXl4G+lgpWaB0Edqetnq6tu3FZhRmcWCsbLqxjvzUeY6mzz4I5Tw3DWhx9u9c7yutvMxtK1tC
ORNBJKcbh81UaS2UMg5U+vD8W+BBHO9A9CfnkVWeBKuLiDNIeWHvgJAOTu8uCvBcWPWuAs7md5Op
03DFpzUNwNt8NvnkKAAQaJyfIrsXt82MZpUTdq9JQ9RAU7VrJO5sYCxHH3rakFwRdGGkSbaCwCR9
rnsBgDovyJw9xC9smYBGWegs0hULHr/KL59mEDNU7z7wn+m/yxo8/NXXPBpRApJlZ7pyvGj04ftA
6kZX1H1rVbaoGynkDOFSMfllRpSo6+Wzh7VxpMu3U9YtjO08usIel4RqNqBGI7AoQwAiug0CdgDJ
mxUr+pZJcCmt4comDLAfv3A7hnfsapjaGAzsc1IoPMIMmB6w3jddxadWX444s+8Ae89cuglGZqcO
+RuwrXoZd1rV2tVJ+mu1nLAmsi7UuMxHloB16LfRaZQdD9J6lZXdub8FQnoARB5TSEGlHsa2ae3F
/S/5FfUG9jihW/NIECjzEZCUFTV8Msm2dvqVVk21sykxiQ7zL+dbnRkot6qlgGtcmVp3EexSh12J
W7CrYVRStkNO+V4cjQy8UNqeofl7o+Qm1Ru0jRfERURZwzCqE1WV1VW3AxYQ2fBgS6VWaXdIzGG5
xHc6XEyozIbN9dAUeYoJ22e5ETI4oxeZPY8qlEiRMoYLDRx8yd0jaHK8Ew6ySRES8fzJcpvmze59
/+oOsMSiraKelWfAhJUypDk6zakeBrRt4K9wzHauhNPHUudo7+pss1Wu+VnyTpXP96rVD30R0g1L
HXJj0HWHT6DttOpBNVYaz+8wSFd6SSq7+CFTptNd9dmWySv4xsbwS1+IZ/cT6r0f3WQ0s2E+Z81Y
FVVUufttJL09dRUsCNYMZ3eBKN8tikveMp85exnrjYsyc1wvDfjy6z8QCzdT+a0qJ38f6NU00T3k
SMqX9kJIV0w2x2pfudnnyP53RAv1Wk2hhs2tNm2m41YgVukgaf4mh8exwOk9zcMEDMx7EELcNaa0
vCYMlW8J/OIthKusPoTa1OuVBYwUcAUnQEdQfBSP7fzzYtic8721wT09FY1c7T4TFe6quGIZSk7k
QiozBjcEtVFK7AKjni7QzO8SJSxP9AV7mtAZuK9f6LxXu8cpy0VcTLkYK7agB/gzRdQebRbybBtz
AbRavPReFMVzjGMSuVY4P3fdBm86TvMIe551Cmi1qSeLtRCFj5pLyQqV4uqTyPzSsW08X4XBhdBM
UpvyAoPis9AXTw4scNG/psEflVHXzH5QxvYw1LgAc4lsru4UUQnqmmhb+DPjWTuwQKujfrNDhibo
cp87b4ymDbIWnwgdO8D0ZpxSHpYnfpZr47i+VtSny3pqUCo10Z4CfUTPfIPwEppQhEwxd3bNbmil
4UNPC4cOMNj0B8RZuL/mNxB036Zg0tSl291LPjpW49Yp8f9aqc8pvdxtijWwsZli5/XblTvvYuky
AYAnwNnuT+9VECW1/gYVnBQlU8JnAP4qeMGTPWzrmUgngZa+j28+9Uq0TAQXn9NToElVpGmkUR7E
roUy1reGf5vQeHAnZ9NwIoIr+37DzQ+v0x13w0jjbTUIguLfEH4r2VwlKEOEJN/8NRZiO0YykW0v
0LswNCsSwUN2N9IQ+8p/ffbeM0k3J9qydT2njVG+t7pozHeSdaPo54ilBMIPOZTqYujhP1PWJAAI
X0oRgS8F1HW0FKeFhlsRJCkeqPqCwPPk8g5wSk3JNlmwOH/zKOhlW+x+RRqao3zUDakX03hHFdgk
vMeeJdm3Lb2JvWanl28dMmNbOvLmbwdhDrLq9kG8CyOENHcfpREIYtf325/06etQ8u/kgUxALgUU
vkiDY4CPo3tm1umE5G6TYT1/OQeEeKflPj/CDy00pTMwWfL12mQfqkAdQE9fEWPft8T16+YXumLc
MV8Q9f7UyhKKqb5wdmNmzDLc09ygxVVo6vZmRgTOjlrzusUrhhW++t7mOW5TqbuxGcvOgNZ2sPp7
YXzPuc1XWQnha15pri/31OF2rH950i96W0m6+BuUWuAVmududEt1EAB7ZlZXUfiguCdftEMU/KZt
NYH3uuuln26mSpGFtF8s1H5jMm/ZexQ+WgUWb5cu67OjnE2/lkpJUKX53DzpYdovESl4lScxyu2t
311CtfTRSPg6eox8Mmjty5YsEJjpuRdwnkRz0MHghZ8kgUAixuF8KyZ+EMdntmmvwqQNpKyRjQWR
TW0YEnHSNdYb5JZPkVaMwCzedvjiDCbTGRBOp/81xhdBTKftr4Kg+I32QUHWRZynVShW5z4VmuXM
MikO+CQnJ+qhGFFzTq9orCgJ+7yfVkSv/A1ACkCOjcyV3+878QLQNfK/ayTHGXRR2quj8s2DxKku
QMtz6KksDx2n4Qu62KWscC5eZ975T+C8l2aVVl6X3Pnqwe5rVlfKM/kRnnZLuUdonbfgntr4xngj
BTCvS6V3zuQO4/YqOu7dY8uPW1s6+RgJWDX7W7Q5ImEpfMwx+23qODI0cxHBmZKhLHjxsI2EbQDP
R41xlehl2tBOt3DS+OFhTBJ8eST/Vahzrf4tjXcSsmMp0iULc1gOVCMQL84v7zlwoRhAGpVKfpgY
0LjGqSzz/Um7nInExdHugyuEsuNWbkaWguGeP41y/vGV1wUvzaANU2FOzSN+t/DsRfS6f528l5e7
WQRR1C/RnlSTF9Xs7DoHLNepgpnij+WAd+Y4ONPRRz6aqUPuOCBl0+qloWlLMJFrRmfooJA/GpaK
Umj4k9wmkrEm/9skpv+K2d072s1Pde6sR8yF5N1ol1Sc8xvyfeOXZYz6zBpWsAnQkMEyEMTAs0uI
LHgUhUyjF0rQKc3QUoEqUACfNHGtaIEtOSzxT4cBkYB6x98XJMkGFsJpHxYlFEqqZ7xuqEidLYho
jPSq09/URkFQev9b5bnsSe3rh6zPi8b5yfq7UEE9rD02tLeAU/VOGfCghzjXPfrzgLqjthoFSKAP
IqKUZ6bLydUmPLfY32MIAPasBPp+GuGogLQk4Q7Q9YWb3BYyMaleZ8cm6x5WD2EjZ+pT5JC1xFl/
IRBfLlObDZKyQkiErQ24rhpeRdss9dioNYWjwwRiNBuITYHm9I8zHBODmfQniiFW6F1ekDu9FNqI
5H5Hci5kuPL2onf71Idep7BEOcmz1pYbSETetnl7lpteGtvXdjfHocQ+jA2s3DmcVL/UOqWq/T3r
85VIoIZYcDp2DAx73MBEpxPzMlFuvCVeC8YuoMZu1D8hbA1tIbr9r03aQkQuV+SEEX01Z/hS1VIN
3zBlCAynNlKrSYrbKDv4F2n01XWmsBnccZE9DBDJvgMkixotdW3pyJV6XwS+qeKlodIUnZqSkIOp
LnnKaajAcjrsA35xDT6XJs4YmzJYu9N51BcFpqUaWb4XsOa+ZNnrSfO2hG2qREuvpy1tTMBEPjnB
Hdbwte1wg/2eLFk8+CnwiIlfcPZ2N1FdQsi+MnUJZACl9fu+5F7zULEe9e37tA744jOphInQXUDb
43/TBv2cZ8gTRq0Q33pSmRdrNETLMgsHlUKK0PPCLRCPDBNlWBK3JpLrpXX9qPv3/Ri1YTfnssmw
I97tnCGC/f3xnzZM6kEsOhgPJkilsefHBOFA68G2zVrtAUnSMH5lbRu4EtvG+/nivbSpmszu3paY
pDYK+J2dneZMNejTI0PmEr++FZ9xApR3A3ojM7T0NLl4an5GQuOcxU3fJTRiyDdkkzettmLDBQm/
4Jrxtl4iHyQo2GznGOBYL3muXPGpM6Uz8/BiKtjw0dVqG9Z0t5R7arusniCwVk1MAqivi2XyUMoB
JSPLZDDDyzGuMjMXXEKv8Ye81GvMfU8ylronEqz8lVvYezoWDOa9BysIoywV3jfbxBObSHd30OUf
1ONSzJPh+nwz0gpLbPn/eVRX42K9SxzWSTZV3bQ9im2hTHb2+HWPrAmComxdqeRhNnYchRwmyueX
LEVwTDprjTlFOvm+ZvOdqjNafFV2GerXgyyhMvrocZReg80JDqISjP78mNySTp4ZkObQ2xJXBw2r
HlU64EV+dEyY8mJsFURM8nYg6OEitm9gCUook6FUJilxOvCxWr7fYngurg873M/+F+y6p46upHTf
fHjA7RKwdsY2h0uuyEJ4DGXpodaBsasQIT721TGjwD9B97zGAW/PWp0lgC690gIWIHQJf2uT/+2f
HAx0XB/KYyj8pXYcOsun7+G8Q4b3cLjgqKFZga2M0uehtFklYq2UfHrmUWCuQ7htGGm/10LAxd/H
tFW5U/ZKu5LZpqf28WckyZoTBnGiZx2z21x3vHUfOUrxeza3vL3IYcNSLCtEQv51nEGEt6uDIA8t
yqSwlf7KUiE8ZYJInWXKsV7lR4xWm/8iG5OvpQtkFFq6zfkEqnqMSFius0pcDBUlg8EoNSzfHlZo
kEDM/4sXzUK6n1FLsNK1rpcdBt+yGzEijQsxtvZ0LYUxmEYKXB63MfffWs2mQxP4Qmf+STfMkjzl
Xr8ponvNOoo3OvO2DuqgnDsLW54DDKdFg+xDmY/MfGpCTEHYP/izzUYs0NE4ISp0LRAsQnb9KFfA
ry+glm9bCaTrOWvaCf4psaieR9A0o+VOEulczGxNx29vQsnQU926fQYnaw15Xsnl8xxzZqf/AlyF
gsfmEBYVQvctfadMMmsodcSczZQZNqZSFu8IN8DLAdlvF4iO3VltU2IsrO+tKUwJlvkJlz60BZEN
DdLlOtHDVcAitHe67K0paM1SxQ3ry+uzBaER4uoKjtyZuhOZHgzUpxS3S1w1upcFFouck2DY/aZe
XaekmHmHzUDh24Ay7oeaPepa64yc5DpG5hyo/sQML+z7sbJ+Y7G6m45yBW0HvyhyQRyhjDqRjL3s
m/sxCkjJ4f9VTIMyDkAuP3IoDa7M3zygxuL7XnVvTWW8jnhiQbELw1oCaUTZUiliHlVRQ8/5V238
Tyxn+abNyC7igMlseM6aU2iRzGnf5Pdmw5gCophDxEDSAjbuA+fJLDsS1E05KeyJnHqNtzzgAYRa
kEebz7mR44LZLN/TdZZqdp+EWsMAx66bdggpy9boddMU7L5YQsA+FU6EJczgnkjQJZmfdZt5h32K
5bdBjfEkZufgxxNVE0uenotv0oxXGrsYQA+2DfMnIn/Vzl1bjVeXnMqdOUN1aMZZitQuX8ALFLUH
5tOY7GC/6Cjqz4rfPGkTmDzlR02JD5+dzmzWXWn3pwJKE6D+rsAvhePuY8wRJZ+xORC9K+CQGx+d
qnqVkuvPo+mD/2KjDxvMyCEelW8/IpBxXvMKMD9bvW1hNogBa8Sr6SIPYTF+BjQY9qa/xA1meIMN
gEkpEU1eWv8zW6r0upfoRCLILHVKQllTu/Z/W67YhsaadvFRICsYvoemtl2FGDuixiiCVgt9ESWt
lyAYrCilzqAwN1Dkr6iuDUD3C7CO++6T65RRvDTYyydWBnfvbKOW9D1sQcO2N1mt7/tFsTcySv8S
/QMueE1EO2W4JqAxmJI8ZQ4DNVpxvYqRqxHSi7vEffvxNiYPiFd0KUb1bMgEjOHDKJ+mzslJnFg8
6vs09yOBC5vXV8vPVZHXWbffykEipDJhmYh8ZAx5lJY0TtCt4zmtuzG7RsOl+arkxE3JS/uGfJiA
KW9Js1h/CufffqHiErDmtz482GuLdxgxSr8zHmNg5oKKT2fv1x4lB0xw45yCv84hkfm3zZnmQL+r
ogGVg7otSGs6QTDp2mBOb224CIAQs1AU9nRyNXyH1kpeXF16Bfz21ARyDVZLO/JPOFvcYXCr7n2q
T1uX2a7vFPbOfvMIG5ClAJsDd26EleVrLvLVbsx7UhhJhF9xNIliN6OE37EVMe9JxXWiEixAM3V1
1l6Api2/hZji3ZcwSanm/Yb2lMKr2p4fdaP4A9QjTeIRvdMe9XHTHAde0FhEUV/Pk5MtMgL3KgO2
M2eNd2nef8ZxG38id976FkD+h7kS779AwCE2rJZbEQFuIwcL6yKBe5uLCrMbeY0jLJ6KJNckxuk8
TpkKBPWEDF1TGfWh/b7CEN1Xv1ETFsdeyIx/AzIFQrxwx+4aehOIjK43eaonrypgB8JJhZgP/Y1Z
+gN5vNGwbMm5jRPBA9jm5kvEy915moxSS97fH+XgEduUw7hJlIcAx3INHK4JQjeTMg0DzCHLRIhS
k+VWEfg//R9DmpfverAbRgx/fCgS9xJ6PVj1TJQtetQIfPMvIkuVAVaPfo7G2bzHc/YO9C7OV1Ja
pXEkWPT3UOia2n99UsKs0HJChvZLaMmDbax+vgwyYUG7BUCyQiBWLfTjflutGwRHA/vjjCBh6udU
sjCrgb3O9X0VZ38ev3uSmCgFZAM/qeY+6FmJIF1wW7WuLt/GV9AMbf4B2wFRSFcRu56zL1lVyn60
w9pxtExUQjN4qShvJ7Ez2jGe5SA/+6FeKLUFrVKL4Xrky4E/1IVs4I43/dl8RLJLId8mqqSqQxHL
Im3Zlob+IjKc4yLp8Ky7wZaIG4404+7zJJKSNpb5SU8ZuPYsZitzswIrZsOCQx1QBgJMVd0mLZUp
KTTbb5UojUGAYBrjDA2e1goGuOpy16nhzbcV7drACPniMnO+4C2xpCQN+hQmpSr4gjO9P6WQrRgn
EKz1ZktZFpFhM8tx8jYCw7kY7kCI0fJ2a5ySWGEbTOx3jLf9k7ZlVE2cL4ExEvqCxwVzPKYUFMit
DutBHy5wQL/qvukqJ6GLhgBTegfNs6qz119dbudRqR2e5+hcqpuyO5iu62JXjCzeLoj/fDHUbQGc
U1CGIy0ONoMQ6gBGvsyPDQoJt1GobYmtW/P4lBN39WN8wUzkdBkwPp5rS8dq7KOZFPNP9F/IHk5V
V80teISOeZ+y3dCY+xLqkqyfsn18wO2AKEEHf4EaKSG+5q9tHYFwzqPju4yBh+A9pfWJZ+oJDhYG
OVi43is5AH3+xJdeUhl8Gcaim5hkZBqU60TMl9bQ5fPLmtXrWAUscrP/bjz/OuNl6F5U0+ETeFnG
sj+7/MOU5DrTYYtrHH94/k7uhV3oP9aPLlH3Lad/0CN9oZFrU4wpwFFgD1y32YxugwfP+hnAcxS7
7fL1deoacjTCX4jpqAPJzGLBYvqG9nJODk8cYIEDbJ/C3gDaGT28zfnZg6EoITRac66lCVN0S3aP
AtWmSeN2wCnS+1/E9wJ10S8/6WnkSVXWOBhXhDO8SHDJknIiXwgnGcd65733mXfuUyvi9A2ThvOp
YS1095GN/gZFZLXi+afK1ajyIypBfOC0FM+OvmMDzMff0MuWFDE0E7awkekOnc95uhsLr3jj9zOe
/wzzsHscnx4DyyDD6xfQR1vPegSEMO8wNtZsFXMliIckFEWHXG+awEyIMpVatiWx5zVYNrDRwktM
ODFDI/K40ix/YobKaztoGo9tQs70rbn4l8WytkJukTlXs6ZbEfKgbH0GkECDtcvf0OTwU9+d5aBO
lsfQ43mbS2b4boBRKi0+R32oD8R3lzlvgQMqBOM9DbukOHEoVeEt49b62VRQu6CKFp0oS9RJ8E9k
ZmuHR651YJSOTy3DtkGlyqT4m9uCtwMbbSLLkcgZGnp4+GC4ST6lWGrAAw+fwJ0bUffdxQuaza74
jS26BaNitZ/NdnFdvAxCdY/wCWCQ8L6QVF65GYsYhhIFGI8KPts3fE5PtHueyUn+Qz/tFhdmKCL1
xbQtKgWpBJWq8Uu+bFfKVaKF8H5GjcEjpU/DUePkNMe8k2AqApum7MJz9h4OQhQ+rbknifSTt7BW
ipKCGnPnMui6gzo13sZR5tWTDBVtMP1k9TPZUoLYGVvWS4CjBicwElom9QXO0SJwsFppEfwVFDsG
zB5Da7uXV/I0UbB+h9DtIY6AeT3DoE4kCL2wGXgIGher7msZIuWUz8LQe9lfoIJFV2SX8gXcyOcA
gm5X5bFxe2X3Iyk9Ra8zfcEAmRa+Dta8N1rQo29Clac1sAGreVqE3H7iupcf0ipPwQkSI34x0Y1Y
mWjHzKxl8dPOdS9K/RZAtL7DzY0s2F9iE2PiTGK+A1mYtzWD4kbzE/XoV5C8ksE1kmDGoGhYKqsD
HU88DtsKFVZvwGU/N2/0LiNdQIezdQpCyMLC/u4I121XRu8yi87OXiqT9ccGSVHAAAINZjD7XFNT
RnDeX4biu8U5aCuu4gXje+tOdIBXw+HwwREP4z6BhIY1EuFlyty04Qt7aExJM8RL5b0LFeyf5F1B
vqjEbyVsxh5Ovqa6Gi68TAohSIHbgKuULo9I5NijUatN+BkjHXLmDuYfXUiTPV0jUgaD7VAopECk
co5x5eRcZO0W3qxJb7wSmO2iCQp1npmhx9rszbpdMU4vGU7ozWLh4iZeBB/nj7tEGiLmjaqcGS9e
+36nM1bglrrjPZOo6qMGmadookzTKlMqCGEuM+f3bHtoSKVgeQ0erYP1VaUMCsb1Y2XoI0tEAEm8
vFHUwJyV2b7wpR2yldOo58M8T/fikOP91AzBwXKNFMd1efmZsjEcpoD+GplUNHcnHtPvWCYryokj
4HUuVVKrcSbTLrE+rURnWgfZrDdK5F9v9UASIFdRcgfnbcdoyMpSLXLqgyRwdWGpMWTotaTgVjhP
vPaJ+yJkN6qYvhY0hOlcx9zd6ua0MH68CXFyeNF8tNm/ZFTZ9VqRykyjPR1aurFtSh88jhsNnjts
lUOBSoeH/a39nDgWp53/f+BHd9Fti5mqFM/VHlRYE7d1Wj9KYT/PyTG7Ej1dBnq6R6xkMEipzr7M
b4zwuOi5lXW/72CvWYIyTg97TwhLH6D5HObxHcDMyHtIdNAce1TBgwUI0CWCp9Qpq3dtUjQr5bEb
wVTJbvtdUevd4t0HtLgT6atcDzpTwNqrvxeL5ETg95PkoZ8Koru8epeiKIWaslfdYauaqTZvjLSQ
szc2PSJZD5gpaGMxNPoqFxHzG5wTkUQpdcasRV12SMrGoDDoIq2B84FVndQ8Ovzh78vWX9s1WNfF
k+2Iym6Do6TPIPoGRMo/KnaIfSQn270uU+TtBmsGjUpnxfI4tVPJeh8D0uap/19nhKbxgg3OaygA
zrnqB2SrFxxefZppsI6z8KkR9Sm81+B1eVNJEpxjDzegC9qlGFj3OnqWvemncw/5EdPy/B6nWY28
VUNuFhb/W1Dz9QnCYWIsRsCfd5yQXAr9ClLLZG1Wr/w31Y+IU3VfWz8MCNFeN0Qrt24Oqx+NGIvu
lTxefNnjzjQ5ocDhbdwaMhqsG39MHYd65ejpXf0x+FeCvbnQ+mg/yanNDc4wNBU5+ksOxMd4fdj3
wV1LIC7kuxmJTXdHhsJYdlqpPVR30Htxv4spiaIMJri8QsXZKS/B3WTAxb6+oJM1UwzPWn6HuZHj
msuOhvbgTll8d439O5IVofOhLoDh0UcLA+bwp2mOJgFoHKq4mie/jEV+lX0fQZXQL29pN3WeUqEV
9gc1hH7QIXLjHtiIIkVDswLtaMQVk9uA9WLI/+lRJgaa5TToT0HPtvM7DyKzwHP3peXZXNsovHvF
K59bxwO/viFgpYNGMD6qCbM5Idc/olsSGCmUBmp5jYgIX1r91K6dw9X+t4kpotHf7QFzMB++a1zr
fnyF8xAgF6xo/ffEmiK3ByFian7x5xD0BQhh+ALWBrSNECw+UQPoPqclPbrXByoVTaMZQm7znRkx
7VWExhF/3ix9UZlKJALgx7V2r3PZ1zSs13uTku3+TCUDZ5GzFWgX8SXtbb7q81tBxG/hv4BbjAoD
pltEfplM9UwVgN/a81rN9CAyDd3zjfp+9ZoQHmp1JJvugGRI5QpV2dm7vH4ZmViZsR0wGc/rdllv
GkQRK0bW/42+dvsyoce9fpD0ymCC11cVqUWVFj/hqdpX7lZ+6t2+4wLKGkS1XnWuoY7OR8jFWZoR
PN+O1x9jMtqkBaqjO1wMTjip3RafqPbiRl4Qx7rZ7+6aNrYlRmwPXBfwVFlHfA4aGJE4NI/UmE60
at4O+s2gsvFePkx6UMwk0MwKMFfUkNQqjjdqlrWYav8rMqHfEKQc/Tb4jOxT8ZyzJ2GSghVUaPSj
5/fNrz8KPvLkucRYghyZQ03KYYz5z6sXPsyDHtpoDbNkyjWiwIQMElRe60YfQ2vHKpCS2TJJTFR2
w0K22jAzaYjuspHJotgo+WxJVxpmO5WgHyqfvW6uVRC1Y6lqPqhdvEEVPYiTLE48ZN7Lvk+aU2qt
DbsUscQhfHY7Vuf8oGbCwqBxWIZTNPc6tdcTPCAdhV9oNHDCidQbG/Q3/WsLP9I/Rp4hSqqzlfRB
kz6n89nZgxpnziJwshFaH7zxjyiO4Q2NxxXWE2msDdnjof0/eA8AjAA4sSIzooXJ2BKZgOv2bchw
4gg8Njz9VxtYfDEi4N7rWGlG3P68U3e4diMF1oGbDewzfe11gtnZBsvwkwImqbSpUH5z7Rnh/Nmf
mtzg7K2YWcaAdp9ntdiHqMP0nD8YWiHpCjt8cWtQEscLqGCAmlinA+4rWA/ppQ2aZW4ghwzf5ov1
lMB36Jk2nyaweO1mzv6J3hvIUHK/wfI5rpDtWCWzX58/l/t2FStFrbuYbtqIsBkVni+Q1V21fJxb
xKk7iky4WylgR7plARAmm1VYGRHA/KXOL4TNKjqFte91S5mq1+UqdSdW/iRXWa01EDS4PSVXzE5A
S66b3wgT9zVzEgoDP+87al0x1X9i+RJua1mS2sPrso6EnvUdos7W4r/P1PvlgxQweNDkumhPYUAn
JfHzmrczum00cHMQkpANk8XIPYVoKTs43hwSFUFF28EriebcGosKJoz+DpdhMlAdXmyRUgm627Xa
6Xf1u6mqXtvWdNYD0H1nrjL8xyHB5AVsIeJxvN2RFXU8t/0lTivohTB3MIC4w6r44M2pV+oZWDgz
T1gcj8sKR5XBUseffSwaFnrJpJhf4y2HrjWVFwzX/4VU8mcxemaOGD+5PNrxuQhNMgZXHUygZsk1
Wp3xEQrKG+iI0sjKt2OgmfGtU7fVoEgTzi9F9xD3ghcBXEDoJiWieZ5vOVnUDlli2IevMNQMGNmt
0wnKe48EkKEStU6EF62ti1RSIKXbfZSQPqTUwRBf+FrudAZejJC0wt7kq9DchDeJZmqBvC4oKnyE
xk+3vqOnw+N51QpWhcfRP8vzXgyJOmmKnHa7lUpU1Yowil72w/c+gmMC5oVVsedxneFM0rpbfEy6
PfSC+8L2kArqTUGNGbNRsLfgfw464d8+ZBaF08lGG90R5hRXpz5e1lmmacX7QYIk6jAXe7Tgpq2i
VaHdHjpAevvdA5ZqejpwcYV2Or76vW7izMZuBGWxZva+FhBpUzRZyIxOlUcdX3TcEZBMBcV6Wq/b
NLB7oMw5qE5XprXsRFzxnBqBqdRSufs/E60uk03UR5+fJLnutQXTbWL+FX6Fmn6KE2PLYiiq5LX8
a0UrDwT1bIWlLB58VlNCni58D3a6K2DjxPxmYw2A/k05MHeNHhC0K3oOVj/WgcoqGmknWbW7NsER
YM2nwc0xImjHI0mhhmJZNGtdsokuBAU5jcWlvK4tnjhleLIH7+oLxyWcThxLzJUeiMmgdR7lQD+I
74NgYXMFysIt2gZyHlw6tBCEPp3b+RAOc0G1ce28mo2eVtVZPv9R88Z3ejYcWt2F7aWS/lJdGppz
WXDBsZwrRGtG+ieQH7htSwUv9/4GSXg4+s70pNF9mVSWOCS8euNF0ea9mtJnZrajsp4oT0ttNqcP
0GvXow5agbVX0EdXk66r+WQB7a8J2TqfzDF+19TTL6i/YMOej9zsKo3pxLfKZb6Nq03rgJt+82//
/NZxZvimHkMuC3BtrLWVCxCv3CRqTPvZCcfGvBFTpDAyEJjEv89ot3nNP+90VVOBsE4+THuka+/d
ED63oKroJJqOHLXSJrcvFG34E9+oynGaUP4GDzZ3IQLCzOA3zhK/Bnm346IO+bQxq30DU8wVl3KR
jrbJJUX0YrxBZq5kvwWDoLnVblyNX82KmVFq/gX8GJg4tbosJTFv8wJnaXBYngYMV/c9DVSMwy1h
SA5r7S56N+DDWHHOj0Y8xUz5eI/IhfjJwbpVk9TPKEZGfjdvlmWFW07LsKFXfdirfhTtsqh7PTTB
n0UnmgEiu5khFPj7zzPkYX2aJ7sgJj/RS80a2r4wdgM4eS5e8dPiWURcPDx3t8Os2gLBdNe+IU2q
K8/0zfO3cpMXzOh4d+TvBrSZCl2J5fY19c+8mTRDDDoOYRJwBrhLreuxX7R9VzTREPYzgm1UNHy3
X+b4NvhoMFtKKHDoWoM49dlmnKpPYlW3huNQPdCkjrMYPy2X+SXVCko/Lj3mBvTN4OCtqp+oEFQb
bSVnRBPU7WuLZiSFkV6KM8IfdM8eBRr6SiVcIMtIT/mzApsIgF84e+9B1ltKgCOKIVI2zuSk7a13
lRxm5CFfErd/wIjsnC8R+nDYQx1kmYZLMdt43SX6S7IoZ1b23alEOE15CN+i7aqV19eYtjj37DYK
JE10eP1y7uO+6mV4MASHKKmcyoGN0qJnp8CQ+mtDDs1dMyYivxciE6wuDdiku7wSRiYvZE0am9R3
3+Am41wR6YlOkW9JSZuoIMpPHy/h1/LBz3B/DfiHrk2R+xS5uteWY83OdlRJ1eeKYYDAeWG2PWBL
J+2S/b546izrkkGr6GZUWw1NGpdelfa8vyDPrTxbe6YQSjS8rAX2TMADgfaS/P5ctk9rkgRXZb94
3TnQYEtsQEm+V3pOBa0gAgAA/n8ZWjKkcGS6Lid9nHsEjr+/sBdB30B4IQ4UyiN/sYmIsxADtcwa
xylQEwJi1if3XfHaH14UFqVa3x7g6GDwqVMBZv6VDD3c1IjhWWI6k2ZP2xBpe/D3IFozMSTiq5RH
JSPqbxgwv9QB8R4okd34efjTXVAwVjiDhZFobXzr9LcTVsaFO5WjKo6DcTCty22/YLnDSK1st1S9
h9EXQqrfTSXWalqeqVggqETY/8bYV3ojtg6biUYknU9uu/q7rbE1afVNuUSSevh4iwyLE6GKoeMY
4uvvXKRiKMt+P4FGltQ00mOHHlfoZfiyfW41QvTDrDeym9H1J0rfTd/qJYBn8a8RwrCzyT+FHAl3
/p/96MefCVAJDFDABKLC/GWiV3366Afclh2F/MESf1XhBQ9WZKe9RxzB0BysfH7JCVQflXDUDMQ+
tUsDRX4WPuRjvPLeEZI4I5Zs/+9o7EP7G7PMWq8ggxZ2gbKhq4tX4aRHnJ9FmffnnQtDMEK0fjr0
dISoMUzPRVjriWKJpBQzgsF8AMcsnW/pESmAvePph8Zi4fPoCm/al4/QQPln3e3ZPsw+G1NdcPlW
qS9CIzFaPx0D4J+n0cdE7PAraNy/UalY3muhbUgOMl72t4HJWC6fYSdKLjod00K8Cux6WoUZgWpE
Q9q9T9IADMME8aAKGJnWNWf0rZ6WIOpP1mE5KrbPd/F1XWRfpfP8y6vuswPULkh7I8+B5BF/udNI
LcuzvitKWFZtTZORlPLOS98efbeFCInxeEkBsrja4ukWB+iwTG8FhjWRREsn4Pg3gwcv+yQLNioz
PDlkV31Xmh9SrprCZykmmXQ4XniUokya/KOgRr6yhw7QoVz0RjGLQmP2tEKRV6he+Fm27i7szK+w
GrasioRmpYs1FEZFx5EgKwX+hoIStH76sHNYAquY+ywxK00J/TTnr0sRN1sjUQBC+CvaVp4cce5z
DUSl9kLUu1MGrpD30w1AK3wa76WZ9sA8MXDwSRNRM3uNLiygbLNiZIUR6shh/S2xMxrsBislyGAL
bAJErTRNNfhnm8y0U3+L7m1omHoR1LIlWJGldbkpNjTJ7UITolSomCAYcxsoa59etzRqsVFKFroA
cjMhmYSL2PoLvVKTfwtRtF7oCz62u7+J2+ieofVyQ5HFCyg4J7cYVXE+S5ylTcDntbQ8kqJlxG1I
6sEj4ftcNTcevCM7yz1VL8UvIyynMlLkqGwCiGY+KLAd3uduZzDRmVPdNMVSHNhRUJFDLzBefxeu
nAzeOvXcT9oNU4ATmc9JmGsTv8h9DRHOl0HDFRK0c9eOc81YU/WsocAxXS0Bd6gvXTlxW7kaTOrv
0eo/AHxwAtzOEcVM3pgkQmOrtyg4xWw+ZD2xVmYrzqpI8sV8pNvgaGg+0iyCfay3sJvKRFhVvpMc
usUiT+TD3uOSmq4PJHO2pdf6eo3ITOKFdQGcHfoa7prv5NEBlDM+UQzXGZxojTJXYU5/GyfEHqJc
/FTzaOBol+LUDXfCBwARF0wp+99E9z3fSU/J2Uu3C+OY9wVuAL0oUnTu6Ooq9AKGtI3DEjN+hmrw
qzIT+S1fe8U7IccagF6Iw6PDADwrfM42LVVYfmrlohbkLwAoqb9m7evjLb/VMMsEwVLcvw8oG/He
1t5t44AVF1+h7TN6ICQwttkkp3IYbPNOFxzv4D8sTuGPaXaOsAo5liDUElBPtbV7HmkysntCwITG
yhejbSbp5L2R9YOiF8D2Ge+0z6ywo4vVB7PI3mFDLII+obApThW1+zaSuCDqoecV2Npzo5hKiw5S
mYUcm0OR/AXpkbHz9gJdh8wWABQMOs0lOor7EUbqhpMA5Rat2BGHym0t4Olc149tJxbe7mDXk+5K
v+zB8LxbNVYURKMPCPCnNbfY75N0JFwCfijwLgkHXlXrn9b7ZCzcxop5P8XEVn8SE8Xvx5IGu1UU
xVn+4laW8SZ5jPKFpBAOC/57uhs9iM3uZil3z40ayDtNIzoATAl0mTK0iHeV9GGVa4JT6btLW0Ks
Oh9XildNEhvQOsG5yNY8DRanKmRnpf1Fpi1Dj5nyAm2KhdzQ97pcH3Xb5M2j1uOOd5xWH3joQG96
rad/zSTiEKxWbgKBuKv/KlM3o781u8lLANWE4MxTnHjQmM4Dt7qNFLOcDF4+Y9VfDqOAdOEli/hy
U/7+AxwLTEfXaTTGup40D0ZXpv/nhPUqPP5QNdmEbV5EY5d1XvNznTga/nc552QEOtQh9TBNcsus
jME9Afp5Cop2zgm2tqqvzaysg79bDvXUK97Ndev+vAOH/l5jB4ad84w27e8rIM+PAH2GcpCoBtCW
55oUdngWL7ZM1fXBc6nLQpXgWku2isU5Ph1ChOQFfqEmiLbb9TPlDfmiI5DP8pyLKRhayJi+bMcS
Bwn3MtFWAfEMHVtUBg9y8eMqGrkUAnqE6l4Y7d+c4e55yf7RWVEr0kvFPXcGFCY/pVpsPRNcTtlO
UvpdTeN6shxN6jikRODDd9BoOzZCA3CSGGeB1zMFJPD5VScnRrXkogLAJWTU7vwx117+TuGXgHs9
OPUVZwL/kYMb9Ry9kAHMYisxrVvfsOu0rr3PNLc3GYgACXE4Fwg8Nlpw7zResvLqpvcsLsIn1l19
kbGUnveBe9WHV7RiuM3fBCODB0TNG9bH/Gjv8NvN+kAwR/4VZhV2sqRIN7kS8r1sDO3IrRgUWEbo
g8SPGTOfxX5+Th5rHBtq2LMEDYoK4sIHNQRY26l1ClStHNYsZmYQaG30vNhotPm1AoSO6oY6S/HR
Fw2UuwEcUH3lX/mOo4opCv5EKD3myzqr7xUvkNUYo4RbIcIF/9YptC/+V6JufXyhVe/JEc3XBlW4
+HENKngfDSqAsilS+vsTfRvNwrcUNb/dnxySV0RnyhT8LRm8gAH6EZaeuILkkVPYuJQGHNb2brmk
OOVDoSgUVXE0SmxZwyiOl4wBPIOXgjyoNCEnIbUIR4ZJdTGM/zibEUVOtTvYmEsb0q838DSKeVft
WBwT9FmOEJEYF7dayWrooYT4CP6BoxcfV1dSDAPZZZ3Fg0JZcrstufxhbKjDqkW6jyAnHHFkO/XG
xnKBPOsPtaMXjFzZImooTPto8lCBn9gLeyO2BPmAniYwsa3vWXPXk3ONPLxCdBtZEnKu7baQHHtI
I8GCEFOY1+eXA2URMD00HlxjPyf8FwL9Ce5SIGZTPJNF8xJEoefCw0xAfuFPuYWWrLPn7ybWUBF0
hPTJK0UHi6Oh/GRtn50dE4ddzEdD4J2MX555JvezFmjPTc0v3d/Od92aFmuJAQ/EDR5UkkzXtxRv
jkBLwqHPsKAwuDqFsZYHYcPoiIA8DodlfJ7JNmrkgUp9PJ/QQ8H6pVhkWsb/6luUXoaXrBKbNUpF
La1mZVpnpUAYBCzMhqEzIxzMgg+LG+YPxZCz7VU0gPhvfH/3KXGFGELuwbaNoCarcF0zr4zwyNu2
Si6XvtDyJUDW2VlpV/Wvn4jVYhtAUsIOt1jNXratZi+Og51u+PYN+H1wIJKVTGadEnZAjJd7Xvfa
hP/1qiLO+JBV0jFIxruKwjbdfAe1OfoM4ah/8SGFh1+SlLuUckvTqvUF2njKHzPDdRlfyJ15b7Sf
2joZJ1esf4MvpcDCcR7IbkK17G/fueAkFdMEcFNw7qmtRsN/fyGxH6PRCQt5YDRXIbas8gKLiMzR
puQJyQZ4x8ezlDqTJQTcQN/M+A+VoCDdJVwnxuhp2GFPJUR3t2pbTPiKRbYnkbwxcuRr93zD6mTL
knQAC7daIfQGPh1vlMJQI0WB7vvgUchjlgWePmPvOVybymejHRFZO1aISQsjc/MDhDEZSXwQg9MI
EBh0TsvHWT12CLtyoz4y7rO195w9NoP2w+ZhYQlfYoSAc5QXcZKaM9hyJrZdDD/dR0HRLmvZ5Cwr
DrbQuZDy6162Cfep3bQjRQMGUWrXtdzYDBpkUYJsxpYlr8wxlws5RKbSCNqtr7Swm4cLe/68cxT5
Vy2Kev+XhOvYAyj8Ybs8zhQ9pq4xKr6DvF74HIKD3Qhsu48e/kVNspexw+dl5nWeHyQht1dasChD
ihbUx7yPK4dgMh6baPOnGBfwSBFlblpZajQASg7eQVylkEW/mNl9rLtu3GU/pQM07HDd76sfloGc
n3nvJG3fnRxvSLi2IlV/Yim7/IZN47+O+xAjrc/MBtS//w1ZqDAi9HYnhmT9HJi4/zFTizuLaY1m
FirnetsAyj5sON2xKLcOxx+YDV6t0WXXuQHgd1Wq6rdlEvt44QlazFz+HfbiS0+1jUvzP1dsssz9
znI4V0xaHBpEPNhWMQe5QRcfprDLZsfEt3RLvXEYyZT2akvjOkYt7GnldYSkJLmIaGT3FHJK9fkW
AxkuawPzn41UM30YEUqAyBmd/LcIEI/YWQAy1l1L+TuCGx8C8N7EGwuZv6ClokTC8HNqDDk7t0WX
QnUdjHlysh5yUII/xknbp/vDHyUoiRLSHXsxy2+TeJLHdrZt91AmKgH833sSfuolrYNobX72OY+z
FW3WpHSX6H+esEJpOCcBTJoUTxJMcVhD/Jnw1UAUGTvo+ivLfmu5ZGdBP/E5f2oe5MnF8Uh89XCF
Ml8l97XrhYl3jmNv5Oc441QIcC7v0qRG3A7AIHeFCKufZAvgjioNO5MHHfiOvh1Ar79tdlL1sdnF
ZJnBjxdhOXtjmK/NXtV5wvQnz+5sqybGxZVwghFXC0/7jtkwSYUZPjAs6ttgh1uxasSB4MeWU/v1
OW55DCAqXqAV6QzNbIvz/A1d5DQRyKrZanEeOzu2bjY4g7lMegmSk+kqnmzN4jBjZ0eivbQD/zv+
9uAy4CuIrFmghN6kNtw69mjm6mBn3ywn5V2q7gelgg32ChX/tG3xql6OvfR0BJd0dXpHcFBAskCo
6T+OgHilpTuwgAlt7GBqUGwdbzEvqWUZ6ECqVLcKKnr+GfhOnApVNqB9Kzz4uvACFBBihWcGUjJw
+XK2VHQO8ETTsawDeMkpZYEl2/0siDJDLf1+FDsQ+nnQJtHsmSEarFeepwbiCJvFhZSdaymB8ic3
CJtyyD7psdw+eFYzdPpZnZcd32VWKmUggKHVC9ANbqDk+4LVRqBL0sl3oTOZDEfga2JTQdhKaGZv
yEtB4LO2Fd467jDowEf5q/EQhLvj0HV+EMpH3l8JV7tKIBfd4AdDFr2iWeOyaYGuvQD+xEGG6+wm
VTRIjuYGJsmF4vWZS7FnR+Pfwaiap0D5u913xYW2KcQQn3/kJzSCQnSDkaqj+6fXHwXNfp6Zc1z2
Bdc/sYF1+fbvbZKiuA9//un0LNfuhYwGWfyQSlfmUUUh6jOLB3wFUPT44VF708iG3aTX2z9vDw9L
hrKYuElSEnSyRqvNYMGpG+MeOdZUf+ApTxzk+ttTT5chPYumhZ8DvyaxdXdi2YUITu6brYjxEgW+
63yJpS77y1ycK8ltp9rtHMNWzgr9yJ4W6fv1K9Thkk+Wrpa1SuXGlyk6m07WJGVjbKoudNviEdO+
fzO+g4cV+tCcLs5EzICyskwAEd6RiOFyU7yvuzANJI09A37feGe97wWwimSHcvISbBTz975RC50q
4RfII9sGVRH93UgggHD3zC/jfcbHw9QqP+n+fHehrlfodsaIDOVQPXMleZqESoaptYeUZcSuGR8e
cgiwglGzkFMzZ9QXvQdSR4YQrTaYToR/fv+n21bvDARfIMI96GTZCecFkNg/Zq7odlTUv5EREHMI
zE2cN6c54M9Zj0ZmZ9v+JuAekKtTU0otUWAMJxDEeVHS3gBeEoHHuzgCVMsXPI0YZz8mD25KtwB+
yWz7WKQp5e3pDakkuenzKg+kfhu6xCBQKo6UHrh8znbaPfsQOY8OTOSoU8/jNZimkLelFPggNTd+
vYZBpAHiJp5KiQPUAI7+DX/bg3tMUrj8IN/USp3q8KO/2/fQ4SsfcddhvgHzT114kCr6ESbL23I2
yspjxD61e8mKwbufb/eyKt5/1GbrQMAONB3RSqq0Nw9HZcNRxF/Yx7uA/0p1Ix6TgM9xT4bt/yJk
ff9FIS8oUS7fWIpC1GpdPclKr1tnQQdCswdC52YeakncaX6obyr6grPdOS4O8tl2SUBe/4qzCqVJ
865laFFHAMYa/4vF8X8gE1/f6azHUqTYdj17H8hVANcgzylKenDxnc12Fk2hDPX/evn8AdfxAmcW
+1ncqGWcX+Spuj7XTsno9cx76aA6YR3TNN9nAXZBrhuR5Pc8dBMaotb1WnX8xGXQPyGjb2XQ0xRn
VLUm+Jt6LFaf/3oJX0g0Sd8Yb7hYulUiKiok/YQHDyOFaWSGK+bqoGF/4CQZovOePs0707fG8RX5
zhpC4l0IQ111ArzLmvRc2jyta2WLnbm9nIvB7WoNF/OQVFPI8TiGKhve+FqVVptd2Dln98JiFtkG
ZHZcCPHHoPmao04JfWH4tyIVsdKTgtGggX7T1dEowePaCzGT9kzZi0rB7FPBwz7FSgQqEKeIphMF
fXaqDDsstFRbmSXg+q4ntSt9nXa+QBmw6CrvmlSax8T1V4z/x+3ukEL4ktFz8jcYI4pEwE8+9lZX
lkUrTYiAM2nhtHA9P6O1Lr7SfGlM9IGsL2ktL6P8ahsPb+59tBGued2P2sZL5IGE94wA6dpRFcXi
eS3shOJjG6YBTTt4xegibo5v6YEQI/bUe6yOCtZioZbILdj1QF/HjXuM98cmf9CTuI0aJNGkpe6Y
L+TNIKhGnoJujRsmhiRGqDyKLFgrzvhKMPAha4SmnjCmg3VPnSGsAb1OrH893aNQsssVGyOLwSpf
xDASEG4jgLR5HdMpeSpV2d4KCYln1zsW9PFT3n9fUYZrqaxg0juV6YNxBwkeLUy0UoKTNVIzCtw1
KweUEIWaZps2WSHsj4M9Gj5evRaKit7uo7+Rc8Eht5r4AJzyZyJHrB2SzmLTN/rARLT14edk3Ixd
M30Bl6ZqesJQdGjdzd7i9hnvbU7yRMjjpGjjEnRoVH/Vzfnm0xYsnB4QX939d4pSFOpTux9y4IZl
fpHET8IqD9RfPYYDxLi8pDUNXEp4kUQio8sY/zmBjSVVRIM4bbJnTKdBavEZaN20AphDDYkBp3WJ
mUTv0lKzFdLpXcLO7C9MBEiiFLhiy9Ikc9d7qWiPdlplRYYH3tJ1v0RTvxeiVon+J3k9xQlQGQQm
xjwABzxRPdn6V7ILm8dT5XLmIq2JH/UuDlQK7wbKO2bwvW4YQb9QlNiQlU/001/v+52yJAdxFj/K
p4Si/czRg1U61j3GoFGL4gj5n3HLr7bcCqbtwQhVKPT6cFzLcusgcZPZc9e/CbF2z+Wu0uFSkRsD
vYpL7JoA8MDVsQaMR1kwj3npDgdYslo6YwYo0eZDmdW9Cou8L9ybRDyTCqdLfq4z06jCapD8mz83
Iq1dkKRsmTWp1aN7//0nN+cfNGFLh5jVXlfef0qvtLeHKKmr7oWe3kwgrjCvuDLy7c4bjnNjMaD4
XEbqXOLSFE1k6jSKszR12hDtwia9vvrDEl0pS0M3yXPUZntE3VEBSm/soAyfXdZfCKwZrjLceaHo
f3Zrh5HHrQdz23SfcGPMeSJP4Ik/7ZoxzLeQRt4yuHBUZ9fxdTupBSf+q+Qx3vzUb7eLa/x1zBGK
Un511zJkdX+U4E6M5v2I7qegU6ZbDKkjgIpJj45kpo8I+VBoIfK520OFOwrK/UXwUJ+2SxyZYyG/
V1VUT6iIA4rylbhPF3ciI2obSAtQlDvD68MYXQVlcG+u8bX394e7CfemR5BOeiFAKoQE8NL+3M3R
vz2fqqxZOPp8movOFNr8t/1mPL0z15F/P65576ehP+Dxt6o7MhQPf+guRkYpPjJh2yHWEN5saU/L
vUWSuWcmPeKvhPO1WavFh8Hxyu3JqD1tEjeAW7SP9nXuM+yM+WEsDZcV1cJJ7VKbNz7CxpEVV5uA
4OHjGl27+CMbQ4cupxBLY0SjTYMzo6YgsVjYh4AWl13vsG952qo3OJjNNxTlqe8BInoMAEYSCMyk
1c0L3J2SINQ3bmABWb0aoKR/U+to+GFzlB8MM7FoYGKkJORl0NR74LZGFHQYZUkyH2Hlvlnfrly4
P+1KAMK9c3/eTNDMSZ6zSY0tz/Lybk7iFr8y3cbukHj8kwiBPgBxGX+7UKfzBUew5XusMoz6qAHK
VlBFBjvfRrWvtRQIJq/KWqw0fAjGU+YT16bkbOVcK7h4LNhryhIhvoXnZdypL6dJKsYpPljcXPAd
FjdziVAbeOlaqKRQb5V4mwmeQr4iB6KH5O8olsWs/JLUWDYKAzyaIOC/l8oIRdfxsyj0TcC14bhF
U56mLaiPtRZ9ScI9VJQd8DFj6uJW832v+R9Z8pPbApTuuY7zyMxJBpJv7XbHQOfhluh/JXGEOIJf
B1nEmUEOFPlQb3bE2yU0OXP7kbCVZn1BPBW+yIFenGcQXOc6BRrBlYbt6BhaA/slaApVfJTu6whm
UoA56IhZW1V3pp7MzO3j5josAbPcfO8Z4YSFy74y5R0cMxXsnFLKyt7V937M/zcLYvJfAiL7Ll78
EjpyKCf8Yb7WvGM1lqtnKzAwyxCuIkoVyGq5YNvSsW7NBwRFuRJJZBwexqz4JTMNzWeeO1EDFAFj
G/uiGOlnN2nTsdLpaePo1uEJPS6u+wAPn8vWGjU1Q1mdUvJMRNXIz5+0CGxR6J2QufAQCJK2Zybb
4BQtK57cWz5NEs+JFjb1/6YCm2CNk9iDDp/NAqe/5FjD/iPbKPtpjPbfdQM/qllIkzvIBct+AKX3
knFAUVjV9dMSwApQPV+F4QqwZexW8O3nzYMfXnerisueOB1tQUA94NW0rQUDaKHwX2BTdcIvmFq2
fADxjMt1DxIkHC96k4T/zZZT+ioPV6HC2xoatC9PUlsyh+Ct5MJVY1o14pe4g8y2ugmPp0w0A5eD
NCqOF/2ceSB6jJ74hHc1YK0T7J9U9P+OAj55lCY2jE1/pmQmJkR0fXLMALakh7k0Hu5FUUb/1IJt
z/AVqVjA2ZpfhfBZtSqN2RGpI+/IDB1T5vLBeSSiGcSKZ0ltzL8SUVmU3uCttRemhSl8pDQ1pgkj
31vCc0pWc2P1kayMxFck7eR1arunXNNHuzJmZMvHzkSRso8O0SqfSKv23bp5b1T+1pwZT6EzUCDE
QZO8QD6CxnWbFzg4ExD0e6xWB8cRSjap8JNjX43SIfvU4OtcUJB7VRpkhDJEkNOE3m/TpV/jLr+C
XFIOWjqRkLjnU3tQ35PqhlztZsmhi30Hj4gZgahAmEDj2PikdD6sFdm7FONSaUCgiFNKJIkCuLUU
3W57Ia0yUPlNLSu3dF1OCk0Wle6UQPDzPTUrvO/OJIwvSJiIs5kL8zMQLgI46cVqRS53o1MyHWT3
n5mMuLS55ntRBj66OQHMWtGJjixilAbnkNKj6+9BkJbn5MHYNbDojZ6xuucLmU5WtdxqnWYWaeYu
TZvxMJd2pELjtO3HW03cLE3eLh/9CmQUK9BqMw7Z38uUKfao4IV2+YGCnAzaRpOX/1uCF3Yudz3Z
1ZU/cM8MH/hWqpto/8qRYeZ12qer87txkpUkcsrqGNN5Oi1diE5+GkdvlDvR4bzHSHtPrmGx1yp4
xOPIpK7ZdT01hdyesTtitpG3CHjoTOL7YjZcA6Uxqcdw1ASxK3kAIKivhmLKt/3sRQ83K0s3tgPm
9Eh/2HRHC8pRu1LI4/zBeTeO9SoI6ATImFuoU+vACrOqEIIZlces0KxUFz1BoqwJoCaQHwIPYxj3
4vy94EYXBz0wm8WOcI/sED8gkQncLJU+LYZSL/e9vYhkIT4tkLrcb8SVNb/W0l3APcUJ2XPwa8gx
e1bXLc2Eb8vB01Y6Pf882NQJjlQUEizScgApiwMNVgj2XW7fX9T33UVWezuGixvN2kU+NXVsiugt
bIT+PpNiz8mbkOM1hgE5MvyVahOl+5lyX3LLREfTcMbYBoT2zLCJCCouFlMrQop071lALec2Q4cr
TwPJapY/RZqUIMO2abKtmp1PeTVwj9AZrc9o5jU0Yyk+YqgrQtael6Qpei5wR9xRdBVqrYbDIqBe
2DjXEDbGKbhrOIl/YImqHnTNA6jmDxisvySa/mzOf8VYSNrm5FblOC0HgbAHfhCtBRRvmHqSWHWc
GQ1zAE1n+rgCOSLQBdd6k2oE1xZ2X3gZQW0ZiXkoA65FDCR6ycrDKnJCWPMnmHFMK/zlERJTUvWS
a7E7+Tqku48weyxt8bDzcYPAUer/8dD5YjE2e3z618fJnzMOTRfuT4AwXyUMpbTBZsxuFVvCuQOB
7DJp7rH8IiuX4p0allyc7mHYoeOfeUKQ6JnODSDK+jbpgZgkGnbYSPEYcvQg1FIYYeg9ZwkCSv4P
1W+0YTVqSUyQ0CuxBXPGbTPYvR/33XrOIe7PdpHjQCW+GHD63BLIjY9Jr2UHcDJFO0P8B5+D2ozd
KpW5E0qeAZqzNgBPeM0an+fZrrpUtkBQGHeKBAg5VHFZlyQalIHQR10YDndWRSNs6DLLnq3ZuvfZ
SO1sV0EMvsUyIJBmM+b3ncpHlgDMskkLxTSPjEcBZ3D/3IiwKYRG7KyrVyuDQyKisCmbnrIyK23o
cr4AWfg8vHKRB6Zdowtpwr4bx8XKDgZpMNXD9uGhMqMui1Bfh1H/3I1YzOw8oR75u3sCgiEX0NW4
XNh6HD21OTpqbtxWGQQTKpBylAR/IoBDTgpuZCy1ZtYTYOPeAtEe4YzXQXCNpiJTYZAFOhjONIdy
U5j6pwCZuquMwrIy1DpmRK4tiidlJTX0u6oX33fKpsP2gLA+ayGnd7z0PHqZMqH1I2DodYrGgiu6
3kB12oojnOcjIAmPF6PvvSXNNqVkrK6IUoE0yDj6dGg986f15wlE/hWjPB/cc2O/fQNjGnKqg+bl
MrcUA32NN1tbUpRGMsfHLQ9GrztE7qHAYSQvJfWIuZeu6l+I8SOaf8VMRnObTTzznlf4EZvrU6oZ
JBVoMHG9CdWwA2M7v0CxhjOpJzOfAI5pJnUOpbNBb82n2SZWv4ov41oi9okwj6g8kzzozV/P5kbB
luIhFFdKxlq/2KJDNa9umfkC6FCiJVR8q8OTk9k964OZrfNds2Bew4yrdUG1+aQGfBAcR1TnD6iO
+GhfoZ9Mw71qfC3ZyGq90E6v/QKyQyyMkZ26monOb9bHNkFvu4juIoQnaBGeixJkxCi5AtvcOBjt
orRWm1q07CZX3A/679TDTk64YM4YIj8JVlskU2QKIhRnGo8Ubzd8XQknc/Y5+tjMW3eqpsyWImv5
7O32XEQBsOiD/wu6hblxWH+obHd9NGxrJJILqXO+d6qeyMLFhOgA3SEAvVTVCm2BWFJEyjShkj5I
O52/fkjmZJpfp5ZA8QAYHhgg5tGzOE2PadXjwWbjYAn5V0MdtlqJN07/eeJKHSgSgWf8Ju1QWQjE
ZXIHXnDseZU01q0GXeMtY/xBPbJkS0vb8f6HR2YiAvAQezOSSk/1udwwLPz9uHPCQJpzZG0Uh7Et
kYL+OLUy7FhU6BhP19JY/x43DHWBqVs+PTDWjMgmz+p/govC1pWylN7RipB+Q2TjZLk5wrH6V7EG
gKfwxEI6Rt8s+hpPsWZRUzo1rdGIsgaLKcYCJP00M12D6AZYW1HUW9HQ/cJmiR/P1dBOnyne81XW
yIoL/vmlktXOej+EviCtVMCk+IzqC0u5tnlZwVYCRDlTm22wSpoG/IGs7CLkjkm29uyouMnESZk2
ZodIbygx55sR6AkRmWZZwhYB3+sDJtK/6bDb4myYv6HMeeoiXUWF1dO2pE91ztQA5tgHU3FSBt6w
ohoIXU4Z/NfNOnd8YKnP0QFckTUv6X410A3Dtln3InkwI88q4+dEF8JATHAFQjV28BxGYwgyMay9
AtPfA9J8GafRh0JDfvoBrkh+XtlY2veEmOoc4R2FF0KrZk5++vIu8XAL1OA93GoM4pnxOFhClgTh
KbIHuEBR8x6A+LHH21dD9A9CP2G1pvMamDZsqBG3RI002wLMmz+U7ftjrjcaTaf7h8ckznV4aTks
EAb+SeKsJwm1OMvdjlatv7JKQ7O2a9KyCj47OgF6XjqkTCcPYxUf88MyVKjPeNpUm++GOggOFm7L
4AFA/XpVopcIGOLxD0Qgqh9DVoslVTjn4PRnMaTH1SCrENUGDk/+rUXzPzJCKMPzBLWe0JKvTE/n
qRWe7d9GUIkmr0pTh84e0v3mxs4qLKHddfyjLF8UJ2Vj6MZUlhNSYlY+Iv6h4TLFAqoY+rt9+jLq
IBUp8QqPTVcnr8GYnQPfEKuWU4jsR4939nkq5EgVJ5TpSrI8giWDAv34jqKZ/JsZE764ynWpUPwG
ZxzgMOSx9U41br9v9PrWET82jxsG/2SLNw7+XmeNQOw2W+oBkHQnwMFYpZAY7u9KkGki6IWpPCxx
HoO+pLGVcMfnxQVx1PPLJbagtZbz+RulmuQWG+dV3YHn861Zqc1UQzjP6Rlx2N8RTiNT6Fk9XMC5
w9TyyLta9v51VhVB3f8/5f1pEqG5nFhGaIMqPL0rdCKX94P9WwL3HdxrXpf8ZSZP0FIkLKO/mdJQ
PTm7rFGiQFrPD0nwAGaQt6Tk/c2qFAz5Z4RI4PEkS1UmKDKvAQpB3ouELYv2PrH0Au+wwh0JcCtu
RbzD/IIeMS/kJdwJCF3rKCWHEFI8ehfe4w4VNGxieF+L46zMPi8WTxNTN954Q2xASqfN58lAOpg8
qlAipodYZLTqHUGB+0AqBzpqnnAKFzWhIzlcPCmZML1YqjNZ4S9hbz7GS64JNcqUq0AyZBckYGYy
OzW40fFvQ1culaZ+xRpwPctk6SOjiSHmU8yUIw6HrtexL6YGNpljhV3C5WXJSwCxtBbmmF0mn/p9
mtorvPBQSpF6gjD19IQyk+9mFdjSB2zk8Q/wgfewmPwL/xDwbx6O8n11kvdZlkxLYaWVYlUl/Dur
Cm75ZWTl7w4cKL3lnVUf1v1mJWYrG7OeVGWnsX7gOHkuKW9lW7oaFmSuz07pdJLVxElJeb55e82w
SMgH//VNpe1gPRcwBl9R8xqj1TrutL/jSxNiZcBYg19nPt4Mx/+r/IIy/92dqzM4bwduN3V5+/GA
Hf66XLrIaw2vNPi9k8FdAOlkrp9tMY32H+vU/Ue9YNyFUdrrYljOfOIn40GdaK5tPH7mcSMjJJSl
JcVu8EmAqVkyxSOsF7/YUHdaNEWxjWeBO1Ifrs5uaB/alJiDIT50rXFpLwr9ReN+OJUTyg1kDy+e
/EtaQI8oxgPSTtqILQ0kBkrkhlDw3r+Me+HKYwjevCGdjzUuU9/KxEIqGAEoAFsd3W67rR8jspRr
LgDnJwGWz5YTwEModOQC7siJBKSvve+lhmFC5NGOBQf66TsYoDClCM4WmtFt64CYfSG86YdFIuZg
QrRoxpUMxLPk/nzvAVDytBPg2O72vBtU/EQDvoI5KMCreScE38ocgfBg8ADAf0llxEi+2f7q54Er
o4oegU6yBOZyYPI4tZRQ/t2b/azGn13by5uHruLrAfyCYXTiw2vACaak6W0xAIsaxnhuaFDyARPH
khAQTo9EYJR9dyRnTk32aCCcq5ETyO6Wb6pcdbe2cEw7gZ/Uaovwp9eNXA9rMyLB1cEVLsDE8Npr
AcqAtJ5QY1a3Jqa8Tl6X52WfFjTF/bIDsdvk5Rf+zulrB83YKNdjtAq0np+ScaKGlNvdhugHBJz4
bEIoF0SXqM55ncd6QWqZ3tRAcS1AXhnQufP7ZIy4nmafaO85D0GwLQDkLq4B9wMDoLkQTlPbOeH1
+FBNeF227J/HlKRwRtIv6c/zdHP8yG8NbKuCBv/oLRu5tV4TY0PzwZKX1C0B6xX5o7YwSyp4pt4V
Y5LQQcPC0zNCaBzNzQd0lrQZk8lTJLqfApBrDSHyWhResE3KCRi50YSUN2kWGybmi9tcoNCCamb0
k6p+FGLq/Jnvkrezrun3K/lOsgkBun1+4UjqSYEYcJzm88HPPPbhQSyJKkz4fHTo9JUINc+VILyB
0OQTNCPf6MEHsmwRaYb8XxzjJ6hRVWoCPP0tGN5NRVKncpDgXrVR0megbmvn0sojKU4fApzoL0Vn
A7zpupvxpD6btnTHWtIFrnYxgUDhPpejJ1Y3Y74MY5DBtqVMpTeBq6vJbGpSjKX0XjLjc8andwiv
GgmT+W8xZBxSXUd2YwM8GkzEyIKzwNOwGbWwLr0cFHX4NWVuTToryifLoBKNL2jvW6cwlPZn8s1Y
z785NoIr7keP2Pb/l98ZAFUzd5hu2Vk2e3a88N5eesOIUkmpMIStuBJidinwefl0vWnad7yqzq1Z
msvytRW22LezxdxRW+kBTP/2t/bW1n+45eBKeByEDb96xvfWySrMkvcRNeUGyvApzUBFBKMhuVH0
HK0RByfNzw1BAkOCnIcyhDuOPBceuremrNIQpYSWfRuwwRGgEjKRT1YJ0z5gwUVywpIBJa2EN/IQ
CPqCGhlyeob/f4hU8lR32gv4mYeEgn6tIT2xJWmSCanDS4ICfPXueZO++Bqsexgj11QhFcREL5ky
DL4W9t0C1CYn98RWrPuqtAWFg95cQm0cw7/6JEERsdMl/g2AO0a6XR0MeFFF4gSKQoPeZ1RwfQN1
9uss7IfLtMCxdXiU7VBmbJWNB4wlGBfWvHyazMcD3FmM4YKq/MKayxmzAR1bdz2xWW75xmg+amjR
cyjWot5aw+XGtRkhT/XE/1w+fItx+04hj0C8ZcayTLRc0eqCa5RFmfcM1jlBagItHsx6kU6fDdIp
rZ3a4eBu1bNBTb+mtG9W3z934/rEZYeGdVGN4TZ2T6+oTW3HEfGozYzBIMiCefD/N0yhqbyQa/Kd
rsCGXw7y7QhqPQMzYAtA6lkrYZYOYsh4/+f1UIdJNk4W/VwIO38g9yM0RiPsDJBmmWQWmvT1jT51
kkVkTQrneEdxLWHjhdSOKkaHAu/M5cH+Wuv+1nfUaAbZMsDExYlqgA53421RduFveQNzGM4Twv70
fw9CIdoOV2i+/ryL7fGDVjWRkg3gMEMke6bqe6l+gYCuqqdrXRRt2hwG+W0K2AqmUqgedGNmTUbL
cxYWG1JNY9w6psM90IHrFoVKphsaiW62iBNq+VTiDAtGSsBhSxcgFIl5EF3TBSyt10nomo8jcaLF
s/+jCDvKjPrRCtpyjPVXtTXYnkqXXWFI8sn72aeyrMzxV4K0pjmOoHvUjbNJkdFqbMtuhVrM8Y64
EWHKFCVpEQ5wHENMLdKIEqraVtXkCtMJLCZuRMWHDzA09Tf0sEVKUQij83K5RJn5BmEXO7IuuNAM
e8L/95jF+GtKZUekx3t+4PPRva4HekopRPgFHhKs/RCtSpzNLc0ZQ7CAm1UuW5YqcFiFKLYKUT22
WaFj4J5T6v7cfcPdIu4VJhf8eHdrCg7K/cminN3pXXmj8YqAHCultirDBqIetoCsHBP0Jpsh9Q72
zHo+xhXUmaOeY0ZpkospPC33ClLMtIlhK767etxATcESDy/qmDpegnaoBobnkWbH8PlTqdbONjau
u3Ty9uQ4tn7DFc+iq+DpASEpEKGGhJtPtOIzjaRHVxEdQHuGH/Y+8Tvpm2NpLrEVDhV+Kj69naFY
fn/TlTqB4QZ3tNL+RvIbTMCszciLJggsLepLzRl2jTKdSC33+Siwu1VK1XYD+foKco70JlhHbh1t
dK8Y5rvZPURu7lxCLn7lBEj6R0jxyZkWhLVZ1MmesRrqv7XiHQGQ6cjgJiUNDF/fJKt1Y9Wy1vzz
FO24PlkGCqY5sURaHxHK9WjFjjOSHJvvLh1q9PxNKIGhljOSmNvyZSc+ORJ4D/rv6PS/wN8pPBrW
CuSo0tt9IgeX7UzL1pSGFa8kaHMCxEw5VeXfx3IU1mxD5V+PWFYuS2wpKSJfQoRFLobqQNPPuRb7
EEAYizq9TIGvMGq74ls2aQ72hbB7fNQN92ktAXXidj8TA6dz9xj5USLVNl9OwRL+9szBzBN2aiVW
hfMFZM9Ha1QkoUufcwVG+Cy1HJNa+x8MdXpe3fl/sBkzmDSVmvm0hrwPO333VZ0jTpuGO6pi5aKv
Cs/7rHEiFw/iuW/mRvhiyHFCW4rlDBCGcMkAz600RQ5qkT+KiWRxV5IpCufxxxI8cZ7ynNKp/oiw
uXP4vvnUW5wAY2WzjTaMWhosRKU3lep8HZnIJtyhPZa8F6njxlY84t7eBHJ+0tZLrBG1ivLqQNE4
3Dd/mozmfzJO7UzHgTsm3Fa38a6qTaj/4EnCYW7g0GbaeymboF/wmTGHb/IplHBbw2kzzbFrIQ28
w+x3QWLZZOR6k2GY76W4We5KR6TKyBu3Urr79iYirGgND55gAC3SDb90PZNeBYE4xmqu8qwJNOWe
lss9qw571lE16CFBbPb9nxvbvkBDrg/4ZLGr2+Lr4X6O/NRBJDTvMx9V+vb3w856ltzQ0/YNyXBd
IBrDkgMS7ErDN0VLv5LqyG5tvtO+4VcQuW/tqPXKfTHumsGOdGOlEi3yNbY8Ni3En/VMqDyrGVAE
3c/08TZWEYpdGEytM1yI4+sTdezsRO3sxYxkP870snU+6PALnsSW+oK3jHQXMl1dT5dh8WDGtCeG
wJWVNiiMXJA3R7tzsFVyFCZoomfDxRaMfBY0XtOvD9g/EyxClTwWxzlOzWx3Qh+rX+iB1d+06YZ8
ZvxVvM5B7ccSW7cbFrgVMWckDpHIv+tOYmT/5xl4HRWwDWdVkUDwJ+zigK3eBK1DgHAMWxDgtyxF
3143nzgqchza1+RdugkW/itqC4cDLkrwwZss+BPxCS/J401mLIqToDRqkzh7Latq3rsL9VBnPEbR
JEW6WevR56ToCu5BdwJhiY6ON3Uhe79QM4SOJsKU2lxRxDQQHwXMjR3iTo1x79GSQPopO6DZBJ5o
NYvKK8zL1XwYp2+UdYG44Go8TzayU/pHuhVgbvmXuDWOSvfZRpBtYFsX4IJEKLb/o2Fi2HlxsAa5
/49sTMY6bNILmnefO6WB/qrF4/i52LeC97p1MYLHMdGisxTARq1yI9NQeAVH97PCZBwJfleO94EA
q+fUBNnjW2wez88XWtALZ6RXBIq27oBoElLt3Ac0Q/vmjNW5dX6IKYK6ecwD7wrgP0SsocbUxLxF
E599d/R6DGnX5TP3wAekVoEI2Vb/SPxg6ZKPKTCWNPsIFVPtn/XDKgv+RyV8wfcxoxYsyoN1PWXE
VZ0bMCisGXpoxj7SVB28kSeinml4il80RlCHoB/xH5zWccktHEw18cLE4Dt+s8DxFKis4zfrMeuT
za74u9gNqUVe6l/C3Pkb/kB4N2y+iw9MupEi1zxPF/NiHosHMtQnUM10pnpFkb7BpCuM+v69cimF
YJB4YLe9YMK6KtPut9jIqW3ZNyeNtaw20YcOJicDCB1pz27q/dutsiMuvgsLLHen5ZTON2ZlVTsL
TXnQ7ZpIj3ub5H4jO1HDlu5ZCBKU3DJUaY9Wy/Nq5NnVQBXDpJGWC2i7T9Z7n0KI7eYfSr8cvwYH
0hFUEQDVz1J+m4ThLzwFGnSpEir0GC49NXnQDYWAeO22LqyoCSVTE54WDZJ9kgHTJpehJjUE/OVf
mWN0FRpuS8OFa3O3PPNCVwDpIqPLL73wWUJtTHoD9g+bDtboUrkqsgqqPoAVnsF5JK1GLW5K02kh
v4OkVwRi6wB6WQzodaUcZqLutksbMR/SK0K5EjABrxBeNu1uUEBr0HV6U2pbVjTJK4LgQKGdhUKi
QKAkd7K/IZXQBef5ByuxE9+zzNFuvhnoipusyq061uEgM3c8JJ8QxiyWw2qUnC7nONuzeDjIpeMH
K8mV8a5TpI9fIXOU5jM4K6tweqn+lKEoaQmzJGwzs+tveHsJ9QdsWCWtC77VFoPKIQqjcPbA+aAd
pugJFEDKUBQ1Z+PrFDg8Vz/3LBQa5h0gX4cJepfW95a34IWTd2U2yB5tn+pqL5GDVf9tivEKg6ty
djqvsEe63op7BKYHLgNUcW9aYFf4PwgkdJxPl4X0calbXySgmhcPXslW8TrdFbPJVgFHu8sTkZYT
U7dM157USUuiY4VVtmbcjSUmmLto+NiwpeXzkOs1Xz2xCt6+DacYz2QNZdh+lB3LVNSFbZViqlgb
FgwBmXFa+tt4VzAG2z7Eh9y/gYXtq0bhnW6lR/gT+eKBFUAvgQofikQJ+1cy+CnGjqj3VVyqOXGh
j1GEgZZtTU2kxc1IBbVNFsNSNhndt8hGqANCgV5pG7YHdzerI8Ftf9aS6EOm8X9EFbhit+rh5JEM
C/ruTwYteAPLMq2n6uSFwTbfNfT6bLFw7jX+PG1F5hr4DQY9p8vtRUGVE80SpZ9d7ylUKbspoG9y
BnVyR1igvuWHRLvVtTKGZbBm+zROKgQIzg6ep6bctv0LeUY8sG+Tj9uWMJXTh97lGxKphwuiAZxa
cvbNl8BSHEnx5v3b+H2LIqiL8bdw1P3kRrCEspmp2Cy/GYHrNaiY2pHT1lY4Ffg3uMAjNY28+qdY
0RCiEmpot7bSuDGX3MQsmq4SSzIhKrEIFi+2ZCNpSDo4NPcZbiyXt6BsfJq8zx7AzIUpAqOd3UDb
uHw9QurT9LEqBEII+oL532Kqhpo3LNvgJGYyfHHprTkQgjOzHRQyR6IcqjGF1x3ANbpRBVPRB/VI
WWi625/Helqfm+K54usH2HZE7xyd7dQ3pdZPQtUot1p9c25iXM7L6TzUSbLrIvnwRhFWFnra5/Fd
wBPO2y4i/oDratTCUBfixT67sCnreG51R7Z3Pghayb+KXZ8IbihuP67t6neW7AwHNN3HWHbVFgG9
TAIoRxsneqwHinJv01/gYAz7I0uNrGTiaB95P3pt6BGpIED1JmlVS6LpCkaJimhriEfyjwPzHLz1
oxO7gDcS0tQ3IRgAL8tU2oPT0yxaLigzhopLXs4yEwiHvMaiLdM4X9yDyo5IIcuYpWYLMfcQ4997
FUaMQelanEtstfQnu+7tbpmfcvxQrL8gv9E74g4FhUgA/DCYwV2k8g8mjKY0pkViUZnfC8YbbZfE
chY2wsO67wOM0fhdOGmog32D0vi6kQ9ziI3629Bd6UfbDEsmidq+SPWs5GCv/ft8hWFYqiRDw2nd
1g6me9Q6o2HhBw/umlTQ075BTtBNKWEbBl3pc5NVi2CRfwCop6uRKDDWtlWdMmOzkiohJ98DU/8E
lcTLNECKt8mPjfdOLXgAPmbz1dITz72wAsiykDPzjCkP9TfudLAT0gb0gdmx+/YKq0q3XASu2xPu
11N7Fh+49/TUukFh2DKszzyUOY2QsM9l0JKquJuIG27Qts1xTclvYtKzDq+35mTooY5Q5QxeEksA
GwQOyuB2Fo9/uULZ/863SncBey9uEKICaJ/igroOBvenoMe3TSmGaMdzknlTJHZ2/U8vWntl2mjT
NzUHF2FT0u9nsBLXHHfDM3+jDb8TgQApzaRzMZKW+bEv7JMZUK4zCp55vhqhfqPr3YvqzVZaQ8is
2oecWCeNrCq91WE0xYek9s/sMNBHc7tHjvXOy4bgbyjcwop7BR6ZH2A0iypn70/8ojfHXNkcFrUI
2rmSeX2vt27T3rP5+KKNk00dph744ZePr338y7/ScSYvhLjKMXQggvMRbzAafDOW7LrYA9qB+GDl
2V8n9q3Bfx/np6huMrlNteOQXoVzPXGQC6LbyFfk5/oBanfZ1vwSOuuWMYU0e6mwLxqlBgHDhski
/fsOMXzjnq/2Eok1koaMQ7ChtI4nf7E6MnW5aG7roud9t/lWvCuoh4uWgFT2YTm/Ezb/xIEr760+
rXFr7agc2y2a3LItD/yYfglCbxeqLCwuT99WCNtBkF+VIR9KIXbFyrvNULw51ZS0docXxKN/zhgc
zoLmTUcx6oNGlR2rjIw4CYDj1KmFGJblbyBYkKyBNYJkwVcW0w5k1TKcUAYpKQiS3wSaLcdeX67O
1Qz2uwpS5+aECJW0IYzmXPLYHlg3KHKMQmgcvbCMHiSgBpqfF/5YE3BbAh40s7zyAnbolcoXdVz1
ra3e1dpuSFp25kOa5SaHqNj7M2cooJDNxD5bQwDQWmrB4YODluybhji34uILvgq0JlNM8PE1y2UF
xLoHoaGagwlQ12lXVg6HorQ+mljaovGdwv7u/EfXMxrD4zQQfm8iBTbx9tyxY2WDItQgGHfDbx+N
uaqFxO8MCjFooBF5b3Sj0fxFt04s7vAStnE1ZKBTIwkUDdAlFP+f8pSmoXt1e7ODdjAu2tcQNc5b
bZ4dqTmAza4wNdHPeLnVd2U0YCFrQ+25a7L7lTDEjHoECaAePr3wRv3aqOlKl9gZpgiF/+LLSxP5
VpBe1cCyGm0YtvsfQWJ8YIpU2vRgqDwScpJ3rLYVRD2U46OIDjIDlvnfADkaXPgI5nu9EnrsttLC
zX5Jh/7ioYl4BnmpHuUxLgjkVeJN5Or5HkSNH/JuRxZrfXxfRyfL1FkoIEB8PtdIgvwLSI/0ukAg
ewSjFwDF5nc2r6xSvhCn+pUCtzYDIMCp4VEw//45yCJXkyOMLV/TMPSv2ENrbJTdVQmKCnEgxeyM
zONI5tb6ep5enFcfWaN8pFAPFDY0R68IMbEmS2cicSeJRBYFVmj2aQyXTyVAHziyuEbLbNZDuXRm
pZ3K7GgnadsfVAoYWGQsCP1o9iwImU4WvRzG+A5cKwPN5kDFZiVQz7iO9HGLxPDZT6QX9zt3hFYW
B2Hj9KMlSoycxAR7hTItjW15yTddmZl9RzcGnogKfATzZGmSP3Nkk4b+qFQwihPQ2FmAxrvVFUZQ
yn96bpK23v0XyB4hmadB0DxS6KsMbVDRdX5PyPEpb4qVe8ANCQ1EEwC1JtjrevBxDd3cVKvxZ8Ev
vmnnD0no9nczehtFFGvS8tkNYc0HRHGo59Lz1YvU6weYqhUSoopeEsBa5WGOEN8Nj76I+qCkiz4n
/wSvm9FD4FXFybC6RT6vgW61dw0YQ/XKSFIe/bHjnn764ru5QGSus2akZ7TkMx9k/5BnL1SscXB4
nWyvx0SuGl6CrnXbA3ETyjHS7gCU2tgY4LQE3dsD/aTgItrHNF88irBmOLcHGWWvfnZNUG59bOnc
Ac63RWsg0WoNaq9jqVbmHb3ynIeK82k2kSKn01h/aYKHKQHBBhKAx0WXq4SUekUWLBR2ocLWW/aq
Trp/yo75nz0juYdn1Vam7uIXTxdg2Wuzky5wTIQUN6eIwE3rw0pUg3upe07RJDJ1D1ZT+kNDgRws
xip6CGH++vBmqfEa3n8Jb/JNmQoniORCGs81F7RnrO5bTyY3jYH2UsRINdJ51++3/QkDfBM1cCnL
xFOh1IzPPa8YFYYE5hjrUqTIDKgAvwgORz52kR40/GABb7lK4tMx/9uHNIklCxWtYQKeX9Ih3SoW
4d/dFVJmMAUEl89LD0T7/9OBc90dK7d/LCxSQ+UJAauZVwmnFEeMq6YZEdFyARNjAZFWmG6Ee+DJ
RhfH5zLvuo80Rdh/T3xIpRHo4Azv4dCYf6mLu9NC/m4RbV0bl4Dats81lQ177+/lF9XVh+IGrHqx
eoeFcldN4V9U2GtZPB7IsWmPY2mbHJY2KQlOwJ2/vb9RFCZEnnouOqsxSFjDqwga71pcYvW4c6uJ
+xwYcZe8GwyTQqJDmqRJPM7V0pFrf2Mmxca85ggxseQAPW1TvFukQfps4v14rC912/UVD+ofIzaT
x0ipBhAL5HF5fzUA1sUg1HXzWMR63bDQkwAMGs5f/mtlT3i+XWAvzdewM4Vhc7uNxjLd1JKEa2r6
Ixb+4vHv/5oSKRRuXH5mrLpwXTi7wYGxwCzl1b+M6zBlLfRfyz3uqu+znFDeK793YHFZFYaoxa9T
Z5IvGJSF9VJP2dRliCCjt46Lb2Zkn9FHorZXBM7mg7eiggQKkzkxFx8zGese06atPkfijum9N8Vz
hChEXXxcWSu195wXVOsGzGICw1R0oi2cd6N9KqcjgWdGWQS/Dy2DhmelzVnWxoc/v0v+Ba5AQWAk
17eRDjNeL5gJx3NTuRq7fT4kWlKaebdLANNc8sBXMBJ7g5XtHZPks8MxA01tIBn7fnK4zn1bMcfO
/xLiP6LfZVgOBytfwRYF17nZMGcbhPNDV4+Qx9kHN0tWyZWK7BYjEImeY9yIs5nfcKCzNbq/cPJx
cxJT+hEQyfvcBPtG8gk6rZtri4anFu4dFY0lr/cuYuvxPB2jnA/dUD36gQu8/B5KrjYJb1igiM2A
tYR+rC+R+1mKX1TfRyoV1xeGE4MK2iWPL+tQG6OyxYd3RwyHHjn33Ca9Ckq7o6kwaYTTly120Xxi
29kP0Xvqpstym8HLeH4ixeRbUM6inVAVEG9NloIbUkdAV/Lfsq6lbCAt3Behq0z6157xz42MT6Bu
WVpMI2Gq9ylMX/ns3RmMbF+Ms+ZfkhwcBejD4wKbnog8k1oZnIe4NDi3zaa2C/CwJx9KTuCBwpnW
xxxidtTjkPqPVdXnB28mmdfd5AhRcBt7Ajfcm40tTPsMR26frSPJWbr0Sfbp2hgYn3vvvbZTFAlx
6/H1BO3k0IU4YjxTpKfs9To28O2H3vfZ/WMRy9yDuM52WaOXH8dR2iyZnOf4RSgP6WmiHng4uQ5S
rvEpQGzGRBFyvJMv/YZm+mpMsL1Pen2R32jhIL7Fcadmmo3NL+OrbvzCxj4OP9hcm7BFTr+HRYQR
pxpWtCQPzDxm0uPzt+9IUdBwlTNiqwOjrLAzBiiswnpdV1P31KuYrkloORL4DfwupADOvbxtFNll
kDfVGPQYmaDnLpz9izJ4AAu+/yikWbZ1Nzm7fgofXno6/Sin7vEv/eWVEr2sGAcJAkukHJQXbDnh
1DmtSoe4mR0YeRxDXHpqJIiCpHxItDtJ6BQD6MmVG4zGQ3v7jjYTDio4ufYZPqaZGH04CQ//Nu63
6EN8BudtiPVfprUDa3waQUCDaPFF8eMZ3QT73gNoHGvz0ZwtgqQH7G9/cGm3q/bIcGnhmOJ5BQu7
dq01fLHDAWU+6DWyxkxMdXeoqWgFBa75VEk4qF4GyVznoe0UbdigPBpG7/44R7DDcCQyU8NdKJGA
ZDAk+sZ4hqsTAh27Q6sLIjTOhjWOHyx3I34417yaMZwSrA8rzgS7YEYZKWj/BWFvcQTFX+UGuKSx
cO8w/gdzERU3Q22O8c0MR/uE7WD8wvVJPLaP7bbGvz58G2JowrZ1miL8BwNfP/DHoWD5z7e6d6s8
RFjh1j4w1hIuenj3K7wHtsfmwfDS9ovnctCdDmW8rLXRD01QnCTFMAFNYB/R7tJfdBb7uNw85jid
6pfuucYQxZ9xrFMo6fAppeekXh+d1pjmR7xM67pD0oy6zOTnRu2TTqFD8irpceNszw9tgLjY+xtC
v2gC3Rwv9yi0Y4fG/0pK7gaCo8naWAr12sTmFRW3/YSSAspr5Wok4NH3N7VdDihGR0pqqW7LcOFK
esi+/XmAhe1iVNj7Fn3t2OlXDiR3/4DtKOCxkcA4JKWawpR823ov8t+I58P9Qtk9ETbMQRzoAXxZ
hi52EIrMajW68V0n1bRCUwWb3dWT/mzJAY/DDI3WRSq7KBv1bo2ahLsxodIgLlNDCw9Jq3rSToTw
B/AnO3DsXL2Fgl+Sv0dbVZ0F0vI4bwoNhDww3JBa/6zErHYySnNBfDuodpMXKwFmsVZ2ojF6GuCn
pm1R5C6uF/uyRj5ppYatkFpPMJHQNmOskS1muBynEb6oNO1s6G1wlYr1XYyWFgiAclcGB9ObiocH
69TMyH1Xp3PFoW4eK+07UKnplTZfOnLdEUzolxmcmuj2xqQeoLsvAVFtCLER7FnnoHRwoUIyl6xJ
Um4aDNsyqsO3eQlxRJd8knvtbEAr/F3AqMS9gByg3qgtFRe0jvX8OW3GiY9tEiatPcfVt7CsV2Hx
ZRqArNGXl1VGKc+ME9EtNe9Fiwmm3PS157b+r3WiWfQflJ/M5QBwt4lDvX8Dk4Ev06aIs4lACvrL
bdjwqW4ZCIZ5+12qoh/IEbhsDo5+X2BEZOUfzjyoDx3pOmKnjDCWKJP4EMhIpWscocCPOcK4y1f8
lKrxJdChA3av6d7e0XjookrgBarST9BhcYMNXirnQB5xzFEr4AjX6EO08z9KQtd1GuBCKDbn4uZ+
iu2f6JIxx3vFvsfLhGeBXrGTmSJKMqCWkS+P1SatefQl/Hgum43YiCE2zOpZsAUWNnKExk/lZSe+
cCLtOVe2PV0jGkf/zuwrqEG3LJt25QDstccIpg/Jv+ccBX/X+laucocw8EOsB+ZSEQq2rEwFa+XQ
VbRM4Bz3tcJ0MvbMoAIzTI4et1CNU+0XMwNVihc8dopA2RdLW8shdCdj1qNKaiwcDFvi0/qIhHla
YmQbCdsEJPGSeM10W+g/0fTSoq7cXH6GJQIhEMFW2AhdDQYdMDViC/7PJv9aOFwvvGxHDoqYBEkV
ZobbtGivYFwQSuVDG8KtCHUI0oFgO/BDIMepmf29JDFLOjSFvRqQXakD+cBQWUBievQcPA+wQmFb
q40vs3ZQX9A6udEpLg9ac1844iccs4M+aSwmPMDgninLEMHr6wDbxWaAyHsaVDUtYLjjgkIG7uRu
LPRh8AaIe4EURvazreiRHc8Zz6XnTFDYpZZlj6aj/N7Vb9+04MRI+YRVVtoiwO/YfOMt9Ze1nJ9E
+ntQnF2u7uJGd3zVgV+WtAJjp2mLI9PGTdosHKfhRPuoTJgNblaTOb3iMuUtBuZXo1tEmaOcULvW
bGrF8hpb5Z8+LlKj+2u9oc8TnljfB57pb3KAO0LtzrbHHPYwBD0YnSpHUiHCqsVZLtGVt8/VDUqb
VEYLf9Mz0mB9n1lZhuDDRm4TCVwmXPzkc0mwhlYlBfwJXUeRl1M48y93L8hZGkS9gByul8NOYHK9
5mL5oCiz44pJwMh4dv6MqSwDpgZeaq0x/C0UDRWEr11mqPT0b0Y16pZiUAlTcjGMwzigNXF5aDJl
Mhwv/Qg3CvWsikhNF9mqAeFKjzqpruN11/GtAVXgqu9N1F6qY6O9Buy9TDZyJsbdQRF9Fke9ao4S
s5+eeBnGbB1GU5uBkYfADDd5RZt73b9a5+ZbaB00c40hG/oI/UUrcUrNpNe/+jmOcc7f7oqVjAHk
JGyHPXwPM1gLrEsiLWT+YYy28gsXBZjoLjOJBxncPCLRHV4kZh9bXRLgB7JHDV9wL4LkDwKxM2AO
0qYKJWZapwzGt9YQg+5vhX7BXDMmvlJKY//B/wezCXCQAqKHN3t0fuOdWFnc5Sbr/I0cuAcYHq0t
vRSDQyA2I9XZxJSXje33l3Q92DLLcuTtLu7Il2W785c2ifiNjaYJOAdDcgK0gN3r2BZ/1UWbqpRp
gbtOFnLFfy/jsqW80XZ1kWfkQgLb8X/9Beo7Zn2eAY+7gsNK0899XKu3MPu5quXmVBkiRCMomOUY
edK/fP3abDP3ZQElwwbNMbVKB/Nvv7IoRQj47THqj122j9L9ayCAb3meHLw4a8M+LFRVs6JAcbbn
pvtboKs7uinYF1ZtKyKzZhK4CNtbe5JVE7K2wljFOpqZu50uGWjnF3fpqm5fGtmZAGtK4AGRYzqZ
HGGITsSpNANnE3RrP5iaHNmbDQXYFZz5QyMCQfbM5V2FHmyvQ1iFdu8qLyc1sEcaWYDmwedOv9vH
Y/vEe2Oo6tHNAhmm5lfTtZTmpWqok7zTHbUOhXuNw8d7ziGn786CvVqAe0FIB44dXc27v6yyegOH
A+MTMle7EA4K/hZyts/pwGkuZqyI8qVwq9/92eR5TapGyY5eoK0YpRZYnw8Z9gK6+ETcVSV9kUp0
uJNPMIHe1wY1HVrpLZjHEuze5/7MVEn3ZsH3YSUCCsxjZz629tozRU57FFmw73LQKYuFm0st6OYd
fVzMg8GLUqdCF/deO2hDtFOUx586iBAqONpXYr8dtqoqzrgwZh7+dZ4DgZ9VVxP8gpHkOf/ryKpA
e7QhSBjy0nO5l9atGgPXDpMN8U4ujQvZ1rpSFh0MDQWeMuui9MzK3XcUz66MZAL3p4uvWVrkIA5R
dn//X/8pd8kpGLLX/3UmJ2uF3Xs1gbaBXw8VQz6auBUSOStmrJTG3IqpMZ0n3+ljM0rZoKvN+jS4
utvNaAnwJXbJXpsvVNBCSYw8N3DX9PlHOU7LS5P0sF7Usu4aq8hDLj3DtSuWhFIUGjxrr7CfUoz6
m9D7cLJVZWSSTTqzeQp2LSst6kh/hPU9wVY2YzPgDf2iGIi1dRQ8CerHzTIbaC/2v3L02jKxDDOC
vuZPKjBpVf6DMAWilBPM67YMylCcocWOhtN9NUEq2YwOSsJTbUrjTFNSKiyebJvoQU8xpV6cQBuj
1VLveYiFFSAUXE8TqtYvQyp4MGzowS8fp8Sgy7h6NFqnWWy8ZCvIk6Do4sAoGdYLwiMCk1+yPI8m
XjUIjmZfSf2M+z827rcH57z3Rmje2mcKUNZ8zsKSyvJxs1Zidvyrg31V2mb5Zfh54XHWfdZGlSZJ
zFqZO3b68iVbJp4/lBKZX6s10Vff0gnmvXUUDJAOssSP2c0nvoqJkPqiI9RrfhperkAIG1jmmAZU
xv6yhnpm+ANRDMmdPI902YXufPx6O8SnhGzhVe/onZan4sUADBL/2oVfYVdFO+k2QzoyT431Mvu0
quzICoXkLG+g9l8b0BRyvS2ZdccxrLKNWV2SH6jsLxZItnzTNC5oM+SB0X+t+Dbhr+0PH/x438kf
VD1r4ghs9Dry9unW9UXAd6AMR/ogNvbTyRIUtr54wmMSHgUMaF3Vk1Q4uxuL0ZDppu/6v7nka+W1
uppF/ZXi3mRJDaP3ecvA1gSolGSIOW3wUzzSD4FgDUo/I2d+SkhOugetDSEjqbsYTw2iBXYZKw6G
bYim5AmfTHBk6fbL2KpVK85IxHRmxDFkBOgzD8eJbkSRitLRa1T/e0l8x33/3q9Swcqpofg7ECDl
KsAXRUZmJGBXWsjXzckBw7YYShwHub5qDNd/PkAUOMzb4oAsmm/tjTLaF9E2+NDBhHR2NqFLAese
mAVgqt87dOpNk5xnnID+e0YeZ9ZrC3AvqsPWqM+cj2wqhKRN9hq7XnMgAM9dF1QRziT5s11YZpWT
aODDb0znH0Oru2jpFj8GxVcFmlp0dsDpPfhIhqf0PNHO+R1OZE6zs/gHN6EAZ3JFxvCgCKzy9SeB
flJHV8ZMLprcS8UC+LYOyELx4WMRoRkSDYWRvcOnrjkqgleFOjab1l9nUGI+Gi0U0BR57vkMjVHh
5bse8LiYiQuH3C7PpoaNqf/pSCWi8w5IMbOyGtSBTr9qxNBhptVtPSvnnUZa+rB0EmT+UJEm/PpH
KZoKWcVPGc8ZPFMtGKnhP4iN4At85BzCJRsrqVGssAkXnaYYaA5+SJPf52BPuuzGBOo24rTyN+yX
ouWPotks2vCtdF8k2yp4ywxWwVnpjRDs49cRWZZfpyJMqzPlLHfYxV9OpQ/BJlxCjaURC7RR6sE1
yOyjGkv2Qih0/c+losGRj+yB7sGrKylZA4FjNAlt9AjG9BJTIwD1XJtXiboyRF7OGyya0e7B5XgC
+JUg6LdYrPX/LDWP7AWcOpjRBBP0cCR+4TJgztk1pRWFibr2FpKHX7itUMtkJiqfByJSoj0A/YFb
9JW6NKdX524B31PsZZS2nIr7D436yJopuaFi7acwOgnvqVWyhMiN16tCWboE9tX0k7mhTVzHyWl4
aSBPmDAKt3HFZO2JMUj2umXjTJx/jpSKsCAaB/BezqyZQck0gZdPEOkB8pVUY0qN5hvIZ9tvf2gj
gzuSujLQWm4Z8XMsSa1K1b4Z0bY8WH9mbzdLBvc7w4uGFlCUVxNoCY13kADUbOe3EFayP+mUCmku
VWkoBQEegtCseFLQPsHWf6HtoIZSqOl+gUL4e64IhVsljnUpA+0IS2a7jdM6uw0fqHzofMxS770d
OR6qIHxHytAdzNGChR5H+mflHLL9Gb9mSL9ot7Qr0HbIwRqoi0MG+HqKrHwdGaDO6PUZedNPFk+p
gfKmZmHPVPR2G9c22tMsmg3Hix7QFGYAcNu1YSsUmuEmD1f0wBkKmYQnsoRTqUOt+9pDKu1ytgZz
s5sRhopoubIqwiGVqs0pkr+KhjUZd+Ph9OiJpJIbHqVH2XXg/axonaEmzJc9jDUZ17mbrfb9g44h
eJbiGw4iw+sgsK0e+p2UbjvFgvgV9fIKI043iMMaawHlg3GlybZA97+H2ddJSUCbPZ/uIXNW2zGd
eX95gQyhmI3WYEivxM08EFw4b5qaVyIc4VQUGnLl5Fpg/ns7Mf0o2YjjdiQ+M9454nmPyRjvpLN3
dFlf3FHAcOgHvTeVHXWME5T7ftDaXmBv8XIxKrCqmWhX/9QRokJVASOVLoNxrCXKuE+ryZTMiwNa
ovZCMukg1nO8K1S0wNUthI4ql+h2HQyO4+KYuDB8/nXZsEEbbL5e3m/p/5B2ejBNDvNIDiqya7bV
sIGXewwZiUc+iJiT87kqCC0kDpbxHnOYankC2bwygTEf2cdlHuodOcMDk/4mlIfkQc2Yd0WnkY63
/wKrCn74yoYPocPSo3x2vS/0wqCwAFYPjN1PcLunoc3NW4nw/ciHdBeuIl4yLo6COIsuCEj9n4fZ
cue+pxgNFgL1128xVdI5wK83wsjHTSgWDDXlTV1cziR0RXLMPvusNDKszYygA7rHqnHxtMwdQD4W
jcSkUtoSlJOhOcD5JXuhvjjPmAXtld9bFAxlLGBXGKuypLty1+5n18VbSbFZmXLjppEDnCUT2esB
NdyWOy2fdsILNJIiMu/ySFa98UU522+9dU++zcBEfuNbuaKE+cqvzDZzrZtRvIxPCxDGGztGRGfZ
jLt1EhN/hj6cYefaBWSrsrzZpywrxq5PR7ED+VC0VfWj1SShd+RIid23UCsRDbdbNmqmZmro68wp
Q2aWnxjUOLrABPRZNhSaRIIlEESxz4EWpI7i3Xa+ZGVOEtfNYjst2p+3lMWMFrQxzwR6vatrWTMd
Rn1wzVLHYdqL9JQv+saXFrzlAOv9tCoF61iE3n/S1J8uLjrVMyJ+VpPBqDKn+dHFoPs4sNn+v0Mi
g7w+q/2pctS9uj9EW87jDTDVWbtahW5LRV90VGUTU4CC4It/YZo7XgTPH2nh8F3l5I37+NewduV/
uRpyFHODPZMPGd7yBOL7YMS6dBNX6g4RvaWxTqt6WKuWwMnzONKmxGJnqU6bNpcanf0XHmXpKY/v
aOtaoVTnLbTA9NVsEM7bQI1f9YqXyv4XwBHliR1+iQTQT7FxvHZdINE3P/YMKXcPK5FJ50dcGpsF
NDpM35Xm2lEJmVUVx21m9BX3rK5eOm7NWQPV+dXPS3ZllurDs9nPU1l1o2DkNiY0kxtjmgmO0hLb
ijFG/b7ZuAezfx5Ge0VUyvdXhloXxrHDZ/MqFJOyfJGVhGyoSDgeN0f86ItSS8cK9C7h4V83BlxW
o094NnQqP/4IISuu06gaNG/oYkn6G3gcWZ479/mMlMmL5I4ChjJ+1t4fhZgZ57QNE0vbz6RX1AFt
4F8szDSZ/F3wOxKmCzg4l5VfIaHoYwGdPj8ac8RJBlcLIYufF9u77o3dMBuXQ19Gnf3G6XxpUTLN
JBx+9GQ5vEEughb31qDwxtLYjJ7KFImcuJkcOODjVzNjJ/5haVjqmr3hnS/aYj3au8qvxkOYc6kP
GVXn0b6I8ZOEXZl1mRBSZymlp8gAyL9gfSRpttbUg1ettwtsPiCFVN4D9ufodbnbi6/lwlcKjCxJ
WHZ6nO3cKZsI2W6RpmopnKnVGKk+y6s6+BbxZegcav0R/caPyCFJLlTyuQVkpklDASzh1pENmTh2
wAQrTT/Cni+UONeGvgRF2VjG3VQQnaIEYh/Bt3lOU095BSgorVlFGjoeXC92Du1L8do9RIFstTKQ
0GV/fsCnv6NLvZesrQRvmwafJ6aHZDA4qRUeoTaj/bXfPlIKN+KlkvAV7jwEQ9sht0kfZVBXfTzB
SEjmrGV6RJyl0XyTOKS7QgMzHX+HOgXxg7z2yZ6EjOtXTLlaqrwTAki/zQ2jKh8p8xYBZWbA+zuG
3ecj75ogKrlhdWOSCOUz5JoORK8BDE5jnNVYKkWuFc3SfLoXJ8fN0fLBCxAcXABBViNxkQyog5GR
JclCOJdTxeY8RhXrLmuV3vmQRuyWnWhUKSTIS0K4yVCeiAVs2Opn692VGKWwHrapovVCzHIYM3ez
5zNbJhRUUYVZsoVfZPLfpBP2+KoIA0VmHvJMKWB0i0vJ8AVpezBdtj24HmHDzD6Ndlk+enXrDK8X
zRq0V8GdAUf9wnRS+bxqN2gLpR9RegLDpecXtcCtFJnCnThceLTKilbNTVS1SXJhkLXtB0qxKfvP
+h6WXSezbi9l6NVHkNmd+QIrdfA/WIdSjgy0j1JYdmH3x9nfoqH87cihwZGXy7Mk3I1QVh9VLXJ8
v3egQZM5bVFZJ5CneF2ATrPURBF7xXy2kA0L2QNWd+cEkF2CunWzI3U8asVBrVXCMk3g8uvEI1GH
GPV8F21zE1ar7/SG7/QuGJn1wC8IGe5gKK9YGShl686oXoGj56rqBn+TTMCxyytk634EVjOXuznS
VHcdrXKDvI6NEFYs7Y9SR3qeL5Jh3J1Ce/jBi+ztbjlwEYSeW4M++/NZHXOrCdj8YmGyEJZHzKzT
a1nrItbGN9hkSL1eJhGiImrY6ujt7dGScQrCa5NJ9/f5myMO27TNsx8dFrc32vh9BcOa/oaBeUcT
ybAdy1sGAZS5jZwMFuM9cxne56S320w0gmu7bhf47oWempS+yoCmKBBE46eAOvCTIHFoVbTiXwEy
UL2EPj45f7a7kU+iMScB5rqwYey6knG+TyLKVqXQ8N9xz6ahWnrpgXxPpT3PogBUAIfNpVDu33fo
Vkce1SYwMF5P0QC/ACDGCwB00wc4PEGw/Og0NdCL1LssndPflT1LIFobexXL7xjE3ukkk/LBfsR0
G0UHuvhf459PPsQh1ImZjJ/lCUHhOdL0oMspir19f53YKCwedB5Rd4OLugDXXPZgknOMKntstAGB
JynRMH3Wm6jmY5VLrHKcjQwOK1IOrfOnbE9e3KeXohxhZ2HblDVBLWI+UaVbabfdqhsfPCpqW9Rf
X1xHjJ6UKyrzZeugyPnJl8VFPiJqgL0BnJx9KGKsv3HsEZRc2dRk+ZGIvcifmloNH6ZuN/AbL35e
PuimtK5JJF6OhufZRW1Tzo9A19r4eO1ew0+DuZx5Wyn6ytIiBCG2pkZL9m4OwJwKgsv9wWOCStKA
u75G8ur/pH4hQW3k1CB6e3GDZCvrOXPjzbPmBiBaGBQcSKP5YkYlSLKKPp4ZUg0t4fowTJNI0da2
xPSPCSuoDWOm75FSuUtgJ5cBn5wrLz1mvWQKfpSrV4Jh10fKnGoiJqk18xBR/G9w5S4mNVh8zO5H
dJBIwjT4XgYaoFcpCvryVNRRiZ3+niV//ARLq3OBr3lMnHF+FQNWv+RSaweTWAUeEPOgFPnveIyw
pVUjzg58cOOdAUsTnctYYAHXeB5cfVRdNGc1hPOLi5Zs2BaMIa+KEXPiyM8huNyt4tp+JqaSdo2m
To3R1KF3qkkVMoJT7riqOqF/fSs6c0+AA+HsXokLkf+8wDH3Oxc+HNNWVrAkyTBCV69D3/YMaBXs
6ola/69guzztsyzm7+v0aNX7uNH9Hu7XdKOmcyB3ekcChnYV3aEPuUuwRizmF2eelRuUFqGShrEB
6+PLlk/ZNcTkeje9v6nMqwOK4UO9uZbCQ+EoCRLvD9EfmNicKYOFJ02ITGDxGdLctnblxrOkzvfj
Z5Kv9aL0YrqGcvqN+MkUnsyXaR1m+Y/9Pl0SlB2xtRCS2g2x9jTPNUhijTJdw7VUOtMCEdcMl5IO
/xaxHO+/x+dRyIMIBetCpoUd26kJiwNKlsYNIbTvpfPOFg5fFZxAfR4Ve/DawYwSXUm5but5eHLj
PhWtPwuNmYX5X/J5Tgj7Ju5eGlHc9eEgJdvaj89LxPtdkOhmd3R+9qhBeGXsMUghtoM3Llj1ZerQ
/1n2PSNgMjoDnRkg9CADd0dbQnN7vj/YEpyX/1OYmgxcR4ktPDn/LYbiQ0sCFb3EQZnasxFkHQkN
0NyWsvY66xKDtp5bEX+mEaPxXSHK4DWK+D5HkT9TKsokYy4FxJKbtya45UwrBQ5kJUJhvmPvyM6R
+wpeF8dsZlosWK3vXr5CuQ82yvXhF0U3tJ7m/JS26cMYOs1YYFD2nSreFUddBzU1e4X33d/eZdlK
gTKdkfoOTnoY9vd8KqkYcgY69z1ysvaHkumDwvp5Yj5TsTva7gzRlnvvA6JpPZHLbE0YQ8TLUEcw
aqlj8I1Cd57daADZRfh9GvQlgM/XqjMinUJF4sKIfv8lxILqx3P1RyIB64WWWsl2+2gATQrSwlDy
QNcx7udyBZCdq9YrR3qo9ycR6KbFq4RlgdeDedwTl58WBasLbDrGqbCjSnmLnya86iWJwW2yBt6U
mlAnKnxRfJuvs1h89IdqiXWufsOBxISRzMQA0+23LLVoYIoB84/6xZBcSju9qWoml3ioMXVh2ILf
AfhlJoXQgeGp5H9IyYrtE381wjWoYljVpQCj01T3HSsLjSKgDf0fdTjyQFisZgITC8s6eCGrXVm7
Tiip2Z15KGQy/aCSJlj4hf0JGc6lpm1I9x4KN4UaTrLvdcLANCbqa1H5mFUVIV4tyYzwldM/VU6X
+At9SL2IKJKEpPKJbaavEKnPfl66GMnHzQzu5pKoFm36wUnInw272fnQzWyyqCqhz4Ysc0j1r0Ce
YFy+Z4vW/I8r6kqWFiIHUCwVOplwQn3kBsB46nx3x598fayRP8HOwXoO6qjrONO7mP7I7ucXmr36
rfafjdSnS7jRLQ4yeEit0UGBNo6YYEW3i7h93yQRsOMJEZk8XPxAmU2X3go96gx9FzBMRMfhGWQp
BiqYCP5dIOJokXZjZ8oT5qrDwS1zaKpH05WNkNvhfGiA460yINGEASfAcgP167A3zMZBsynV283k
3qsxvb8PFvq9lCra1EnoALa8M/R1Ely54U8E2SOtlVLSfA0QY1IuFe99FUqn8ms7bbOeA7jo9sNt
65REAMSzs+CHneXFLzUrepRXOyWtxA2OsrMPecgCYyWnLEFyJpB7ukR3lw9b6oZaoFuNIae0L/hn
OLwhNj+YJuJqeCD95s69xejxV2dC2w6MZ2sBHPhAs3c4pCfBOqRfHciQUlUfYML2tqoTifAsYtyE
zTaKw0eYj2oW6WwKBFOaMVNA3ni9ofFDQJCSPuqRNHdsG2o7u1Ia2Ji3i2qII89soiB8v2ctxFZl
OUbkVDAAjcDy482k51ab3jB6rVfr5yaFjGVROIWxTFq3BqtfqboKAJGlKxCpao7DTbXbPBNCS7IF
waypy2+yVF27e8QnE5TSf0EYz1pJWNtRM00mTF7pn0ZxThLqbzZYdP7+qDLUiulwTOTTtlG6zovf
+d3jDvCRc/m3RTBZ5alR7vEfD+9uIErTJmxLWedqUo6iqKP0czoYqf1Tsuo8diFnwsi7Bh6rlKlw
hhLntegdz77wdLWgCNJLg2nI3PkWcCFO/ikenlvkjVxAkqxi+gEN1qYLjB62GPIDmn9sSjChK/tQ
cupLzxeK2hcnix4lWIenEGhfLzYQG3SsN6fDAT6PObwKEhQDS7Erm8haqt0sWNNyu3G/DK7LidvN
9bNwDa1TZMxbSnP5cGkBZ5GT1OVHNDOlm8VV7RAm3pGG3sEPF4bn6Ujmfi4tioT84XOhbakDiWCi
wjS2WmOyObMHVEJzH2Nw9Y/etn4ozcFYm9sTiTyTwhrWW4daZ9HDjVu3Itv3t+eK2RTmK3DJAvhD
HawYQSnSdrQFlQNxw5YByUs6Y/G1FCj828IwBKB55ySNzrxMhMkfV8AaI82Zkd3ir/5WYdf8J24p
xLnb5P/IE/z1Hm/yMPcoBM04ww3bgmWQGIK+jF4ZLROcAJuuJf6uxXCHSXo8oMGI7UgvIg4LGJuQ
qlAL7engjAKq49R55tCO5V8upnUdGmtP5eFUkH59gvmW1mzYbM6ahzPahfNpu52uFzk0NmtcamJC
RpG3tgs9iDcMwcGPRBmM+rUfkfE6tZTa5cU3GRxg/whzGL0JYPAv31nmRUgkiuSn7qvH5wUyD+K3
7J62iD/0iznkGLFW6FkLf3tR2epJeBs02rYNvX/qkX668P3xiCulOOnGc6Lea9esQJfa6n8v31Rk
sjjY+/Fb5AMSzZnnjkRGXwywZYlKybaxHRoO+lgtsHi/7QfccPOYFVMIWJJElW/xUwUBKYd6j9kW
y5nS0X8doXsWMqyG/b3SN3jkHCTswa2Acbi8FmKcLJQI1EgCnQATveT9dOSZTFQ3tX67hSm2O68p
6jkoX/fCvg2/XLdbfVogtla08PNJJZUpuf7Yu/xXM6NbC0/fvAQGp4Td2cEFZkbGYTaCxXkDSLWP
qqxqHPU08HdX2f8EjcMVcHuX4RumSY1c0G8KHYXauMnLC6+Lyvu8dFHuFm6etEwtBrVmJHRomvW4
b6Mqcx5Wq2ScTYAfbDMHELFOHz/7F8jumldATPL7rBdFN2TumPQk1ZMO6Lmizhd1tes+obpiI6Wh
vzGUf3BvlPKmpAwxN17FOXIDXNEwvZ8sLyKyJi8+A2GG0tS6QBO4MGw/dds0yuF78pGw8aO/XPZz
LpNPx+R5TdG2Gb1stEB5DVAf/eWM2FdrDGEEb+eiadBBSWZbrz16n6BqRK+p03/tdEI6oYIeXaz5
EdlG7wWapf5H5WA/cM6CKAX7/cyio2lGkDIRzq/cEq4lWBtZN/5lG6uS9QqfvoxvQY2h+ZUvHRRu
LN8rSks9IAz8FvJ7cxMydEe5jfRH3IYPVL4OJ7U7mI1V8j3HOZwo97pI5aWJcrD5LBjOYNzZRoTJ
P+VC/6EHCk1dAbwIHrOCKEsN4yG+lr7B2QNr7vCZBujtAMP70tXqP4Oe0Ykvsllx8Lgzn38cy2tl
0i8bCSejY7b+BI/eGq0snshsXZ0/a1mr6IqnSjw/3ruSlbMt4Byjex2tmtkKkRRs160X+HBI9RNR
WYcEwzMbhULg7/2KQ+eL3U5dlUNI6l6BpTEPiQMlJ7SyLwxyxF9rOIPScUHhERk0/0wNBBnUM41R
/U9fQQt6Dd6F4NXlUMjicbyqFpcpxoGb2Q9cO5R3hkV9IkzbF7aO0oXUGkXEoQquCQ6QK0XXpcwt
RcNHsde5GcS+rSfvEkVS1nQA55kAz4h8MsnFQn2pEGXd6iecQJ2AclVRgdbxYTe0xFtq5+XvMs22
O19mcRSRc9V5sBQEeU1eb9QFzSPWXle2GkMhTvKzmJAJsELLaXpkg6pmhg+tfE5elmCQ9yOU9Mzm
Zqtz59Ktk1KatyFaQjjVLa8J0+fbdHIXYvVoZlKZFBrVRrfrcUMSme8m8x67DcqVFttu6XcPxHkr
SHmcjaq6zaVyn9TIrVzfKUw9lhDMa35SyGm7EkDGVGBNeczEyzHCuV+yQf8FfgGRCHbElPzdy07g
ZPHgYUwjh1GkIJAS8JymdXhQVMQc8scifULhjAh4tmEyzJ06//x4Dp7nzx0AXED2RW/VTex7GsUo
nLM3ALN7fEDFVV1mt1AeFA4dguqw/bPVCdBPif8nW9ov2V5IGKBSnONBl8MHEL02pE0WUjsUl8oF
SaXVc4nPeC4anour5gjq3Hv/vJdy6I4O7b2QN2J25B3rWVYfjm26wS6mfuRiCSiXF7kU8+sKTRJI
7Q2zVIg5l0eHy47dNDOvaki4LOBq2bq2tZZ1psKEfL9lghH5iv4xUlMxzEx1VlKUYAOG3Q7npGDA
5p8oqPU4ZHHuloPp6TkzEiWq1iZJeHqLTuVYeeIMcuTL/Gx2YKzBxn1xaNV4V6juYutGoscdYt4s
93Gaq3egHu5zayDr+UbIFnksI6eU63q33uTf9ilywaj0V6KC34laIqwJwbKRtQRp/uQt2a+wQhuH
Av1ZDG2xJ65qVvhkuh7FNWK5YmnEvzs50QuXFHm4Eff9oNqyaoi2ZucplLBVxrvZ6rATQNamiurH
Udo6oN9u2xy7sDsaHCJ21ViVpQcsMElnjcf4YCCQ0aV8oBVH44Rj4ODi6wYr5lDBsePq/AM60tLk
EVa90ql623AvoF8I5pMpqrS1j8Z9yNIQsP8yABeigSonHPRraTzt0m6dlCRseoYt5toXp578/KKm
StZ07cRXpdn/oj1pO+tTlBwC+O8S1ol6hT+P3tDq9jprKSQMH/4s5AAwDx3It3Kvz0dDaIqNglKo
A6G2E3FXTgru1xXIH9peZAvFbm/7gvT67G50p7UthRBY36H/FrBM4RuOjwoLUSSYlIFVMIGqRqXb
sEW8SU4fsnKYLTlaotCjfulhm/S+jWmFnQ0HC2qM3xzgPKZSq5GEzLHezvsttnSCp/VvDQXAvwAs
KeVKt22N7Vq380RwrVD3d3fPXAdZ53IjMS78AomjazVfESzatYfVfinsVrkEIGwgdvA+mvLPXISA
GAsnKzrRTED9+mr96HPxCywb7iNC14W/m0fGeQ3DSb+MMfR9C1p8uw7xp2prC6B3uDi8F62knbzp
dZl00Oh9hy1Vcu1hI00JQqm7bM+sOoIoUlZxM2Y1e2FC7kGTcUg2VdkAQJDt5OUHQYWXibpgaUfS
SGtF/hW2oq/zuxsvVEIY/CElmD2yCGTVwTggRUSw+qEV0LdIHRZAGn/ZHeNmrso9VrZLScK/By8u
AU+O77b0mcy4N19UaFNWMi8vdvQEcJPPu8UcPHcsmLkTqNdl8j3ylWglJWIHvDT/rRE5ExN7xTGz
BoBXX9u4sEsrR8oVCKMdH8bLnVeLfMaLUBOSLxYBRuZUjSsH1GuIHX6Jdxd9IdMo4fVILE2HX04L
0B2y11sksaVKr1oqzjykyz5s2dlECWmEaZjl5fGXV66HAC0/7ypLIckDGr//cXGEArG7Z/7Zka+R
0aL47hS0jILP01oDnk13XT8LTHfNja6GCu88ahClSPPv17L+xq5/QCfY5P8B9dGM6L0yZ4YnAsTq
Uvr5WM/ZM5EYip7MwuGKW6j0oBdWBWcnuSBhgAPq4Xd+izuLzMQgcdPx/Os7/G8y1BJqTJdUmfBu
zY2fTNENEV7V030UQK/paRiN+lXp4+YAkx+X6YL4oqwbj8xKuPWrm5TrL64PzhxPn7YY4+3EPmJD
zqB4k7LVHr2nDGyvdOh2i9HpyULXVbTibTPoddcFV3EDTYBjOqChsaVSzy5toTlWx8alC38AaYrf
6YeAj43GLZFV2OLzrM2JN4p+2i77iGsYlmtUsK4k8Yt2cTdQZhLgLHx4QHziFdCYs/geLrrRloRd
sOHGwl+GuJC5HlFrMA0g4a3lf+sp5V7jlAdAWVm+9YNiABsxQ0icQYL8d4JrM0wBhVVBbubZZacj
ZL1fOQcBQekO+EAB0mbg9D6XlVLOwrQyZIfQRY93bzEjG9WeyZFiYaWqrktsVrpCks9JMAkxbQQv
zEsOSNuAWuhjQc39sIKpz23/Pi9ZQcc1zKKdOHP99nBEm1oUpdT67akiFhy69kj+2KbUspebHLd+
Lttk73h/pmjmdfmD/HDAcoITp09kfHHtO493d57FfKU4PYrchMyf4mtzWGNPcXdNz/SR+29L23xT
3hR9unKQqgsXbGm7PHY6/r/iqEMPUGCiodq8k5ZF0f8uuOCqZ/gXciHrBGelyruWSIBZuTu3tAUO
b89Mcb6pvTHtJcLblqrnA+w+gnCXlibI6skpXpxTJ72HeWdpyHm49oVBCwf5dx5fdXddhcKtYW1H
ANpGRzA7q18GuHz3Vd2NsNGPGwxGpMGZBr3iP4VzMD99FIgtZEshYN0zSY6NH+pCFNHgFGCj16+s
YGvTNx5r9yddce6VyDhYlbkSs668duoEAzh2vfSGy9KJqqxTrQIHmfiPRoFJTmft8t4si0fFScFB
2mgl6PTTGIQw3HDp5+ARv/mcWAF+GpMvYwwveF6t8Esd/7LJ5NwmFdRKRW8qcLgRktL1eWK44RhG
Gf8Yo9yTK7tqxepF8IkF+8aXTHlA7A7gVVLdfW7z9Tw/Sl8CvPJIRkC4jx8XUdjgpmyzpixvhcLa
22tbqByYvA0wFQFfSyatO0IJEm8/vUNUuvpcXpSF7o+d9A+aUJ/nkeEeaGeA+pyw7RSwGClwHBmo
n3S5+R4HoTtzpPZgizlm35hFMVvUHoFySGbU8G1BjWofqSPQ9aBhJSRN/bfCyyszhUfOpHP2rjML
w1pTmXksTnqoSRP/AJB8TN220lTap4SAaFGgtSJ6+ADTcRwDvLX/chXOQ9GbOt4dS0BlZuz47R24
vQmrxHATkQAG/4qQBzPt06Ny56FBHjOpIYXpfcQFZ7rKjHdLIwRwVziSaoBmSNepAE/T9GmNQjdZ
05pQ6HM7m+FtH02K5xQKvDbqEOa82jpC9SDuVnVTnl/uG3SSl/4lRtLXl+0lcqj20oU7ITFADCk/
MZaPoOO8jVtg5sAMKS71vqR1OV9YBBdzLQsnyJcR8LjJIpR2VFdXu9CEjeIYMWUwnz2yuUCP+6Zs
KhzN28PO3oLW6z/Hnhm8+eAINLiVyCwbY+jdUbTxlgvBW8vJHP7W+O5Xi7bPXhibLHK6MPFiSQEr
6Ef5kUZ4M/sgYyCcM1KojwRoAUOAEHfvflUN8wMo0e74WxjyBj52hijXc2gJBKr7+1eSXTj931yu
yHPu+WiNj4Ah4XCD8NDlejUbNks0kN4LU7ZzY8fY3hwadz2XU4DWHQs3bfObhrdtZ3A10AzNnzdV
6Z2yVEXjOPqtceQbyVHbyS21UHgC0U0sF6tHfDfhFrVKPCKgJSKhtDOzmZ8giZOH8XMLSESvuTlW
nDVV+imve34kqLVE738Nho7nC3GXAv0Q8/mkjo1QK/t5EcauLeVBm89opZiT97d4NsfA+/3Ijt3z
g1k7ZxxcofDJBCadaJmwpDlNHCThz9YVlRTvqOAps2VSeBcnjqIc2OsQLVcfG8A1wayEdIM1U4ih
VkgJB8jM9mAawFQgSqiunlZVgNQn3BksTK9Wp3RxF2ToQ6r9tHn9KIppsuxN4R9O5Z8vG5CmDrM2
hrxzNQbR5SdBWkCON7WXymMwNucE3ESbFisdlghN1sQ75cffWv5tYZYRfHGSl8T4unTcYNrPQbbe
+XS19/A4NDT3aenVjcPkM4VA2g0nnXp1FlP2peCy6xThs9F2aDJoMIW93lIUBTE+rGqULgV/atD9
brmOED9Of887Ot88LBVmBdUpzsufXIrTzS/Ui063IIZrwz4lrKTB6rAflJq8EAILw2IrHaNtn9w8
Emmll4WM6u7jbwBnScrHKS1vzaOvn02X1oZ2K1C+qPGzpErwqGLTxNDAECyuL6I72TNuIcNOLPMy
NC3YT09CsNjRj1tlsftK/OtoPS514fcs2y2QGSRYu8jHraC1rvKTpLJKmEeJlGmNq0crx+mkFhcO
sWkBj7aVLoihACYAc5DcK0fSJAgEWfQOLPofZAAL4I1o9QYWddJllJJnsG/k1MG8r2stXCcAMQ8p
GvPzMSJuKvl5VLDEQheam/4R0vwy0H3QM1b3yZeknDDwY/ZDYKhPmY+1f36o2tCq8zhcAOIq0tbT
PYClEVcOoucTM+9rOEDHBqJNrQsUHIvJttHaMVHI6gbOt91VL8gCVedcVQX7wOWdC5yYyIi+FeP/
fYfyauNj5GHqm7kvNhNWBlFRLf5a3ENYC3bae2XgLhXkzuWuMTkQ45IGl5Ij492o5Re0xdvboRYm
BvOkWS/Y0fCuwsMDoHh/bUY4RGPDR81AmY24IoaUf+lCA85MC94dR6NU8rWh9U8+jv2uN0yDcMGb
sx9zRip5lSOnk55i9v9tmy+swO+2f32vwOTA7IQ3k2GM57K2cGJDgfkpwJALz9fYf9UiLiQt1wr1
X0Lpdl20QdyeJlgm4kdEzfxaWYqvLsqw9fRFCxuLUmc6tKJhNc1yaJfuMgvUeHPuZ+9uDKrsMVL1
t/PVYKqY2A2YB0/CTSySlubFAL35GhgY0nAReo/Gt8jyr0+8DdLfCCbVdFUHoARxkfLZzrH9LuG0
YWY5u0nkypYrdKGWdK+DKm+mWtodgTZ6SMzqF0FyWnEwMKMqI4nY9q0YJ/+eUGCtDgMOowxlrx9A
/Yewj2HQnNE0EimZiC8NarR0Vt/ivS1Valkew+5ZwZxtSC1/68Dm3CVCU0dwp3XBGREIVIsouzYr
bSb8QqClCFstJQvUUiABF46tE/baHXycnCmbRImOwCuYnd5b84v0pTsyTecDryU4uUZpNf+LFV0z
xWbX7t7YOqAPnS5eAMTKiQElGa6xCxa0dSrHvnk/S8mP+J9VbL6Rqh0mQG2F2Y9N2w10/+9o45Me
3Z0G4l3LjDEUEKUv+/4sICIspo4RRdcbjuTTL2eXSMXCtdjb7Q9PBFufF8tMyQdDIg14y1w+B5+n
g9naa2VGmLl0loQliQ5c7kkYet5A7Gml3ToVHBsTAaSEKb74ddXxOju1LEhZ4xXz4qbVOIuvBl//
p9jOUahxFKh2SpPXPVZrfkH7mkNuVyJBqvyNrM2rYIV11Vbha0Ki/Sp2hOBOOlYtfdH2DquAT6vy
L0GjZVgVvf4YN7NWsyWYrQCkJPVQR9i/Dz0+gVQyuNpmkqjw6ulpTFx6CmSma+3Ww6rlxO8Sa7Lv
WcgqG2rM6qJKNt/8/KTVtIFTUdMXuqkVRzWMNRYpAAB/pimyB3scaZiiUe1ESnwh/i+DeHZKVWz8
YyKYzSMto+A4PYfBQ6kgCHIJVn8bBvMuH5maf1nSowUmvmt+96jvicwAXtq1RJydmmNq8FfsUtJ0
MPssENr3jfS7iinNyFPa8NIww67nyrzGPrhrC8Bx+BylSkTuwImJ6QVRBOJyfQV6jJrxPYBAL6+L
0Tk1K17B+s76B4ED3vVkyDaY8GhTfX1rASa9iJIdeuGH+TsdFAV43urEMRUt5q+2vIaMyb5dyBzs
H00NtjC0771Rnt3Avg8cMUafyUeUEDvHPIrIarcyk4iauiQ4e8Shbs57kYZiTdULsEIRSrQbFUgL
5EhiRuqj4z4xg1EvoIv1R3pTz/+WQP41lJ1bhnjXyu1AL31qB4yithlhUgODU9xt+6HC1sNWcaIm
28bWf6+elTAc5AQVmxfqt2ob3FsIhFZ7bKmtZZ5X1BMyKSXGjrYb99A5o1K0w577Q+pQWEzeSgOV
ps8NCc9/DpT/gj0JbEXhdgUOsXEQiwCBHO6kO/LNTPQhGpZkmGkTTZJHDBDGyTi2K3CIesEwuFq0
YTavRyjg99xfC7KAnask4N60ENEq3Ubc0+SVyyWYp6EjlyDUYrlzfFYc1ZccZ87IQWjCrRXXdn/9
5U6nQi1zmcPXBcR+AlkM3/puB4ntDT0LCH1crVwY9OTM9mJn+CqDzqS7AqI1abBFtHTQXM0VfoS1
/Jt7IpGb+gjqGUZeoJYYY1EiQVq9LiU2c8iVaa3cuXvEQoU705weuwau9upu3Aj6XB0u3ANBObnz
kl4qiFkcv/qRB09/Yty45ZlU47miTFTK4DPqzsd2h02nlBm3uGNGzbW1SAFnSZ9KN6nKhkIMRekw
y6XRz6ZNbg+wC4yC+NohEYGiGzNxOe8Tdy5VwgpgUz0Zi8e7QCxTePlKIO2h8FMvEiU3JBKFo+Cs
PLC2U9qAuH59lbKv72FmnAGcaKj2fBHCTZIHqd683cfd19G0Dy4JdHuaXLeBFHCFib4ZcivpYbyi
2k3fhDW+XeKf1gol/uVwIG+nmEwoo/AGSLdqLFHaOpfUE4D9dLWQTQNL2BFRXg1DhubblcH1+woZ
6kobPuj8kyCHf9Zftp1Pceso6IkGPQ1MsAFIT4cw+E7EJh5A3w/rGiSY5LkEWgmK4UskywgvYdTy
jP2PH0DPlcW5ZbOFHZeI6/NIzZ2HZnL/tXtnxQa0+CAnYTVNG74odu8vOdo0iPRdDrEuJcBNtr3F
H6uo3qWtEP0oZc85Nfl86vqvzvYtvjZO4eEeFwA8GjMRxeYkrO7y2XmORYPno/WwtcqMBTUSdCt6
+ZFFXIIrfuxLnLYhnLqO0UHH/+IRu37t4GH39Y512zpyL4nr+jAXqxc5hxmldGD6Kno2SyJZBvqP
8DPPRGs6xAIyq6AAFXPmZc1t7LnFtT3mOUe5JnnwqdR7iZowEt3bKiIrnFHe9JX9p7jwhL+ptnSc
uQgIpWeA1RCvv6QsD+2d8YhSCVV6zxQKLeD7b/RkJ/oiaz3DdxwGgM6mH618i6HGKZg0oAKwGN84
q7AH0Lgqadziaw6qdNERHt98S5vXbeAtPXsE9eldbAJ4OrvUY53U6iBhLtJ9d3uemH+P215qC8MG
f2YvR6EsIsDPwSHkuwP+DWNaahpXBsC2y22koFPeRNe2naMzmVo+mEU+4PxO3exU/cyvxD/45yvc
5v9AB5XSZC3+lPUWcg58BX38TfivTvVsGI5BYr84BSxnZ6MC2SdEV4WvDh5d5Q8MEIUcWBz/frIn
FBGSiPm0M0Sn9benCQFdblXiKvypFR2GBFnhxgX17O3OSYDT66rb2lhhtPtb3uQx2cTCcuLE+tmc
iQ3dIasLk5G1ze4OW6WoJRnv+1dU0rGRgY5a1rTLAzthBJPcDIe53nBQchSMVS844aEL/Yf1mwV0
KrfaHNjNKo7gxRW+6EXpTKtH4fWgVZTbWoon5QoIz6pPnLpBc45Hii3DCGdM5/ws1dcOmQr+5ngE
V9lgDwQtR+McuFDg2/5tsqg3D1k/UKfIg4PUtj/JaOWoELa6B/Gj3zHG6mzQT21YGEX/Z7X9gwH/
BCJ0jpOOHhsvkJWgYPI1747U99+1H+xYLARj8SLnhU4rji3hTHWF67mmYWFtoqThfV/YSFDsySlu
ZQzIAyytf/DsquECLDAqu9VS8FtgVHEGgfHbpWPEQKjHalFjaVySb0iRy2qBSsYLxawz0SQsPB+b
jULzZkQllDVWNYPVLGLUDNKDl8hlZA7qheYXYlSSqBkQXXi2oxuWRGJcxOdvIPRzBinrkdeIKj9+
2hHK9Wf5RqXiMRMPGOxUl2gsqyWkfwEF7IIIvdzpoy3XVjDjPvPd1j2wB9O0F10iXJ1gijJV/a+U
zzC32xle5h4xZpS3bU/4/ocQHcVYGALlokZ14ZTwmyfOjuBVUM1kf3PCQ1MQ+Mrja881hip/rB8i
lqE9iFJROCdmFnE6EdrMTfZCqlHhyj2SzKfKHozthXpEH9iaAFGLZb9Pt2ZakIOW19m3JPZGdOCo
oohUbH9JTx00WCkm+LXtI4s9xZJNPNEF1pvFRXk/k/a27ZezN8bzmRq+NC5FYE8S9d48VuZXja2g
kRVDIV/PRV//D1iviQt6/Mbk3oIrhcu7pR+2MkwyjcnWzsIH8TirtEl8jNrInPRUIrfA8DDqa1Jt
UwLSdWiEbkDhnw6650DxnzYI9h+MsKsX3gCdCiXwxtqJr/6TiTDCbqfcPhNJ7C41a4jwIuNnGXVa
vehoO7LtbhGX+twz6bpw1OlGK6eiYKO7Pjb9ZD3lvEfe2rSKhtG2ZkoPSf+03TreqnM933xQh1K5
C3i/argjKeT7RTwVB7tdZK/3emfoLw7bsoWtKNml4+J0xHO2FwmCuJepy9bv0fqdet0Y8Kk/BvVa
CV1SC5NRmSTtpbbVbxnHok/Dl83jk+X7K4MJL1E/K5cZqa9ArSRNdaA20TIdGcES4XLRiZRcw+li
e39Uip6uePtApJ3mFX8JQEtFl65MMGgR8jaieZweoR2F3bzvvRlTysefQfXsrZ1Evu9sHnCfe/2E
o5a+H3+Ogg2uWBKsqx8MlgJfZ0QnBqPswTCjSx+RDYK+46D5J4/JQEM5Cq+s6ZWbrVtsDhfwLrDx
EVN5HBpraEqKw467XGYv2AzgcMT5XYw3mpiGu+4rrFIikbgaV2so5c25PMvF8ztKrgphP8AmyV1E
A+BRgHkbe2pvCQDZ4HFWnFOTpDmpyufWPb2m8sTDLpRMl2jz5YcxzimSbBKFPnxsS2D8DuX/NAaS
OshomaCGxDGxma8XJeGSAcuW1uTbLb83YaNexqskbE5scq8ZZzmITo0aOQrPbtqgpsKdX7PTeLBA
a0uUTv85eqjdwXqhdl1VSzsdj64/aqaEqg2AjjeFCNaIElBgujnxzk+lx3vPQTJPK3U8BF1nhUk0
1Hknas3b83ap2vScw8Mfh6hMrVbZ7+TpWA0JxhYVn66lj3s99egrogqjNrz3rMFYABZHaemrJre0
FJlTY+6FYzemUYLBz3ouvoWnAtckU3XXi2akm2Z0WuBbhGh4FU5CIg+vn/n683wh5gwyX2xPyQ9Z
QIoTCb3rAnuzuOmmTv2bpSOVgMI+OIb84F4pd426yEKpkfMVBCcGs+Stu3yVp/Ajd1Jw2gJiJuQr
C94fTtfGPcKDt8pEvaC+94Kb5fKOnRw3A7wnYJg+t5rzoddi5pCBitVMM7jN+8BCIwkB7327bH6o
s6DEevY+HoTW9QnIT10pURWvDmm9T12yvC/7N36ceEyYC14G3pt/luweEFrrKK4/AyXnnVQ3N9tY
swbyMlklNn6H2t0Xa/KENy41kXMelOQYTb0g1a96oL1PPX4cN2b8gwjdz42HZRekDx8ggcMRMWNq
UGWrB8N/UKMylh1/zSHuDXsbTeAQBQCNNCcoPGOqAFXPRBA1JKndobj0zFvogxGqU+Uh+cdk3jwk
pLo6YWeoo5xpaR951DE2s00jtKKkJO1pjC7yP2RlMewXuMxvouJFVkEVrdnZhpqLsJHmQ707YN2/
HipulNo+ll8kmhZ3felC9Xf52/ckZ0297zwLWzPYvsGfBYCjSttStMG70quu8WKk7RfbbCdu7bRe
IFK+Tdifvt1rXoYsreZ5AKsSfJ6XHFxtmC07ExeXKyAIgmIlWugbpcobAZul402sLZvIgaq7nHYI
uh2n7b1WNzPEQVSYbE0q7bL0Ea4RSJVV/7ysghUwjh5VZVeixqTdc+1YgMNpz62DRG5GEbfaVqPt
KsUAdloRM/Zd+PHdcykWX90EJiaIvDX8HaJlXNmSi+mUgFtGpRckNHGzTABgR1rVnmpi2o7D5IXl
LZDHXlA2gUIfPYXLbq68WubVn5ciz2MxqNoTQd/jDv/rDNOm/J62w27YzZgDkJY0O8XLwa3C1+To
IeKmOb5oRHTiekQFwk45oGsLcaHVxqNcy2Htl+bCkjmdWNtdPJrqrPeJkEgQ6S7fegVaXPdYfTjP
np9HB1hEB/CwxAQULAhDFZX6+knn1DXzrXN+GVJtOeQqvUoC2S1QxG2TVSHXF/t8Y1wv8nmDAu16
R0weMaXjNQI/JTbvyB6WtI1tuQ+9yw6bJYpj7V9z3huW0zanPaZMHDok4SeqafsQClRIu93u5/7b
X4ijrTojgN5Lh03beC6miK+K0P/JQMKhk/wzBz+ojwx4tClFcu3N+gC3e9ucDr0XuKg2a058+odU
QlqAkiE0vpsSom1MbLdC84CzuH1oDeuHqMN8zsQivg82VkPrUr9NiI5u5LkKBkMESnxZj7wzKntG
iT/p8DBgF2/UgGfocqFrWYCINVsni8D8OZGNQFFHtj5iHQr2u7rdvTHnQWC4coCZ2MbfWblDG9zZ
cJymthKYIz8ypLa57O9jyFV1XekS/L0vOn7t//WH6X8PLThA6V1sA9CZiAqGmuJs4zoB7OQkRPHS
xX1V2YRt4u1C+YfFK/9FkREPW2cOlFNcVu2qeSa2tFZJo3ltplVN6nazbcf9ZVFPocECPg6ioAII
1ZyoyugH6CXE4izvMiWurNX7WejM0xBKrZBcquotKZbgXtdch54ypVSjXi1la/g+NyrI1xmjmrsd
bIluZgXmEdIdezfyY3FwrOOW0oYZuFWIFG5SMhHuiCvxcmxyccNeink97oUmRRDW1O/V9u5rPmaK
z7Sag/fGvtkMIqkNuR/5+8D0lu0laZy6cjgvexJbGiqNlDcjBCEgwu0Wk0uoHItFj/T5A96baYfr
AHmYzLDl13bKSKP8iAQk1EprTTvK5q56ywsCQw3Eiwz8oEwQ4ZQAeHTIYjV1TaQrZGWGU6jX8Iy6
Lk0dXwpE8AUs5DY/U/YJ7VGVDTW5cBEyoElB5WMPPFZ/PFgNPFlX96cmhB1yH8NRAxnUlXY5JUgx
IEtWjEhuiQLqngL09RG+rrzrH7ZK817XXIc9zN2gKP7pAXF6aHvEazgIKDiyQNzgizFTw4XIUhgy
K1VGIG/tYZgBn6EWtnyLzbOYAszMzKU3epIynaQt/uD7sl4ggKDWLhLeCy15itWUxnc4dIF2QzJs
qGM8OyAN6bcu9YhrfCc2wcWoO9PQQ0JMPc6f3EiHSi/9yJctlI7EvnyKiXyXrQeDXMdw+e5T5N9S
0ArV80zu4bgS8bu57WIsPihfxXI1n6DyYC5qNDgCa/oIoUhGvrpvWsuaCGN+d1Pw7wKh3ZojmmX/
JRHy0s4OdizLOG34gmsasJGT7GV3Z7NEi9HyymymQEOH6oxy3ExB9Re3zz1VwH8CYjUJnxm3oxF7
+aUSnNCoqT+ADe7VEyKiyHm81MgbBsWXuhJj1Y+yPS/iNepl9GIx5LdI2qvKkFWwM+0t0G2MbgiZ
US6GJNDscDcEpjXHEApIse17gKbFfP2OIHDIOG64cOnzAtQ6vVZknRvQx26+Qpa2N31DKoqtEvBJ
eOVBEhEq1wMq39i51b0fbCWpF0GJfbqDo81s9GaWHM1FWpvrTmooDInbv/QDzuzFvHIcZxBaU5VM
eXzbVIbRuSS8DROG+r5hwtS8AEVr5VDTpuHNZyq/+rn0MswcX0mMYTKmFV3jduIC+sXZIas+hzpk
UlIRcbEJb4peK4QMVau7f/LUKnp7P+6MAwHUsWg5T1nHY8bMkXrbgMTs+vPQQFSfsA0ptwisCAQf
XjBz2JRMV5tdHX4eFl4CuIOeWySRi+fOcmZmAv3h154xihLstMGDapZEWS/OcxlD/qDgomB218Lf
vakNLyhlDLdfvK1wT2pN3Go87urZQ7QtGT7bCUbcXf6rNk/iG7biWmqVG4HTRCdt/8qcYlT7PN5z
68S5aS/dIl/xSA7QtlkZu+/gJfz2e8fXul2JwA25UzOgomRIpJCJNIH0eF2EQCGbvqUT/R8RL6Bd
pdmwQlkHBiBMxZP/xzoUOZnDAsUj5ae8LRGCQ284aaJK7NzClgCeP83beSDr7WikNCGZqldtp06i
8Wz6dcNNAIa1gZmIWgRITIb6+9o2H2okLC1uOKnhddfMSIUV6+1X9UkFbUPrBVpa7Z4JXi5nXTX7
y+ELqMe6AY1SE2gUWtlkxkQxv4U89E3Sk5RYHZieOEEKktNaY5UNOfLfVObJ11oYsSruR6MlJdNB
eG2hY79WhoUbTmaX7ADTt7tK1WdnLkm5il/bhON0g8aART+Wddr+SvLKK0nTiGPq48dnFRQe9jYH
wSxl7ubkxTVKR5VtT03iaOBfN8BRLBpXiu/1LwcmnifcILbH51+viiCrkopCdxa9eZX2rLh8nJhd
Ru8sWElpzRwNXYPuhCt002ppXBZjBMnf03/Z8WHqkRpIxYelKaBabMf9h8veWCkHm0nrbLmTf9+/
t41Q95/Onq+ZX3Ob33abtLFxyIhBxCJejYYk9fNLjk6IudD9ULAys/wJOZtObv28+YlfpoAGYZkX
H5QbzMfY9dbuln98VMA3PQN4UgRM0xibZEkSMwyKpT4MxhrMlQd6yAeAZuqrVx+XEVb4U01aJ8ZB
piYEhDLB1xXpZQ9kZ5Np0uuM7t6X6RvOhk7G3ixU5brhukb+NP1MmVGNbgSbfHsKAaPCjDfS/oxn
A7b4W63L4qEctJBFcpMMZZIoj6Xj3kTKioxUlr5QMbMGCPurEHMQfAGOshFzM7oKyC1mh4remm+D
NrYfOdkWnKgs34jyMn1dSyXtnqkSTHwS4mqRY2ezRayLL7xws13kc+wL17E+unmSonSm9gemi5Yn
Tvxv3UbiRoRWTJGEXXRSkamCGKxand5EF6uzeCAP69Nyrt9v938JJAiUq5vAuXO8A5JlErirMyhA
Ja8UKneAj43Twc9LCH+bZDp+39X0YIfPcnBstB62yuSxhR7XIbLOW4Ot4fNh80HXyY2JwViPkR7s
79361b0joo77aIAru9jSoMBN+STM7DDC+TY97oEbsCqwYSKFBpW8Coapy90UAqvMjqp6K00GBzoe
ved1ceCI+RS6yQpb30JaFYIJ5LLiNSiTKbRK+msOXcGhDLo7hJEAUdN/frLtwjXac2jlLRUV3FH/
WgW4Gkm7mLmKt1O4U+HAAG/ilT6mTNpG7jh9i7HW9uTeafw6vW591UEzxwg99lMlvBpLaN4QziDX
VPr7o7H15tPnWIHtDsCXOPe88YMo+HtzOHL8KqwV7uNoaDRQeVKMsongVu/rUlb3s2nvk4gVQBBz
LVLvovhSm0bL1C3emOg/rR4Rkeimza2fZVq1465XdfYjnmGixKi6aPnHpIoSTuWuiUrD0coQJqUT
46sSQZYtUqsdtfgCEWfj52WjV0UUrWs5Zo+de3t0vw832jQ8vX/DcRDrC2f0WPbLO6UHOkEIKTMj
HsRkWZLSQywFpw9ZqB3oRgEiClNb76hQht4resm7XEBZNNh9ehAjjxnsJ9eFgp6c7K+yPjZXI+Og
/HNT7BH8Bn+C3T9SalgjWjLpXaL+g2zZgJhl1fBATSA3aTRMXfs5n7AuK9Nqz7IfJPftJu6HA0mf
fJnuHSMHkd5javfmlEnYTAiDwD6K8C6UB/ePzEIvYYMxUlGWh/62Zgc7HbLTdwwK8bLJ0Pd5MslS
nF435epToyUcJBs7KLPTety7pOaQYLZ0uGkZdxdsOYiIjRv9HbXwBEn8sSt5HwsE5Ta9JzBPPT6L
H3w43n8vlVcKdaLe39QhC+DNw6lX4S7sMaOppDXYnl2nPr+gMRWX3hRux4/i64mRD3kE3cvKsWpu
lb2xAMjW6vjzIHAV1HVN/3R4Q6OtaUcYeFGUkLRq6zkAJ9iKv0zGEHig9k/9k/ItgEXVxc1r8JgY
Sl1iCDvhh1q0Kx22yu8Ywolo6+5PPRff1623PKKNdlSQHcoeVdBbfQM+40v3/NXEkkr7Y5Ws8+VT
by+NmQaE3ut7rS6PWsDEdQFSNh3kcLyOB5pA6lubposvJRtJPg4JlH6gpBI0eN4NH8EpJ0de3dZV
jDODvXqbY3o/ZHrJWOHDTERh6tV8ChETEoIeHjH67DNyh51Q42VC3Vlyz2jDePHDXnHQ34unC9ZC
7N3LNoAoTxAj1LCUpLlKbc/XHJ0Yv3KvD2g3790R1AD3f1PDRT2jNL9NrmhOqHmg0mdaKqv7oo0R
IiBX7bE2DxC75vSKfrCnzz1kMZsQgXrnoS/WCdQbZxZtMcITVru++vYv5r4FRep1DuX4ATxN1sa1
gkzYT9epb7DFumJCddCQNLsDOe/yatCLD6tdmlkksLzn3g2PRDgzV6GP8mPPTRysa68dpIWM0fGS
N8FwGaswQDo0ST1mbO1DdjaQEeuJS4RDNtQhk1XQ4ozFDm+kxTtmdiEsQHXRW3hzJBu/LRrSwlh2
ImhVU0kWjLAbKwD2qqV1glYJSEZhB2966UvqS8CExDW/LhZqeDvhvqQe7WNoHY6qjO16kaadsEtW
4xrAk4UkrMrlsyhP2o0LY2t5wncKjobuRDFVrMAog8t6lwVNKQG2yfcL6t/tbmlq+oQzlMqqQ+B4
xK5P27Ze3rZci/7jKd+BU0lvPX4lQhbcym5RuzJPnDtnwGk3hCEsEPAOT57PfpKJTdiCncFM6xs2
0ckfO292tGbq4cwDZmWJsNNrUXm9w+GMobgaLEE3oeQfkt6UDQeZ0UvVPytsH9v4h2XP95cLplFr
yhHGAOzXax14M2WbYdr/K4SVAsH63WTDZggrQOGg6myT7w8ryCcfITSRryFu9d72JmO9JURQFR3v
qfDKN1Xe+HwzTchLFofrCLHG11cGSqw//XdFCkZKPYoM9HAnpVa16eheUn1CvCJr1MVJ7QVvERPo
Ge5jg0asNOpU+Rn1vOWH+2BYe5YPb2ZkE5BLru4vdUP6M0QqyvdvaMbU4F8YEyq/v2w7xb7pqqSv
wJ68NTJKNm36KnScg2ss8Maa5MQmO5yzbWYO1VpW7CIjNHEbvCzH2wEQw8YrLpYIiKwwb+xPfC8A
/8XNkhKkUID1cSOMMqSToYGZHasYClPLBFWqXLTNOxx8OfxzGtKkwBxANUzkWP1OLBQkrvmvReRk
aCEVT62QkR2vCNHNqVmEF45tWYUlYLQbCHNTb+d5kxMk2c4R4pUbDphMU6vvxNDlQDGT9ellqFsC
w12YIC+mKOSKdiQJPzO51SFBzGMD+c+s2gFbEXjkn0cfXZWkNgu4lFXaXgX2X51DRHqwvs4RjrKg
URn7UVRw+O+cKqBKX9sxUSeZobqJL6a9lP27R1M9LgQ2TkTlh+ykT++UZP5jkkQMzzuktJ9UExYy
YEZpifgqq7DWq+2W9bVWUOjo8AeXvuXCODssroLPIMawKi483vPxar7eqFsncq1/K1dBXo9IIY1t
CvAB8osVO7FpL9iTmN/a5mB4b7ZrnpI4VSuivlO3BwX8bFdfPoT8vFeJpZn/EZMWKbkuItqSizFE
nopdC0iuSWFotjNBZ9dw4u7kFb2aRHyF7UkDym7pR7C87dk+ta3njxCXCU3WlEvnJO5z+HM73Zyu
hAqB3rX9EdoqoDL9JYwarMSigNGkxgV7sWVo083+ZAVRGsCK4Vv4517nJf4TgaTf7WV5fp7NdVNh
yCtctjksMn/9Tcv0yYUCQR7a9wr0Wa0OWN8ukQJI+cEGv6mlwXsnNcNnCMNocuPcCwu/Yy8TmxJ1
tBOy+jaHZAvQcbCdFw8LHoGf2x1KbhwtOT4jXflztjvQ30q16yWbOovixsnlw/Pclahbze/Kp8Vk
qSKmHyOtRxrkCOI4rbtM4gPKPylRWG83b3+6sroeMxiv+zKR6mqRbAlfCyPOiMRs7gy3h+P6zgvT
DNealsjw7EQb5a7u9MLzubUw+xNhyWrHWsfg6jY3GIu1iKPXkAtAVBkC7u0UlzaoNhqs6mwVMYlS
ew3t82yaJ3W0Ux1yLa7WlUcXbYugMiiCkJdULtMR9uqO6aghTtdeyU5J0ZPtbg8e9oO4QRlA11qz
kzWmTT4vkTvqoMaWhTSdHG+ABZncd9uQYv44wNu+k8P1zliyGJSDS9fevoH4+prXef9tzheyqMCl
pzbECMY3FHWJQnRIAqfNeg+DnQ7ZZi6JEFiinMdR8VvpMpacHvzQoLVeSn60bA+GoaZHl4bVYyIZ
Z4NPfBi6li610GxaKZDYu/4kupwTQHKWB89pqSvxQnDUZ3sSzz+4pXX/gefny1WKRCBJUktGnTQ+
i+HuBZ9G32EGI3r6ZgZUKqax2uCIqJpH/cRLcwUnw2VVxVSRCtkug4lTDxzo1+tf0UTECcdf3Zil
lm9B1ztuiCtz50Ft/obYD0geRbSC1mPLMtp+zOhcBjoI1qjoT4huqQ7brOo0MUjlvd1qtdp3qwMx
p7ZO7mgLJD9ZiqrJ7S+4uARmNHU243FRF4U5jO3rA+ukbBvXps69R+80UykV066Lcss8OAx8ztxP
kVv6+1R/OE9bDGgMPhjbRWxlB4RbwSTHE9VGXRHzIxEcIlAWesdLgRO9hYbN7dp4BvPaZAFgu/so
UHDsMlxN895Oog+7cfNzOZsOp4nY0eIVkBRwIz1p5BqCee+LfQpOivUdIm6x/7g/qStaMMsfgxTs
vxyCnc+6k5HRCG94igj/2eIKl21DjS6jZSdiBOOXqvmDJe1sxyGzPnl2p7sSDP+K41d4DAtSIxXM
catVAV2WlMs1S060EHFVgC0xXXSsuCw76bza7Ligf9hCuEm2PQZH6VN9lHc+GSfjmU3/ZdMw7dA/
V+OECv2qWykz9cDCSZ/Gggk5ZLWFbIvJ2y5mzH5zBnuuPSeV03SoENEvPUS1Xd+pAPpsNTEIyxsB
a0lt1wmulzCNOO4rPWWNNmlb3FDMkqns8XjciAQKRC6/zRlfypUITZWG+R0bzFszQSb6/EPlcbuz
Zmn6RcZGb3JO0/GUpupnilxhcxq7qJNn+7BVveVHQWT5YDIs1Pjy8SLeQjqxxTX3Nqjk7ZY5eg1l
YBtH/rw04Ef8Sgmz2lFzph/FJFKxlD7B5RxmPZAn9u66kGO3OpemxQ95tCgB01Q+WUg6qFUCvuo2
jeTLGUKLrXMOqYVClqF4kVqappj/RJPPwp0Xej5r+zmHAFJvsejiviTCusr/aF/KTzBM+yOqTLK5
S7/g7E56BSbIVhw7Kd+KjVkIbpBu+HCu798vfnneeDbEp+rCWCFv8mUthYNUPelJVMB1iQag44Db
ltKScC3Zx2H7z/CURPGphPTK3FmEneNAjjLFpNNdCRaEQGc0/KYw6YeBZQttkl+faT9vu9pXzhQ5
FUEWMKrd/zaYyL19FrX/N+2Zwi8t0lyo405p75WxUDt/zh8zIaYvl3k4V+rmZFxYGv8O/ARVPtGh
Itd+4JBsoV/uSPV23tVt/bcW1Bsc+PvmMhER0XRRpwm+MyP4gipL3nOTgONHes9xKyDl97byTIGH
nNyqsW9fQEltAbGpQBYY5XgqvYRh5QQVRQpTbcSZiywg/0YPIlAg9Q+bNZW6xEWqQbXsuBWlPYMj
bC1LqHDdNAx6wWkvAJEsW1gqFTCCalNyxYusx3zPEnBAKenBS0HTopa0BgnLLB2o+VLQlq3cf0bZ
g9H21SjkFoucF+eggaLoPpcpTAesxAYU7ypfUx8w6/AbH8po+M6VmDvyr2gOOnzWI3Eu/nBzpAWY
UcygWBdhNbiRfLGXnTKebzlh59D2D36Ylopd/uH6IOEu7IbNc/vyvndLxNArMIoEi0b72HanCh8Y
pCm69fSDkBfV53aA09ibe0o2UvI9PxDe+efP3szx3aMyYXNgjKPrD9uexBkjvB3VnpDgQcFLZl8M
UsQ7tgMvBaZc+IKoK9jY/tFMnJPPdFe8LUQQZME6SsZnz26ApLcDJ9zAmcxLuAaBOMNfF1U3pC4J
jGH3Y86FHQ5Z8CgRefWJg1IRDHDUWR1KsQd6QZnZfza1wKhA/+LP7j4oZmz8So1awiIUfEUz9hta
TQHxQH9SSlemfW4blF8xeTaz7DCx8L3E2NUgC0YjlDztFF6OwzpRA3cCYeOvCsUU0LC8tRLRxKQz
O9iHwqYIKUtkko7NGkaKUri+4cYyNtv/1nQwmNq8pVWsGD+hrirjMYGf0glEbicLhQMAv+lTK0a/
H34LJRGbgt1KUUFin2o/2Xy2pE9bKJsHogWYreH9XgGdMpuly2FjHx6rYf5XmGa6YVj1VVHL2hzB
iXuLEkr6A+fuTzdamGgM9ariMYWLrFMqYHY8+4hAo+XfrM3TcMcSLWTpJQo0DS7rZxrZEkhvLYnO
vSTIcexHqzeYF8X4z0dRLy1mGeSQD21I+2ilD1UAYMwhiBOwlvOcB2yK9QZNvwnpJoUTurfb/2Gx
o6wdQbitwoP1EFuFVWHlfvR78HRBMeD4UXUVvVMQvB5u4OMiAkMiFtkTeTn1nq2/fy46fFTlo+60
LLIIfVycgNY7gEmv0ruUMkIbOU0jM/S2WcMAnwQgVAmo+FEVxT/v9X1YO3W2b8NybBkjBhOojNEU
TH4S614OYmj7dh9EhEgW0ROMQGdoaG/g+1Cn2dJN3A2+xMtyTnTI0qnig4s1gUVlSB7NA4ixQOU3
erQXNj3/Xkl9LTZ7t3GYRbsObgHhnYxElK6v0Zu3pSxH59BlW8AsCSQwAlIEkO4iskwLgHaN+ujH
ut8y3/HmXpg4jUDX4Z0nBEd848qpxskOHKSvOGmvFopDLO8f37SX4Yk/jxz1Q9GcNr+z7AeMEnuA
sgqiLwJ6ZwYhtqLGHox41INSr8+6FWt9F6BjIAyRp/95rBwjD0k7CNIvbyYGE/LsOCoGygsFC2Mi
sB74BSu3345DaEJjpkGkZUJ98rfRGsATl5lSlqk38BVY9Dw0j0vs5STi6e64HPZxyyzGd5905jAT
lRGveQ5T+Fo4JZr6dkK5P5JS2E9opMEgP2q44c7HsYrqSUZDwu2TnwBSiiaNUtoloF2K7CZSrXP0
t1wogchWf7PBum3KPPogiaMl25sAwr5LCxLFNwuCz3yDd9B3s2vurc3HbvHfQ/jPsEPw7JIBSD9b
x4Mjgw4DaZEZ4WLUPTpu2hQq1o97QxpkHzLqrFR9zwNWnFZXc/qOSyQLdsDE4H5aJncVrohbOK70
ffKrnd8jQTlj6t7Oc7FN4DB00ebgu2p4eJGCz3dSJ+zNZtL1aRKtRfNmvSneVI/T1beF/bFxXy/y
KwMBi6+3pF++Jm7EpUk0ZDP74UOEpGjGPb7yPSu6mWXJb0IPYRMrLv2Cgd8KMcwrJ6aMczNVq7wb
bI1eU4HgaSiK1ZBo2U7/UY0habS/IE4KuFoQUWmm71TPue0FVlR31IwZ6upiNkIdGSB4nNNPP3Vy
+gWZsxzxD5PUpktHqN5OL7weFN+sMMt6pT/iHe9/h8UYtRoYCqtK+r6qwxhO3UlXZwhPvpa3+8wL
F5LgTw+TACH1h4AA2KHcQdbM5tLvYcxUxdfXH4jbJWD+S5VHLd413bQPIm3OgaSbF6xOTjX1iRyr
fT1v45w89pWRs6YLaVt4LJZRVZk161ff+w3FSIxhRKVqondCu+lpwAvUbKw9xa38YT4eyAGIK69l
VTnfDPQtoIh5ocOJU2RTiFVEccs4kvXi/MVJ7sXfBL0l1mt2gGsp7OK7nCeVK6CgYbCeQVtNdlPo
bVgM8VnkCXYM4MF8RkrFywQ8WZZBgnN4EmTi0+frVxJabp1miwCP1TZfbT50gPxe2O2lJAdY1y3k
PuB7bi0zpywybrMq0sn4w+2VcbeGSGmAZ2gHOVg30e8GvLzuzJoxWJVhXD1p3jdEGmxeKqW3v7hl
fE9unNXRk6vF92SrRhHSPKwFYNtAul+9rDoL+vbbGe51pkry8AqABhFgQ5LmRJYsUvL3o+hjHwF6
saZTiPAeatK3Bn4PWUD2ccwfY2RIGE9arh6WwL3VK5mqpTgB8qdq31QMVm/+WE+oeD90eGDF3sJS
x8mhBByRtWcUG8oqyfiBVOiw1QqJ7p/hCpnCp723a0lEhQrWhKUitllNAe8l+LVGCF2klAJj0SK9
BsgYf2ZWI6a35f/ryncqvGYG+xPnn9DA6PHXBJoWmIz9PtwKnf8duMoeBsI9eXQ7RwJLiq68zaqz
lJj7ffhGMe2/4Q89orJpi0BkSjP7OJEZ8DTUXlW9q/NHyjVKab0Nc2qngvaHQ0iI3MKLON63YQiy
z2oMRPVXWbb6R8jiERRjd3mC/bKoRfjyuOXSsFfsIuoFa0o9L3Ad0NzINErzjVRyY8oyZrNjmzqj
rQb5G8PWqVp4zhE6gyLMFjD7Yj1jv2CBDmjM86+GSJ7Cu64haKKEJfvIldrPUSQL+NncY3811Zh0
/edKNmajtVb2oazDDBbuIFq7OIoS9HNeSk1x9ZDMwvsOmPya/Ns8G7Wsqu1mjkpBQDNjUH8/Wwl2
SDb1b44yI3ikML/opac0uqkSda6+jvxweeqHOWgU0LHiey6yfCv2QpFxPlULSuZ3behI47uY+R9u
7/ZXBNVldse1wBkw9VBpvzSYgGAQFP5NX/tFMLihP4mmZIOWds1YkAPB7Mk0ir41EEo/SNeyo4go
6e2ELF7YSf1ZKrDYGLxv6VD1RjqoDXQKTXayx46Mc5y3p4Sb9xlYLvk0AOvByETIbMchf4GMIUH7
frL7j8r+SLg/Q69KLx9qwWTwnthExTguLUtpc2RFM4aF2AI+GfroTnXpJY8vcJv0uJEm6YeQE2zp
E0vVxbwiqKdjmQ2r4MdgNCDmtjMIQ6wMXUzqjlCXW45K3xKQSXSCdnqf+Dxs0GfiMPlpnB6W1Mlu
NizS1EchuopeOBdIXySNnH8BI7JiX/T1Ws/YGl4LRmiPMdL8hGmSn1BuzCf+KrpoQd5Qocf92ohI
g5TsTIMJEpuOaaIiMTcbgefpj7NiZZptrS5BmTIL1SGJAxIN5w2U6Tyx0qXnxiIbkhiHwz9L5q7f
4dke7y4eXYQBaAsygl/nhE4vAL9aQPDxwrdyONr425HO8tky84R4qWJgpyS7x1cs84sb14qfTKdi
Q4sTkY4Q2uE5wiS8Veasldv6px2S+EDS1HVKPujY2bNUbBxq79x1m4LDtLB6QXo2ug/n6MxWzDt6
Or/zHKOzny39oIQavyVrY7nu36GdvTqwJSGDT5fgjDvMvHX+07x7tMK1z56iMeLIPMwDnY5GlDIo
3VgqMTBzLsLYib9ToXCH6+211qz+417vy7Z9GC68l6o9KZgHQNonHukj72xOqeYwdaBlAjOnDSBP
jFUaZZUL17Db3g4pvG/o7fGJ5Hm25wFh/kTcEh276LVgawxpEptodjvX1xo8zaE5ZkbjCyEwgV6r
lapjU7gQzZQ57H27Z9Y8inVTxw61oTjIHKSz1UY/0YlkyOt44l4kSNW3R+mbQzwYtb6QRQRL5plu
Sbb3tsHSapQOSRyr9FpOCAkS2rMtygZWtaXBat2yTjTU+MIsZFpZASB82pmNXsq9bJokkv12gBdB
r10ii2ZvmGYLxtJ/meTNQIik+L+JBmypMoNLSXN4DZpFOh1ueRP7SBMAt1VljJ1LkMrrZCGxL96S
w1qwuSw+gFxkTe4Cv3DAoNaJ2mJubYUXNrvsCBWHHqdoVr2SqIDJ7a5NFuDA6+dlrmH0z4WevcKu
3ZsrHoPTAM+oqZg/pPx9uu1yiuT6gc1p2BzdPNlBmSYFG5AvhU92HoY1+0Lckb0ACSOExl8HY74F
OjBudTZpuEp/CeecvnQ+3UqtUfGzaMUlxxSQk47gm9Sug2icTRsfxugOPfT/atO3UMhSC0NS5Xrj
K6Q9MbOJ+ImEvqTD844H4kUvbFv8wAbq0WFWGJUCAOagX2K8ssg187vGitkfTlOGzHIwH9099epE
1ms7RMuGtbIQEB+CcQRnIc8GcXhIVT1S1rFCagaYuuuU6W7RQD1GQqc3fnWi8dAc+NURY3bUYJnX
N1OmBcCuExNbbIEL/72ittSmRKkuQrODLEiv1fjjiyQNHqmBPalL8A69VNaAaKYE4083cbdDDhCw
tJw27PVsOUoPutstRDEP5fk/0/hLl+ciJ065FGJ/gJRXBklL3A8L+XpdQGfhtynyLkHrrlqWvTHY
NrIDeCNfyIXHjex/waSG0Rk02sq9LcIdRSZfxdB5w1sLv5G1t+Fch3khuTHKbK8v/SQKRvRJS8rQ
hzHxAXy5YyqgNWc5S1XVYbP7IQ0Oi/7YUQxNpRKeQz4e1LzKPBbkoMEjgF5AHfj9L+ZYiJZmVvLh
9pDjyx9Ers1TDQDQUOJ2AiTySsZu/vIcm62EEStOizNeM53vXAnp5wu61IfhYzY0qu6czOitapj2
D19FwEo6dYlQxwvV76xnWlG2tBe5gtDsDHUyfKMXzSyNojvqiP6JjO5byYWgQwaBrGJx5EzJoTKL
yepXVaA/nHVx2Z72TOBH9eoTJUykRCwu2UrsnPcuEL4d/JPyTQtwvvPckOYY0SiW/v/wvdemyQTp
D7C/9OB/pg7AfcHIvIyxvRNTGYnHM28WQl49RqEp1r78UJEAYltLXsmAwtwlMrUDNF7rDSmx8dTj
Tb59PSic+7nx0VYQuxX7fYzUtzVow5VHNP7CXDlxRFsGaSJ5Nb9aNKye7eyDBbelI+stZ0LUxLFw
vvjetuzaNmrzv94fCSgYq4tWC4nP5+Fk9SjBYUTEFkIm7W9R684UmCMNV9LItLhriSWTuNbLzXsm
iiGTgJOlWIxf8iWeE5hgHpWBz0h9/x7ckymbsxk+iNyTPA+DOM25d6Ve/uyO5y9mCdoGV6w/nBon
f5S2vDu6XnPUHArGSWN7Cq9jEyOLy+1kzh9TNvo9i2IlXCoyC6ZUhOCA6LV4jvzcLvlkHjZwOEx+
MHWf4Z3vH/k8EtJCM/pv3LVi3Zj7rCswspwYtE3G71CH3R5wXDfpM5jgOKgELkAsS3p0UblLgy4E
QhGy99T/FNq1G1rQvODnobInsf8RkxRU4EFGryyVKQbHnSYHQWQzgmXCZCtrypyJzKyvyT1IpAFX
OOnxC59KIPRqkI0dv3qqxllR+BDvsOnDo8ct5RzSc+3FMiE92Vti0+TNjr/UTYBoYYGq1JQbJAwK
01ZloKR4It5J8pVkAX6sWbystFq3rznwnEDGCkwV+yoWMh/aERHFwrIRPnWTBaDvDLHN/aBcpE6Q
E5M/lw97xbuD4ZBf96WiulStxH32HDUFqBSGHt2rv8yjO9Z0KjdCl9W3BuzAi8jFSsilELEv6aTN
6H1xAedlYRTR6cM/jQ3qQ+SfgP7+6gRivkPsuKm6iVQdr9j4soFUFhu2W/wV9Z8DLibONSUV6lVE
db16/rnVFjCstDMX6490zQVBidETJKM3Ad+0u+cEyLYJvhYtU9D36Qk9WztG1Mk5/9NJ1tvqIudK
bWCZv5vCPlADsVVr2BOz+ob9yDlxfa+mVywsvOjurDpAiK8JJtH5kgiyb+kfANUMvlan3mceJSkf
70gxdfUzE+3C9Rc3zYGxNEupLrPYkVJJc9WGxYryLw/w98NgCJuFlY3u+Twjq0va5jCc/aT9e6Ty
dvQpCUQBo7G3T1fRY9NokMEs3PAnd0m+72JUxTSUQl7pdrb27XdTBhLX4goGgTT41DLNUeMDTY68
dZOiCFuME3r0E9vp60BwtVMSKrP5o0xp5ZgmrmFPBACsVSnGK7AW6JAt9xEptLu7kjMR5zsqe0gW
v+rZP1BMoZoEfDSkTeeEkgnVUMRCgZiSYvyv1UCp6r5CawngWShjiY6hAjuMwoCs41ULLrWJ6HJ7
WnOEc19Oa+r9jFvdqoK+8elS/JGnaRnpWd4jZgNWaGbEMADe2E3uolI4M75y8XjzOe0WkevsVR62
/aCfLWJooceV/Hf1248qhvMXFkPCE42T0XDWSR1yT1LZ/qsEIhj3AxRwzdbKRdATTTb7UgTTOTAu
y9PJFUHqCRqqf6s408R+KWHfII274vuaWZbdD4WRaB/thqAy6o8911PMXn1RB45UY/iBf3emzubY
lsEQnhnVwlDI+jZ7C5QEA+smpY79QW4QQLnkO8Yg+Hc3vF9xXVrZPUNKKohxmbIXZkK7fAFjJ9lQ
NM4mpLqzLixN7gTz6Xjbk45XvpMj6rZX7UgJvpcfmNd9kt7LEinHwPdJMPtMBgDTnhuHdQC4atvO
9JCZWjdwxTtd6Adnu65LUk5xXy/XXN7uMU3+OYTV76qumwcE5xNXLzZYvfRls0+snxOxs0R64W+K
wDMTm4n1W/9WeHais5PbTWXsZIhTsD74tWgOuQl87j8gzOM/nwdqShWuv1dFUSjFLiF2zV6V30S3
utr7ykpKebxvRS3pAXFFPhyl+qgXIV/Z0Yydf/8t7A9Qy67IvCisuBWig2WufMuc+FJ531Gc+v5K
NHEZZMIldPauYwmdTu7szjCjWrAIR0d40OgDDFNpIXyz2YLIrOlvAoL5CJwriPgGNrkp5nI3CfP6
TvOROJaZQWepajIkJK2vFhsxCEBRHOOBgpxpvHp5uPe+wu46nvr0a6qxGGMOBhizR6INkCe0BUCO
TjD9QzPNzdfn9yyHY/gedr/ij2CkhMQ/P2NOquICiwqdUUS7NEADAEe7+7dgNn7wf8Ykt5e5LRxN
TrH/TVx2NosHX+Jdm7SJJj2238hC5NdebrzfpfzrzGEKeVOeIwKCwJZLLNKfXriO8WysL3fHPOTR
Cd7xLiqAWjJUyKT+hhOvYiYvobwEO3/UdNAcmm0OHx15C7F0dXVMdYnlfLJ5BZTMlof4o/21ZHUB
JcFtos7ptv8SfFlJOny5maxb43tPLp8D3fvagcfYM2vwvVqEnqdbBhAETCpRp9mg6iW7c6Nc3KYN
xZrYYe1locysbq4h0IVyxRgVQV893P/ebRvum0LoH1diJ1sV4+OSIezcJUJIuLK9YL52qsk9rvwv
ZaGGtPU9oR+laFMAJga/cnELOideNL9nr7pyYb7M0D3t5ocaTBuwclCYYDAmvWxAZmI/ICJ1gJj/
9+WbPcod/3UncHZ6U+Iuq3D2dCrE7s0crd+OrCss7d2dVIt6AAw1tmwhwkl7+iBdEjHBAjks+XH6
D++RNLUi1fZlkk8yYuuKBuoYk6gU0LC8yM2Yadz9gmnLChgaBUrQTZYUORsiXVG6jkFwBfaHwmce
a/O+wIdt7DjgtuMEarBUf1DptonDG9giyTrz2otIdr/KXEa9CHVd9PwJ5oIHnlOcqgs9ikVhz7Qi
Zz5oli7UQ0r/Ha+GzX8NQqAm0OTUNi/euRLeFe4wPJL3DbCtYrX+x3VurVKz1RPN9mw89agR+8Jw
kDFccPqGIzI62U6V7RnXvetDYcuMoILocSEMyT359C3XeSZJYRVzYcf0tX4FvyQM6+Vvoe01Z7SJ
eaCxVo8SC+Jy6kpzybx1emYvVluvjpL7u53QvaUdBh+D/iFSrqKu0EJVkRQN4kmMhDno5HHGN5iq
b0bwvyr6K9UldVhETFplGcD89YBila2lmEeYaTpaXlm781gNJbg1yoSmjpNMAIuJ5iXaE3rXH9Ck
TtbuaTNYeyK4ydKywyac2O3M+5DNOr99OPEA9Kg93kv01U8TEkMj7Xs6RD3ZQLy9vjgiMVysEMBg
lyt3h+X7NLXHsPM7s4/bDQ/di+LjdwkxLsL31qRQeDecuphj3bbeloUvstQNbBZdtH9pQso39h7l
RfsKp2eVdZ3tEVpGRVbyDIDus3SvrPgE5WMIu8WdWknRnxygM59R2WuojlWp2XdX0FMzU8ifQtJq
iz4i7/56TLF1C0Xj6tlPyYpT5M2Rjvb4XsXwg7ouFZBo/f+7LsQFRDnuC9qewUleJCpK77P/cNxm
TEmIHn/iNl18SCBrqW85zwKf71EXEBkTHD5YC3rFRtUkl+nSJuSqV29GH5mrzmhbMiMsG+pLVq2T
MfjX6p8qrgcQ3gzJY+aGf94ILGCBPdwN6y4r/M5mvBbX/4coJNJSNY0askXS99/u4uWHQ8jJwcZh
ZWA/VWWCnRLcPqIEY733NDzGrudXhlhqle9RY6ReKhV0jHTczJ240t8OTTfYLUCNwMaTrx4KE4FK
pe2BDPnhZkRvghqdeBuyjPDZ2XecpRQND19fGZhEa3CbZI9JBS97jS1i+octcWCCcEThuHaFkbv8
YcPoQ38N0rXsYeLf85qSnv+xzb94bQ6mRBCIrkCsV+n3705WX9wfVR7XIb2IftULYht49AGGJT1n
6H4839trq/9YSd1rZ3ns8WMsKZqqMXT18H+htArCMiE+JXjCuwgcgGfhoQrh4bKPGjmW72mhOz5X
GjjGhsk6eewgWoTHZHDbUQeDiNiWMYAahUEy4ed4aUCXX/5E5/xcqOkQZKJjYkUFsbK+kwizyz79
osIOQLtU2bqRz7Ufh7xOLre18IqXWJKXD5Uo7YWMS9GsFJW6WKE1SlGxPpDacJPdl6ofJBZFIcCe
CjnPnJSVYWU5G75pwoZIWLB3tBOevN7VZdLjcat/M5FD+d2tipPqQgJqGUv/IrFkSSFGXwIsQwrR
HZjmrrMylY7ixh3hBVEEteJny2tQba7GhIO+DDFOH55OKsQ0pCYlT5qQWiojIT1xOCs/S0Q3Rgq1
5r6dbvGslaeHgFYGBSDlk+jeEZJ/9e1EdBAOUntQGZyMTNBmvuxH2UUuP8wmubPZZb8zJPOD0+wd
xLR7hD8bjO07+EtKnZchdLXMxwQY3wgVzeWQ6QnrVoMqCJbtUR6IRUTvCPk/FxJYbJOPHPk6hlV8
wa+GHwYj6DaNLAa+2mMmGUaXdv3BMn7avLC3fJDjbo0HsCCsH8f8fPDdwpey64BZ8RyPOuLPcIBR
rkg++8UC5u5HDl7/TZSzrzwzK+Du6xdNuqU9yjkyPCy4N+uCefqrQMxBxM4BxPLzahaQQgcHcLlF
izRm6Lvp7vAfQLIGzvPrRpDmDVakt/O00c2oZg6rLvmrfiOU7ZAkH0WivpibTXP9j2U7iR95uVgQ
N0vWNuOSeQIDl/uBNa5LfqUwoV9dqiAcEQL77jvEQTsKhqjznipkAk4/tIZFyMBiXuyF9tXKe5fn
A2zVD84WcW69WeVZ5y4hoVzIlm4Zppz9waTuz/S+umqhcUMfqSn7D2GW8z+R165QC0SXQhPhdtbI
zF0XyaisyPhKQvszT9T8fD1dTvusWhisDKsmLt5imoOix9069S33sJ+xaIApgCTSiHENYK99I/pz
rBhCVuN2HCaUCmlJbuFgWg603DlNTLu2EmWhhqQcGJKQuyYto9RBPNSLgWlRQgo38zmLsZt5e6hV
masZY7mVx3LMDQOuNaF4y7N0D+FbmcPWb88t2LgtQDaZG0p/ZKaTbtpyiIV8kCvOOARy6oyJtpa/
0Mgl6CnEThNbkAWX4h0RgOMiU56XRuLoNUO48o/SOp6FlGEe50mC5HRrg6nNUs6MHAxfO8K5eq+S
ekcHnNYJ/JZkryUiQ9ToRRW0LGkcMsG/p9fSM2de5EIL5LznUYuh+/zKN8GPgixx4tN8vMnPKUx0
oWopmIHkmeYPYPFWNP49gQRKud/lTHujFK/WFJkY7qeRigZO29uOTMOEoJP1U7XNtiFOKcdbFUHC
PrnfPbtZjDqqhiFpQ7i9068jxpjkNdLuUAuGfwIVb3301vMDR1H5fGMZoaOnpdREUMc9vIN6fXsH
kFyYhgw8etPOoqyyXPr/frYbuzzc8O4QlyOmjnL3GqhT1USAoObwHDQ2tCXHN4bE7YXhuwSbJwBx
1mhdWGKUS3Y594EXdcwTl6FyLxtfP+H67ZdRld2hI8MDVNn5o5tuUpXT2626pNJAifACAaXqsozu
xq3F3w+I2RjXXm/CeXpkLEIMX3d1RaY1X42ijwLKIvhBYgGM8u6/1XcMKAS8NC6CxbaZIux0Y9Zy
UDttEbnjFiAJ9HTdLIptnQj/nr++gCzwDZFtTAFPOqq5FzrX3Uz85jX9RnTu6fhAu+WT+KpHzT0/
B/MItHXvHwe8pzNGsMimc85z2AGVAHxj+O0BVonubppfDFhmOU/6a4accw4AWcXTnVntR8T4oklr
MQReke3ZGLVYB71Kr57us6TDQotZO8V5lc1jRGg9KLTKmpTCRHxVWEFHjhZ4m3Z4j0tUzvrlH0Gp
+d5rCnNftJEMRtllHjRzuCNxkEvJgyTIFx8AaSi6k2WQIf3HdHqjOjZg8733d0+dF2bLGTbi5zmm
RYR4VaTsYt66HfNmDWDQhRHsRru+lpCpFIZ/tlvrr7Vp7YcHDtvZZ4EkpF+GiaKoGSRFn4drQx0z
hzgeJ1eabBaASUdzjwKyEE4wPxP+PyrjmBT+TG1QMKu5+WCezc+8PLjvO8XSfNM1kMUt/IX0siUs
cZ9zak6GCutD6P+wZQZnx281ZC7/54s22F7KnZLtvXQ6IIlEy7+FTnP87th70Pw1rxbcUZmF/Nno
DUGAwu0PaEWjp7k8kopDtFRTEmkDH869/mxrdj2/t4l2pnliiaIEzDMTpc6VqNzRwWNd2ivjBo7K
+uz4VpsVIejyaNZ1zSmeLm0EbGrVzJ/v6yJaP4BW6GC1G6MMBBQlj14QsTwW900Mj567cBzBTG8i
fm19J6+ltx/kNGZzzlYF9+wxfbRb/f5Nngr/r0Mmwm30IUdgakyOSBKdT6vXaSWayMbOjxTDdQVF
7DeYSXpxB5DmFKn0oUjsU9zgXqAT7B82sW84GiY4AwpBx+B+LPPqfVHu7hA0ncNlg2VN77MZGW5k
JckVuW9SJqdAiMC3ryUblfIfg3BflCPsMp5eigG04S7x5nyisnBEWbK1rs8tMYfzKqoSupsH44gd
CJaw6eTCGP29/5eL6g6ML/XF/8wUPZOSxt1HL5pxNblhd+0TEPT30lHa+hfIDBJo49Ljwb/krW2s
p1X2lcd8fGr0lCHV0K1nxVhZ7J2MO1G/BOjWNzeK4s5loEIBmrmtKeo2RnwzEQfjsy0WHyNCSw2J
ErNIcTV3rRnKBnxhb2Molq7muMo5icbkw6Gtq8ckTTPwT0Me3aUt7kYp9wQCGmch2XaDRiBZBVNb
Z8AnuD6oEDON/LKpH7I2/jqIJ/fkuKzwNdqpI+EaeuyiT1GVMLpiAyfuiMuGG6DwMKQCGLBCLj21
kEwzhSrFakO3WareaLp3RmeVRpRTH2f5Ati0V2lO1fe+pfzVCZW6qMNOoSrHADFHI1xFl/XtyOyh
t1YnM7H3Af3t0MI+bgUFchTw+Pv+q+hVGq5NPDGpAmGmixNZwjCX7bdJHcjkpT8LjJnsfCHBPAQ3
UVi0xn/T69ppscEdc5x+mj2fxLuqG9gGMnNn6M/p4YW4BOR5KfI/S/oJImOlqzxNjfXMw17hcTzp
7CjTjZg8bsAjN90xo/OBxbB3XlEISzA47YhYTYPSng19fDMi/JBMtATTLlJpMUOm0qrT+wxj4Gzj
h4tTkUIypr802YKfz0V+xshZjTmQkOsSnfTrQcBq7jhkvFs5OMmAe+jco9HoLGRXMUBMU/MP9Bk4
BmWHdeUtPHhQxBylxXhib+rMClLiTEpLDAfQIBYkUNh6347xlmaoo+Wa66hK4do82vDPIWys/tHL
hl3R+6oUvJnGu1L3zUxU2hq6IQjp0Cvib9LB9dCR87fxw4Ddj1JxrIblFR17QdWfaGIi8Tuo9Vmi
glrOm4vAh5MkNBIbusDWZqiBtf97RI7+GV4EQbTR+h6jNzXh4qOXHuM/2Lt+Fm6g45hdb+cLVt88
9RSsi3p6cH17N6e8reuJRXXBYhCXdywXEPD/vc+84qJXcZyPUUkGJ6x38/F0//GgBNX4dfru9q53
ab4GchF91+kPDKm+8UdeaKYDBd5WFIcO0HuPrBXi4NQWoifRnXttFnSlk42E/esB/+Vv6uL3gJda
NdqSypgAtFKKE6N2ZmYsb/sfJ8+iJEsRR7iiq2P2G9BBYRv7eS59aO7FMlU6YxbZsbP5IiI6soF2
1bQmP+zn3Q7DXH0WFT9F6izTRunG4K1fruYK3SFuQ3b4c7hzbeKC7W8EtuHkAc0rgC5zceEXxfTa
0YkQX8H5fgm3LrTYplc1d73CJFvLGak/fpuQNR0k5XhIkHZ8x0JU0LiQwEQYnG323YNf3ti1MUuH
zlXNpNu1pKTP6tg6+adyg2Ejq6DdttmTgw0rZS9kkGTe4JNwiyQbfQNANu207a3pDDDOhvqp5yDp
/pHQdDtT/hqIp5ekdyNpWyD5fPzr4F+3VWMOxtR07myCY83UI6CfnBZk7RZn5ZKm1MYPk1hnAl+b
iJwwW54GxlIFQrSWmj93JHCoSGIQ0XUus6CTF4msR+F0OsPDnH7b0x9N1Ya6nnllS7nEDvc4wl0f
ymnMEv8YzN7Z7mCUU2A/FQDBW6d7EqlJkB7hvv2xZ8Nlqp/oSPc/I3/wHHk+l/yLv4JGciB3TOOk
Q2mM+DMOGppt/S4tlLKlVF0maj72S6qs8NlZzfYIYd2v6Uidak3GlDk9Z2EIbB0Bw3uT7xaRDY5t
JFgZAxrITIpv/ZwH1urJmln8aGSmNCd5tP4MDRg/lgW6TXOk1PKWoYuZQ2FFXhw0xOKnf2Y7Zpds
VK5FwPcYSQPXOtrRQ10CjvFRBafxmUaXa5zFzPdC/+K6SJmhhZDHAew/Uj7RRsRlzpCV60wBdrUL
nnN46i14n8RX6EHGtHfV0u4OTuHMstfSJwkAjTHkyTKR53QFlp/BZhFjneBEF49tTW9cmhRpXhFx
8NhFIkjVjRrcIYXj+x3M25+6mgD+5s37IZ97F02WrOFhFFI9fLFAGl4HlV/2TDm2EP7A/4iVgzm8
or8QYevZVdBhnnOa0vGmMXa4LxLMr/LH8DeuVuE05HFTD+jIIXZhbTSZXWojyNNztCtKSGvZrX8P
tSxsJkBB7UNtALbFN1VyN2ghHFUMVjBX6yCSP9INet+NpdtK0GMMzT2Y2jbeXmQzh4WOechefLYv
88Ai1jkERdSOrtqYtMTFf/bujAmsEyiWbkmVU3XYYg59QbvEJiTeXTNTGqQ+uJJr0czvrU5UMfcF
ydNkL5KU/+O5IEJAYbRA5oYUX/BG/kk3difS6pJ2NrkDLvSp6vS8IqqS5cL+4dRzIFUEy6xe9AXi
XBCSoXo5um32TYYrMwx92h3OoDrKnm9Igpw1S8MfLBEEDlgnt32xP3g5+sRN6sp/qklkokv4eZI7
JecronXvhbIquBEWphvWG23L7j/Gl2eSbRyvrMkxn3NTIqymfVYVsmm8x7KCXcLydwXa8xw+CLpD
N2NHk1EvFWBDk+41les8cylymtLpB32uXlFh8USTRkIRWA2IwIBHqmiRAOGG9z5b9jznM2LVmcX3
xasMonJ+V9dC13bFYdRXqG1dp5DFZHtusd8F/AeuQejnbVVX1dyCfv1YCPJqpsr6ky1yy9h/aLj7
CCW7qKmk8sNLD8+ZSUXBLgtCyhpIv87IvNh3XlkfnkPaBCSqpIr2ZcH2pr8nwHq3b5J2poFADeAm
xNhoN0/f96f2fKOIguXnjXo+65zPyGbtVVkY2xB6ra/gGOhXZQbwlmVq7lesiTUs/kBLVXMPlFcy
WK6uWQODgYyqlq42GiY7nZkdLKTGr4Myi0brtqBj5yPL5BSomuakek4at2JdtjM1r60jWtERVJYF
hugHf7k0PmVcWohCwBh2fQ4F4Cycm5jOY8R/rK9Lki1N4n6+OWoU1HaqFFJrWxgxwdFH/B7t4EEu
4FuMOl3FIzkMbeTGyO2pn+Ha0HoLo1kicVXjkgj7wI1ZEiHaOzdtORG6WjM6sYDRKlwNKKMc16SY
8OymkoieHru4PZ0W4qBF8K6MvulgXejn0Jk9G37i+uBIn9ERqZ/A23uvJGcx/xyeoxngrQQHCmu7
fBB6TxCvUObssaSnVK6BwRdezZrwwVTb+Mnw0XQg2TpT/LiMeHLRelE+p2FSLZ+CiiUZfY9YUmuO
P5eCfUimJ32pkN82WMt+yyX8pDj8C6tzyEEB8AH3xRwLwmN56uc3saN6kE40WNBSf8MV+L66s2PI
Xo1N2s+0q1Eoyv6kH+xdgjpjMLlkh+btOaPEF7LpACscNvl3aKL9uYGWDxou08UkX3Ogn3DqyFH5
pjvTG+7n0bO6saKOXrYaaapklFhpBLqO3XLnF5siHoi9kuNSviQnYCx2JunEyeJWw0u2JvBSgex/
ooJ1b9EtST/aaq7xKh3YGWyWtPB//I1ZICiIJCeTv9YNu8EWjZ5pEmkcfMZNyF6zHFF7tSagfZnr
rQZuwhiTXN9JRDMirEnWzDGooahYwwoGRoFKEnmYfoEpGAqx+tPAakeSHZmkXsxTYUL57DXLJsmF
/GGkveEL5WQrBMm7XsCbyfdfw0KhzujJFEOdB15DWANr3fPm7RrK/DrPLbRI6H3fYkULYcQ+0B5o
mkR3bLSk//FtiSnXxWo9nbqCvnFABP7YknN+YnAiQIL7sz5A49V56eYbCNQZEQWFT66v0pmoPXaU
IkxoXoQMS1f2CBkyue+516yAxHboSzdKtsXE4wBpHeK8BOfVCNZUu7YpN5Bx09vu2IKCXIqyPKYL
Oym5igQA4cHwFqh1UUYJNS9UYPtOY1AWgIOsd1bl2XKSOFQlvqkYNiChR9bjJhpWPihITjFLb1jY
Lpsi9p15REzvD47oh7vl1VEXLdNFlZZDbZGsBvNAixKDS8M3386q354oEXVdvkDjl7hNTARlYBAl
UtZrUZks97kvmdq7qKgxl8r9pEm2VLxQtG2k9sqIgtiQ2g9gn5FQ+bbBj16EVUpRnNakUyuclDdE
IpBrSMzMsFnTg19NXrOzW/pbuZw84gIPAh7dUYY7qgb5R+aFhwAuS/gqRqWEZYKgK3XktVS6Mr6r
X6FxjaNISDd5bHMJDF4YPZV3ILo33vcbIvSKOsoEKla3nDIhBiqmiUIxTL6zQkXvyIe2/VpedmMX
vBERikT9lzanNsyjLFSJfK+gRQjchUepyDWEeey02t7ondU5aWEgm5kR19oR8yzpQ4HxqXIJqVmP
NVHh6NUUbFYXtKUEK5iq2rlSwODWPFueOxNZUycayY9PthvPs8k8g9rVz6Pw5DDbgalrk6Sla8NV
wViRiKbIc+NnKoHQfWDBXorvYWq68QB/qk5kiizESh70t58pLPMxYI7XwA7BRyIJ17nvc07H9/Yv
M6D7QWcja3+OsLkTVtl/VjDZy1ZWvNwNaz7LE/kRzfFp5ydNZWUwPgKb7GykdGCR6D8fiVT1korP
84+cILZGrn3pTqljOP+QbDDZW+3yOsI3bB8btQjvOjFUSTjm3D/W1LQsAuH4MWM3tzQUi3POlbYD
5+rdJZX1/I6WA0oFW1BnGZvyY+ZBuTBbUt9Er5Z/VcrjqXRRCtBEYtRxsOI/HUYUUgnj0VnZL4TD
827ugriOuhdCWnX6R+QvmuAp2IHhwYJphf/Lry0C6MLMKVLUBV90pvXyFkLks2B6QYE7Fv6Rwxzi
9OPJFXeia96HDQKZ7s0rWXHYYPNPBEEflfOpSwfr+q33R7gh5dIM9Ktlz5vV0S7GDdPmcxv+289J
OvfWjlhXPhpZLVmN8pd7hXa5A0cR2Fc6QStuLQrzr9nLl4zUdqR9LCziarRs2ShAcD23RZLmwZRX
yWO/PxaJczfXBgrfMa6BhGB3qYE/Qi58pdmh3fv5UNGGlg3eusCZusXdJlCUdNVV0lzYWt4eis9h
Q8E/mXVuJdMW3Nqcr+15rYDXwykXZiAWrhU4noPePOVX2dsMHfe285g24Llk/VXMp/IkXIxNM6zN
EWOMgr/izG8dbBFcIjcagiSrhmBvMWxz/PM8g++00XYXKK7FCX0dE75nSfnSx/P6R5F4hfcORAa0
JTf93JXLaJjBHnr2QprSA3YTET+gQ26ADF+yHnz0RPOeHh+Cn733JoVnHXx/lmS8RGD7mRWOQ9uh
CHBTHxuNyEFZd2+kSFQoH5GDCCzYjkH6vbKIckRDUHaSrT8nk3Zhvzzio73NsEmEJ5iFavH37ILh
lz3jf2m+EoFtZXcUlpQceQQ5WLa6g0YWbOJTzojjZx/GR8bEmb1iA9sjz7JapNNUw4NSX4ysmkgK
r9zhQgmA0Qz3naZ0MGpI7skQIZeCvQeBaLjYhcJ5nvFQj/rsDXzbIZ3Ig2RNc3Yz7ZBvgpPAr3Sy
pSc3bTWabuUWpD+njB/mrTN+qZJLYlD12R6C8voDyxcoTbv9N35sz7EeTVLlelxPJxHTaqs77LHt
qtvMW20dnSiNJX8qbXS+UBi2Kq2mIieY70O6fCmxMz9cY84byyYvSgE4hNrM+i2RpPaUDpzUnxGY
GuWkOgMgsnXYJJ/kFTgPkvpFWMhiemTr7yqUUVD35hp/zX6sUXDd4UzUu/ouVcOGNF0KK1DPz/G2
4b9SrvDa8qr+nWeosBbNHt0xGqchExVzV4UUQB3F77MnnBd1a7+o/qnpN8dF8UZZPkXBPRhMQf7l
g7ur4ot/5OTJ6uafJb7+WMIjuZHfyl6TpxikTy5a5Kl5SI0+XGeMMhhhgCIDurdQ1pcPanqEho12
4l622AMAZInbHghq/7X8kHw1o1N6/LWxcRj6hEhPz1W3Rf5lW9qGSaqdnSMFyju79q4Nx+lQZb6f
3QwEM1Q0/nyiE6xSm8lRSSBGc2POqU+Q+wYYazNAajbNjSt0nPlhSQcOwf2O7CDsdtmntxLMpJyD
AjahPuAkCvUa0tO8KzOg3Si2g+DaNJ5v6eG+1W09ziUqXB9fUI1jgLsW0YV2Sap+Z69o+wjjF4sR
Cr0LllLmt4Im1sHiJAJDpa7sJo470mqB4w0HzUWjmnlA4GEYcgMptC/H7jUUMWgzqoYRojQsmbsU
b1wSaisfJ+VVsdrUTjio6ThG/OMc4fkJr0buV6/HKYpCf9rKoHyLUxZqRkpr25dNH0PCtR2FYz9e
Te1Y8z1dqHw1JIGz0+RQyKVZNdgQfXa/0NgZxaEYr6bcBp1gpay2amSs4vYxrcHljWrQpsbyhYDQ
MolPn9kblcjymzXNtempYBUT7i0OcYbjbKhNr30/sEtHuCFI67OS29fI5EfQsWsCFLjdSFNgY7vA
radc7AlOmcXf/h1ggFuMi0taAiO/cK94V+M1HgrArkDeJmSLClEuuuKZEAR21O+umilE5LfwThG3
FBTih7bwDSFwxOrATzoml41VBwu76d2dyNN1j7LlZYnTIYLuvpypPKFwStLnIxZZYbk8iq9T4YwF
Wdbq1Le09bFM96KY3JADZcVVllpIpsQPz5GF3gbJTBOr4Z9o0DZ2oO4DYReCGTwLztxw5pkpxjow
a8VpLfezDDGypQhwr2iI7FCDTILiaEfpVoGHJA9/FObGbnjfXbxYsqWfOFAhGYmGha/fwhy2GDBI
bwS4rhsxol9qxJWRUhmKDoQgFh41yDrOfsPQsetVvpsy6OLPMJjOApgk0zrcP0wWmmSvwUg8Kq3z
NZ/55DC5r/bLOcAFNGa1h5s43sFMO2oScwr+NFwgarfDz2ycaf4dRGlW2kWUeB/Xf6iZQa2dJcYQ
yrE81jDyDojgu09GewIJBdjGtB/fdjsNfcMRZLw/3gckgLjoMJdpcQhR+8RjbjUI66fjFKnH7gu1
LuraHfoOUG7Imxwq3lT/WYhRnBzJGZqdkqo0O00BLfrdoGacBWyyM5SiD3ezpgqvVreZgi0cjM1s
6FFyq2SbjlaF2nCgDLxxvvzYNB+i5kTBcCB+zlA9OEsfoYr5pOQ2rmR3ojDbCywnd4hfSPIQ1NU/
hRIYQtW8htYVBSSKstFdZnFhtBbpJWOe6C9BQ8AvvnLcooW4T93Ij3EaQHt5zeQ/ved+K/d5LtNp
R9AwD0emNIL70o6vSkw+XULxdPyT2K/GRlwl92ckTg/NjSlCIT0imxvSCkDobNAzG0qHatX+BvJY
7dBC0dzYVKX6E8aQNUVu700wBPpVmwwMUw6sa5mSqtSc9FDm54nc+Mxu0vlz/FaFjuq8LrXbHY9D
ahn+66f2pTgkGA8aTC2Uc7sIL3VYt330G5rpiuSp2QkFI65VgRdLFlly8/RXs6/3+WF0JDLMgVzR
2TNNZiDkVjGGbhRXkmrMje5r2p11S28uVQeEvXsQ8P/u2Wl/1TcTXwVK2EHi0KbQCaqS4vkzHGIc
l9P7Twzay7xRglj+jEYL8hgkZIN2YRK9H2SijSmTvBQgligsAhT7YeplVVEy5/0KPjwedgD/EBHc
gUzrdxS9fD222DYTrHyttF18RTqXimp+ACzqv+KHWNE4VncjJxRSWnFPZHaOkynEl9Ik6rX9Pb+9
0zUD7lLhgHuSKLPhnYbZxnRc1zPoKYjC20ybtUzSsWyJ3iH9SOhD2P1PYl8S4qqEl4505VkFN8tw
uBV0zMkU+b1EOZsEB9q88J4ZrGY4gST+ECa3vKfgUic/Cfq+0SimiMAA5FNPl0RMe3f/MwOalmKf
/3zKL6XGHpX7bLPLcE80TzR2sh4POjpVueZl3g/cz+WCRFNxupC+rvckf/l1bjYScIE9TypIugAh
hViApQi0blWGhbQYYGq05xviWr66EGScs0NmAWgAixv978Pd5ZP/jm8eh0mJkXL2Q9CK0n08qcbv
9E+YhbZ8i6uTG+rJ6FfADIqZJQpMugL6Wu7qTY3EJbVw/wo8BVLPTbrmmaKhybvqDu1BaPArzAwx
FiHQxjnjYRHpI2UdyUq0whgp94wPHWi3gIg2laXzdl+U0SZm1EYr2YZbM9gw8VQD9DqV2LJ9ygnz
LrwJLWTXDwpzDKtiKM7GHLpI6jTDkmWiv2ZBgLmiTb1OfOTYE8Qem8TGap789dWYdNaCYhMxOHrv
SgMLTdGZP7sUT6pDJjo1GTEOd0jaPbDCDQA2YzO3PYvf1FwtwrU9At1pHtyzqJXhkdHmb8HTrEp1
Oq2tlKvCRLXAhh1DiFaOV4gRgNRpI07SP64dpT+fggH612UnC40MlpDUgW+PcFYtvU08DPlPTqML
en+/LysJ9o2tvVaYZuzfoDpANvmdTKt2rnBECgSCddQnbxnnu0j9BazYNVIaazWyfC9k84Q4Lo9k
X/hH7KfTJO1EjQIUK1MSJl0+qXdqheRzqG/1IjKmIVzLFBHFQyxge2sqR91zymEPtFx5FcW9ybXp
1TRmldimxlI1qW+liigkDFHLrJ2Np2XJ2ar2qH+h46m34iQ1SXWdyMmY5EuHvdNzczZBvXb6PxKK
rEiyY3XxTawuGij/6j3/bav3CUKhBDjdyHHo8JaWTEkgAhWUyuedOmqYTZm9xgSCB6Of9vSTiGyt
/ljjz7s9zm3UBvkeieknugfePgNAFZgw+mU3u1EEH6jnrkvSnENTiWM4qkvIo2AFecYNmHkIwaqM
jYeq+7+KtTMOVBGPfgZcvv9W2sKg1dJaXsz7gZLnwHrKTTiytklfDVro8SeBXPkWl2eWI3QOY2Yh
xid/vUuyA+Cd2io9XhhoCmfje//T9nxQj9i8JpLBcyUB1OHNmYBLxyLaw6xbkfuOSyx8lQA5W0Rk
G0Af4RuVLA+gKRpc28i0yunIFRAS59UEGcib/A1aZ3WniQxdCPn1U14sINY8/FiS1+yXGOhLaDc9
hqdzZ36nNnLaKlreTB/5GwXltnTnLGw20f1LcugIuHF5dREpsEj/CEfeUEQ1PhclOCcKhzCgUVds
r2RePRBfoTxWoS6bIlK44bs67xjOi9GLeqNq1KctcmpMTsqCH/pOKu3vUbzY8dBgCjU7bzKWXAKn
DLG2Jow0LCpZtnMng/+JJBvXf4JZqBFbbxwYBf6SRvEhLxL2BMAqXBxP8afnGVj3kwAk2DM1Y6ds
oFREmUm2AclrBLmctAPoccoAjnw0z1RzerQY/G/eBtrQCdUAUQ3vWXl1iade34U3RUqcW1DYfiTV
D+rSLnzaT1dBlVO3Em4KigoiShteLQ9TgNe5mA1YvbaYgV6+5yP0ommExguYutiUQt9MGoe7ICKQ
uUu7ABn/rj/HTM8MlCwYluBY/F3AfGJr2P0/BTcBF24VFRkzHzp7ct/eCyrsPB2RW+nbe1xwMGJ+
FNo3ZZoBNfAUkuCxEiIS7G4fbrkb8uZFl1j8ANsgGrRmtwmd9J7b45IzZ/e5jgwwJGBHz6Qap1Sz
qJF6kltMXsoMmFR6kaI4r1ZQ1vmyCPYEecZYDpl0XCu5lP9Bnwew9anhj8Oeutn++VuDjENghC42
v97PIcDwY/0GQUPcz81F3shXbbtJUjFXr2biBTWnEa0wFozv8HsgsblI+ef333eSA0rI525tX+ST
LeHVUzfoT+x7s3NCsuB1+02KlI659injKJekm1Y6QfejRY1Jb0cvxtH1I4kA2eFBHAt8E6i+w2az
x1jRmFVSAiqmibrhuRe4LdyjS1WsHfh/q5aT/eDWqflulsqdNfj1ZH5k1KOfU41ZDekPfqaQUKXR
0UXDU5p0b0LXvno+9+b3ga2oZpAQDhFvqW6RwiyZSX7pVKF0U6ZGPUf8mMMIu42gZv0G461ooucA
Bss9ilJQA2d8vlvgl9TZvwbb5LXiUhBxXODdkur4JvOIpNaeosdvQcVNB3XstixawlbPGnFbPin4
dHcneI6fKhNdwccyKkShxGIJUKEaJcoDM14UuLQ7XRsN1g0wCcWe99/QUkV4ellqwDjzzJEAOCbW
KzHDd8G/1apoJV78oAD2O7efSRZbFf4yl71TkTACYzosO+c/1MJl3XbqaOF/qy3JfkCwEwgck1/H
l9siqzw5Y3dXA0Kgi8/EDJc3vuXTnWrF0unMaII28ifiYCLclXL9APbUOSJemM1uAcMbxxfxdQZE
zrE3gu2ozPD/3LNjrcF6zlmzKkpfyx9rmi8rOM5ocresngdHtoW7tYCVhDO79fE6A/VnBhlcaWgU
kFqbte2fAimapf1tq+veQM7lsaqCyg+57I10GTcyjjqvKOLy2WH36vTfF2pCWeZvAo6vWoixOMf+
0qLiGUp2woqHEteWw91hssErmx+BEgNIev8RKnKmJ+K96Pmy/cZasNr/j9/23YZRoNd8mZC0GMU1
xz444J7Hqnx5MAa60zM0/viVm50wsZT4bSFx/7rF3UyIggQQtXzxdztyT/k3PhbLtO/Y5y7pbymY
ipheRy0zjpM2OWkivrLkznXxB9xG+23Uc21AiH0CnXXjpoiPKC0nSh6NrRS7t+9/mLHL/cEWxpVF
peXMRwc+Dzl4iLbQynzGPb3aCumB1lLQCV+gOBHG+7uq9f8HmvA0Pbv8wwzNO2zleBI8pKNOvIVO
7nQzwBxpPsDAc//2mF1B+uEwkFIh1CBMFw4wEyXPOtlOzBCFUw2jqvlmqAQSAFXVhZYP8zWUzSJJ
FiWc3Ucs5HkETe1TusKE5eMw7IHKFKo3wdOzZzbVYf+PrlxpE66+fVecF4xLpdWhf2H510UFF4RA
+LXDT522QemImsftRXojDVmCZ1z+z4RDLjIjpI6wA+cOXVUIzZjtWMC6BhuTuPvgbb0CjcLf1ZBa
Idur3HXuCRIcuqbgZsFl7YMStjenYsF40556nbo2xZwsqmbWZHMwzRmVZX5IEwsAbi8YnYPV/Alx
GygAJ0oA1hjJVsZ96VDqR0+W0bfCg2OQkvWFbcpL9AklTADugOy6o4Y/LMla7Kzp9Hcy3Gz/srkG
NZYbLJAwL+zrU5lLg+0xWxVj5w9AJO+Nj66PYBXCyW4gqSjHJcFE/mG48R/yQVZdGmKLl8ouEZNP
cST0hLUbRsdEWTkKxvmxydUrAIygJZHRY/FR73bHUqobiCJZqi5ezT/vqJrrO63JcXXAZBdYRYUf
gDkg7RPr9jqMEZQL0/RYAlhhzrbFmz+/eRiz3HqiU4d8Y4hmRTp/mVKMBjqn0wtUEbRtoA1eprNL
ATMaJoi92dLFSB2935oxKPPlhrxyka0DOIbBtl6mEaDxFz7szoX9PlwDiQt8xVQbVgaTfYZZJnBF
DTlwK3KRg0jLkViQqekc40ZE9EVqDfVo/5R27Pl9YM6IV5UZM25YAtUk0EcqmcR+xRh+uVfezEkD
Ve98o1z/td7lTnLx7Wiu2txG0lpsa9DX/IHJQDTK2CiaF57aNiuGi1kj6jQbdlI0EcGhpiBqPKQI
TmTpjPkO8pTBK4X4LTMQtGerD5FrGpFGcRIyaawGjU+C/HPddFS9tqnYaKuXLZdV6kHXsQJMDgbB
Zx11Z7Ud3jCoAz49MyexUzZjkA1YrxCjUgUPGBV6Ysd+RmhFa/atM1IV4VkvSzVjza5KLMJuLVSB
8ZqZmSX315+gmEI5X9xSfvTp1UPHCvXdsRsT7//ZU0ZUKQq0T1JiAGbF6IPXhHuFCQ3mUy+Y0UTa
wKmQeddXGTQeRu0PSsN0/g7hTmDJA8OaW//5ywPaDYOi128fAQQBONmqBnWWWPKFa03TYEQsHVVf
AIqXJEbp3mpis/W1Tkv9lSjdjRIVR9kpHDYL8TQQ7hr12GOJ/5YW1uybFONgzH8a4CveyBV9gt4t
3OdTR5+aJyF9H3LLolR9IT4NTH5UqDJ9oth8Bt0ZX7WVu1U4qX97aMMgQMyPA4OWsCJkxqnjDSHc
IVGLTGUpAfm6hTlvxD8k5FKOwqzWTlFIy1Kj359Y7mUBoo4Yd8zb+lB2tT2CiaQlb4X4E7CLoLR1
dpy/K5Gh9uHoUW0VsIrsBTqWpUbeCWfd309qGAuixZQDmFmNPTFj8dPZubU237SQRDbuJRm8HH4P
SAstzH04KeXktEkUgUXEajPERM99zRSee3qoo4SxfJ4zmQ6iyP7Yw6QwbIQSpaovzdzyFgDOL6t8
wuBuMAumgxG5b6c6mThP3K6OnEOpv6ag14Z6L7FUGz9fwYASapYgRbyfEymbKuo6bI/Fs+76dlcs
vthHy0Z7sEIADYVq+LtAE4zsFkKGyvU3aPVfJ80sjvq8ncMAhOgfRucSykb+RPIyiG04tWM1usqv
umwln1oI3evOECKJyG29HdaiGNvi0QUB8JlmRvDUFgTVTGO5pdz1zbfSfv27Z4I5fv4FkmTCmFa5
km8/psQdMjmYA+VJE9CQq5XPXHSU3QBM5gi1TSr+CvWyrU6fMsI8MU5NOi1veVR7rrcgXuE8VGAL
r5/Phtqug1dRKZO39hVtfJ4qmROulNq5754PAn4/4PJcpAGwLg9j8tV53yMa1QAY/2c4B1mIySIP
L5/Fp0p3MgnCSE5tmMSmAwDFCnNeQz2MHZjq7BQesg7MEumWKmyt9XCs9DNIsmnXfg0ncuBYDqG+
nwMth1q/dj9onX5gcYTBesGUGgo04ZvALzoRaN4jdTuFZ5qQasI3dd84XtjS0fZeWeWCjDKRRa1t
JHGFvbcClmXgNLYTUjPY1pR5UynbD3Srimhi2kPqa9mJDcmy6OfX0T/d6twCikmMHWnoIUM8o5Wf
C8UCzd0wdMjv6dkXcF3d6acCsFjfuosXyHU10bR5fN+FC9gh6AziBAjgLdN7whU/72Jlw5Cz2GC2
DQkhyVmdy/dyLuPrh8mf8h9ytmzBLv77wial6HGvZCV+rH/HtN48JlWjr0Jyp2RqxvuHXA/wAoU9
rwoxu2DeFCazBhfbftNc/YiDPV++IuxWEZ4O/NZ7MnzvUYhHDTgY6YrdOEbTHtjveC7Zr+b9peTO
9wMXBafQkonYF6b5oGdsFzw/Zfa854nNJLaVJ78/9xP8ewzWWcZdD40mWefdc5htF8AfDcyvHgC1
ebNR+Q5k0I7Wk8BBppdeeglcijI0IPfUBbWB/RPpzP6ycovV511Wavk+INpOL3tmvbsgrs8lsyke
eQ2W7w6igYT9NVh6iw7Cg72eQj7LVtXRDT/GsXxX65ROoaIB1VxxOiYEhF3KLlUq+QVUhTe8kIrn
7IxLv886xrdB7sJUxVNQMra1sgfrEd/0nXzhrgn1SVDPqTI8MWnRBddI+v0CCof1/ak2De9YnNc6
rmt85zCYeyn60Su+i8lLCaw6O/lZmSi1m3nRtbwucBst6vV+sHWjgD4SzB0yz2i4KbR013lHD1/v
FjTQKGUXWMIzx5mhKmAvkOP+pOqKbmrC+rCCBVx62Gc2tHp5EMB9dESQ8knUmnkk+AiSw+ewdnly
Ff8FD4aVEeMbE6VcXYZcKq8GETD2bpTi6hCTyPeE1iQyoLGfn3riPfQSuym6HrC0SD6F3zuksKrP
kVAefTBJl2GWitJI1c6J4Z5HRwz1OupT8ClYqp9xbWIXw1o+7iKsiaqPQHtMxAF8gRDrYmBKxEaG
YpYOjarp04783lMmPooNMKV7NkpgEfzdmCOWMCJJ8TVGq+1jlPEcbw5wLra7MLA5XloKplX9gQO/
LiQUYSIFu9YI6gU5xrBtJFpG3QXYvcs5mn2ZJTq2V0qfpmrp2TmK+v/NeCiGXomi8bz8vlxz5vej
44TwnHVGu2Tn4sspe3QQBVzTV3y47Lrb53nwbXQ1SxpGKmo1MdD7iLkvZNnxe2Kb2kmyDAAOPGLI
K3YsZTtTolVy8FXIcvMzr9i7bOPwFBJwwB0NtHR1mb9OEyiKhhAHUdSSaRStVNSCCpKNZjGl1DDq
bBQxjBnR54fYk2WztEdqaY6EFpVOXweaPbkHEelKu/In5i2eJYNjXs2wUZHfEWsixATCMvJtPNM8
yxNy3XFx2LcvkCJbA2M7BIzOCSJfa320YlgSvlRihKVQnOtPqG7ruAngk/2bUIc3/I3Pyh/sDXrf
TRV9SQ1prRbSG1wTs0RRSdSoS2oXin95lKprU1vJTRhJNSYZjNOyR/08w+xdoigUlFBvaFssn0X8
/KOcBIRY+0OtC/zvn5Chnxjdieo0AfrCwJBPwPHV9ia+m35QmWpIOZSAa9z72Wpxw+VRpv0d/K+2
GB7U1KvAb+khOtyTng/YtFBeb3xgY5UPN5W8FdlWHxemF+tm2UserK2h48WW6vQDQb+flZ+DRLQL
v+XxDAnRBowp7Ymg2WcbKNEQSgmDX4HLh/ZNQVT35icbaKUT4o8WaVqgz+/rQ51tx8qYr6nIVHip
LlcpX/BAz2fRpGWVfx58TlvFrXfBWlKMPc4CRq5RZ55d/ItTMVSIoV0hjBAHQwh/SBx+8eUHeigu
R8BrwXqKuwz/ay29tkZ4vmHwsSDjyRn4fedgXLnNCiFVdVO/iEGYBnZIv35Mar1e8Yv74gnlFnsY
T5pVvJ5rM4lS6xAadSFIxEq7dOu4h/VMKmsvZ0GTaWNNHVpSstFP7ouGZD4TgGx+zlfyEobvTGYP
bt4dUeCoGZIpbtlVVH7ZRnoknnfwJq13hmX0wwoNSby6rkCyPteN1CbS0LedrZFeLdsq8ZELW8Xp
yZshZxRSSGl25pU/h+MIFE+VAtOMAEqh6o14LEbEqm2/pnhk62UQoKtboqmrqQ0ygRGa70KwLc4H
Lpt+2N7brfJZiYFxggsEm3A/nvLjuP2T2s0JtFbUg2zEuuK6kUAxxrSvEU5WKYd0dPCdGHuGJglE
jxuDj4Y4PWVLtTcpI4SxDhdrEmhQT0wIoxIiqC0yicwlQD5rQFrx7hSZ7UhOTxNzgCuSlHjolF6I
yJIBgRHZ+4+tKKqyH7fcwUJWMU5vp5ZvxXKwQxc59VZKyjMDLNHUmoOW09ovoyPjeE9tOzECFPqp
v5FzrNQXNqL+cz5WhEK1jBfEufWWRbVsGwJrJA1mvrM2iBCy7U6PTH1L49kMn7cABE4KSuF9Lmqx
c8O4+NJY92eJFIF6G1trfi1vCfZv7onXG3+MFSP1XVX+nHHCRHKQnBmAqTSPmVgK3666iV/yGHHI
NLF5oBFaXolvFe0mSm1Q7wzTosnp2a6vhKKAVuOF/Zzx+QVqAF3jtp3seg5SG4DS2BVFtwQhllJ+
XzceZRhR9ijbxLwfS3l6KsTg33vj3n8cfgHswJ0gqgZrxfX0feBpbi2937eKealMJLO8Bg0waEsW
YE7NBF6aGAp0In3IVkYBzr6rWpye1j35vvNO/ie5hqiD4+ZUF5jtHGreev1AoMLe6R2DneXb7dFm
n841TRAsiptlcI+kSc4om+GF0hYtkP1B5dnAVUIYmTrFptuwXBSmg3YU/HieDTW0m6FPzrO5jqow
LgW+9low8q9vBH431fe0nGxZZgVOp+Sb+6RC3oPo4/xRR4NA5V/Qg/qDoFFOPLniOMjYgFJwgfsP
S/cwKuxhRCq0mXgmvh+qMroFcjpQhHhOhUEjatb5pyR8SzuARedA68zxB6ZJgKiCVgP14QszolLG
jdBL87gvV+UTRPOwfj8my4kx04ljSKgdvCEvDZoM7dsuN8jfnVDoGQJHqp7BabjL21JzIFvW2tOK
C5YJIc/eGrf/vP74Z/+BPF2R5aQPFzR/5AMJ5A/W2nzcBpz1Qwri0eNcpmziAgnZfsa1YNinhGH4
JzVcHqtoIh70z+E4au86XeDHZEYwGu/WgFpVTiy/rOkrvtD7mBVNrI62tMzxbsIh+zQo3PizclUE
c/bQmAWTonbzfWoEL7cjLHfWBT6GCzmiRO3JlOkiPNNjRVwteq3x3dNegaDCeo9Q8VKSn7rT7v1x
Zu69/QSlwW7Ppp6zn6zmvIyypCQGhKqdVOwx8tth9fdA0U9eN8fwHXqbu101dKOGG9BKSwmFeve6
7ES5B0ZMVBdr0QcdTKA0+6MDAr4lRxU5SVBfVUmphvb9b6HxapEJsoaINmlYtPrPZlB8R6A/sia+
OWP0FF4ZGgGYcahsKC1eh+K4aOH+UEGDy49cjjKnwkF8VWSEqn6imcbk10s9cHjLWcLUFJSKziER
FQ4l2loe20hjjyK2PD+UJedMEP0IH34KAUuLTo/awWs3GXddxNJB/IYvCqxsSuqW1S3Y/QS7MEdY
AmWsmnUJAe583Gx9EyyF6dZTYaR5c++dFwo8xCkU0PBMUCXVXUlWvWyp2fFWSocZoM1chLWVGqwM
kkm0degrN91M/HYV/qDls231dAeWKljCPNhs+f0ebnmOoJrj58Qb1x2Budh7n9qarpVsgUeljLvu
z6RstFtdxrKGNfXj23yvg1V5cQljLi117VvQIAzxvnlCryuVPLhNfKeO4/OTdISNpFppG1IGRqmO
RzHznUTPHOS7xeGrsuXHqMDu+2f4+IR+j17kxeZQTs6Yj8icNiyxn8At4KZu4IjD+un1SOkqpod1
5oprBEsbbi9ylde1fEun230Pxn9YsaZIhW3Jl5b3xLYQScLf+jJ1RIPLgzcfVSH5/rmm3Ai8boZW
rEAj8Rp9Y/ZAXCfhPAZkgHrygUDIlNsy9quVTncYu0zWuXhtLUUh0wYX7ffKkdGslH6zEoR/cd//
Ynut91dSXQTrMbsXA3XfGGDFb5mSivCoF7K++MdGmJbZBurmyC6fAMzPppCrxONl0TLrdvOXjGb+
6LxA0DC+3BycZY3aIvitLB4LfmdAlvaHWG7cGe0r4PIJk9BVBF7v5KAYto+BJGcB6GVKQTchJcwz
xnOiQ74fHYxJrT50UImuhqTXfdEwFEwJ1Or0HNRB2RcUchJ0CE8/r9YY0w7PcGPeSRvB98SYmWFH
NOcllva+RMVddcagkFn3nyj60L64j7cq/zBMEfQaWofYZLP6WeaEgigWa0w5tCKmGJkUeI8CVzSk
eSzOBWEfu8wIKiaUPN+/H9buAHlDbHNXQkY24i+s1oDJO9vK2a4KGJ37wvji/Osnx+y7yJ4U0rr2
BWTfnzLksDyxjGYrDwtjDdcL2pIFR6GSL1EKiee0Ia4pOJRb4js1n0pA9+kk5LEhC344il/4gSbA
9gG9GkSN9nJhtLgFChUDMCeufub/fR7fXBohTlnWjbO73Le4xO1pEFEzNGARUHcVwjkam3iradKh
AiUg5JShQUqEdZCJzgduwLmFW5r0s8mO9HxTw//GXdDhc9bjzuVnHHFhpKlgpCOxWVS6JQTkkI6L
scnYjt2T5bDLe+rY1yrcNqrIVOzKMRVyC7t+YX91z1KGQBatzl61zis2k4egSm7XAiJc6SDWX7PW
ORApbzHAS/VJE35im/G8InVGdVqyMtDKtx27+EkA/djoOSGo7JutvJuUIOtazDQmxCdfBOUby1r2
eEZFsb4j1KSj5azJgDT6VhayUB2nQ1ejBlpdOXtB3ou0fMktGgsK6Zyaq65wLDlUjCitbMPG5qCu
dJWDmvQ4sm0uKl82Yi+nAwnPxsLax8zxBKQ0nkZ9BpwegljalhnrkibK8rqWJLPyAPsXwNsZhJIB
z/TnWQw8OYkwNemXzF40KM/s/niFma/LVuwTW8OHj6vhbaJjzp6fRPAiNuAI1RWQOYGggaZrviNR
RoW4eO/kBjD5AxrxlpQwKXMmr+Db8zZnhr3QL2zu9Qav+/Dd5I0gCAk2GzYgc9nkpUVSzxVd1ebO
BSQpQSrPutEfoW9WvdSi66DPNpQ5ugyFW8XdBUyNnwcIPBWeWpah9653bOPle8HyhJEoFE3xnyED
v0PIMd1GkycTeTSoIyely8HFb1mV7T2MJY1i79l8s9i4lfjtKnCvRFOy0y93ffiHSLwHG45Foo4e
czE1EUbD5G8aV0gEUXhUb15D489TcuVXu8KhnqvNcU8SaKsrz5byfU7njVeA+qFheKDH1zxW7eID
GaTQHcFomPIBJNrh6oxZFdA66WkMW27g1sRU0c4Bs9tIehlfaiEdNRPAy3U4i2RX6X5IrNhxW7KI
4jhAuSHRSIsZOXAz44a0h4UfBdI86auTwhe0AmdPM95QSBrSoyelO9bZrxjIlgzN2rjqBOXhKtNc
naRlMEqdOIQjjF92yA/7X1BXGycXsrTK1Epi5wSjncTLtyvXJeXJFYsSf4vZsfIuwMsuPBWYQqBh
38ogPD+9vyRt2Pr3vxRdn6SdEu0OCB/5vpBAvQEENMUv3YUxX/6UE6hvheUnwuOA2Yvz5T0bQlYq
jhjBK5pD4ZkRqKAdVrtwKrJIzwyLz2xJ9/LsUsbKBLiXfCmz92hDmFhxbSpCI0C6o02/O6JaQoV1
l+4X3H8STy518llBAu4Kx5z1Rleka5zBBWBh2xFeZr0fLEAytmS/tXl/Sgxpn2Hdcf++CBn+RKRX
M40f/NgyQ0cTahYVjD6s8jczEvMTdNfNzOcCCQ0FigMBfzNPMmPA/N74vs/OK0/1EOwf12Zh1p3q
4ZhmMnHbpe1ytZ+/mbD87JJQ7LxSX10doYPaO9BpsNPDdDmndb+XeE9D+a6MpmqPsNfaPNhqxO2F
BqtYzxJ8eWhBT/cs07xO/radhDdfF+KGJzinTmGVN+w2kSLTvu1PLgvJNDQJmkGMaCCywynycjdU
dv+lHPDcUJMbdfyJsLZ3AmgWV109ReAwNQz0fUGxgE6cHleYGtAMIAhOWxmlYtYsb/67TFqtcCGM
Mi7qA/RvGlDXX0sukwRrCLbIHcyvfX6GMVVJBhl2LlD8BJqcx5idvjIW4ZEZ/qJyXw1ZuxgI4iNy
CX1ZZTDAyMnUAERtR5wfftUivuYwPfBo14MhffjBY2C4H25sSwiltR/q5SX9AiQI/IhfINuuKT8U
3TZmmhW1rtUbqgeGzF3KopH5WKXL0IDJEYDrMKK14CGHqjEQw5CH+8oMlDlY+zs1yqqk/gVLR5qY
ihGCaoIa+AGYPlaVtCLDxGeI1F4qxvCMv/gWDFJYA7ZcH/aGC65Tt0PtasxpkN4+Q9PyLK2/nNgC
t30eJgcUR1SE4KFr/mmeAoDS9DRNqwsw6AFd2tDiu5xODFw0ZsbWq5z8wA0tkZuMFDQzRv+p0wsf
d/9AvzOpKNMbnfujVMXAlgS0eN6LHmxH+Mi9sszjuyIu9amPUkFRsShxKUCQLiNN8zP9aV6F8Kxf
1cwWRGZVCJuFExEPv0RBACuxW+7PD5ZQODjyrLXE8xijkKnQ+OKfjuHEhIDDuvl7ONk3B7FeRa9F
q6fQKjWg1j0SZBZ+1uhuliiFBy1CYCE3XvoTJ41Y9l4st91f9xcsiuwcv4wzUHXKzU0Rxl7x6pud
lb2pNes1NSC7SLfTLH2B7OyGbRjbssO9w89/jBHZXOvuytqdpr32TM3IArwmHwLwGLuiuM8iR9ap
184cB62bais2rBpwYWGla9/jWPH3m5Pc3ebSxzXf1xvJFoq5iNkE3OvNdsYWT4AAN/ZpL3U9lhDt
pxXBQGyWppxoGs3pE7MfagSYOkOzD2pHHlb+i7fEjUM7TqjBejTvD5f9RAzhK1BIEkSx2X/4o0NW
wPUpERCOHCT1MZQXM2N5A5JNjiEPsEj8pUc44dKkcLJQJjE1V+TSlHVmzvTfbAq1PnKzUy9vCvUB
SzrXwV0CiUh51aQz6F7BSjyh4xtocOWJ9K8GKLu9XaXMcy1mvTfCMri0jQikeDvOAGkcpSOBZE9w
UAIS/uM66hv6XOVlJCjVkGihl5vj+HQSYXmA8ScfDehDDn0M790DvRwZTmXZgNTh7MwVcVF3ZYPO
JR2Tw3Bq+CHiZviD3ydwyYZhHVCYNWyxYRD3GUeO0X7eLF+BbxyLsSZXn7QgOEdtowOY5Vw8gnL4
gO4knkREivf2Jzs6Vy/rSUXy1KR6ObwkAnJ9w4Xnx1DQBMW3Wwuw2Qv0KUqsGJBq4inxeLtY/XkX
AM84HUA0RBw57nvaeSaNrb9115xK0p7OIpnnCVBtJKXEVSRqnW7Lg7dX2Qst783Bl1w/QFAKcDmx
gZ4wYPhikWgSrFufAZSalLlLk070wh3oBV8hh2GDZOudswcuXaDgdhJenHRIkfK0a1Hzn9x57Llc
Y7ob2wbjvCk2xE6cLVqCNugZVR4QmYDluVPftIajUiQq9eE0GMG/q9sVZUttLYWw16f/6meCA/i+
+TigmySbvgot15BX1R0v80t9N7LHfRHKFKGSboJjKvbP0aGahZvy6vniAzw7Od+cU+3mXmAFY7uj
uXG3N8+0SNZg8LM2Xc7rGUwO5USXf3MfwScs+mLJ2TQrGty+fWkyRq1UEDPi8OzoqoMz7sj9T3cg
l7cHdn+iEzYvTyG5Tt6LZ3vNHaS9X0SqCFOe4/EpHZIWc2e3OXj07laucLfQqaT1lMoHK7ozxZDY
Xm+WzXJKDHsoeRY2SRnHXqrXxuytgFwLylS2v2R7J4ZHWZcQBCBpd1wpUyxKtjkE+q5OAdQnItD7
zUHRAO/lLFcyrVODKMGvMOWBr3klYBjk1/jNGjq5YVngUxT1D0UoCHrMa+C3xMUM9hrDGnxpVAQy
zRN9eZLR7AHBQ6KYaf098TOoYaGzagVt3OC6fmeM+a5Y9YUNxl5N6HQBYL1iZgOxMC5Ge5GwxCmp
vhEdq6YV5lmKQ6648uGcsmctRJYSz8jqbg0IiRhz0pKqK1Jtw54wswEPMuogrzdhHKScTYVmWFds
DG1s1pwn02Fu46aXfVCRDelXUpPtnP+gMmyULiQYJ4QpArsrxRnikqbHjJH3YjQ8mT1csXZumUmH
Lq8JY+YJgvsrKpZDB3ejzbFI88KFzRPow/+pk5gLhYlzW4y33BUgxBmp55pqWxm9o/+cCGLD6oTO
7cnU++GJ8tUdlGKC3zTs1fhLOHfyvaw3pBuN+OViE7uXtHhd9SKp8XCIFn0tc9u1o4p98zJhNgDz
CwHFBuvAGRT+p5g3dtcwBMzHE/RzCvYNRjetELfAAi6zjWjPqOCXJ/ztQEfPAm3ConftDNv3h1pV
1DkvZzENK/9AnC7xUxpdRLtzlo46Va4KvSl4qvCikwuJSHsW111UXoZ+ZXem66ErUv/WeZj9e4jF
kEhdJgkDs2gHulHWv+bsCdkKjvkrJ3Yt1wUz+/i29clAn/QV9SK+jqO9QFHmunUdWVu1Egh4F8ju
A8nM6xoo+vjEFrnAItEVR+4xvpBCs+Vp1+7zvoGBuVZQKgyKJfwKr6DNWing+yWzwXHcQJ2JbAup
YRVgfyDukb2OnfI467iE29ELziTJSABH4Ghz02Z/lbDdoYQTVO5CEjzWKtmeyPBGCIv8GRCw3a/L
pSoB3Ugr3IQj17IZcqV5x9uKmelIfcpe65UcyLPo/cJpFaiOCh4q/wbRO6nxEsQBAHovvZqhrtsC
VoD5xketazABQf1KKq4o8FgdpHRW0Zw9f6frQE9d8DSv9NNRpH4dPx0nw0+vqjvP9OSjP3d17p8S
t/Q05rCQTictLk8Y/SljcH/n7JqARR9ueHkFfOL91n30xGm3gMyPxj6+uhHPYJAJs1UaEI9enILV
4rLhG4hZrd1P523C4ZgiuoexKaK6fHahxtFhCpTbk3VzfOxIC+eU50hH34DMo5asd6o22zCecHgJ
AVJD6ULo4GbH5KFI9FWE5snEXkzn30rf4dAVRtmPJL4neEFfmnqTuBhwLd8HmqtZ55dlVcGy1b2F
0Fv+SjizLE5a1E/Woncj8bRCebk8ugAXfHg3vxpUhmufTOLKmV/H2h7MuUrW4VBt6SkaL6rKAU0k
zcU6YyEAReB66F+muOMcmv99xUAS5GDJIN8+tF+PPZWM/5H6/SCoIlyJtIXE1cOmQMy7Iqkbnx7b
Z+nzQZFd4MSGgd3DEuDgeB5N37yheVaOJ74yzo71UqoAVdBNUM+sf+EY+ONhV0RtWf28JAHHqnO6
p4njJoSmxNM8VvTHygNXk813z55S3a6Dr6EEZFLnP63inkJM+TU8BG2I13AlXFLeSOJcYDxW9TTR
jlxU25mPAsDThd4JyxxKaIhf67IzD/LSKT6X51V3Eh5YGPldO5AsJeVSEOO6YR54SuqpIwd1TA6Z
noq6zunnqlyAVlauhlKhui98kh4AsU8u02rGDc8Qp7lXgE2ZXLEQbU3kUB+lrn8KINuScbTUcGXt
OgcfMphFu9l0CoJw+fABqVO8MdSVtGFpUQ/+VlTbWy68H69drz0StZnuMxXlLX/jTp0JSzC1Iv26
Hd32pYao6XsCfVrMDPTWbkU+VRgShz3OS4uI6p4oxvdloLOBAlv4X8CA3ZPxaAKViBwQIXs8FFvZ
9UvdRUETP0cfvZTCJCIS9wk+jbzQH3050Uz8hFs0J52oK1Co7/E9z981QvX9hyOhFsNdLGzqS09B
jcK0g7NGC5onMMxxfFvspuNdTAVX/d9K64XulkjJaIMEq3gdm1f4/Dw9XgrlyId1qxJE+dYpirPw
Wy+J5MYQxKmPz9BjQ1mLvllb9tBhLsYvMFZPq8S1JJTsVt6/iRw2dAXmLNTLv8VPLi8RA064e7SG
3yf5XpNFE6iOMSj4mdK0ipeYvdUTUc1diNrqP+SJN083hjyUp1XkSlHv7DLaT9sBy0o78SDtN/S6
PeVB7XN2Ds6QGwVOEybEpnHrrzbEwi4vYRleo9w0J4mk1beMhykEskkdU/HcId90VR6p1SSF1qNk
+IndQtbGD///iWTIxUgp5WsdFEdRVEvWGfmanZYkYI4iKw74AK3+fvngLc3dvW8xqT+0lEtPi+e8
fwXQ5XZ0tSKedxsQHHMDZfELZl4kHhSKW/EZnw/MvitxJ1e58b2QAEREe7zBj9fNlyuOKNgDUTtq
KKGYTVJinUKat6Mcs2AsecAeHdvzhILIcD+m6v+mcuDY6I1I3nuYb+zkzQ93n3vpE/YxqoOLDXhA
Vvvi8hnLbCbuy/BUMWoHZ48wIjKJXArYUbJPy7aKUeF6/oARHB15qfEGzzDaVi92IINVShOKHpvI
t1XUoNX5pAd8f9gctLpeIMYkxc1sMyWYtgg0RHZWL3Z6adCj72dGLbs0PkWMKVaNjdwCjTKhYdDk
n7gvZ2C8uW5k+3ClNCaSZ32sJkoeQuM4uByBsKeWnrtiayazLxLS/b1Og2dxFI1HKhBlsVlf9NAb
l/FM8WT3MaWkSxJGAXnZKENzIx9g2rJrflOMbAaL7fRtSl04y66CR7caTj5vg9J8S2UXnfnbzqwR
m0L9ZW2tdMPITH5EMAzug/MHk8NEV+0EZ9BLXmg8ghW87vHjorLUOENWw08VlPS+qeXua8sxm4P4
h0Xw9PSznPbEyIXlOGH6ojnACW7zBB11gfci2t03jCOZZ13wQjnpmxNO9mAvRqyrDMDvIcA+t4Wb
wtFuh+tHAHqsOX1R7NoiaagXg7qXqLgUVm/sKdoxF2zfwhIDs2J6r6dpO7oPKSR3YvgQefyusFjL
InWnlAxPgMmvKAM5jPSJgP5nhA4GLKvvF5nFNi3uik+vNFWBTMoz/4oP2qnlZBYEp8zgUlIqx7uT
srfmGHTWwaBLtpBtMgo5WX8EmzfW+S/V3dqL0HtyeIQhpNA4fVND/tc7j7BWyZw/uP618sO81HR5
7Wkj0F4RPsNYWvM1xkAPkLsS5sIzi+OQX67kFdp3z3DT3+n3b6v00pQ2oLOffx9N+ZEVwXTVqJHH
kujNy2BIW0m9PkP1g/GeT+aTLV5BBbe3+W1f0+AKmvmsJdCtZXQLmLRS/h9ZETWv3FLqnlFEpmoD
qaF8eJy6/vvuTiCzL0M/mcUqgD4vSHMNlNKjiOgBrJk/BaybR5STYiaiRNDLUEVZLu+TGM/hQJW9
s9IUB4O6J1ok1pzlHZT08m8lREnAx4rrUN8PJ5uJX6YgwZLW5L4w7nYOIMtf3OUNx3bWGXMoI+GW
mQAvmr84VtE1F6GUPC39AAR0nHumb3TKy5ArPFW4bHrdsalw6aew9Cv5wBr3ohv5pxqNIFFVBXQF
cHkCoi2L3ggWTv5kA9wLrB0N4J8SWmgDmCTgPhiHPZojgr5oq5vM0IuJpGDbcnrTCB29Fl1xqDGy
Re2CbWXA0/s5UJeM60Dp12TKDOFw6ERIUbwhK7dZzCpT1tiyNvcxYDAEzKe3s8eVow7tqZ/c5tjU
h5TCj4UER6KJtUoS6FONAywoOJr4qlPJTRCSOX6UpKRtjvUaIvkD970cPMoGf1z4ivFD/XLX0che
GkgkBsKnNV9Gi7o1Y/nUVq5HNuX9N7hQdvnqTAfYbcxJ2WcCsOurX9fGj02C9vVmWEbUS65gHqKB
c3XVX6iD3LYFNBGGWYrlyZYRzcxbCyWbg7113p/hzyK7Ri0qOXwMY2mM9x7CKP2BmJsN3Gn98/7S
gMfKU6lBvJl0CVN00fW8CvsMnvNlizEQLcsJH6Dv20oc6tGle+auk/2xPGJK0Z4OAbdbz7g2Kq7Y
fMTQ3tWIBrYxNwqdlUD6gKPMuO4tNxkRPLLCw9OOp40bUs4ZuHyD225yVkSEbugASR+CnhP/KMgs
X6t2m0kPEHSNLezqaeKwkX0MqSslRsZRQyeNsHadW+b8NpPLY/heYOb7ukhJIWAieYqiWSFGR7sl
qcD+Og6Ux8v7eI414Z1rHZWGWSVuZaJASPyL0jZ2HmQc0UbeM70cXkyJrZlSthRoeu0UlrbHsKTB
+/fq7SIUke3rKSYgL4t78Ns8PAf1C4rhYJTD2nMQmOCuyqPUhQJigRBfiLF46IyAACNX/adPAEJ8
EPPJibrgJFIokvHOLKwFU2m2LSj2ySNp1ZKeBaL2Uu2Kadxw4ykYLtFi0UuoCj+rzAmwJyVJdxgd
OSfNlaUeFCXvVd64NUteXEtzAwqSm9MQAfvuOr0Gs3p5vRHndCwy+Oo+mnVAXzHIqhrze8KeKkvs
+ycVtL8iItlMnpX4TVc9RtN78qubTh7mYKqh663/kkIpkPBUTxwB73p7GWCJUYbdJRus0ynaEEce
+OTK/oe7PR8gVz5O1W41qdMaGs2s/EU2wA1GYkt+MpS/bBAyiN2+5Ycn4Y3wiPAreqlQKHAYtYKp
XCpZqpviqbTCj1/4OUb5hPdm1FyDst2RlKE9FFPxN9XOnjHlGo2ElOQqAwbVdv+B969PX0k3d+IJ
DY/htaajWBTwLUxTFRCAu9WQmvtIjNP/ib0PiXoWXdOT5WZ/TDlm3gpT6PVR2WnQBDRgpz72ejyC
BcxBaYpIZCM/e1SX9dnQJxu+6sX2f0N3fOXUt+m0DxjpTBXIfga40yLC4p2gfKfR9aMsxu1Q0QzY
kSy+QdH91xMjLFHTC7GCFGoCq59mRNH97SyVPviQGyofMJKRgCS66HNV0Q44a+ZO++GeawSFgcYk
eCx3b2tlSjqRCXjDjKhNi9C73dg+VHCblX00HlOmg/1vgqzLD0rT7cQMLa2Cl85T44PSiWnyu41h
sXt0CLFO4EMwH3Gp0/ZKRsht9WuWEqFyg5GAOyyRLVTHC7etoaXBsNNCeqjkotk+URkJqbUw7WCl
4/EU2e5Mu6lMkSY49jCZQwp4LNEZPi/1yQYV8qqsLRacmtkVYQ23kJnejUnlx6XxSiGV7DxH7Pj8
RNjOLRNvIKFytegKaLfeuXCAucTIhVd+vjOwcURTovHrz96LMpz79Oe7SaYQNaaNThfRC2vc/nje
sEHV8iaZsQJGydew335IF7Sj4PbFDPQVYgiW0yox6XsQlOacSOowy2dYv5gHhLaBcEWB8pNNhN47
JJuJh8tMsG5+HCeGMmOCpUV4CYIf+v/51Wl6JMRjTmUIQdJBmO193xdzXvWsmMFBZFRyIQZViEd9
mdQkqV6S/01s3tKxDXjAChhoqN9Da2oRfEPeNi3wsiTAi9KZmiFGSuFpsyFIGYaqQEk9msCrwmeA
0qEQZ06J2Ew/LpKmdHzsWd7iX3CmwcggpUpQisdcoqY5ma4F/LbYaCh6d1a+F8mvgAlfzWEzDgH1
3POFHwoL4kKDF0bVwf8aAY/jYm82Vw7waFXT9b0rwZtzoombUaOElpDxJLpdQ+bWzRVvKSjC4wHf
djRemaxMZGzTJct4EAY/SSSYb8Oo2CnvWYVBCJTLRqzNpJnr8mJ4XGX4/o0F/C9okSMFjUtbqNkf
UIhwugBTRpuDpRWHlhRNwO71CbcWYoXC8G1K+s3Yfq+U2uRcYgyogI7hprElU+NjZ1GAg6yVWuiD
yOC+0CCw88ypD7cUQWCQNCT70C2lEnBJiZA2YwnxHI+p8hDehS8NHgkekSTL2O7HZHh8/lxRsNEt
EKWydH3vxzI+Ev7Pu7RG4UDqyL7X6OJ9CQo81J3BEimDvheM9p9lWCT+k1s/ndksShFN31OXYVGj
46Av4xX0n3KwCbIIZJk+wC8JWwyrUO4r1WBtw4wYUlaiopzMbyYoSEc7USuE+WD+26MqPr0EroPj
QPA+jS70AxfKDCD1O8zTwVWPVCvAoKK8jBY3LXlzRTBnVNpmPYVN7UBWCZNdVCW7izX304vRTQ81
mcGKQFPap68r31iEY+iJO9G9S41o6/cXwRPVnSVL2hmOYkiFLomvZ4JUdRLErD8q1n+BKyh9cqk1
OIa4KQudKmf++WtoIY/OAsSKbe6agT9W7deGj8Le333sMBw2xGAQgBMttpgL9zGiWO48lA60S1JK
8rEseAjYShA2J0viney5Q0srBQFjH5Pn1Z91YZqIDTdNifbkKq6d40fj1qc+1TxUlC3l1Ivcl0/I
SzG5YwWL2KWO8uCQj98BvpKjPcZ68UErs7N3p171+GyEtAQCSiglwoG6R4rvzPbBIVp7LQfbGemu
tG+Z7AOzbsde3qfNZljuN+5uTEP3zn2B4CYYRuYArx6uQZMInquPRhF+SfdOuW6136DFk4wSdIib
eeHgT8PmkcvzvVn6Petzw5zk1Lifen+45bn8feadZyEaoMLkcIG2W8+BXr+YjANUbJb6/FDm2jeA
nOdTlNmartlIqsS/I57P6PIG53VuRmR1GukvwvRwZiNjrlbPFippT3i1YZe1/Ce0sfyhvfT6TuSi
ezpDLfmrau92d2V8S+PaiLdtNFcxu5dlGirce2dKy9/Z4+Z0RFTXrneZr/8qjhvHzwMtmY399Cc+
+ue7zeq/TCTYvxeCJAo9S62ipx9pg9YT8JaLyadpMcbC5JZLLLcxsJ/E/Jo6FVf3KlZSJZoUy+Rr
rqoPyCJlrRWHX1nPKqxpDkIDpWTybwGVyD6bmefC4xCcP1xGAo6dDMcpJA486EKTyBXwaAZOHv+3
eYIJ25AtFP9Z1ESr2nRuM/gUrWQbO74TW7Aro4ACFSoiCvVTzxt78sHlHNyjlShjnEVxpp3Cqgtg
gRbwpKjARFDUHcCbgdt0O+8/kcg2uJNeI/H9jNotiE9Xw93r2YqQIOqEnAQXdoyJnZ/wUdsSbFfP
UxZ45SEacX+kEhwVrbjWi2xTImR2WN65D0hRg2FI4dYIu2vD6tuZ48cHFP5+DDObfzsGmUM7QUTV
UD+7lgp9yIXFBMdKj7FjctCoicZt8Ci1Lr1hvL63pu1+lRRBb6gwCyMx4kNBV6cY6KxVYLrR2KbC
4x/whxauOzxRqCS6DEnfz1dWimiHHu6cb5vdY7luyfkKm8FQTbYjPYgVyNWZX0dXxKEQd1yEAGel
ZAj/o6GwfNgRNzRcpoYwcKX9RwbWD5vNursOzdHoBsbs/Tng+chidVm7FVgv7xFgUMzUxocMWWQF
RY7AiJ4gM8cRUSfwHyejSB3AMyhe39f4jS6V/FYyDUgFZw4U/E2cIPRsJMXE6mqxhma1n0z/zn8K
EvlhAIxus55vtEf/OdF4/ax+8eiYq9BcLdGwPBIm7giHFiO1d/QTvSY1P2TTXX8IADsnT4r7CmQF
wdqyUwGeAK77ohK+2cpgjYppKhKZFTlEkepZn+7ddipVq7Pg7yCrZD4VA3UB/1lSKMYMrFhftuA0
V9b9M7GbLnAMru7xF/JXwep3ZTIaUuXzXOZEqyumdL8tW7BI4//3uQ9sH1XXXjzgdMafulijf2k4
oKsmqz/Q58DmlAobK2wHP2Sv8hFY8OIhRvLgght7hlHiDlkRUpoNpgtdLtMkSDOTP/a7KefKT2qb
Js59Ifdp68bno/1KTtc8uMojsrZKtVIHh05RU2opCK8q2BtzdEC/ZstpxyyN/dDl9qyB3aSIk3ec
t7ulLxITlQhZD0kpkWnWWlc1hBEg8utj4k1v+qdiKGNR/4J3JS3/4w8GYKd6AP2eGphIWzWD2tSB
LsJ5p09LnQaPXIARqs/KZBCmx0rHfLV2y1VGreYlVinOHSEXK5qOS8AyuVrsQbNZMPXOCFh59faw
GnxqmVWxnltCR3On75b+lCc7+97rYytznhM+SBzkuHKQ5SxsLw7hUUbdGMmthZZkjlq4ZMUua/Uo
MLP9U7tou8duLQNczBUJuyr3KLQ+r+7DJ2YX8nGZGneHdbu3XZ/1RNCUpcqx/a+b10MG0cH9zkih
As6ZYTny8iQq8IUvScHK3mXILL8mKOijZnYgCzsmUEeEfWTfGgGWTMjqXcxAcCVYXY5LKb6uEWD8
EK+o3ipTAC9h2MxEckvj5arBR4L6zS9CaLypHPh4zD+7QbEGAZ5EoDW1ABoMBTYZFvhJiyB6Gffq
yYC3qpRzdMz0BLtO6p8K/ByCJFlgvg+XHH5xwExFBq3aEsVMhMSlfLPRQJF8Vfzi20FtKsbtKzSp
NeX3k5AISAqcnt4E692ONlyfs44v1fTiPS5FpAK3ncnvvuiwlPbjLRwfELJbh1MClJ/Ce0LTVAzn
tXqUDElkx2IahdlGxmONG3bytX+Etm3lL7954eIcWY46AksC/PG9uByrDQPdGoUvQ3Sc3vBsu2s4
uM3/r/JTMo2/kASlg4HeE0jyAOmVWQ/CnsYWpHy+9GRmWGGVQaBodmyzxF+fhJ8fFTjIVxLT295n
9c1GwjFdT7/xi3E+MLX+u7XFTayJFMWfKZBp/Z/Wo0w2pr3GJThNipjH1gj8GVmb7DQHecDZ9eaJ
UQFBv06NLMvnZsYVfjDHMOq/Lioipe9bT/49+iK7ZternzKNDDUUF+phc+NZWyg0iP1ZLmFDwkAR
I688wxIaDJ3XV391MZS2JIUvVpG5H6KfZfVN2HpgvH5lFkGY9YlTeCYNdauA3mRgvojCLAZUPy2p
/aH9wtHB0AyXEyjA8PPEG/8tUBRLfTqbOEJC4F8V/5bim8++7L20RtpDpyxap36ZGwXVClMYB7ro
WUYyVi6N+RH6KJeTuu8pk+/gVR7dbU6sPI7RxVvuL5F0ehhwNp2mP9d/xtpv+gsHO6B6BMFcEnUn
7KiLFOgBo71d6w2kTtKTGK7Ek72UNupuIWjnpjljFUgo7WbRBmrhmewqfjByY6NQ1Emno6PDFJoR
aDqHZPn82UHsznzgl03JIKYaiS8dAl00kODVUMHZg1OAKbxQ+yvktel9YV3Ci3tXvqDSxGFqZ6np
23fRa/qT3YdSI6Tx1rvHA0Ri3uQM20aGrGBHtn5i1MTR6SDKJUFQCqJMxq20mm/+nynFm11tPpRZ
MDBKS0AdgE3wZ2ekpq5eT15cMePlqizHto9guMxQqOE9Dmo2HNJQEJvsDphr4WtXJSExUkBknCKE
ky+VB1AJAAZdf3e+RBIYMANJZkvabdh6V0wfJQzXi65ofRWC/xzclhE1JOpzr5A9hXGfAFE2pyQN
DNthRBPSghbRwfG8gPhcxyz+KSL7fMZxFxpUIpWjCQH0yUbUbMv7F5cfrYAicVnbh0CVlHYqk3n7
Ums7uEd6zERgwNtWfYapupXFoNQElB3dMB0dC1t4vZG3DglrKRKaD9rf77O3coV3wK2krOuJTUQV
TfgyjQatObcPZuesPYnwQg+xI/n4kuR4gTmfn2U9jBVuenaIGNOCdyQ8Yd8a/lGdNs83GZ5bsGGW
eWRd7iB/8MtGXHe/DY6iXN3bw+vw81PqNgm9hDFKtL0zwfECINYLfUfQ7kJ3hB6jxTUDGusCFdkL
MiuIc7h3cBa7jEw0V45+4KfU/wbF5YNneaC8yTBrWbWdsU99zZgDCNcfciBhgdjBBR3HNGsnAlhh
YisGHAZboRl0OfTTpA5+7sFdrXhUEvfiQIX5n4GNb40f8vszwrWCtNVu3J55rWQ3J4VNQqjVX6sj
f8B9uYifSxyQeeN2Z2sEHooOpAkBQeZDH07MHox1F5eiMtHhJ7tYOakcFeqnjT4qvyV+JGpalfo7
p67P7oBNgWl7wVpycaOqMCGl2eEiNZrgcbTQnst1diRzTdlaNSKZF7EfExtBvShx4oyye8xfC1mH
+Xzy9SWO6PYIz1YHHhZGPGBxnJvpXJggIG3Ir1xK+DUpX7kJmVRWGcUIBO1nM2WVW86PYhl6lKTH
zq1afN2GtKQ/0T02dDmv2rze2lG9jp6WGo2SbUosDeFPmLLOVZLcQT1MDzoEc5UOD3ajVhZrCM74
L11gCKy8TprHDF2d82J2nXvbZIlPkUqENg5itqFabAHAh4hzjB1do2vfvPrEtc3kxZAFPMi3sc+z
2KWQt8QoZRM2gLhR0LpfBIPxe5b0Q5hVK15qdzPWZtEjFSWn+g+XUnTktNiNWwqUzV4AcuWcoVf0
tZKvsgi24DlUanDLdOFWUOo2SD8L0l9bROs/a/p8n5KaXZRBHqy9sjcmV8zgpeM1v5BUzDpgyrz5
DxgG+y/QmUMa//Lb8hsHAoaDdB1goeBJ0xp8ngSsrj70IUZ9vL5tytp3xlaWsSmf7fiKTNvcxVhm
Jnmi3FgOkCwNAzKU4TS35Hdbya0GdjgOPA2Losaz6RzA1D8DAxLscTp2hvSlvqEDpLkG9s/lXUoe
1SHob54O66T7FtC9O11HSLY7QoZbqyjtbaHtIF8RZ3tYAATXYEurxZrxykE94uR2RyaSWIWP99SR
KplvhS7jxEFtC0OddH9Id1Ui+TouEBSocgeCVuZ+WHGySRsyf+Mxw6D6N+aYXF7kBAFBY/y1Qzyr
bjLbUxCzoQDFig4O1qXKTD/Tp7rr1QYSa9Dc+93ktzY6WhDz8gOMDtII+Br/47RKZjF7mH3TgIFF
OItZ8HbIh63jFx9SpRaxNDQeN17ffePRZuWUEZkTGXSfkfkOiZyJ45LCspgngU+zmLllVq0A2yoU
GAvkTwN82BN/ulgHpr/jSggc8UYMVTRNiNRjCLA51QrFbHGU51KmKFMAmjYLfo3avdBd2tpbFwFP
hq1ygDUPHDncdLCn8YwK3kqqhuPPwl9h+yLQKzBFTVSeJ16UuYeTWmIRMPbqV6Dc7N+hcxmHpxls
n2q5ki24REfbmgU4wK4ZVPh27vk+vGzbxH9WlQoQlAs4H+p85fqQ7sWHP62xUpXNGYQq49KLiIwi
FhjBzICmY8gKWYCu1qcSccbP0wAoyFI1H6vc1Jxa3m5oSOW5zPpAw3zvdbDUhddVyJeexxfcydh/
XTRI2maqMbo1PcfHbVKPGriXFtXFPRQeNzqKahuyhbrlxiGZ2DvkSUBbOzOJtiKXKe/A8BXSmFTM
K7S8H+9dejqhx6vzHwMSpFBdQLD8les7jWjTs05JTMhfKEHRxl/pR17KeEohFByDuKAMLYKJY019
BlA9KiXpf10s9B7itZ+3MyAKig7J2/+Y2lr5aKJXVgNWWpA64D5b5CpmeDhGXDRXGOaYr1hA1x49
NV4dreoVsFRHBkRaFr5wRsWkIDdvxyCI2JPJRlr8bKHNGKxp5EhPBH41fIoGfIWmYiTmFPapqlC+
T7C6wZXIGXZhNdgHCRewlRq76cEvwmbCl1hNAeyb5yjrkAJaMtjaWSa4cexfRR2yQl0h6a6vdIao
+t+h4QUQtippDrTEIiphCd/v30fkCflUMqDLvyBEgr87nXb8E5e+up8Xn50D28XERj81GAZ2hy/L
Qq4I0zseGhDjhmpFhZb3w2rp36aNabTnpdy0Dwv+j4Gm6SoijaGzfF4z81160Mbo1naYUnpfeQ4v
y1BwWGW9QhaaLwdcvwFq4UwqxZDsPWl6tmWxHCsvj488hRrIsEijx9xhbQ8qhmxuHBBqFX401HMs
NwcZh1H2Ues5jdLNzVIMljB2i/9DWBqVCJvEpsYePBtcNWcRq+Spc1VJGM9b5Enaan/piaHQ5UAN
mTJaJ4Ta/ft/zA5WV7U8VSVZWT1VDaEshYcf40c4YhmE5mYmZsmouHAN0hr/c2p6juHiQCSJn6VI
HCIjNrSnCDui1CKDFSPXZf0D0S/FmOtpAuB49KfNGQJutjZubwbvOiSCr3ehlTM1X9DYXuuHurh4
nYfU+TFXVagmuRL6DBAuqXlcfrj4NDvtDEqgxh/7sVDpteDLG3P66AJTsKansfc/ydzwJjRfmZ2m
d58JTHCvGagh7Upp52obaBJubAqwD2g1nNLGOw6msKPJa9bTQzrCJol8NL80fetUMUdh96T+lnVD
miPrJtprGu0cDB23MxTOtL+0vZ3Y1crhxjl1KAQMOZ4OXq9uJqIeIkHgvc+EZHhJIyVlFqEKgV4B
pbqXe4Q8C96IrwZn4kjH2xhufzaywHxS6stUHz8sgAZzXtRYIte3QKmrihzgZcamiIkQxqDeKC1z
R1B4KwRaaqsTDViN7rTL+euI9aASNXsnr/iXQgsfc/8NvBoogdQFlJKFhRqgd7jR0No+MbwsuNar
Zd6Io/Vr9Va+K+IRSEfArSZ8VfsFVJOYUYw9sb3r2s4YXfO5gJydCv+qxs72oHnnwuv6ETDZFvIa
YKz4355csU2/Z9tOPCP2rE0f3xNhbDmzilK0TdpehTAARWmiK3VG+Nn6I/AIUFN1NI5vIA7sDmu4
IfCoyqUdhcSZaPwgYG1c940ogsvrm16mUTXqpNrEuI0f8rwBJCLDDhtTKAIplHcFOcJq98S/j405
PvltgEa/1GW2MM/4IbyLDxRCu849abDNvlARNPkW1n8u3zTmUmsgKvVs/5KHQyr2ZxhaVl2JhrYm
s+OQrMdRnIGus0AsmvDDksuujuSZLz/mCpLdvfsf4TFSSLWyNS6pmIz7w5exoHuTkIgYObz6vXtl
4A/8C6cUXBHve2W5Z/1UveSfBIWjS+EZUz0Cmyn+tbN1WtSPNyVHBz1bCxRMw/658t+bCVOYFYUe
i0ONzNhKtrWObkEJ604rJ9DcZNZo4+QrjETIaj/7xSK+uFaqjUANgpJcAnurz0Aw4pEgT/jUiESx
1hlyq8l9XHEAJteEFIXIwA5QQaGTGx4+ivqu0ElLe3V4tMQqY27DLFQzIho1ga8Xo0DXJWiJovrh
mOttRD0DAEY1JY+EUzuAnp6vATCLk0+4C5nUdfZIZ/eQNn/yjtgr++1Qoo7sfYp+5yh0l/L3WHNP
Pyrykb4f2BO79lCrA8RQX/MYOkJNhGVJI3nfzBcBll9RSvPVU7A0GnyXfkA8qalIAZyTbujwCFxX
QwjdfOC8obQjW7Fsal8rzp9TcRQ10hWyKv5HwjSZkRAoq+77UAbrHZamONmPrGumsxcLIbIsIgkR
B7+I5ZK33nC6aOCY2GLs51pvmpi5N16glDpt3W16KkOOB1LFvYgWugGqN9/xiDXCC6Zmel24gueI
xZlhwzoSQpHMjQg7RvJbiQ51GArgYpmMwh5o6EGe+Bh8zHPaWdTLg0hiIQ1r476LRxHGqxu56QFw
/LQ8zzYngOUSbKTv7Oual+2CtyHuptXY7tBYvi+Y3pel/FcIbMcqCbKHEGTU1gQ4fa0kE52muwK/
EvespTDGtJd856Y3OGiiz5TWfdPIoo9ATyNCEIAM4a3qR3D+ZfQynurjdSVV2TYOZtKwWO1hT/GB
2+/MI0RWFTE0dae9ffS6cH1wRWpksrZumkU6dDfs6JdREuZT80xk9a7KS3WCVKwrJ/lgn+05w1bf
9sb+qWYnNPVqZUWN06dYUSysqP83SMrIKHcPRSAMco2bP+Ix9474Yia/8TxL/7sB2795HZD6Cn8Z
FqENW5apQop8iavafPDXSzuM1JzIb8jB8wCXEWfzfXPIfdd8XqieGrVRkW7kMAJaAbNAtkbUc9SZ
n9z5h9xHCqtlq340jPSp0mMOo9Sd+NjphXlWskbyHXA+L2Zq02XqUT1ZjNve0uemntsi36LY+rQt
Zg4tmnLYapzE2K+UFl2lZMEzCTdcW2Cs/OdnOEDxXCUckR1B3cLUScihRj4yTKOa0zm82IquiKfJ
BR4Xzzf6Mlz3surt+wYBDKG+yG7sT9nHSuXiUQ7obN4J/VfWcu0jfeKaulMb2UWhSiEl8OzzwctA
bo4EPrbCfackpus9t2DlRHgtwc2K5/PghMI2q/AV1TWQfQI6Yh38vFeRERysy9lz4N7kvtRiQGY0
ix0lfUCLUnKXsx7GpM4/SzhQTtmzWKka8IZ+EVBkT8eSqm2uPnoq9DXhLq28eo8YtfPSD9ADvCi4
CbAjSYm9cfC7wtB10o8VhwKeL+/3c/BYg1jOAlLwwb6mglhMliH0mGm7g0YgYhKnUibczYVf3Cc6
Gr0d9QrYTV1JnscQF67nPjyGF7uy+YCYnlaElRkaRNrMoBqkJk5EaGqr+fly9qKzgpQX/xbKtnQA
MS2VO7hYgsJe/0fQtj4l1iAy3uGo0JNTETWC7+qm6J+MnUKS4rbJ457/XziGuAaPy+PiyoExoqeG
YNyIoXjn926jyOp/7TxjncKLYh7bZsK6G3W855L5k4oKLn59atJZsFzpKlrW45aAmgkg6x8rQlPQ
w1IdoxQadJQ/OPSeHCKJvHScGNHSiKO2rjx3kZfAEoYBHAJi2OcYG+pqV3R+Oqrr7hA7zKL/n0RO
yjroFtkZSfaKkMVqIOmdWy7zZngnedy+F5eafpCmh7jkJdZkgEEX7mIFGQMjZOuOAkop+NYkj8MS
vBlUxT+2xEShjm5aMFJ+ZMVnq1B7uJbTDpxMvoZTmDhzBUQKPRwHEZ8BJhYTKiw9WHisQCUYPRYd
SXg53RNIJf6hvam/PpiPx0+v0rT0q52TPk6sez1e+fyqHthNfjwB6hlsPrVC4d03kDFyBdFUSqgb
2fV7a5CVmZOcbsw6y1euvwjGlRUPKoEvSPjzaQOpLSj6P23YkYMveZCrMrGAgXy5wnRqtYW1o+sb
1+PNx3dEEuluZPDz5+zTF6b2ddlTXt4toudLpn6jmrT6DmFwXrzJylRss9agtrxrzTpAO39EY8/Z
jTbhmxEPjM5BRiELpN7PoZxK+qk8IgNmuwy/i9kzlekJV2VQ24NOsrV0gxgN6JXFVM6wBrFL4Ubm
UIams6Ykwu8OctnZac1LFrcUuvOdApov870+ixch9metcv1zqs2YwRE55Jl1Is3OfO/zOUH1z8dc
omzeDF0GNyfvouWU2MSA1nf/218c4laQcKNiAPF7V257ZP1uarv9BqKzQVHUNIt+GbHqekv3ktxq
dyXR/km8cSRFqiLbNqbRvBEVJL3cOVJaObRTue4HjKnFTDoze1UWcWNatoa/iNa5v4nhmQVJmKRV
jsw5kVEY5B27VKln+1U/lfkMvLiEEUilQu+XHCXF+eeHaEI16scmxDKg6dFBjk/rqigajFMMe0Rw
knRXU/ieIxVvcO+p1xiMKaeJGFMUGh8BaqcLKSg9DtIFrBnjivEwgL3eBolAp3wN0N12Ww0wAfTM
Fw77YYtp20ikyI2nqe+B8t+EdDqO9ETo/zEg24bJqdO9TgRuQuIZB/PSVH8rWvPB2Pdss5lwKott
n37A3b+bCZn4Eto+2pfN9VKYLvT0m+R8RvzGnOR8Te69WZ47PfmvwLzArAPTIhXY3F7nJUUGOmFg
0oW1b75lVUUPyRRNMx+W7Na5Wx+reVDC6RpyJWKo63wkttCGU6RiFP6+HdmPScGJBAfThXZNG5oJ
Z20WO1OYtC8k9BW3zwfE6W3/71NJdKcIBF5i6wR0IietK1pPYdqqJ2g8hN3TJQeMBIirI+CiPUVC
xn3se5CQUiXPBjKNww0s7WVZSI2jp1wSkIkDFIDVNYRREUIjvsEaZhz5PZi4bAFDhTHZxo+hYKQ9
ZufYWV8hBcmE2KHgntRzKdEAs2dYyqqtN0BzsOxtI7lTTX4rPrLS1u55uvQm7WEBiLRC4qpfYFFZ
V+3idH2evSM4lMtI24i1SI9Kgb779l5VFmFwTBluvNi65e1QGevKkQI6JeHn1K4lnukWu9+H4OxV
rbi+XdmGN1gbKicxSHPSPbTrIVS+zOJ75jzhTLURWmYK6ocZmMmPC0lb1kEqySwn0faDQmKOgnho
RHH5qm0l333fn3WqM/cPwI8U1Frm/2Lrb2CWbCXdZGl7RAW3x/6wjTeP2PhSbXxVNm3lcw3XBOCG
u6AdhW0X5R+DKXMRfN7lGzf7jBSqIzcdTq7BtuZDPNpmsUF0IswjrQOILhKQM48O5jqizU0febYK
A7Ai57Bl34qWQ+QuxktpW9ddLZKkcXolb35cC8VShSKfeEKiTkN4f+ZF0IjRCkcHmes7KwMKG9Za
VF31LTLVuvEYvvJtHFJlo7/6xgTLnagAzGvnn3HsXzgByv8iNJ9Jf8Bg4AtypJLh7N6+o+OVriF6
fXzqULPZeZ+K6W6jf+2CxsBfJLGj23xE6pid6poUwYksb4+pvo/DtlNsw6WPvzHUdDZX2DJscpaW
xZz9S6WyOk19X6qCHKwOJhRHzZT28pPDHeef/j7Tknx9O0IDCiMImkAkDECNhRZ0ZeU40z3nUdp3
FY/C461gcrBY+20R6eQR0LkcOfN/0IBB5Tan/ix0EZtPbfPdDYB8pLkrM2hC2n8QVjGVg/BlwAFi
uY1WqNQzTf+zR7nzK4TICW09Vyjwgl8wp/tAHmMhNOkcmiokomCR0NDzNDeTkC5ifC0UEZUSkUCL
mW96nPyLCIPYcPpfRQG/gYE8TPRWTQYgbotB5FFN1zQwGxFduM8jSLhJTeZHATmcGQDFHgqgazJv
YS8GANwl9ht9ljsZj1m6w3LZP/EbqKdMMu7dxeEpN7Ks1Q19pwR97wtCyaCjs3/spkajElNWWoLD
fwTVGmaPzxHUdjoljKv9PvS7HgwXecJPcbRmuI4+NAec21WxLov1S7xV0vXNGI02tPWvXqp/sRg0
iNCnPplaDDKY/y7Qlo2S6Fq3XY1K5lR6FGvDlnUzBU+Oh3yRU/PS4yrgqdq8S9FpG8tFLgP11XM0
+NKzEbCZLZIFga3rRkz0uZ4CCyADX4Hd/I9aL1CY8Cz84cm4Z8ZYnaNeqgmMA9BImsZWLG4P25R6
ZFi/rTotOba5cGuoSPdVjO54TCsNNol/ADQ8h5EMZE3qN4oECMsekRcp/c5MY2VvNUts5hiDJt9a
zk7Re1TTSanTBr8y4kAGm2CcOtawaVbrv2wgPOY/4fAxFTajcCBS5fsXOKShrBSTBMvALN351VTx
DcOaLZZG7xdBkdXHiMnRm7urVHJFPlc3/Q0x6wqoztJOrxwuBxdRcOcOHWgk6VKlfLRnGlY+qRzN
I3gOCYFjaSTXbiUvy6DRgKroFynQy8aQLRshAtYVYfhmLa/Dudzv0S70ODzOrt7H1LmaW1elKqwh
XXlwYIspJkdj12JwxnEjpNAB0nVVX7OeXOZCEbFCXh5zBBE88WsQ4ZMCAKZ9oCSVTwdYHSHSFFEQ
BLWiOxFjzuXKMBnd6QYdUPAwDm5+NRfueah7VHd+VoqbQIz7VOpbs/zU78yvp2lReBDjX772bTp+
q+PDsvPBnKvbNhQ8QlPW3cj706G1oxgKifHSzx7dEuAplJTiLBEVpBKhOJOvnpIN0xJ16cxBCR+s
AVK0G03PoWYRC/s0jSw0pD0kbSIXN/9Rv0D/kzKkHDitsOX3EI7BbrWl+RP+wn3Fj1HEdpFyQCDN
VVDR04RyRBoZ00krJ8ttqjLMilQLQaDCKlQnQHMAFZmXaKpAYjBkFnvCZ1Ol/dh3m2C3gRsOxSDy
TDpOjePMQhAxVRDtv1nlK5WceYGn8VK3otg1qYZGcHaDKKxi1Bzbp9P5Fzm6pCIdmXY9btTXKrgz
Rt7UcPhMoz8EFuXnp3fxrppyo8S2co10A72E775/nqAssf8rrZ42IUxAUIJPVOCa2zr/6qnlKIo7
vvFTAG+LyGmUhA0s/+wo3DkTq2VD9ueES5gy+ZDy0dJcEfSW2KbOlVgkaD1hCe3zlvcEXvkXNDQn
KQy3MQAKcHx68EnYia0SJyWdMoJKQDz9dL7DCpsTMgEMiv+ihg3m1FYkSZdCQHV2hFiZRSegAXmZ
XBFTJTGuJv+NpsTlkJWHhc0SPOxTrhLZaQgcWDQ4ZycqcJ5tkqipdWazKQNgz4TE/FFh8MjEC9w3
CLmzbbmFaPtfmgyhZGfmqfexpWY0OpUGq7BGJ0CB2DpugcIeNElDY9imdrNomUQ/7B9F2QnRna4w
StK8+uVotP0U6qoLX9cRobuOp4mKweHfVJKqNoDXYkeFSYBZ5khLhMJF+JxoHZnSHbJ52GW6xhJV
2+ZWGutY3yDxc5ltbyYjDa70UJSTcMFtkoFbTUGh0X2yzYGDq/JfsQQRnLoHbgskPbRHZoWLoiQH
mvRt5Davy8St48GunvlhvKuRWlQspM4nkuh+y7I87b23jiylyIDdg0vf6w4adlmxHLm6echxvIsQ
S0uvFfhHR0CNDLwPMTzDAni1XkoCd9DIHk6mGxNxo3ShFeAQ2FziO8drvqtc3yToKqtDutfxFZ5b
LenJsOoMiO29rkM+HPzofw7kg2213+i4esUOY83t+5TojLVZ+UtUFl1uPwRgci7MkCtllrc4kysy
xVvPfP3G8PqvPvwPHEhpu0KHuEgE85nP77YNASin2ztccqQ2oUdcDfOf5M3vrIhqmEniVZd2JQOJ
FR2bVVxAJSlhRTxBCqQoQvVkvJEPCoiugKilAy69/FQaxsGogzI6P0LygJYm10FUBlssotdhzmeC
4d00ltcca8VgMF4uchx7NBci7UyHUvap1iWm144KrlfAwtyJEFq9Q5/Bgx2hbSyeXpnNKuZH0pd9
tOSpYHZgspD9Iq5HM9Iz68v+2eMmYDinAmjwxFLDw6FJiVuZZ41FMRl9mj0ABLoxwFITHH0WRSdH
vxn6Gaq9H3eFhzqJZhb5ZXcLs7ktfUU6edT2wQi+oZgVjXINHgTpcGXKXYlse6X03nXYtHuchbAe
iKXxd9xK7G1m7spX6Hma4C1H/SDb0y8ikQuhSN4fk0CFQxR7tz8XF1/7Jrp4hMNGybqcrhuPvjxh
GwxH+cOhYfkZPSIsPtbTjdpW9TnxZslGbcBOQFSewXUekLPV8K4bogqaIs04I5Kcq6wyk08om0jK
xt3NHcyf79v0SvpgNCbe/FXjjPMISNrXi1VyoE/IxAhYB+BUUuXxI55DlSp9khMfU7x3HauZyCTe
UUkeycRir4HlIPFFhM6EJtnpf5bpJSoYSpXkmsquf7+J0PjcmR6chxbs6WXNBrnpfxL2WHy0So3c
3zS7YLGmRGzWajdyilulard2pIS/sHBS4HJ+w30hueAq3q0hTFywPv3O9pQw86dPrKtOzCHA3Lf+
V+fXkxbkwcmqBUBEDsMuWa6expQCjZAbHgM0PFqCSnk4V5YwWpAZ9oF+Fn/A1cJZcJ/ML7fj1HMX
90lXpSqEgMQwGweYzAWWiZKCxKaYjZe3zT6bPfMMv9kT79qS0KSQQmOxhpaCGKxo8f0Xp9PTYiwo
der7reycQYkE26G8wB5OnooNU23pVaS9qtU+tT2y22S7i3E4oA28dhxsHOAxfB1Fk6lTUzRt6sgu
oeRdQ5USgG+73FpuQ+y9eXGzEMt1TI4oojaqHnWuFuvSV2hvLP3XI19Lf8UuW1G68fgWA4NnmqDU
q/0HjDxJSRw5ygG58n76BDqLyOtrM1edI9kQorf+gCh3Pbb0snAAG5m89gouMYeVQ83EoVgj/tX2
rXWL/fR4cS2K5xpa0cqDC2MRtnbe3yAzolFRuCgiK91TDlQonnuG/GmPzfW4ict/Lig6ut5QY+zt
phddJ3BHOujaNGDF5pLP2HGe+8k2qeC3BtQvTMH7TgXfE1pKRdfI2uVwHBBNSJLCw6OYGvr1xhXI
csbiC6nc5DDPtWEc5pbLvNHiEi84ixANPYrnC7KWn0h7nesuffFQJ8FFFFtJgATYul4tXtJPbcRQ
i+kEfjLKy7z5xmKVpEgJae0e999QWOtwkuxkyvEZw34Ks1xMW0DSSf3I0qYSn8zxM5jxqyymv8aA
I+S1PbUWbVBpxtsyPtdwlD0PkV0xjRA0B5bAQIzqV+eG0I3S5mXoYhVeTfsM2CLuQ6r1WnvYNZLL
UjLNpjcyhV3RbV9+S6cs88VYBXVpAQNK8BdWA8bpaAItzPWV/l0eZh0GP5+WP6hWBtqpFLzLafdb
rRfBOnbbyL7offt66G9I/K/DyTKTExSzN/PmsK+/bVO/L96CdPE+IG9zFkIUanm0Ci5yL5XSIeoT
vLVhtcuJqKGhfrmTLVR/ha6mHnKbJDSox7NCB6CI8qhC98m88oX0GXLOkCrvNB6oPow9HC0Mwitz
skzPKWqG9yz6W/uOprWzgHcCa5asbhJi27YuYjqgzF4bUAK5aeFn7/cuVUjrYpX5ia1OLSZFcWeA
k2n8ZtZdFMY73WJsASl+wnOGVjma7thyltKok7cfzGx3ELzgJnIoGNB0JliXJFQ1C5viR3Wdn/Pw
0MXZpHp/8rWeLT9pqFXA6HHUHP3hfrcufMV5KrbIa2+lAVdW13tqn3Zvop2qY/Uy+tYQDH6lQxpe
CvuwqnNuHq59LUs9uYjA3lit09SS1MT0C34NRlDjssDgTfuSBj4rzEoBy0IrNzFKVvD3VyiK6ZPm
EpNwfLv/nAEzRvYUSOsmXsXPaKSTfaoADeYhOGXU5ZTWRHLBWsR6PzJyA17EbAooE+Slujo/SlaP
wVAWNVri2GM5SJlQSB0jMIj/xPCRunP8WwTBnCrS2WW5HVZsqCZpA2rx351k0f4y6+mGyB0u/qcI
8amK0od12UChKuWBMaWNCT9GbYoeDzAEvW1U/1nVIkX6c4qI9TIn6DGg3nPG6vYmTt9MYsv4Cl0f
7j+2GNUBbz/24y5XgcgZgs895MNk0GvZ7Dj0kjD5F/ngjP3J4AXOxpkIxkQGMzauckUYliIdO9lj
JQoTPsiZLD4V/YYTXAgNHKNDwjMnA2pRtwi+lzGIhJ2Bgeuj30UNJ12maNIxPAhAdUSHrc8PVKIV
fR7/WbIWe9UdHqH+7bwys3ijsXdgICHNyAtd1XvXGUEm5/ctDMj+2xxBJSYJ9X/MWu9BLeh0Vi5o
mBBVKZxSVrUngwNxQDa/ueD48C2MmETA+5PoSVoRfd1OLDLz++vT+DtFxXoyeZave1nJUNutzgeV
YpEI3LNVucSSVUl43fRohRe8+hCtqJqXLrz8JFvznBy/uei9kZqiNxT0c9uEmtQjJzafkoEsvlG2
I2E5JjicwCawMloazXXrFKKawqMfR5edUe+k0oHP+1S9s24p2wXlGm3AlbNOV0pPkXiK3AeJGBJR
BAvVnn2PMYXmTITLnwQOX1NLmEtLn736VYYGiPx0hMKLShv9j1d4yeC0vdgyvx34kJJvlYYPKDe3
hNP4n6r5FdlQsYNWIL8Ab6vdEQT90rfUZEWk5UvZMtKsuo0lqlvkrlXGkZroKCZVBIuEicQj8jtJ
GkY0pOk0wWdcWtoUPhiugU7DG4n2S21n1asNfr/OC7mGn1rodco47GaLZzRgIUGTY+ui0h7GmrAr
TXl9QsjJDyiCrf0qe31p3Ksn/2Ir6huZwrWlC9FSz/jzX8uMcUmqIW1lvY4G0U8mZi6HzHNRvx1Q
2rtRThXhBZAla4f0coWT2aOyaA4fpBSoszKIbNRpff7g/OXSVLAKnJOQ+EcziML9QwUXpGzgZMT1
STOmVQ0ZUP0mZxabQz3d/tltDoPwJVtW3cJi2w49NJsY0QOw+d5yPEe1QT/bVWBeDFe/bLWZ0YUZ
UZKoha697Qn8s+3x+IMQxq2Oph9Sp4peicmhU5BUKd9kUliUyXHlY/8HkKMlzG5aoeDejuTQUbI/
0sN3/u+D4SIDsLcYyVgGx8AEUpB6IonMxoe01cDP63CUCz12lEkavjv8LsHEYEpx7G4qcb2DBqlE
cvcoV3s6MFHPTk621uIyM6IVg1ssJPhT0GpoQhCRigzw8nDgx3i7T25xO0dhyd+rJvuA7EnxZJae
oDEPVQtZfHkagxp7XgPKZoXuTYMdpc84XTD8Q1Q6hnDIzvDlk5wcI10i58WD6kyA5EHVwwCkXS/+
Nky6y6f5hoxtoQOsP1lGYhIw7jvedj94Ducl2AYTYtzOj6/lpYGYU+rcoFZysypyARAoBACBuvhj
wK7Qu1tIxOcKZdtvHO2ETBaCNgntm17/iLTQtsuLQoWeBStsILNaYYDElupCCQa05js8Uj9Yl8Hq
zvDa4T/RBYzganTL6lsS/3rPO/zMRAtmMIPU5S7+CKIbZcYMkvsS3NbvTfGeaWDXtjEBxa67xZ5P
4OJXjb4+5pQdTIEOW3K2K+u88dSIEN2Nab1aA+qq9iVoFyE/U5KNmcGAK9n8PqOgMWKdQVBnFlnk
iX5QLmDK7TiKb602DeCY6bVhOu8DXidFT8KmbScM5xa+X87v1kGrU2b3dudGYCpax5VrhSunn1oM
2Y6X/qfkHwbIZehfrtCc7hDJrxNqpNQczk+Z0BphuQkH/lWW1skAXJe1wrISU2GjbjjOs80rQbFN
d62ZwgCckQSep6h4laZpjXuKS9XZQTAZHAwQM8VIt2grX+qFJ0VDtireCkrFOR7YIUFbs5aJ6idA
YqM/KOHqQ5/xuMui+jU4st4bd8HTdveVq9JDeFhj4SVTvBxb13lpsidWdjaXFTSxwWn6Fj+2w9YB
yy+H14OoM+8t+y8uYZ7Dm6hkgWJU2zQfY/4J6SRd0ZUH8YyNwIYoQj+rRCRbtPivdBe3f/AaNSGe
kNypeTlnw/oVLwTcBrxl300WuevWpxxrzfHjk2oOJ48gDymiA7hgRxBVq/55/YNgL3no7aoyuYc8
/wk8+xCyGcqwOptZq1oJPndZBwkFDzBLAIDFo/X8PZYv2gPRQHs0LjIHdTzrwSwzTZ8LBbKCHXa3
EsW0VB01M+jm0UNj6wKTPYRHekWdNfFA0+NLWQIWqyGmdBpNggbT00qg+oT0fbYiEtgbiHzTF1yI
HhaZScVUMebeqBE6dO6wT7cKQwnLe3zj/Ezbf21rCbu+7lbP4S2Y8bmZYKdQBVPXp0ejnE6sZWtL
lPldYzlVhBFLyjEWhHZlYtEe3E/aUZBtLb3zLlquQ9X6O8DKbtY6cs3N0QFa6HKZQr7vWKxDnZbb
5OcZDOmoJpejzenCAGfHMdjJm33Cbg3sXW1P3TZP++iKiMMognuuyjKp59s0c1iG/aGaetxiPDva
uOWyrgO9RVNqhA5t6gFTOrK6Z/nHdF0sFdRi63nJjD83PRDmxtU7HwEL3kL4QZYpSdBc+xuE7NLD
gKGI80KszAe1fDbrDG0rh2gbYjaUq4fbGlU71vsYTXryOnrBPV+0WoRFGH2Nr7cCYd0fI2DAfP6t
gB5zCxfrv47RBL/0KVcYDubS5ZEdSs7Tj60v77dePj+VvLpU9es5uEl/xOhh5oSWoHUpsxEVYEHZ
hkA/+X3/mYUQynSUwxwM++lvlIS+Hh1/u//x/RGJWr7r4H8UlaP0KQtuvwIcoZeFYGpMoXjwUSAI
EY/Ns+8WoQfwSAn8bzpTQfV4KfwtfjtaBEJ3OhwSFuzvSepbrtSuSlJc8hybqH6t80jfQbzq9KQH
n5W0gfLYuhTIBXotBJMibae4EONUqRRgdBwD6Dp5kRc70JbPMEREMv5jwMtQZ0BF406lKFa9JgXV
PMM7CzrtP3J43h70TjajQOjxgbLsDyFLlFfrO2QyPF94qeBJs7toTMOuluWf8ZSJPQu5l55XehM2
7wCIaxVnQ2h2WOAVYO7eYSNhWXk9uzYRS87vvbg/pSIzvJOZXzPKhHQDqUG+0p+oq5Zyq33E5ujQ
a9SiuI58EkpHk+8vqvTk2SxK3/nw0vNzbC/miZgTYkewLIsJdt19ZiZqrFRuYsB3P2LN1jndyUEA
VWB9RdrRNR5gg3Q14uybOI9m+nsYaGgEbmp0VmOE+Mkn+cMzgT1liZth3b9LA/BByNLN5Dp1TM+G
VNHaJxAM34OqrMJxbZI4Q/cAuXVh27sUw4fNnwicGfC6Ad2n15a7xdu3aLM6hDIGFdSy82yfUfMg
8cfKgU5SYW13SXYZgEQZqpsYFMsjsh+30rn/S/m35aHqip6Ii//VBVMN9CENQU0xkQ+h+DLPJ4xl
KTn90FyxlWC0ckXEWE+dmcbs9aws5otMVJfb+zxk7gnr839H4ZOK0WsRxo2ha6z9yuJ1hFk7dzK+
JJvDY+PNrde+GvBtn5fstkAkPEf26U929ffqMxmjd/QGsBnGV/NtIUBacVq6FXCoiW00gKWbeBM5
wcRMYLmvUR0qI/avaYpB618NYX497VnWDyyDboz5R3V8epsfJaHzzMZv3h82OY0AvQ7zJZFLQ9bi
4J580wlagCGDkyhsbIvFN3OKWliEDoU/1eAUDPFOhKatUCLweHymzBmkRUsYbQaFiMpsQ+lAKMF8
nWVrep/HmiYFic39dbKfaxDphGvbm2mhzoI9st8KT3xbBa+KkxEo1T8XFtZM3nTchtt/AEgp5dRV
pzziG9XGNTZl2drzgl1Z0sHjts+JYW6ruXL5f01qNsEqAvzqV+lGLs6KGWkPuDtfrxtN/CMmotpu
pSZKm9amJ7y0hOAW3FS1nyLPnaMgaGlhgnB9UJ3LOrDP3LeTw7Q6M+TtGoZYV4J/rmFnT68VRCwZ
czInWSDpIEGLjLei6oQ3rQxu7SOjQYpO18bDybeYJp6FoTkb+VJpYi5fqtnXg5IqL6jpFcPSFz0u
GqFSoIaxirZRCHuCDCjdHAKBUvZgnUpbZpPdPiuqrbghrnWCtfd3hx8N/GUZmtlJi90eEuARF2QL
7X3ZL9PHBgPl6Kxl99d+RVnYzbtlK+dXxpVDbz9JBN1rEX4Bd59bCh06MrpZ0fjqmqIQ3j2JGuEo
9MOQDnpBubXv0R5sH28wJGBPPFXMq7+lZjcKCc+PL/GgWz4qlXvfIM0BVP+/iZ0eJ3LGyazDA7le
BrQMI5jUUjxGZorvd4yzh3EgRVDIUuuaKaaoET/iw8MW4ahzQdjQbLNSmcEV+weyTqo1QZbSEhyS
cl9XSLD/RtM4qnp6xkSomBsOsVGkc6G1fHQYoYh4Y87N1pK9tvz5WRY3SwP/U0Ywjzg6xQLnb87i
655dr7JVWNY8/OlhQlvBKSJwMu/dSkY8w7563GHdy3a4JJrrPJOw0t1sXc5dcJwwAYTTjD3V8ZoN
wzUqZ1F0m8wTwaFzxG1FJfOusulZRxNjTCxu8CcAExcJWGjSzzt68CiZNmcN7h7gBGyzxL7yOwZi
Lrb2EtCIs2ykAxGV5l2d2BJKUTRa8BJd7G5NYLEiwHuPJFFlPiN6HSwN+KBk4qDgu0mgP3ZoAvbE
NNYxV3B3FMWC7p9hdqrwaAfLf6XYheCUXA2RidsfyZZDcTEvwWWFRjW38HM4Uz0c5eCnZ6fBJuDC
h8e30HaOnym8m0//3mXTj+f0LtNm4WE7Kk3T4U0ZdyjhHWV2ZoLCE5prp2tahlZyOghMWb18z8I3
VqLqvOaUZg1vwuStnnzmyIO8HK+UKNgFEV+dyKLwD7A2ezm1VKgdVHOsqSP9L1FPMSX8wwTX+hSf
nZFqZ9LFVjxUyXIi9K1JiV7Ajk5ju0dTBBRrs3LVGFTo3KBkgMOreYYlvsIiwzetmFKSWKfkm6Jq
pJ1ZYa4opMGAB8HUb/VNPeHNA5NdNve0K97g92QhU7W4/3YAghEdQIG4eJ3/OXKETSf43utvq84Q
KztLCBKZJyB6Wqu9wljLRCfcWikSpgLnfqPxGB0F66m3dBdDXzKGx7UfDmi7h0Nqb7iOtpTLZJz3
TyCfJFKPXjh0DahnvYWLd8wuVu2jMc5Ulju3LxUXfNV6hGpuPTS6rP3M+5badDfBLVT2AFPPjsUa
fVWdXKZ2Rwk1cN6IEpTW5X1Gb6qcfrp6RiVZ34RCjIWitYFoD8HO2ZeA5ttTRQtKEK2LuznzKLiL
/ELmLzDs63n549tVHH9xWVt81be77ZYOE+obcFqNuYngFSW8IKe5kffAQWtCk3g/MAf8Z/GV/UNm
k+BPVv69ida1vUWP7HXVo/k6jWsxDYbW/D7siJP3zFqJYXePBOQ3djvWWzJkvZv9lT8l0wQ4nvk1
YbWhivXjXYHVxOWa5FaOaUWRjJqUMDGT0WgSJ/Y6Ovmn3SFXj79UjG5JxJ3UP4o3KDThBHouF4ue
16AryGoiKgsC7wTDcTtQSbmgll8f1XRe50UUYTgkjpBHL3jbbo79QuDVFFHpAU4L5psn2AR97xEq
vFKmb+LU7IuFcaZEcxsnYjCroNm7YUzPhh5G/QYDZBA2tgQkKphNQ/IpsaLveG3IrLkn2S7a7x/v
zwkcQoMA4xpPVE6RGif3NAaFnb5ruxg5aHybbIw9stePKnjWit91j66KDkqLJN9RHnPalr7+YA2I
TIZFMPyrAUdqhWKR4mCloxHOEYo4AT0fIAerGIgwZpjILmr/RG56AlkowQKQg3Ju3MS0i/AJqeyM
O3NgIXfHzylkJHFR8A5mTTaCWlnAQ9NkWbIuTo872Pum/cMpoo9zHQ/TzbJ4uWVabhmAbqLZ8Mj2
hnpzpKgSl0tv89xQIvSltfDHu14Jn1t1AKKxl5dNaKpdAGejeX/YXCWPH+I504yEcKnqwWr+wvfy
SE6MuOfVIgai2XSlzhh2O4zd20+8Wb8uwTM5p2QCrwKvCvIUbXKF0YzD5c7kDPSVr0tq3SZ648va
ah9ztIZnGB1155qi9wGglf/AqfM5CKvyZ58gZECWUoUSg9O03sBNt9xJzOpgxPxExB/B3aPZncyO
q84NAG5fzTPwSbCPkuAYqiMJCpxvqPYvav0thAi/orl44mUMl4Xhv2S/ylHnxMK5lY+TZzrp79GA
egu/MteiDW6UVsxPraIIl2+NaXs9y55LUrwPN3Du8w4aKAvjgTnbX7O0hD00h8D85Mzyc8/RJ3ic
EPaweUWiWlJjy4u2Jn+vX/SxGe0u4dYKCxuJRxgDaIYJphtSDaY17D2sZ/1l+Dxy4Ab0Q3xK54gQ
6Y3BCuDbdssIcuaX+aipSsKqjuiKabyD7IFFwJdJDdqtWI9Z0faggPJzod9o0eDVWQybxNCF0JTI
v7P4m48GrWRmWfz0rWq078X2JMNil4uh46iEq/Hm2UOLzfzF7fhXFiv2WQFDF5Qq4pJXX8wMgqOz
CuU0p3jGFCv+Y5C+nD3KswRQAi2jOg5xwcJkS5vRPVX56s8z0DEmcy4UsB6fTjlaxJOO9xlhJPHo
AHaYy6KTOJWp+oIHvw0BwrRaFe/U6meuFFa6xSBMFTaqpz9jrJ7jCfi0Ect33R7DbVSQXn1ReHG7
/siEqTq0wUlfx/ZMBwuHED6Erppro7+m/LtKYv4QgJMEAFhh0yg9idLmQriAt+XWv2ZqYW9COZOd
tsDNSipV0EYcpVEB3vrZweNV1arnaupO2OSZleWo/j2Weev6EaXK89CMjui+PwtNLBl4mN2fPh2k
3Yi+5GmL3L562YZKGru0xpDrMgECVq2atr7zqi82t8DSLh5ADdd9TYohnSBHiia+8ACcClsgq/x3
uY+4vb8ZA4RVe3sgooQEErR1oWC0svRWMu9/9DH0Y+1VwpQ5+Es9KaFrqWGjslVOFBrIygUZT4rJ
keJTnhhGGLPjJLh5/SLX+h/WPVjtm7ZZaSMCgeg9vQI2LdzbQjPz8bHdQy82NQwINMzd6W3rDQzA
VnRH1VTTlKVya8+46ouVq4tR0r6i9nBtoDEyAQHGkPQ8X17ZEsP6VRjw3Gh4b4gt01L6q3flZNIZ
nidcyIgLiUGfKfXreReyR8LGJBrligc9IbmKTQeqU8ADpuIZIA3+bA/kmEIBZTZdOS8Ta5Vijtl8
cJoetlpy67lDnVsJnrI5zgkx8/OjfHNemV93PxvJcg2Xo6TeOURX82KAiC8DrkilFHYysgVoHDtG
WL4Ne2OtJZIpvkzmzOwUi8Rwiiip0ezz694k7/HXcEpy6y47tRRnnI0y7PJobjmWTu17+6Rbthzl
W64G9Oz99E0QioEeDfJZMbtFIxzbQLJ0EbrD3hKHxSvrcqUMACRJZOWwLO7Qcn3W18ruRCmyRFVe
Bt2tyEobpm/tHNK5ZJfOatYVxLPf0ofAXVOxwRHw3Qdw8BSYOE/wgfYCXBrwPNpKrUw/SSO6b9p+
MaGCj0ofZQTug+w3YXuxSxZnPHtxazCBfWjXUe6BWa11TQRStI0cMntorA28kXqXQHs2mvjB1dPX
iHkfbpbQ9TUmTqRhqPFK9VKqCCCRVCk/4SQM/JyldnE1FlETyzLfSm6v7xN6cn6tNimQsUUQfG6i
dEqNemn4qatNXV4w17YEbjIdJAZkyBPpr0T+4gQNiHOXRPHQxDLixc/U+wwSRpC9fdKvynsTmxUf
FnLpCtXXQH7BCgAAN+u3g41DCEs7Odo9Sgh/SaMGn046HSaaA0cXVqe18+33iBfZtyRHz2gVHf0I
BoNC5QwzD1pLTC0a3WZEgeJB/G6TLz5vjSrX6Ku8WFwTW5i9AesI8rR0ezcQVJr3Ndjfwb/Axsen
mku3teL4f/C19LNaISK7SqZIMtgr38G7GTQSlAGlGB6VgkMtotEdyuLBReBRIS5wfBump/1F6bHT
Z6Z0BAubWwAF8k7Nlv26nL7PkwaahekI2IpAfU4gDCTMH6qHvM+q1Udu/jOh7OTlq9Uevzi1midq
1sG5LEgtXdrCgIRdmh2QSKDJ74eGdnhMleKil6n6HKC4tw8qSq1GiIM7yJracLaVzX/xlsyvtTcl
OXU8yJZG5K7xChTTGqBxBgZfxQBGUXNixsNo7MSKdyA3EkFO2OmxcRCIDW79NiTyQ8/XCSu79Xhl
BO3yMXH1aybeOGaG+N/RSSTNH5WSsEsOf0ViQhpZAPwfwYlUvtaErNSFqfagOlN66N+vZT4pYOeh
d12szTFfz3LmrhZoRr3BqrYmYYifYahMwGz69PsV0r8pnPhsdU8HY3MuHNQtHBqjsljH7zIqg4e2
m/uFJpinpaIdifxkOXwGDXWIOUovbpYnBbm4mufloLbpLdBK8zD/64w98/pNi8ivHfNNsT7iEtS6
noxfTIxTxUdz4CtKasDs+ghlWo6A601qprWD4OwPswsLP6idz22bHIOZs5oKbxDEROzHICKE4ubs
Oss0WLfd2Y5BW06xYxtcpharmy1v9G8S4fPk3KTzPfmzpTAkmxdxGPQOUW6AqOhzeqXscvM77jHH
2FAdzFOL6DDulFVQA6A41H8il/CjwgDOGHtovYFDllUUEqhESJNNUP9+flXmjiJS+iU7AiCT/PfX
PE3HGkKAGXXIBmwkWzE+Yk1ixmZMLOPvgf7iPtbkRikH7rhTs0FFbWK7xGpElyqMzg7YumZNddM6
iWHXUWq91HgzrqxePg+xdaAASuvpRpLcmmP3slVA83C+ELksa4TsT8MnapHk09g3k+GEYeGtWEwF
N6lCQlvU0dL+Tlk89pH13C8//9zm8jRRwD03EJ2C+MTbfkaTLBjjP7Hsbg9qWhksY8R5C4g5J4Z6
Y50Ltj/vaDHnVhJ+9ON+bR4OXb9/S3MPHOCKyq60V6rUU3vyq3ToRjtzZ6ZjzamZdIwLgquCUMvE
gFGJwgdEE5R/8MgN1vh7wQt6sCuNrGJ+RFhS3haK/OHWAU9sYDs/8qiICzNRoeB6Z7Iw5S+0Hxh8
p2b7DraNi+gebfVXTeoxW8gjSEXdPFX4wKB5OWNsFUHfBKP8kmezn9D3IN2VQrWQYQAUXC96xG3m
hMzGxFK+hD7K7PlZ0MUuhWtoJZUtlazLV+DhkFlxZEuxU2bg+yvOhNX6xbUx5QxcudbBIN76fDa0
1Yxh2Ks9jc6s/BBT6HQzpbEK0WbyWfGnlWAAXVGIfofaEdoc1e9c2bHrEUsZjp7YGFmzeBYwbCk2
Bx2y5rs8ofNerNx7XKXKopBiVlDFBPkKEoPq9Fm021YF/KyhTDnnuK4aF09K9rd9+6qAKRXeA8ut
g3+jX5oYsXdKVpNWYPr+xwvGgpu/93T4w6iulcSf20F08b52I5HvQTodzXGcjKfPq/73nmRRr87Y
0qYArAfglgLgn8mIb5e/6hlov2yAaVsU63J97dMPUFKPtPHCSjcsiNwIiURuFOyxtPgSVluDVL0F
aFOriwNzqh+7p/tzdAAGr0/ElKrSn4b8S+1XE4g52Ci1+2BRHs2SafUbDPca5dsFvGc2wVjctqVP
iqQvOjZPPLI9tqTnna83pdtGsjdUtN1DPd9nP4vdOLyySEFjo/Egitul69EgRnym0CvYWC8JLvhd
9nfMglstYKuaF4cXHvQrmQ6CzrzCt8Gki8SY/VYyxDW5SpkkD+zAmr7/ZxMTquaEmRQqUam6BcST
3mFnCQcnPetVeljhtnq2l3H82q20Q7cRFpcFkGoua20DFcJ/NA0DiJCNrhXOJtAtSnP7Ft6Mgieq
0PJHcCu6wAwMRqsB9h/If8y8hztzM8/f9jr+qcry//0sGm5VxvDMIoexaIOYABrDb679AnV83Zkt
9BseiSckwhqCVG1coQXUg4kSAr4fxl+k66uXlWelKw+4WvFdKOLGpiACRpY4S7Xi9nrxqsJjn2yF
c3qzxMkOPJJi5jDOVY36zPwvhB37E/UI1LuEF24kfL2U4H8xeMtAKCPt3X5/xX07nRNGXROQgMki
RMXpUOTt86cngfA0TZFtDNyiRJzq2QeY1v4ksaFrbhuboejXQY3A2A1ArGSeuIRFXA5ImrM8b4iS
uBCebdoVwtsGr/bwUy2pUinH4EIi+qzwg4wcAQT4mvYSPRCjNk2uSfeXo8UwRw5mpBdnvF0OBHyo
L49kEuGRqTfr9kCwxrAlgzPICBjQSWnGpSJZsduuRlFFTLcfrAE3c+jAOhvWl9vlHBdLe6Tq6XZa
jmztv0Zrcr5T0uv981dMPbBjoUqDapB1HL3fcLAJ0rinrIxaNESQ5f6rQTKadtH5PsYYeZq2Ppdy
s6A3g7+u8ZKJxqYLb+16WZis3ooVzYXrAq5kvDyBU8OelGlZUROtwaJXnBFhERov2JT3VrM0nl5x
LJouA+/eFX3NikTaYtMkF1lj0AeUMnbwvAZlEO7ZnyIThev3K14txtlIJ5ij7HRNjKC4QbRIjH6K
L9JxQX4xi/cqr3EVaiRoUsjMRu8QDtYZBcG6GPqX8U7GeIf80VC45HdgZTcY4SbL7HGKydwRw3mi
aSUZ/g8SAKlUpmz2Ivvs7z8D30vA7j1ThB0/ZxeAckn7hxzjxL/oQWfnxws/bR+wO1gUg2yqHl9G
3S5v0Cv0h0SNP7n4XIiJkEspxFBexdEw2rLVF+XAWZdx0Jdbcv/dK3vGNyyxJk6CUCHGZ3Kgzg8o
3ysq05jSr4EiNmIJOMpBHfCoclFTWPwaOQGqDIgkfVzR6gdX6O1WSUT16OYnXwHUf4BrodkktbvR
Y3UtVZPiNFAUt37liUlFGEi2TxaIr7hsBRRRU/g4B5Uv9+it2sLO58vsou6p6nzWzojQqOwHcu0d
B9C65Xv+7segF6P70FLS7VJWoGZCfdmZHOfZyc/cEIj/kXj2B5d6AsFnFEIz2+wAuBmrnKsToiuX
d07SiyLJX1SVluA3EdHBornJCIgLyztndjBOmcxM9rMJDUuvB2jTBdONFjWnrJrXKsZoV0mLBr2p
GXyynHj+2ACE+nvZZ6RSAgMcIr7Q7owRlE1aUNucRd7mawrzN8AiFMpRBf6mAjYNjKHfGvv99BWt
8oTbRc6PLQIK1VWPu8R6jH2rxR0lvxXDhtaiKb4/Zz2UikkiiiqsLsaHKhzgkbpm/W4mDoeGJsyn
0+40FY/5t5Yt8UuFPWYGvURr5YJShZX4y2Q5hxVSjpEv7WPm/x7AcZF5Y5vRUo0D5M7jrTZeNPGn
txFoZh7J93cgYLjFXpHGe9+dhb1dszT5nd6yWnhcO3p/05L+mgFSrL5dkcdkyU2OOVawog2KIhGl
TycV6M0+jEa3fwVoa4BaTx/ADkfuDuAs6Uz6kNCf7Grw1IM7UMxcFLbeJhJu++j0kpfhY5jnIu4z
VmegRYE+WFgP8b/eEtK+8xVTeRcHXIdQdPwzDW4VGhfg5njqfOcZepvrzBOk57BWgOZM5Y4F6qoV
rtu42pby3uQmWL1WIbrgsudK+0R+zB7BNb7YtSoHkLh6H6Rf/+8JIGtNOkii9rWmq4ELaVcWzpDC
EpTy8IkL3Gy+MJFePmeq1ypzCum+PN3gHgWxkMTVoIrT2tSJgCV8kAQU2TYlvDax8hiqRFplcs3l
rc9Z0Zs2FN8cqkVlpPxd9L7ECo0YtL8cxKdwXDiZLh03MD0qLL9/epKVuDH/R9jZO7WA3NXHsRbb
Z/Px+5Sa/fDdGxIxdc+jOdoN4KVVI3EP4huLxSoiNcWonQegjpDNISnN+FT/HPA7druDp/7KW9SX
PYpFreBFZjq2mp9sLc5IUyopHYHOTYc0yymv9Uso2pgvNI/khnpyxdRKx3V+HJ+DwxcIfxFqoDnb
OV9HS09rh7atE+gTfvEXfCdWwPMBstAPybkpJ+BERCaFt1YJbFKT/V5um0DAbBc7mBxM9kO1SrNX
HtOnfO12t42m+Ahrr/XzXj1+5Tgg9BqiMIS+fOMijdkQflBaUBVm1o0uf+F0F6nN0AjPR7Y8MDQ+
hydpv5yIC9Rr02fYdXAnV/AO7j5383WF0EeLrwq849dvRpBOZwZJPf5U4fW5wq2rI5I2aLrH4ghV
/POiFUsbnjkpeW025xQfVU9Djd3yDOXqSBLTxHTnW1ZgP9nJ4EdC4621C7CT/T0At7NokaR2yeKl
pQ1rP3oT4kqXxY+JJWoSjqtIe7XBQDCqJRzq5sHYd6C8cr2i6J9tOaUHIe8wQS2jK6mrF411ObLB
Yf1K1fpBA6QNRrYpV0xFH/mIoxQ4jLO1f9JE8g7Cn2GK3O9SWVBchZ9l1OaZhLMVXz4pGooKKrlK
j2cWfl8QSOfV3BzMhpI2jbPpVrByS4ZFzXDoBaxJTJ2vo6BSPjimTx0l8tYwRRcjF2GvRhkZjd3O
jqzMAVff2odYBw0/o6s3RtG9rm5VLZ6pZc99/KtmpWkLb7qcPF0Q++IwTLi/OTye9r7P6bOY7wVY
lt7n5tJEsP9JFI/9z8uKmZynpr8MQFhv1HBG/2WEUH3OTX4qNdV+ThNK+33ndCyJefwDsBB9W2dX
W150yLqwwIjUShmYGffzYCrhEIWqVaaLmr29brz/IS/b40sNFBza+ahQk1c9cWWAGW0cdM7eawmL
2ZLYNUtV/TzNM8BZLqUJjTLh0oycaU1IeQwYtkxFmL6Sc5MxIaqjOj01sV546j787DbIoFOdSjlT
tmFu/6Y/VFcUbUpJm8samF9dVCQINMQa2bearGZYWCb597vCc0sKk8oe1WLZI+jMfJPoJ2npSAOZ
BDvf15OlRxnqsYzOCQfWm3brqxQWvi0a179xqJ8mu0IrKkWZsd+x3yq074gB45o1YMqQkfBntZtl
hGetElg2I8G7GOCAsSvyyD42QnLp4QZZAguH/kTNGzqzr4HFztAroEpt1e6VRuiJmkjxUz93jR9N
oQs1KZ6JmDGcYs7aRRdEWzFyrI9lgYZu8h99vhAi9zb5W37PP7UBnPUF2V1pPQghCRLIuOu6Txqe
E4bLu2wbyEehGaWUQ3vYdmawaFBipjYzVVGC6VEMiadWQav6MIUaS/DuE5nxlmUyl0cFC9AHZ5OW
YFe/IW7VOToqhFFdSLHOTko3/yf+GS9XOutG5/4eApX+gAi80I4YQVspw+6Jz3+fkPKsy/TcibBn
x17C/dmVm5n0tfdhUqE7JqfU6DZ0QmLwsDYaK/iilifNpHtotRiDDaa6N5RSxakrPK5fwhpSgUzg
tgN6RINJGUVGnTVO2bECDEscBS7eg9MdqubdCVko7oP5Wu0cFyWDCyNI41OsLXSTzXEfXTrcPk/V
mI3JPk0w05vnaXSAaMjkU6ao+w7o5w3Qml91XuN6L6SqVdcJGODqSk5KxMUa5NMRGVJiCbZ+2gL6
y2EUlXYDy9dpZxp70z+2gQ1t5zQBAZY3k0bOOsM8bF0UaeD5wPvOo52uxhsToggayVT03Lud21Ns
QSASWg5aRIFNVzYzke1zy4++cRlXF4hLYnwIuq/tE2e/vRwBp+asnF2XTzQu22mAenQRa099LME4
XXWTqK8wn7cpfRaHo5vvHmNNdJNsOXM//c12o3dNqVDsXrNqLBnJ79pMiz4HX/b4LSCsVdJH0AJK
x8N9X0oqqbyVJ7oEgRvMK2SP+AHFfF3DnOE0I6iwnPC9gJnGt8CFkX/P8fBu+Ct0U1qpAm+TYBr1
BrZNltV9P0CyPzh4TXcoxtg3KRvP1UeEjhqFdOWks+tFV72edU3GXJIozya3c/ELb9ysHZcRw3kP
kkwJ+Zzl1UZSf0T6c1yA+xdT8SxvlP3Hqd6adV8TiUFAGzTk2D5CvhpF6OQLVyY6s22O4fXwOEBj
ohckJCt9eJODfuokE3E3g5WsJ8HQgxUn0goIuFg/NiGYNA15Q3MMAFKnv+pVsKbRRLmMjTnyCIN3
vR/3gxLy+ZDlJ/Zg2LLjcLj61GMJWUg/EZPWqLZYdrpkAg31yRN8f7UxwbOEbiOcSLStqV/MIOxZ
9H1mDF8B4CGGxM6ElTFeq023y5AV8w5S2V4v70XsRp+kb2gc2WrVcA4KsMYvj21gqsW8g9DLKLJP
nMH2AzFD+dYNfC8tnzfu6g7BsgYr9RVQtlg2QFAvWivO2CQWPp39QDezZ2At2VArlbZpq38rNoPb
u0z+AFqHxJU2W1vm8z8KngNcPTT9mWX693XxOgLfHLoHZvRTcQR4u8wnnkC910sYd6usqLekxa8T
8wjZIJvMyEWskDg4qxZHkRimgnr+ZSzWAFJ6+AThrTSUlFCCup8pqK0iYnT9x285INHu+mOJ9WPM
1FEpW8IGnk/hNYKkXlwlxEl4nIJYaW6j+/zleJC84XYB0B1b+oWevaWdaw88EX3/jPiDTQvaFlxn
aGPipa2iWGVf/hcg5ZXRad+jKX8i2g8dMWko893mY46oGDdIqMxOwt6dh1iRQmTEeoWhJ6j7La+D
QjfKS5chgjUTu79SoXiyqHS5LHLaaKgr3ecZJs65hf95BLigxLsMkeApyQ82zKW/XdirPL1FDjIj
/6n/ypER1mASqqCi6g1M01xG0OM4ab51dAFovCrAnL8kJgl5mZTBykP/4h80yrOr7d0GHJo4Ib1O
2gDJJus/46Vtfkon0h6ogC4tkFH0DYDZcP9YyUMJbkrizCRhycBTykdtWQuIWIHMTtLW7V0n/U6d
ynBZj5rzXbYt8Xnfca+JkpJKkGDbg8pyNbtfCxlfeMqh1r5IhpcEZ5M70k62rdIsG3SWUfYqaYnu
q7r+byTspdDhsUqFe/Q83XJ74NrK01ms6dv7m+MEnPip7P7WtirAnFXXEQzReqYbA2VOcSg8AxS7
hTvZpFDiEdAc/cvL21G7Nm0fvk5VIbM6I4CVHu22TT4KUXfGOmOaTfeN/L0Po7F2hUToaSx9H5Qv
2zLnPowxWWBpdPDJeDjhSHUByBkTkZjcr8w2ovLJyfPgngpYEQ3zIPXabc1NRjSFFJz/FD1LizxO
ZIUxAOnGPg5Op4jCr+K0A6h8TD+nC436LNvZIeonTjWHEb+8q5e+wUOCZ4E6sCrf/MvaxX3kWHvm
WzflTDXMP2F+x0tVzFh1nbFK7im56jgfi1TPa/E0JGnrlyq0WWe+LiIeSwGg9dqgezwlCcCnSq5l
xsi/2v7vfBpgktJz5lh27kVRx+8bc+70MkdvbjOS7g87unSl64NEnI4K+NAFzPTYhmazUMPi05Hw
S2I9+r9tLU7NBl5agOYRfC/XANRgJfEoEdrHvOCBREgqyFUlBxQMAq7cOuVi7rsEBFGL9dJP+QbA
+QnKWDewD1QcW0Bz4bxR6MgCzens+ezdfw6+SGwarEKrW0OgbOD9NbUg0wnMVK92FlXy0TtNrgZV
6Ii3j8w43gfzjSvgHtU7KUAtK/AXNhW1xVcS+meucPEZswenI8riZ1WJ8zFj22m0NU9lQaiT4o3t
REtZ7Z/BTh3JDuORmqCHcJBZQlFJDZSQuOw1NcI/v+LxLF53gcuFoFK03aeCVIFWROlkETzc/ssG
pKJso9VokFLlHsju6r2ZPNSAQH7u1hZ1vjt1s4KNIIzpqMGw91xIVGBaQIAO2nEZVxOgpBH2eKfp
dPSHDJZFFSKY/W3pByVrCSeBgQ3WpsKfgaIwN9H7MpThgErStEQFJWEGFAL15EPIWZ2t4eN3uhVR
KnGKc5KfTAgkOJBQz49o+a0tmweXk3/sJoh/+/MBGLPJLE4mEWa2xkiAxvOa5NAJQF2uHnARcy7q
4p2Xs543smNv9xyNwWRnmaMwE3iYSjOCqBAUEfbQ5xCe5dddeZQyej4d1ipfUSYIXYSzBgPNKEDS
8jkmWOmcINqmCJW7eS6VzdFmpgx7UX/TqpAWALt9Sj1+I0TpCcmtKSwLMoes//+klWfJB4SZko3t
UQRBQrhaG6pKMHdHuhs/ntPdt0RP7WVmbvwGQvfGKh/loXMwWiT4uYuxGVVjXb0BgF6AVFwF9AfX
eLax51/qU4UHVOPQLZu/Sl4N9XHg9D8Z8trjwZjW7vPFxDND7+aFfNmefVVkTmU09TzYvKvib4d/
FAN+etXJS2K93lZr6C7rJ2QFLv0w3d73lv+mU8cRp25I/efWlYaxSz2NpvO5bbnVq5zpxXZPpG2C
jmFxgyAXSzPYbqps1IsGuBT6SQi87D4+WSvxOmklRyqQzQLI8huqIQ6j00lViZds+rPTnUYkiXVm
3jhDmdLpY7yxEYkJh2mLD9e4Zh2RXtVCYjwrCsO997uk6B01a6s1gXAJs+FUMLj3PAVkbddNiys4
C2PrGgV5lHgthFC6mm5hsAhTN8ofH73NP2AlOzmCFGJYAXwGIpy4jtP9OtSJQl2tz2ZMHGsMCZeG
FAUDgoHjkMgUvGPwGtpOQsG4GlY/2aJXY7mJ5HiikuEHNtKjv2SaKwQSQcYXJfYtyW4DHol85b+0
E1QfDWTZw3DydLlpjaWI7JHwxFgSBcN2UrmjwF9kLObWZnLSJAWXmkG6PFWO6l9PURY9Yx37ih73
nRvdFseBlNf1eo8RPDANzBhH0Sa9QqrIlx2h1Q8+zCONCu1pZ3pSVHJEPrzOAM1L4r/KS57Mh+va
9bUt4EJYr2nL8B11ICTMavGuVPEnny1TCfX83PT8xlVYn/jXMgJiyQ0kg3S/CMVhUqkqvgdILrcy
F0CFYNO9N0FeQyLPhP++XK92fUwuIRZdA8ppeC9OfNzPsTg4y4LEliJteS2NL4I9wNxtve6oJiTs
dvODkjDBftfr1WQrBVjcFbDAo6aG6OtquOGkmz/vyIVCx1QTJKXXxHytSQ4xCmKyxL0CDDqFAYBO
RZQAYfbO/rBa4LCOiOzYXwZc5tp7u+SjzFio1BZ3kkWfZuegstnMQaJyv+jaMVV40cpfVyIQ62Zt
k1MkUP++krVh4VIrDjFjVJseoph5XVHg8sLW9GGlrChR68/vOwZL/iBY7zAUN23JadrWQE0A6Vud
S7tRo+HNcfwFFyptDFZi3p5AI3KJo1fwXUz7DK9QUkBvmjlpKl1sdj/K85aYOPxbFzezO/w9yCW6
KUVGEhpKpjouVYBBNnqviMYkw64uGaipnd5hM+szKMNhsP6+sGY2AQ9fmAPqfJowchiKJVIgI9t0
vZfcCvo4vPKstzu434xN6dv9HBhdjWYHwTIjLVtMmRUmiKA/gHNeXO8isY7Q+d/rL4+jnlLukjkv
+8Y+xwsmlB8fRMiFlVj9bnAT4CEibLf/I6PkZweYMwzvimPLlu60PI+s+8sis61ljJDx1AuzZ3ak
N2Oj97FWtrkw06S8nwo/e4yCssca6ZJHqZ5vbInypJkfYhqoaEWGQ+qHEm5KDh0K0+lvQNm3+rJ9
kUJwds4pM37y1/QJaO9ZWmHE9gT0sn7iU0TfTRtu67A8/bXgKMJP3MBOHs8A4PzRh7lSee2dI9zs
xjTkR5bhaJsR2No4p0RCigMERUO0LDbMCBGO7PgX1qhCHsdSkDFSscu28tBW17hDPhXbpyuIBkTs
RJyjpvYhfwkPwZYBcF7Zbp2V0JyOsZI74pGX+hzwzAfDtYqilYgzCWSjWgFWJxgGNwa8GEHtw+2M
SgANlZD+9brgrQcGAi8sakAXyW8M43Ak/TN9ChZXC2l4ylM+VexFtqdTTcABJpz58QmixEJs3Pt6
ajLTgoEiPsRsOr4UdjvpmSMYzipbtzJdhEJkqp816WkAxLS5JIPLKpIUSzxogQlarX8nqA4R9Wp/
p9nOESvPE1uokmNUAfNCjglgnouivpvpCvAREfHImprnAqqAYB15maqua+klbTUcNiinA1u7l63G
Qa2sOWnj+XPns8yZ/v5adq6Fx8y0ChjAJ5oJ6LwQjpWbieCGh7GAsQBye22t53bdbiAvw9uUxOL/
+CK8+kWOciz3nAa0BvIK51M5cSvELSjaeocL0qPq7gSDsX6SfypuSPQMkozpBqBGecB9aaH1pJ9m
E72iiOkVip6EeBp5d078fDEwhggjeDW6Eb9pfYgotygdmEyAtLPOdFQjsafzApsGg+O50FjRTJua
nexC+LTPWnWYgVYSHdwbP/ZRxQQY7xrWVaJNGlpE0Bdl/VPYydtpY/SacMpErUVBy2Rf2aNP/9lJ
gdWZac2ndZUitlSTlqY0YHTVxS10JD1H2wmJektMAfOpBPJkpDyz9crkzkPPkUcqInHM6Cqzq+gS
LMT59xXRY+JPlI96NMBdISjEGQ00wemKEe1N5GVsVWmW3j20oM816mpVVlx1cLbsoXPWxybPsEKe
T9p8DVkoknZIHMLlXcpkAtHcCTBzm9BAtv3vd7Hit7iGceWgjL4O9C+pnQrtzx7flh4/MfoMfbsK
G7jdbYTGZBrntcKDQ151NRNhgNuk2V4z+VWX232tVPn7KyIPVdRgj5Hm2gLLF68t7bR8DXlkRWgB
hK2C8Ccz1McaAo3Z61Idn4GxNVNyDxjsEwp0hvZRmVI4SkBCO9OyYGfn633dpLjanYdAKOp0dvV0
02PFAdf2pkt6EP1XJgQf+V+Qfhrs61YFuCxWbC+X3ow7alcRl+uKRPzpn1GkBQeJxTBCivAtoukw
0YwveHdDEKAIrcKNY+QUVlslQOfelJ+Y1o/YX7+DnWqxj/fV7jbhW23hvOvAaqnddZ5s6VXgTbHk
L0Nsq4LuT8dIEZ4x7jApgt2yIDcpCBBooVEy/h9yqGYhaJcXER9hugSQ0/8ydtwKcZQILHfPWjEC
+s9zOfE9M/5A/i+hLLy40OjpLgr7O+e7WVDdTmkahsdz2QTCIBUqgCwOJSThSWttDBPg1FVaWAx1
B8DsMv+ac0GKNJUbcyPYD3QDmWxbQGvvkrYSycvGT3++AS+KKDLfe/6dCwzUb4x/mZ3HlI/LKVlq
X35Oim0Ndfvj5IX9wFATVIEKARsQBe/qrIryZW/oT6KzRWNHpeeIixUEUSlUdX3B6rn8gu19uAN8
3VFkQdqnQrR0eg9g7qcyfWQ2NgomPKsZUoV961ndiT4ajy/u2A8XS6ovyw1feNAELoTEpoP6nx8E
QQwYmjBXx03kZyGIM4mr+LkPuC+E4/psrAFNS+Qysgv9/5XUkQS0zp1Ys16E2ry3SZ00YRKvkNOJ
iI9fNDRbM4p0KD0X/6PHIPHghRe4FXEZ7RwWMBjq79ipR3uNy4TZj0uWnyOPXxjd5diNFgC2EMWJ
IDozzPiA3XqzbnwqKjveJxx3mAHGI8sQJjIZ9UcxXWQJQAD1mmH5ArOesYMQwcgj1rwudhsdFYD4
rDBmfgpCCfL+Ygtko6u8YSbaZIWON7zT10KlUjciAPzb7rtUZNHDtZsE+NNHMuT6sChNwQ/cwlbu
bbxa7F5e07FVgUXjCX8kLmndgJtJzoUi6Anx7Yg18sAXxjN13kF6Hc/0b7KuS1kcj2wSEpwK5a29
cIWfhrA/Pqn4UeSrTq/DFVNJrt6u1VtGGOQDanT5Z2ucb2hQmAODfd63XQwE14magF4d7AlX/YDU
JdTh0RJ9JfqaWSdMQRynVX1g1hBe5vgRxbMRx7vdZyuxPG0bxrASmeTsO0avXaml/GB7sbsDNpjH
hE+N9Hu63ejVejhcMk//y0y3aTDhjfa4dF8r+bDlJkzd9OQFY022RXHJnpq0lBlCRAyuAIJ8Pgha
Y/kBKFlzbotj5LHf/Dt/ja67Frh6PWLhZvVyt5E3x1lrvP1AQ8r6fw25vFrgKDcGCSmB+/vllOiO
Ypg3Ou+jkw4nVabn4tcKo9rD/XlKw1rJx4y+7dizuEknS2DYClpis3S+yr4sh9tlz4M7RfkLDtkT
U+VXM4vlX8LISYgAMAPM8VTPzDXJdKPgnr60OKuLadTP/dQNi2Yg7fgO1x9Yd5EAwVMScuhwKZ+a
WJ9lNXGxCcjRcTgGdP6PakXAFh6gsLBIhedegeNF/xCLul2jnKE0cHw8ATpB5r8bl1+AkzMh0x0N
f64GRyODPJlJv28ykZ4TeVbga8tL1h/8IfErLQGwCWIxp3PJV4mUnytUR6tQLIVWffBs97ss6UAY
Koae5+7nib9erVyMHLnNS8LexF6boMLo7n4+XyQpMJs6MLXvGFU8qKTp6UQkFbqiKXX4jRMMFyDI
j9jzX/KpVaN8t6r4Wwfu/bYNeQU8KqMVSO6U6qMBsxe6NDiuCLFDA8fwzJgE9nE08AeYjxOEJjdj
HsG+5G7QY0a/uUCOXX/tPhGVAe/JjxI7jxShnToHOK4MULtyszXnt3wD3DzSDk6Bft/8Uz2DY60H
JAAKhK0eKEo9yD1cE8h77tWiMDHbWCULs5A5dsP4D6Yx2iCCh8YBqoPltLWb1iBaUq4GxKi1tfZJ
tyEzhlGoYQAV0aKyyxMacZSFyCKBZz+OvSZlrupv15CgTz792zstVDacoRrAcheaKqcxh74AxAga
GtgntmqA0kA7rk1b/jgM5uQIAFtaAoMomAM05Ai+GaTXSw0XReFqmvhgffcTzmWzYEd6wx4eWrtf
awSKf82Q5fXVDpDBh4na2quE0lMqxs1s6ln+hnNzDbqHP7R2WIfelDrMppYBlPFQDA30ehgp+l38
89g7aUlVxGhB/dHA6x+rcqOLienfBJ0FSXbbUjxwlSGILuq+L/t8FZWlfE97aSZbgmnKx3ibsC5S
WLMS/XD0cSpsTYI2aRR1tb2w6g+Nz2BmyEfnSojBIwIkcN/dt9yqeubCK41c8wMtfoK5P8GrlDRO
IsGUfz8EIIuRtbvIxc2A0JST67V5GO5LcT122WXifEXhbyPIgp1qj5zMhjs7TY5v7vuRUNu1ihqx
J5g4qBft5ONb+oFQleCdwvBIyq0zPJvp3ezNwipYi6t1HW03kcHVo/Vpp1wtd9EPdq9uhdtvtJa0
7sJrj6MOYbDRejPBlirJzDC7/f92+QDUfy6ConRJ+2BPcbr6I9wIa8vASvwPmsqzpHpNFtmyFtl+
SZoNf1wsAMJJLT7MIJOdBmw5r7UAQxfb+o2E0fm9jy3MwG0sT/zPhvq3pX765X8NT68olkHXuq3H
RGexY/dD8pQuBPRw9BFU2utBgSitR2eyN9Wtqse4t91zIX208WjdPZ3NPCie/VWsKLTFitG5bYDa
kLaCjFIkswWteCiGlj8qCn5EGvZFhdRe4YjsPO191LGwhRkKGOIzlKsvdhETPJK2PPe2uAun6sta
k4rq/1IctwnUW9CK19qkagjdddRUuV6FKwylIPyitVt0i5Ok337xrzXAnvOj516UL254rykLHpEG
E/o0WYuvBSne75e5A2yNWwIkNPhJKKCNgla9LhCZU1Ai3x8chYEk7q2yjuxXZA9t2Lj3QYtI/mH1
OG+7GtU8ApnpJiNlqUWemzxP6cyqWvoqF2YS4e38sXAOMKJKdMYpk1Nh7xw1DBRoG5joXtp2mPcL
H5lCVeAjuoRMhHNdUVt/Fta6xfs9ceJ6M3glVjqvIs4CZW1Op7LAHy802i6ap6rVc/fEyWwZ4anu
GSC7jpgG5DmWYl8gYCcCS1xNOH8xZYMp8ffgamRYeeupuY+ykVQNQa5R/rDv8LwckvuhLGuOSSMH
3k5Fk3LLcebW6x3ivdA3MUHaonwuQxtAkbCzgXqXgpkCPA88urU8ZzzC+OUhvPR6N1Ix0I56/vAY
bOUImdjRKk6bJqgTlJNskleoCjuDbDSLIyPp+s8bduOVi1QxDI+apo8/NYRCUm77x/K7pch0YRu4
QrEB3AWCM7lNBFpy+Tu8tBYjV3A6yLEi83vZmV+8PkuNoLfiNuIBexnRP47wovEZPrW4gdklypMS
HbNCbzOawjtKfk/Jo/kiAaDv6cc56fuYPoE/vArsSplAUgQq4S8TCyWDIIjAUlzLimyPS1MEy/gr
/kBH9OWyvO8D+b4ELrif3eZvsb7bVNZV0r+AMxS6rlqCsDepvG7YHgGBFk42j2XqOj1dRgMPAOre
g7/dmkDbQ6fSRqP6tdegSdP3NPhqupdOmiNEhe8dBJN6k8Rw+kl2ZazF6sqBsRnlwbQuCxxBsPXT
Md70lH9egzEK5AQcvAsiZjBV2GZ2t+dKg5LIKbYJpRnpaOB/bgPe5EbKeGEABW+/IN9/HOhGqovZ
StYSPD+wyW/MuOl7xK4xx69CcitufvQME1g7TQA1KBj91TUHJNoyqLicb96T2F4ly+6bkF1NGgwx
WsgTI/85RLN80HuegoDzpyGQZOMjpe2Bopj+KZ7WkGRcrmB5ixEtrnZXaW63yxh/M756h4tJ+esj
U2HzDAxZGchCrFNeG9j8DzEjgchKwVi+00dUEZDybWTTZGBrKCj+DJvqr5ahVH+I7d/SQKob3Aiz
wnqpgc6u+kbyOsCvIYbvAPu9IBWr7LFdQVhTxi2gFkPd3zM8uGD+3xlJC3Mw4T78DKPF0eW3qMDS
c3MqP/MykpWPB2C4EN829SmIhu5z0eHWOwA790r436GzL1Ml18f0hy2/ybg80uT+2xk4DXRsjdSO
b9p5CElG0Ib7LPcw2kIkFaczJSTimqfUeqXmPhXHG4QBaQhP6WsN51tadg084Eq1LzblwAaPg5fr
IllCz4RB0C0ooukzEvi5A5R9bb7aSt+pmGoFMvBDizeqFSpVrCGWmA7Y01L4mSIqzWNgHOHYDbBg
oYTHVgg5q4nAjB9V79YFaPKAfY+ZwuMGWjvPSCQMyQqxkoIDLG4KCS/FFPZxA7JEZxe5xNCKDJb/
PaMRaBo9yPn7Ee8mRVyf3gvY2tenxRbTKENQByGJ5KRf5ehibvYrqrmcGfq5V2XmEy+jenDxaNZ0
uk9ivyFU3PB6sgpG+UTDtQzhqpdMirQ9t0M2PHcRI2I8Dz/POeGcgZuV/OjDFECC/EowTlBlYzqD
1j1/nO1OxWSi4+W6YQB+O8dabVpjd7Aj+ZBpXgSg+x3d73gf+Tx13AFAswZrtcf+8mHqDl723CVU
HCcZHYY6KO25vPKTvDYZw2lCeDw6D/IIwsvA7lD5Fz6VLV4nIKhyIpoBuVDllKUK83sL0uyKEJq2
sD/PRC+Ug2W7JMoG8NiLfgL0LC0HKyv47loSAGaXSvO73wBMXIHqMX4NIQJ5OUibj4HKxthq9PTJ
+PIuZa/oFGKILHAUG8NPn5T5BGuwu4e6E4OQs7kG2t/jPCYjjx5O+3zPGHvM/VE77NtgeJifQfpO
3q4GFxh2LonnXuE3v2OGIL8w0NKmh+d4ulv4GWbwSlWaFqXtojEHro92YOuwy8zDzT2j135SNNu7
2wD1I5uunxsAdc/wnRrUnJ6bpjZTngtDPg3ak0ZM6lvweq5Q1/NXPmWZiNQ211O2p/LloCVfV24U
Fjw+V+8OvIUwFFANnqAOjhx2xk1dPf/yQZk5Gx1HVR1xDkrqujnCzriVsjjvJQOaPKfpwpxEj/2X
dRC7TKLlbzR+pKWF9I6uVrvTJsjJdaG2RtcimnYqtRNwemIiS4hW2XvPxAM5VyaAgnZF5JouConh
OtbFAd5FBY1MWaGFtd7OiBjeTcv7UFpt00OtBrZul3m/kKuEfyOIlcc62yB9wBDtz2FeDekG7men
b/bEvdv/gNM4pOnAZOOUPkqc4pEohbrqesAjvFxNE5Av6kJqPwHEHBH6Gw2qOINe0dkxhdb3HRVc
A9pXOibTUF+HPK4wdhg32dn4WjPD/gbGnfeJ+x0kiz0Q4fZDjrir/TF4zh5Q7SyL40EZZ+Zg9lI9
LWn8PxuttuEgge0dmuKlH4KY5XPH9Sgk3uF0Swo0RFQD1IG/IH7nLL9kxrjSR6vyVkK7qObFTgFv
SOVuheDJmewXsM78U96qCM/6FcuJKZ/YTzj1/meZmCZ7RErW0jCuYxQBtSQuF+D5pwTjNthOnuRr
MPuZ4qX59KuwPqwo1oE8FuBk9c99kDmCXFcqVPR/Ul0IFUSUCkpvq40mYff0wWOPpAYmy+6xgRZs
geQ553imNZ8yU86mq6Wr/45MBbxlLUpZfuGT8zUzRDEzj9tSulnLKetQ8aXtSMULtUia/nJpb20C
Izlk+YXzAAGXqQ7t1BobBfHr4lh9SER7VD9Ik22jeTie++2NGRLoKPdt+eZkGkkvG262Mv7kTDea
tK08ofuKrPe5XvcuVtU0e8O3/9l8VNK54kEElhpsipaxHqEuHuY37ybwUFAxCwhEiANRDgqm4Ki7
Nv8ILG+UvvSBZHKr8Vg2m3dCxHDS+26ohe+EyBbZXPtGMXpDn7ESgHQkhvH6nBAAZxg2xno5J4qF
3ZRn4kKibjKvqOrCr8vNOf4iYl6+c47hnLxjkUdARPjNG1/E4nTyWb88CWmo/ttgeiz5ryDZKWXt
QVu0uVjMd/Ec/ESru6OL+CrCQ0eikhVtHKb1yYQcLaaRq76ypuMnd6gAAYuRXxcsOaGxUQkqBNr8
AYF/I3NoCA4unEh7ECfN0piIXMqyH9C4dIhkMEsFIrlOJKTmzeGO4FwCdgW0uPqnMAjUDyz4Czaa
HL35z4TNBrtzoOrlgb6DqOPxQCEWHFTgoVWoyPva/KoJjtkjWIlOitaF3gdc1pqSTYiVlashoxLW
zyQjzVeBk6l4RNOAf6syaJGDYpOS/g9QIxcfeOp48Uo0sfsC55LcLx9pr6MWPKgwF9JmDl/LpVVv
gKsN1h7CEjhwvlPQz1LeC3pbRLDGKgvUSv6H/w/PpdrrodovHFWbvHQn35Ye39Ha5QYqinECtdA+
StZ/7h/pfv45Fa93kzrUc/2MrnBTubycJZ5InqhjZRpHtN/co+l9s0YtaRbL8h0OPnapaFpQAdfU
RcY2xr7aN/Rnykh1fw3Qjx3R9795V9Js0baLygNT4kB3beCnk7vrW8w/LE5nBagbcNldUVDIZu1O
G/DjC38SiU5z2maRU3bx5WZI/JAK7xaHGHTtBRmejzDi3mTRAX2xgwakk0LtDXWImSjuVLA4d5d+
OcV/91VADiq7vhkpIDFu6T6uSwM6mWcLmh/3/dTC2ZIPmG9TrtojXF/QaLIiidilzDTQN6pSxMgT
UyTZpyzrpmwkeZUpCKdB2O5oTF5ZznOFRdcmHz+N4Wy/oVQjhPCsNF0IzWlhsbkoVbklm/1BuDFZ
7WrhTon9YnqH3qM9Jor7wrRO+/Bv7TR0L2pMN3LZriFCkL9rkhW0nrjzDf7qDoZp19saaU3Xc1IT
+TYtcJjkFBfbIT4izbx0rohmNtMzSQza050vHs0VrQswQOAXodK2XKhxM4Uoaw1e94esB2vJCV03
NwSbgpJ8iGfAM1Tr+EaLAlRgs9DUtlLMSR78qOMVbbJaJmJmukT6GefC2naHFk1/grATmWRlRiBx
QfeyfbDo2ho4ZGXSUY9uOvmPON3CduO8JC2TTEVuf3C8vNsvmVRWeC8rFxlmhU3rWgqnb+pYDptA
sVtxkCnaJEQ/h6xUYwbshVRUtlnWGS3FEEoPb/VuzRVodCIXZkXklZVvH/qlwXLRDCVLnMSNGmKs
w+G7DHxSRIl5/IkB/dJ6DVdIlUzzeHuCO4PXsdlGhV4Pp+KSy2WbKx7dIYAGIQ7PGebqst+uCyg3
0Sh9OMkE7hlCarH6Tgqcy2ihG1ExABG6QniwW3zUFBpg/JFugdQpwnCB3qIQMPYZ5Spw0dD7t2xZ
gMetoyP+m+AjeRYpc4F7YwEHm677tLjhNdwDyYnxzxSC5z3qMdBCxErKeNpTvIwzhWZLL1Eyjx08
SMpCEPqVqz6REacqrhBUtbsTajsmUOvUzR/xTcK1E+11NjuhPsUnMi2ydVtir9ORQbA8HLuK3uyv
4X1YX+N3aPx4u7Sxp/W89Npf2QiIEKwRHGmygbSke+jg0gkJXCryvx1slQleTU8LfdvFaphUp3je
wzlDp9Bd2D1yXLeTY9yavcaurhe1FuP1dji7zy+87VoFAwKr6QN9IZ8klQ61qH+n0IDu5rUm223c
7LxJiFzfbfE+CtV3sAL8tJV05xoaVVvhqw0r/QCOalAzcNAWQzjAxVLZfqnm6qGEW7WeR/zpLAXP
uzF+a9sz8y1jsIz4ysrflDssE3O5P3QvZFGXCOSfO+ZEDl6+82DC5ypNEE8Uyvp+r7/u/WkkHOIq
EienqYFQEfun47XSAbmRjq4OzFlL14Sd2b4QgvyHMVDXcUSRjVhONXiOs8P/HkFDXm3P5Pmfa3Ey
jfp92bjKXJOnVMLpsMvKbwbrlS9IcYhmVlDr3qpgCNiC0LBNkuP5wg5QfgsAZBcCJJ535wQ1rks3
ePiv2mkG1KMF3Os4YeaJ4d5//zbyOTzq7QIhwpC235HGuY2gSaGNFodKNgf0iuGpxuFkAo4388lM
kbLMZjfjlQ8ma/A7RZTLmgKGyNoK24UGZQaZ7QHpOnHRttdtEL/v42UMPCaTkBzmGamFvdAh8lM6
uvkuZEraDjYnmJm1hB4LoACn3G5DCIXCq9miKNXyGKPTxOHbEJfg7834KxQCzc3OdFtkxEfKUOsR
3rNkuzVm7LzXDzzWB3Q3l+3sNkPUOrluFxxiwdZ9VteeLiKQj1x+QtTiMh3DiKoh6JgAHgcawU2T
PbnIirFUl+MugiLyNHkTBvrN8wrPQ0vgPPE1i8tCp6PdQE/gBwFu8Asuj42GynosMxyMBAkGNMLK
A7ovTpyZ5+7a8sGCuP7sXXz4lCCo/Y4VaRvUjx1Alh0rCk7e38zYYLzgy7Ga9/KZNFctvR9Wq5GM
EW3VHUFVrqJ6e+dnRrL/E7PmuMmZ8bFm43dk6pcESHeco/DvSy37r74leyl3aR+oiXjxQ8VY+S0w
Sgq4PeXxDuU98vA+c/WxzhD4jopDffnzKdbwchnVP/OttKgWTheBvYtWUmcXMEF4ECSRLH9177A+
OD2Z304qlzGo0X3kMWbi8FosfQ77e/XGQ13vKIWeeiW6aPghvhfCVWHwfV1wOLUG7WpkIiX3v5XX
P2adGtxM1GitfjcRHIrao2FUUFIa93HjNwGMSvRkQt6wZisO2TbqhLiUveop1FewCTulvHPODDfo
ecSNFanUvwlvZqhPGVMSOYbzswvi0EIPB383HOICfWI7jvs/bDahHNW/COwkRKWmXHZlGexIONjK
jOTeyKQyTnZk5+wLOR/R3SzoRuc5MjOG5hJb9wgVk8+kBBxW8sx6UqUra5+3dqgvTo3uP96jMlnc
yEUqyVAuuYRF4qACDvhvRchxesyTTF9wyMO1fDx09jmPitNgwBm0J1g6sHPWm/hIj+n3nqDb10bt
w7f6TizumeMQuutq6pY2SUIdlOyaZhjSzc56yJYXXEmkdzZTx68lHKaVyrSVwX4DtLVVDe1vNmRj
FDmSq4gGWnTP/4tYZwG1UQS+t4kxupdIPEoSUQNi0D8fYgVLL05NhMPWhPe6y9mWlQYg0eGfZN6z
UH06TgFw8BKGP4f1LS/VG+QilK4/1DMvLL9sDf/7s9Fy6BQsTvzlcbH+UkiEFbJkIsRV0IrLWWZs
qNZEn1ZKKneSfsLYCutR4rkmk1NOi1dOvpsua5d7mAZ8NmdUNwo5hGx/ZGYu/X67CIg77LbyaVsC
i7qtZzaT/ED0FglSRYq0OeACFw3ahqPRNioS4UAn0nKqGvfwEpXgQt0Nuj6RAI23jJspR2FEsPKp
qUNZk6z1oeQs7zo8IxBST4DVisEpx/lPy8d+2Q8vvb5WX9RmGpYa4SC48t9QaOX0xGCK0Nk1kqI2
jy6qZOVms6IylwzQ0STRK4ozCM6tJHc5eJwZ4aFZluJ4XeohNefNED+bAxG+qcQytUzSJv3gB77z
yuwktAB0oaQckWuQPpFmKu35XaZjoO91kxJtHdT7KZF3OcZApgQ4s04IyogMVSgwjP7q8M1fQUm/
A+s45ZLk9tAr/iH4a0JnBL2Yf2Wofmk2ZHcUoU6anT3tyeG+tLRpipkgc5U6UeoMna0oUXS0WABw
ial46j2OHHnLDieiqObwiI13NwmCnrIqeWXxpmj2eKbzrHnpuJvBEyyoiMI3rsP6bZSq5WL5DOMU
zY6OD9wklReE48LdjzalVr2axDog50YJoi1EQNR5NUorRB3xdRJMfo4aLrq7VpGsET9m39u6A+V4
cEEhLQCQH7FUCl7+gc+6s1ji3K12idz5z5LA/8xNMIN1ctwV74KN6zS8+kEobncbThW3qv4P7QI3
si0lcfXCbxqWi4pg9mwyuKrllJcuKl1rYKmj23T23vhduKGEFdfBc/DvnkbVVc87UlRdglTwriTx
DA39iTN0dMhRUvHL6JSDfwP92feLiLiEDG7wE9jLNzo7B9tFcYovetSZdz1yf+4PqX/fHp4dEwea
g+l8fsScJoYuWYzu0lOMz15wqVjJgc5V4cuxCiS2xTgLdy9RMPmaFFV1fv7dK2oJbfSDu9pieuT+
0K+aKWc06HdHXSe1AFfgof4mvGYHV8dxLIh8LRPFO/SGG3YxgnyFBHAnmh4P5kF7gLMEwi4glP1S
NvvAZhGbAoblq3AHmZ/tJHoAzJt/rliNXF+6PsxfNUIEghIsJoF7RyH2zTrI1Bb6Gk+OYrJQgfvJ
ct9DhWAx4yYbVtJzjDjLaebJ2V19kTdlzSwIW4ujD3lgA531kmC67kWjNHr192oZHmw/56w8U54W
+OnTkq5dVkaV5j+xx2lJGnlSJop7ymq3h0x+A9aWG0IBKQjrUrBhpS75LUAtKM3VLWaA4ITeaist
tRnlwmft44wjp8P16kM8g0HQqDWLQtgw834g6pBhgf+Eo64YZXy+JFj0gbIrlSefc5faTzmJlzrX
BmxW7f7GHi97IJmZmlVrv4pJr6F5sSmjMSVR8bVBFGFWjx4861uuJsHmYVvQdNRf8rWmx1UED77k
+Q2wL6TJHQNSNQrurHEss7ziMNm8QgJC7pPwL7+LUblEkl8LcHlkJu4Xu0xMsNLD228ByotJtxhG
Pd1sF5mEKmWep7wfFMZWk3Gatpo1MGQ7klLbhvWc7vRLqygyPpIGUHTDwduoWtQI1oJ30wms2wyD
9FfyvWs0W8zHuAFPrfPa0pZP6f9WpvMb0ppCB2BT3jHajS1xliXjmxMzG9SxzTSuKajRo87oe5vI
V98rz8u9t7TQKkJuOwjNC3h6L3a16gfwwhFKgA0vSMDAffpI3s9BJP3GNgui1dX19Vfoc5saeFHB
OEQLnb7dDoQyCAoCLw2DtcXYVpmgznt3udgLksv/dR/x8cY2LHXCL6AR7wfgD8r6oyfiEc0jjoxX
nujbnC6Gnf+XLDlU8GR5tYG0WKIJXNJ0Eo2BZKHIpZW3tGYTZgonJvMqFKPpnqvD91+n8WCAadAj
H2UUHkghuCy454Sac5z7cp8Qn82KG7VpOE7TgOsN0P2StzeHSkSa2ESOQkdOxOc6zIhLK3d7sbSx
R4dGVJhGy0ww8T8+rqV9GLa1vWXyliLs+jYr8Bjpw9wF8vH8wH8PYozVbX/cpjZgEGNt7fgY8QOS
7xVEoOgL3z3OufVqeXGQxzxlY6/8ux4zkdsn+PpKr630vTwJSuJWnVhWL3uJKFPH7b4SANiUfAA7
r2tm6H7DSODK54OAb8IAvopMxdVZphCAE1Vo1dodZHM5mWJUtqy1oGrxHuh/ZujDZvkhY7K4/95K
JrGUVrEo5+V5G+eVdCgZLuvvV0WDS7ZJT7I4175MQsJJeGKnbFjl9ErJlEEIF9DAgLeaSdTUZ50p
vzNHTXpBJCD6jlMpvzZMhGppdutXzskTZsUU33iDkfxw0VcJlH5DuTGjZQTTu1arnLrsgv5Gdv2p
54VB6925nC04+OhC1rRAGM8YyVSohmA2UPY6l48pytVT5ozRrpGwI+Y1bf+5hwmprFG28sIJxfIJ
vF84dpBd9j12K385iNSu/GKkmHlCxSN0AEZ1Ts+F5MjirfN36dbJEGCo19avXo9uqtHCwnK6W5zX
PxAq992AnfCSvNji8ITEjOgZKyZZKp7XKeiPtQ9Q/Myzp/d9pa609ojuM9C62NvLyA0z9K3gMsrF
TbJCqkr6y+kqaXTWENvtlYfYyzL/UbNhAnrqf0GU6Y4xD+jH5ry8lhWWm/O4mhvQrgfoeoh5SZC1
a7odmHYuQzu3VupoJDj9M34Tduu2vo0RuVahzS5fpAmTG9KLXbNNZhkmtjkje6Yu5AFAyivViPm5
1WZwqa/ouS7a4nT4tl6aBl9KR/0j/5h3oPfvji3i/p2Tl/efBCxnwJt/QrPF1YYuRsXEv8OSUfVz
X1VT9r9k/KzH3bpwFYJdF+PbtdYduNnrwVXjeyYB+/ULmSWK2P/HnU80l4iAvZoJDdgn49COFC7K
i0MhmoCDt+oAwqhF3pQx1Ofwl1puH6xesxFKPdan4IEUdJSwMGVIaZZGj0KeAv8mV6ilBUTABvLi
fRcNkUfY6SXjHYnPGkdxtkc2/VJkbiNyJ79x/1lVrP6FcspNSe6d6U5sAbBjZRUleQy9wwy1Vedz
2yXWtH9U+N+Aezs8zcJLJFbl92nyZ+MpXT55qvyFMpYq035hUrwPHgVE4n+nSfPMJl2S4s33oc9p
/YEixLgRDn8phv5y/vVro+VbXCQyiavh24580IBNSoh28UXydQKIs694Q5+Z8AkBwXOnyxTrTG5z
VGiipQqBS8P0wHPvV62/zAOsqG74EHd3ku7pZBngascWJz6BtFttaha16fYPHhwjdnPKHzu8xRQl
hQFm0D9wdpFRT7T4vlLUM90wyt5bGPU1/v2jT3DNLrGl9yZjAnbTN9sWKtVBCXN+ZBY+8cMaNYIZ
eD09nvTSoN46omNHEg7qiynNOx+QlC5Litw/UwrSfiuYPfnEXuZXeEJ4rx0w81pK6hU0ENq82Ksc
55xs2Mvvu47mfyfBTFjCLLeRTTdS2DHkdmKaetFrJ/ygpCwSBxJHt5mINVccQWe7U5GTmlXow6lZ
rqGVcV/R+hnTTkpAdZo9ubONjeE6/iratHh6HsiqA7Qmf8XWG9wbz8Oy/UUf4OQR5WopYMS1YEYE
qb1l50LaBdj+RQ/RqdOn+yBDudNWIMlKDrpwwfBZXSuqPMhC6JXpd3btGRJskKdz/QujSt4CNd0t
+MMc6eEqZTHmHEwvSwupVeF5h4ulmIBIc34WFUa6ooGz5rQLnsN0TSCQSTs+Hyqrxew53EP1EDoK
EFD2cV7I2OcNxdRSoObsFM2TZQHWZ9Jh/uqrUYS+9QAUcCIXHsuiwi/pxrb463xtccG+LeAlyoXo
zZVb8WwgVjRsV3kh+ZCYwu956Gxw+HSm0HP0re5GhW1FypaiCky5S2tf5CaTTNzWcrgFCJUCn5it
qo0KvMMFC3hYN4006NqOg0cV3Ko7i5pZXcjMmIjEsVayi2Y0VYqvOHfRPyRtZaUiF4jJYVDcxoxP
mAx7NrJzCQXP3xjZ//+YXHpMk46qmzUG3SxWe4soU+y299Hhq/Jd0GzeJMZXau5pJXc83XPrh7SX
moOGmoIc1PHzJgUsJmCQhny6s8Ua81toc0c8URA6zLlTfU7wEBGAnJBsEt/G7+NFX/eZcJJ0xlSp
ys8+rp9migta1gwLw71yBjRmTZClZZjcXN/U4JVBFzVzr14WW1UgMqcPw4E1KdFpqRNRWyRgjDch
EaXUbiRo1ATDYEFXEAAkenlnx2+WoGbg7omwhhcYtIoNQ8AZvl3H3ZzYpP/CA6r4+B2JrhRJdCQ2
pH6Kf+HsTfUFsOusVPtiOzDtPuWKM/9bZ77iybkMuNih5CRZHjDgeaG9g/UmQiDN0pn+Ly6mnl/O
dnIdEeOOchr2nxJO1RSGwoyClqcy+5WEUttQWhCqqKeeZtGf56sA/UII2Mj7n8OCIsY+cNmcN7u6
BwlOpArQyJVLehXV0clLKEpeli5X7k52+zzEGgPi2mbwTJfHZ1AidUacihL14y60cO5NvEo+e0te
kNRgtRUfDDxbCrYpeEmukb1JQ+lobPXbcyKo/0s9+msbJFVasj50fgUOxMlWyUIvXyxmHnmlr7rS
BzuFtK0nbYDtSkrUEgFhGRBP49H7H1gQOOI9WNb2P3A6D96+Yvou/OJeA+yewMe5icN4nKWkTYc/
TsEKHnlyIx07eE3Yb5z5+NFmLH6K/Oarq5kZjrTg2Cg57jllFZglveTRzUjPLn/L/L8EQkbiaatq
4pHV+D+iRTZFxL00I+5lbJCFGwQcUQNBPFowRMi91PyPOUnHyllREYhF4YrJf7cUcPWgU+KD0eWq
0injaipIePWecJTfJcskVQNN7DCk5ddVEl64siVwAppWCJ72WlCpq8GSy4AhyBYwkuk8dEANbyLV
JqCKT8fJIFKHmKBc7RihU/5+2JgXYfGQwUYv2YLqA99k2kQ/OFT2DCqOX0VIgZ0eIZhriEEpgeA5
xOmqr6PNC2eMJPHFePxVqewuxYdbthKFktd4y6rlq/V7O0z5CtZ/C5CauTDm5pn71UM+WVTJwdE9
LI2kCAUyr7eQxVEQk0/+TUhQU+SbSTzXoMoyKoveBOOJsTEgCWRVStYTIA6klB9bgB5jcu0G2p+h
gaEewSfpb5P4VWVLIs4A6AhMSsmVl0bxEQSbQPAmz5btNDoX47SGFMndsFMc2RR8JOlUG2Z7/gMG
IkxuzLy59rkXjy1FPVsISu4rDGesMZXyOrXhoZ2maFQMbpjwSD2yMlixN1eBC2MxJz+hpzLppKX6
thrUFvRnYfw614T9ryC/vACEYVjHUepjqCXJqcGPDqU27YgNoaaa0AIHnQ/QxgRX82Uv7YQqECyH
+VpYwqVLoVJnc6g9GoZT/viYhcaBpisnVdvV8t3ewvRIIHpLxkAXnzruRS3rZMBTTBPwatRwE+0a
GIr84C7JIJUsfuokV3j0lfKvMYJ1FV0wP2EhopZ8onGWSjDSKIdsmoiL8xpzoRyc1d1ZZq/ymBcD
PcFWIPFuWJ6UOY1ThbioYylfM66MvKRFVDkMhANPzMfZleKWELF7c47vxxIDhj6V97rm2tIvZj0F
I9033q7ez0g6wMtenWaXunPG8NRSgen7gK+GZKn2JNTiTTARsJn62xPbOeVJaT0CUWgQFY2j8JiU
kGL3uJtiOK+DCA2FZJS3+9aozsptPojOlxD5ZvR9VszNAx01TzAibawiyTVUA6P+gP04GoVEMTpE
CkOdy/34AjCzS3XnE/SWaKMEkjo1BqoMbMysNMHu9h1K7rbXyD3nxpHI6YPkc123vDnXbN/6ingR
PIK8uB0XFeuUYwcQiLfNju0k5YnthYglE+th3FrDWjmTtCN0zBVR/Gaj50kXqPlG2V5oGN8l6SJg
i4DmsKmV3EvaCU9TtuoOSwCwl8wjdTCUqnFQMpetGnBARe58zgxtsHHl8jwCQNaGRBlHbS52SrPT
/q1y50Hv21r7BxzI+gjqpLZrgMk+kEafRUzI+z/0Xh3HT+jBxLkQtQ8c6UBdQRBx0yGRqbtSvNT9
bZnN3d/1rgGEIbg489XepIMUQRpdloQrdZ7bGUyVVCzbnijfQ6WsNjH6nIIGigSEFYuSqXErkcEa
rycEmRr1Kw0krUJaS21KkTca2z1n/8pMMlrR+s6RoFh4ttgFGltf52o/aFqUDE8lEfiU6sFyTjn4
83hAHQ8QGSidKxVveGdtJ05FU/I0poxmrmMJkCg0TkbdwIblvxD3BdQgiliGeKO/p1iaTsup0TOY
p6J1yBCUOx6Xa3NR/TU2kTTC1fE67D4FJgggRq+FTZQb9tVYUI9Z9CH/NQIKtrGQTLp0LFOqVQAP
WUXU4ZNIL9I5L1dwkpFRJMAkvjKzy355BsLidvBFjB5QvQNctYlLRx4C6ce7AolNFj4fPVBMSeoN
NOkg448CKQQOHE7cIHaoJ9TqiBeY57f/whTYwMBvkwOHPnao+hPaySrlH/xbxU/7sBjlo1ED2kta
Bv2N2ZmO2cqBM5MSOaC/h18sF4VtacioYqa/l05AGHyEkT6ptKg1GZWpp2LsDKzPbO0DXkO5WQAG
A/4LS9QZ7osUKof7W386C8+61Ptb7IIqu2Rj5c6et+AuXuEWmMEL29Zzl8fPjVn7Xk+zSnOkgaHm
VSkaYx9JzpL96JKK3A1gSUL+lbrDDb7EBFv8zB/oD7HzAxDZCC/Zku22hva5ixovCiTK/0HV8Vy2
7oiWAv44ryUF3C5kdsxCyRb5sJPoRx/an+m4hlb5X63+9+/SiXoSQq2aeu/cEsgwx1b3KbWRVa2/
00MmMSYimkCCcwsjLABRQYa6UcUExPwBUt1gXUkEVxY8b8WMAFoH+/NTdTduLK3GOXPlEkKDwNdC
UY9pbh3mVwzpY2gsEUDSp8HZWfa6L47xWPbEyTc+UmOA1A+FlGJxeBFhsOXP6qH22D09HtUuzL6A
ZZ1oxOzMOnTgbzouWzzxhu5l0hsNTW2XMsnvTMua2oL2TqJ+BMwbR6AYHszcQTq1g/4bz4iecr1t
eQVco9OFyfj1I2Op5iw1fuMoOrQfTWvlHC9rpui5BeTTO3eeTTElXlpBuA4lHThYOsGdMn340o+0
rVVnnWgV88R5OBMg7BNSTTw16TT4nohtCGNCgd0FEdA/rXkJdnVMb7Nz+Qa8waIYIsXprUUKggP8
btv/iQjsXtrOGzC08nVdhreUpfRdacZSNnl4xYpfy6aAt1yCUnCAzeAUtxFSbJntoUiOvZp5kl8h
K5YRofWP2gsc4+3rZQhOWwrSg++JXPfgcAuelVcJYwkpHnyj/N0Y9KbC2xD1se9FTiysREb2b0cm
58vb52AdljaerD7mf4mJyrsmuoGbZ9rB9YOYW5rB7mN95FdpHBCYSS+6/UbFPYEgeCtn729X6JOb
MMiMFKHcQZnhRf14csf3lQvomSd8yYnSFQj7aWb9u+z22/wXHRqYnHRtK1r56634YLT5q4IaFDpo
hC3erhsmhIxo6jKzQmCrUu/NwQdrbaCsAxTTnQXWJAQwP5w63kxF5VDZnUVopJ3rS+IP+8U1sv+i
NlCR1U1ZqZQoA2G4qLJX3nPwUvp/msiQYj1PPT4Lhw7lHpoDK1QSOyPeJi6FjhibMRZeyiZJfK1w
Ij9AvSp2kbnK09k+FNjS7BQoXci5eqV1EM6SzPdRcZ0v4E/2pjx/Nq0i4FLLv6lMRpVjEf4j8yyG
+OLqksS2nu1cnZgj5FzWnWn6jxrwePDZvLWqfbbbmckDOp9Z4QfOubcI9aLSKJR/MOBGPA3grw07
XhpR5gDphfhzshiCJhRIZpNUljTNXg/kB++uUpjT3O+8CsxmYRSLBTwuwsd+ikMWcK7ljAFK2yQs
OaKQwX3hhqxjgqfPFRrzFAKi69Ad+Jz93Hq3VNaSIx4SWLLZrQB5PaosLFmkalPEZvs5yzo8p0fV
eXyDxrHR4xgB5A9l4kbVj646izTMXyFa17viPNm0s9tYZ97DlakRMpVSICYuCfbN++ACYbI6XgyS
8ESTAIsgWnsMLO8nY3UuqFfZUZevqnx5EXvkgQ852QxcFD8gyFOsC9/EvUMqW5QQB4Mkfe0cFto9
RZWoTNdJSbHLI8WplRLL+ymMJPMqIJBLEE/dNRDsCMdh5fLvhtyutNTa1Hici6uWRCHmCOUDxK4U
KG7H4K4c2uMZuTahH6XURd3asdC30OS2BPfRZfmXlLUAcy6PLXfiTQQsXXoGrqzPrTTbZrQGC+4A
cEKPJenvo/E/cSiXDBFHrACNSo8GOxdxdkyCAdJBEIYE0J8SPjnD/ANDN3tFAiv+wZ2lC97B7bLz
dhE0kPCIy5DryJb1B0cXbhVrdlXU4fobVUTQg8O5TKnZAkiErZCIZvSuP7EAyJm7KhXqP3jCBJ0a
MT9+yK/TzDAK3glFSZ6HFLNEMAB5fXaCUT2SPW27w7PKsKZhs7H6Xv/DUz9cisGFlEPLnwtvwGms
bqYn94mgXNPfX9ut6p4TQdOeW6+lM2kXBwKdXcdPvHuKN5/p0IwleyhSD4W2RnVx/HIwIf8Nqfrw
EPq3ELrNoKNFek2YFRZsDL3E9VkpNwoX2GHpTCITUtnFyABflXuQkxJcJtJDvhNu8ESQXeDGhrdF
ubKajM+FejrjjWj0GLzb4JIDccKccWYgMCXR0QPIQxtycyblPUm80DJ+KYD5e54AvCIHkDD6LNwz
kl3kxMuk9DP4nOjtrDeX2bzU2u7DFsAVrjw5A6sJ8AhHyjeQDMAuwOcsqtOQjL8EISd0bdga+QOs
v6pvWWose+SiNVwq3znfMBa876ZFAbGI4IeS+/GADkuRr+ZHkdFEJZu/YCYnmY/tIQWxBJzwzaKS
/ojW7IqYtqcbteiMNONAQ5VYYhjP2PciO7LX3c7tds0zNO9/gskpyWCFmMQBGd6oDDp0FvgEFalt
42cGLQ6/oomXwoja0PEHr8SRQajkoY21iK3tP+/TsMvIIXdGVnNa8dpFLqx4bk/340BYT3DOiNZf
aUDSOi30bkUppLX0gHqLCwnBQ0j0Yoq21D+6ZEUoNppEBAGBHaF2YZqTPGQkN5qaQUS3/wqWG+tA
mlmfoau7mxULLyEALB3pZU5t25s6aQyZzQT7S0Ee491K6Dh/RhTZGMbA1OhZkj5FcSWqWBl52/q6
bKv4jbi67D45nDUFdfwkeMHsV8EUPN9Bs120Xcu8np7N40kmw3pFH0imxEb+WNDE92kAAEqphJj+
LUt2CxmETWrtEMo1ugXT21bkpTHHD3rEGTvMoK9z3jhccAdEYbAV1mztZ5fJ9+/t1zIOFrLbgyDG
iDdecOd7/lok3uZKBXAcNjgQ4w+ukQyb6JB7hiWa6IkOaojuWHOtT18HeUnVUFASVXjUWOGnNs3t
eqKlHLPZxZYsFogMzIEqA6n98dAXiaPQd1ZsW41dReRnh1T3I9DZKYG6V5yIIHVnd80XptN+He0H
aslaQ4LG08G8REDUIBUbhz1e+4z4iUqE8haazxpEFP1xzKEUdGd6Wp9T5ib6oIsS04/mHb7IUBbp
wMn08yGFtWiH4h+in96hPeiyiJQoXivQ33DnNmD0J0bKatnVva943W4E3CP2PxA+nNbMXH/ivBOe
3MwrJ/f7tAOJ1k790q7jSAnhzHM3GbkSaZghJfcwiT+Lmm6++qIEVYKHh2GXsHAXc9wrRIEPz8tD
RPOgx0+cuVaAu8UGSNYSPCzvrBYnWsFsMpz4XuP9oASwNmp4TxR5om17dRV3Wm0daghUVzDjv+FW
h9Dszor07JzlABHPuBDpQrFDGEuJ3q4Q2ZaMFFc6LaIQNdoGMtG1VOpJtp8rQP9eYV8wEQkBQNXd
nUJi9th8N2fbwE9PtmewhKX2QkMQR+Qwj/c1ehgbuQv0tJhwyl7hieuNqcU0R+Qd0vQ2IYuoamo/
C86AeCr6qrdFonMXCu0XeOMZLGlcD5B+vh4QP9PBeoHqn10Ho+D4ENBGBjeCaAo1h8w6D5PCqwAd
liuV3oVeTw0IHS/dlAs65w5DHH2jaAxfJhKae7nQQAGio3tuzYd2QbXlWbVGOpl8VecQp2hOf7EO
6bVuFS25wjda5ToQfKRYr6FLVDy76hxyFmibDtvqEhj4H2wjzN6vAx81F5q6SV9R4b6CLz+Yd9Ir
Q5Cdgt1znz8xI4wi3T0dSCEEVeoYH32FltK4kpvkuDx+ji5G6+W8hx74CIzmuPuBJzZ2UsTv9hLV
mX8p6XwmNQ4Cfi1AAEyHkQJcalAr1fC1xdNxOvBKjsfCmxB4AHhPBdWM6Y9JSJBy96xCrwSI9KTe
QC04+d69Qz/UDbzLmBWF19IqZcRPE96ahHuMc8SWe6j2HNJV6IunFLickhYYNqkeF5maV8vlVRTv
3SSoxA8mWqcbjnIDwXms5wk9Thn4sLDXBDmmDjBskbFhOkj9sdJ0hAYv0syGl96GXYjs+YLzgWBk
gmF+MIe+zZutt4vigNfHCkSfkwELhcDrz3S795mPzwmd1PaFRCnqDC2P82ZW1jVtm4pXxeUB/NFf
1NVh7o3JhKGkG4yZcT3xz7s81/Q7Cn8CK4WCGeyeqBXSQP299RTPsv19/0hWRWPp/LSyLEqd7ND2
ndMz//Pj8OCsd5E62ep+AQcoTfDHGIq3gntAIpM1d5VqdrHPQdVhvGcH3q1HMUF1U6Owk8/raZr+
P9r1CY4MTbtYFdefRhT4MgI5Ga1U0IF/7rn7wEfGghDHymcJIjDVUz9+3AM+OnHoErYYUX3unSaa
4bzjhnmC53+bn5ywKUCEbDDt1R1YZl91DsjxJQkLTG9i1IRoqyA8VIdhe3PeZiwL9CZS9GaEtQaL
7oKPgZSOACbENBODneHQ8xJcyB82ZJiGRJJ/kq4a8YrySa4wE6sAiA72HmX5ZyYFuDekI7CZD3fh
AT/nXAkBsGRul09wR8h+4F5JprIK70wdWVvVtp0rHwmjMf8InpKJeE73RBXuq6vbM/HFCNawlqwr
BNpqb5tVMC9CXR6hs+X7eqIEiHsPmRwRIkjx3jZt5covt1mJ6wTWBhvYbL3Z6zEE75ZFFdOO0qsv
urGRqn12ZGR5dUMUwCecCoR4noBtE4AGBKJMn1aF4Ah+tAh6YhOTC/Bv2ajJIT+iNJk611mb7G5T
pXWTB1QiVrRQlHIwH73Tm+zhBAJgn7xxV7rNpZlnY1LLVmcjbu2d8re94XkR6Z6QnQMp3HlKgvCt
ZiLz2vTlARNY7opmX0REmu1bPFvfKEqBTLRomyOMAom8fVWybleklBAp21Xh7tAnMaF9HcNYZRA7
8zu4JoBNj0q0mvoq1mAj1XzYseJOClpqVTFQds3wdJYL0F9u0ybbAr5B1nZ7mb2KGZ+bOqCDI7oI
L3+C+NK0MQwQD0TgoSeByvgSn40BAxTuf0E7cylylEE95Zx8Q16OvtiENf3efQg2cM402oyl63XW
wjXZXY8TFwXE9WaUf5Ij/7fYxYfSO4yiJ+k6QSj9bdJkPJ68+tIHL/WNOPivKwDhgbJU5dxApCCq
EYVH/D4pTBBYWuzbk0RRq/MOOMDtsyIrDtineyM9BlZsRyGBKKh88AxaTXYKiIMIaMzBTGA7jp+T
hhLoP92fimJyZEls8ZXg98/dUV8QxCLc6m+QbmZ3edp1Fuu3XV45s6sNgI3EiZm9jDC6dnhrAUIV
KnuaRawco2ivWh8nRV86ZZZWoIPeihGbFNWZ8mR6DjvEnotM+jty43Ns6q80+r7/GOn/wXvPT2uG
49tkzqSzRJuyGdWyrSBacSUeuyMUt+jFTH+6fg3V+eHMpnwfms0ZlYnqnNZTTXug6VS7+a3l1AEz
I3wZVsnanOlJf0r/K3FRsOQqhp9fQWay4aZjJJB3vIOh/6qTCafbPdJWfQyzTPLizkKTY0CXmop9
z/UaO6yf74olMJQgeySl9pqUb7zCehLTrBp90aWTUrfgSZk7be2Qnr7dU0yf6BpDTdRi9Ir+7SyG
IgXDs4Gz+rMEQd6kn5wVb53Yo6ZNBh90X99s8QO8u1Buoc6XL9UdPAv/Z5HQX+1fSvNbI6gnDBKL
LbKb7W4exRuKnvemX3gGguYJO/J3ggnW4Qo0Q7C5OVYgwl4jNJjS8biNzziVaDOBEZIYCL8T1Af+
OJvgFcxqyXHjMURPrgkeK66ye0et6UFQ/Vu2BimwRK4s2KPAqVsT4jWLWvT0PdUxluyvwcXA3TwN
pdpxFk6fuZ/ndmqtMRVUv7DD30CxmgD8HJinXh1txRU0M6zFbpeK9PdCuv9V2J3UnYUVUTdWGEbI
Sju9kG8Z/Dg8eXZ/qpmLe5+hwmsgSnS3G1eHw8/B9V21Bj6H9OWjlg8GH4uznaySRXpTWvOsMcb5
HpeF0DYwIIcy4qKaxeCICF538u2dYPDNLE57FTHbZTTbkqpGll5sb++c3E9iN8RCPazf4+wcNrRQ
jzxuPJ99o2CGWOtgXZ6EDGGh7AqPGYeomppAXFsLrEBX4Yu3VAHz19fKsPGPcqsfssmoZ7yaWzM4
3dz916bA8qN0fvJ00uHBra1c1LICElGL9Ss/83dzRGO92n5X8j05k248weHUnxJzmHK4VjAXC13V
/FWLGWTZ57yXV4E6dnj49lNocZhsZadZeOn/KS6NAylq1Df3iS5Ds/23wd8OyCpw88p5IfihKtZg
Trg1XQKUN/de1c5C39lKdjdrQiG/yRrqIKnXpBVdyZ3XaVgj8M2uFCwpiiBLEO1WAs5YAKuvLUcC
5MmN/BJnLqV/HRtPYGjWmqQTSr0pt7THFPkK2uIQkHUH+lXQ55h8eQc0v8nuO91+izqFgpkUPgqQ
2ANxBGnhp33FLQ+5Vs9RWMuMUcAC4CwKc+MjpfMpmoJIkh3d88eNrtsBcB6b8Xdm7dSTem/MqlRm
qjTwrLUWxKh/DPstDDc3WapqIva1viLLVb9hu4TL6CyleB+L7dNZabmlrFOueN8WIPoJBvivCnly
nkwrqCel0a+fqYkBFza7DPYBegnII8yMci5RNP7DWY4KyqIMO28cA3hAfMM94inbjMactml20AN9
f5iujJYQpR3qS7kY8pDYQjOFK5evyIdjcCw25ijzH98TCqGUs1zGD3cni7X+Tyccq/OHXk/urZW4
4lmTds9xY/3PhlBKlXJVDQ9H67uy2zFZx70FbJPhto8JrnKL9kqnU76M2LiDuxdvKrF17lJjA6jL
WJ7HOyeLNskk6I0vYpcCuvgTxypDwgAUJBQ/AvLTrNXp9AGF4K/d2V6NTXij9v0amtYPqRMUjHck
9beKChzTbHZyA4aB2aKcrHmMOMPcJSYA5ASDJz5lyNMOHmHa5ZlgFO0O8pcsAyuU7s1mRlDOxqp0
zjXcpsi3EE3VXH9lmMRsO0jYvs9RqpJ39ad+FRowhtr4c6dvypcjwhWiANDDmFGqWpw4LV2i0h4y
WJxu7RZGhEAtXcfvbmtB3Lu3aC9VjQGD+OgDvpeImIJI8mXoVFNnZl4aZ7YpRR30WfStgUKWWn88
JSwm4mKohB2SNzbitS+ajZi7/ZWfO57OPtRIcxy5LFBbjtD1ONQz+TVxwHojtvPxPhPGsO903kdp
loeNZ7qpH3bflYm6Lk/ly1zU/prnQqKpFz2TbByfb2SQuboJPbSGS0M0GoywlcbnIRFUizBSXxNM
zqbTfdJHs60kx6qUQ1fxgzoJiDDS3+n6kuig8S/7cm2rlkPLtKLpwDa0IbiXupRhZSPnbMWTDRxp
Ws5BgAC73iDpXkI8w2tX1vis3VY5SzSr+lInjiY524qR+qPzwBMitAjvPzdU4h8VdNIJQNfZpu0r
2gwr0tV9CBPFk5rp9BXAYY6BBhbr0H+d5Ll68Erz/vfh/FgM3yG09gfZdzubPaw2PvAZHNE3QJta
FviRKzUEPkGbmJhEv4tl8bkVAacHx+XyKYhtVWWHjJbfaPYWHyspW6uGd/mflCktZX/T0zdebMAw
+V6WOz8hnpGrA6MnvS4fhrJEnw9dfzprQsucvHGuJUKSM3a41+Uo6VIuQlMFCqEppUTlwzfIKduh
P/ES70lFJ0SBS2x2gykXpTDXVRoExm3TbofeZICqdOO0MY7CYD2+d49JlI2XN14mC8x8E0qXlZuk
tLSXdehCu2cjCiKjkHLFanCmyvzOOGv52iZjp7DhpwhPkXIvonqnht9ovShcC3Tq1lCrVK02pNYS
NRqDmLEhBd9/GlrzZjz/x/sK27Iw5FeygMsPKErZo87nrRCvDsdpjM96NES7c6c38J611d1Cc78S
ps3gSJaBAfVq8z4vtDiqmkewa7Mg9h7L4dBGvIyOQfk5eCMLUEojGCweexIvsY1eEUjjQA2aRn10
CtAZK+oe6u1ryTN5ujtKUolKPF6VeUrqjZfO2nOCBj8VvkDBwBdV1oDzVcLt0oHlAK9Z+xRe3D1P
CYuRWC0tnGb0uRBzzXmgtY/Taq/s75dtMkX68FTd2uYWfsejf2N33KK3W4quY+ETJIMhuY7nXaJ6
8i+uniB0lbp8CWOXKMRNHBnu7V6ZAeWqqutaKYHqkbZv272Oi471jqWnpxTKUW08Ov7W+2qRuaqx
KsjJFBGozKtUEnRxFH7uCijRpyZg8/vwfNhsKWEzNBfvLaZK4RyeDEs94crZx5ombjW4KD4M4pbj
ANOhsqc42br2ysdZkF2B3bgMp3TSNAAkzMCrK7s8F0a+QrcL74A1OkS+VWteAQ5xpff/xMYVmqrH
L/hyL+NUFzyQGgRUG/XpbAyJFOvPV33Lsf9OL4E+0C9uhcqo1/9d1xOBkAhSKqlmTp79LhFEnG9x
MxSQCjdnusnzItC6RhinpShFMUDBvpxulJ2fxIHUN8TjFMBCdunlDULmK/MPwh6NLml74tK/Ti7e
/lXWF8BS6FtR19+vYVfMh8ZxlPuF+OLy18nGpGeXBoXi6rCTCQmp9Pv8TtncUKw8+vEpwo6Z5Vjf
uOENAX9MOIg6O6Uw606z0oTHZHfHINFArSNyQZOHKXe+yPFe1ubntAPZ7HNUF+mw/+GO1yy/Ia79
7Xl+h9Gyvd2IOgNYN9fmOkXOOlYFzxrYxNa3kOT18GSakDFq41zbjb2NdsKIjyStMGcPc64zKDG1
76vHME016O32JYwPiDr9mJkYTOnBvGxgARla8pYhMUrc9G1QhfOE9bIlNEvS+O/hP5HHeE9kLB0y
Xn7LKAikuFnI+y0J3KdxDqZ2JpRRsrzLxEJ+Xk6m1EjSzCSKDWZs6oFdiiFLBtzrYQD1mbjkX0iK
Jmc7xMN+KxegqKu3J7fzqpBUA9NUhCRWHl6I7LKkj/y1o/CAfTW4a1Mpilb6sXRENmAQW6DpmllS
Vjhznbrd5F1ZTZQ9uBSl/G2nhTXqNOhBwFt+zBC9xt0lFv8K9zgNXCgVtVW9jwWex+nzHZ5ImgFU
DeRKMrWfxRstKlxDIK+bMFGrIK0bycriaKzLZ7oOiC+7E3y3PQda+mqy/jkTWcZYMwuEvnUk0fWx
uRGuunvJxWKvfttSRj7mWSjwQ+OMJVRrEvqe+K0t49/HFye446ivXW2EWI1fqDSMxsI6IHlMuOpF
/jWuo5gOlRfmFk9Y0CO/TdEyXrD7skmppo3/uLydrqhVRXdOi2/3aD2SyIjN9fvoLjWdsQqkBrzs
m3TujSUzGWR808cw7l+de0Y2mxva4CVQLqN04K/4MD0uiPa8oECOWeJZJ+GAD4pqF4eqPBPj2ImC
13OtcmqksCwMi/r5pxBTNHRjnOFSe3BTj6kQLhz5y23ufQwk0Dh3emnRoHorz5nrMRZLxDpCVIpG
p+aT+cyj3A+CJ+qrZqlamZ/ozyWw5eVd8BFf1uV4nuenxhnpIfgHVP8erg6yRk8iuwSW3H7GGeD1
DiZ7yk3jNkyrExYGCHyD0X01jciszByOXVhK9PlLW/0oOjVBZ/GdtzlupvjW7nuI19o9Kn0QeQLe
Pzn8Yhp/BkPXu3E4jgw9lLTbQSDgfH01U0gcy6wNWyo1ftM0qQBg6L0MFTazi/nJD8RK6NHnN9AM
V4a7d1YLI3yNwjRn5+zRDtNGEN9rG881Lk9x+sbCEydRVRN2TuBImOPoc+PcS5ZpUjTQvBAUljPp
2PZruT1lWKxcEyb1LrKHJ+qqKxQfGE9iVLLOJ8eCxpiv6TioueblcU8w0KSL/eM+j5lo/Y1zOk0b
yk9WiNvjDbRVubezMAieTAHOCdZKAs9XS96PbUhR1TLGY4P3gnxlK1DOvEyFzB9utrzhDZxAO7jC
BzxQ4nw5HEWs1U6xgSX9ZNiznJhmK679mvbMstxvcBWXgehZfH7JIPK0mo2l1l0iiEmfO9+tMNCU
CUNXcme3yk5muuOhsw2Hj8Mk2z93fcasP/xwcf9fHYkKQWURqkdS2ymzAp48Eu8Pd/KYaOghHcau
Kngb2dtp9Y4l0jEpPwYn1BJmBcX9E4dGMkYxHY2WXnITyONb5hNcMzjRYscO4XLTD9TvLN9LDbJy
YcdoUv050EAAuRZfCTgldgWOQxCaJa3goT+WNnS3cXXj39+7eNS7RAw6UoneuScVcbASoeRLOFQM
exwAisKu+JNArXcioAVv1LyifnnZmyI5cXshG7OcQi/GAkO0ugj2eJKyh5UzYAdne7UT125qv+FA
cpxj7Ow+1z8BrQBU6AR306HVI6ErY6ibHTi98OUmDcvnTo1Ns3ZTb/aJMOReHZawsWLEQH9r/wMG
VOT4uV9eGYnmLbLJ1z29NnGxBY8pjdd8XC/tJI/uEYR3uz7EvMLoDwPVaYTjMJegqAWvH3lu2hC/
+JFcOVgkeXjxQx6Nk6H4FbbmvctwfCWHBNCiuxCmzHD7lbiVlc9Ke2zkW43nxpRgPInYQsyWBESz
m8AmRgVaj/HsgtSOQP0WVagwMpxriczDWtFjkQArEA5Cs6QKnCdaeNt27HCFJJhAlR2Z21Rvfqtm
jXhxf8v5yAsfAEuDv1CiBY+9yQ1nm4CRYWKz9xEy0mBwtdtZUSFInW29fed3Nzt/5WO0iJx4E/AL
nsWxjDWQ8jjIUFQyToRMW0fanP7toGOIjx/Q5Y8EKhHLRCa48oV8m2L+mnTB8imIQh3fzSA8QUcR
88AtMdbaDi5E1ZxG15tosZ7w8w3mS0Pds8a2oKZsElnWLpsUFJUrOTbrxKEC5pe4RFaO9NW+Loch
wKgoB/RVfQw9u0x4EtpzlzvklWywb/GxNTkJtFYg+aVooeqVNl/D+p26/wSYreke9rF1cSDe3dJ0
05VMyaoVAipysxEktmK889I67s5GjJCTlHcABcEjAdBbdJxFhYDFImuR2RG0OtKU8pojHEmb3bVo
k6k8m6EOVwd45PYiJBloSQrQn/7E3QSkhkwgh1tvMMipnfbBAmbNT2R3GrfbT5zc9k/m5A+/3rIk
t4mNjSKwvs6NrrALnQfcosjh82m8gQRgaMXA9EKv5KUW5i9bxVBwBI3k/0/vx5kd91XCB91O07sw
dlMGUm+8Zxmm0WrxO8UYDivrMy7Sqc64IRWF75TycFwA5FVyxDJj+GTekdPxl3Hxeso8maHs0pOO
CpApCMMJfmxoVd2RXpQ6Nw0PuHjVwvBWKamZ49DBUD8F2BvoeJYJtdE4f8mzR83TMAcIXAtRvII5
qwkSw+5CaUviqXIGHTb7aXWy0iCf6sFkY7ihY2u//4e1bgED6ItNTyylge4xTm++jCuBoFAHSiBa
7Wub3JQiLF1jDPR3EiqpXpk2hk6gjLrjKl7F76KT3PRVVDxBhTnKFMOd/gCB1QYBHTIFkHhd/h0A
RrwLeWCAwsV8daI92QCU9z0/iZ8sscQ1/fHuJ/qAdLE4VkCXWFw6y4aqAEOfaefhfz3hRjtgc3mZ
0p5TkAqkMj86xwbcMlER+HUfj3YMZTJv/dYFyWndvzHTD/Qn7FakYWiJFP4ONS+vIKUW6mjQ5Ibk
Ib47AeXKK9mhaz+sTQPdqLSp8BYasXhB5KNO5cbqnWhsJcp9pA6FoiEewlt0/xTSOK5fSY6ai37Z
cS9RF106zr2F6XT/beiZrbpWGk72JVKvoQrS+CVeXE288f5ebdFJaz141Ri0CvKrVevediwDogll
ZpYcXPxtyLch3YbocLD5MtmudduawjFPVKkOF2bi1sYdIPqF34/wZkKeI5n2/v5rgzJRzn2AZ8L0
ngayCmrXpYAzvRIVAb1QESJC1eGw4D84M4BMSycI/b2UwPvsbcGofNk7GUQ+fYq7OiFKlAl+1yXG
dEydLGAcmAYlvu63Nj1a26j10u6M8GQmOro6lDi4oRif+7/LRbkeGgeJB0SQwL9f947i1BvRJoF/
N2p/XDZxOpcqvMshbCJF4RJNwrif2n1lfQhu+PFIYFUTMPDfX2yGryVSzR4fEvE5jH/ar91oRzm+
LrU6b4rkE7YZ/wjzyV2SuXZnYJw7JYw6YifaN2lmn7tqXE+bP+WuNl+8SE1InuUH1Nm+hCfva6sQ
VP6DsD8EovaiWcrjiJR/FMtu0/RH1fA7K3kGA4dcbb/ON/fjHNaFTs3eOlvYxnFnY6GqcAz9gM7U
oYo12GGMp2tkk99N+l+84q66vOKl/LiaDRfVzeXqPPioj0eeEIENOSDwVrSwU9Mefox9ZXNxWOK7
yWrbZGixD5eBZS8Db9KwZukv0Lr3v/ue+BPPgIQ+NFfDT150yO+S+s8t6j3v2480PIHwvgbKZHl5
UegUDX/XTkqFHArGP5gGFgvZ3XNwuVbKPIIr1ewSewhOz0ckjghP+ZWsTDo2bcubX4wdH68SRZmC
/wLrCyfBkORm2Lmc25TX+O7oQkcfmjnieBwUw1SzUVY9k+fRQWWi3dcQhJpKOOHMQ5Kq0z20toiH
FeovEawEXfQkNhUWB5XjLJUzmcgvHy6wxxoPo7I0EOPOoe0M82Rn+taGqcCW+7pn5PoK1Q/hemuo
OsEdAdKmeNn+bzdaOdIw7D9R94NGVn5IdJfIURBhjQG3j63VwVLESX3DLQqfZtG/jZyxrAOhbG94
j63oJDo2p2DsdtWch/WZZOS2MdIIJvscqGTL/cnVlEt95tzTPy2T6W1DC+arQwzl3HszzizezPJx
WGEijSB2csJw4zznXk1g/kqp0BORCgbrQiAsSJ3VnWhlD10Sxv6e4C7QCr4zZVEJTLZEp+oMdu90
3QwIoav6FeJfzAyDhHsCLD6uDSacfdFhezQrO5SDKyMQvb028crYsY8eZfcF1Ds/niJTAc2tBocT
s2lJ0SjFaw6RUhkpGlU8m6wpx0MZtLg8k0MGS1OJYS+X8OGHkWnUDlHXyZbCsIAPaUHpMn/Z3nVI
6IavPXgokBL4ar9SgobufpOIIGdpK5Yk0CVueslPHOOn1pCCxKvpCQ5GJb+YQZqwToYQTXcf8JhW
ttKWOrZRLixMXKrbq2FT+xLhpRjjU/p9Ac67HwKmUV5xAa3sg0eGcdMVR8oS9js6yiyEmKfQF8c6
0/jUTj3UPhzq/xnvZBGvXxbRTBupcvmpZM9V8eq3xPoQannvjfJst28tO1GZFpKlNuZbTc5qrIhw
5c2Qoso/fxtCisc740giKn7fR9fCtPU9p4Jjv8AdpuiaX9zRZY5208Lfx5z/5+f2p9BYoGxDOBtQ
hgu6MleB+IEOYyksTeiyguoK/7WjGEbdb0Fj85+xskAK9jF1NILe3mj/GgcPaHbnnvWSIa9u3B7b
zoMhQLqIew7dnTNMIUGODemGPSgA7i8z6Et4lYgbkm4lk9T1xbXz3MkeqwCkUtVed2JfCVGms7cN
yooaytjh3JX5uBwAG2mFz2en6u/NXC0JSn7kUWzEugCS7nVEmrRl3ZAMfULiKA9QC2S4yPXfBzGu
zaNaaKXs3ErAj4CUMYe8vojwDh+C+6G8Ohux5mFOAOa6V9yHk4dL4ezfHYnOeJcK9noAoM35DYET
lt8ncQydcQmY2laa1GUC/M8Zk4kmL4A14RrOHlQ4rFyjQSJZH203pfz8atS7IjNGW0j00Az8UkTR
N10jr6+WrwJYfKaVkcutdUWrvOlkBtCTyOHkhlR+AnNkWH3yxtnjEZV/XQ9W7irdn0wvMh25BaPE
kk0RxafF/je6+7sXiW9G1tJkol0zoToyGGbb9anONCft9G74q9+fcoZ2/4JJztScfrD+dXxHw9SF
Tqqg6I/5JNAeW6QrMtQ4ijUZiSP0B3ovWH66DcM+J38p6/ca64cfucuUYD/TqPCpylyQH7JOidzv
ELKMWqle2ejnovZvI0B/uL3C4HcLdI/kzHPyTZj263UKMuwXrwDWNyI5eVbMaEo+xntGqkxmyPNI
tgE9YKxEHVUYLifbm2/p1s9osMDvzRJx7OlH/zPCAPphDylIEwHeeEnIClWoigX+yEt4s8dXbS7b
4jotFoHdUTzBQyAtPLMc4GtW5cqJ4KVjGb3VKSyh/ysbKgcSfbN7pfmsWgS9eJEOfcijAwfm3JE0
ZMo9T7b5mHS3sk4TC5B99qOpwr9tzENR9MRI8VmOsVW5fyi/6Vt3HcC/Gq0aUsM7A8B+ZbxLIcG0
jftMZDoUTOxY9iKfQNe688FAvZ4Vgy3mcAKGSy2jAV2FCAeOeOBCFmy2BZw81PDzTkJVQrbFk4SA
z7F3oejbQEnu3XYBNO5bILIgp160cBpEyQ0gBKNYoGH7A64Kmc1Sh48kjSDlx+bsIJjUATDJBQln
ce/ip6AJcFwiMJLJ9G/EepulFWhZ1VfSKITkrFF9LUNIWmNn9LIhNEaa2S0MSGsVH0xPla9JM5nM
P64HTUKeJllSx9w+0+DyWNj82Xt3YEimku6wwzFIdGUWS3wVb7MNXl7bZYXB7CR86137Ub6siYLE
NtDfaDUE8hAAjIiVSYjkNB03yJT3u6+fRVZpid1wLkoMW8hi0VsCbjiThuV7xXfMYNZ//OrSHog8
fjicC5+ltCQf/xJ8drWKGQUTbR711SvSYE7rWC+zy/e6txozkMdAAgpmEM8MGhanllvK2AxG+3uP
45El8dhFlnWEA6R+oReReViaK/ZkYIlj38WuW72Vsi3QhO/GtAURnIkyJCDJ49HtxmihhzzES6Jb
Ix1Szo3lpIuxZiiBdqYC2Fax3+gRflJHYK/OZhfO2jOLSryGgfS9cNCUZQa378p3TgGsXBgCM1D1
q8PV9NC6ygYWb5fm1Brq8puilPan3OgKnPeZTv6mmgyN1MpsaPmB523Qqz3DMBuNX3kTOJaFnrvk
mjyOco1TOSqmun7Yr3SZAvQn0sNQqy37UV6PDiiFEBVDB6XXYh0E8no7lUxt6ADAmtbRbc3gS7NI
LmDq2dpNEx4dfSRNH4xqcx6siMF6OG6nBLNE9Jq+9wVLSW0caymU8vgMJzF0cToxs/tfhxBL7wTZ
N6jWO/G9bV4xPBGE2YNFxmmFoXb+xOhk6vGpl8cxcIonAuaT4v3DhOCSS3FHlAN4TejvmZzpGmc7
ht9yMhqUd5SVawsAkv21G2RxIrb8cTmQlP8VR+NCBO2Z3f00ijLBmVPvAxhtNAF79BFSrVGvWz0+
4nTIN/5dE6Ne1gaimCf2LP6zHJqs6MF5aDj70QXtlYtLHOprh+vc+AwVWvD10q13DToSiOHGof7W
TgWAj9LwNvloB05QuXdWfsrRU2JaEqTNCxt6RRdm3Zo657jHH4BCmHah/J2p5GbuKo8UCMCf9veS
YIfBIFyAHpzuUsWlKzNExiT4UNDpmRi4xhStOf27vuX3LfEu6FbyV+z6miOu5sGvLka1Boj196Yp
R94/RwGzLvvV2DDrMBgOBRnJoX+pZA2AH64wnRtyZkyty5uPKHehqR1DRQI7W8HMzkP9T9+b78n3
xtf9RS0AyCHtKmI573Idk5hz8atwN+kG29VnW6uwWlj3N6oJBuAeBbzwDm8KTLSu0qoh28Enc/f2
bJoFeh8kBs/aNxJvK/CfuDRBFhPkEivNrzfKSjTx7Mpa7LlHF/CFzA9rrtla76HuQchmSdKW6Yul
T8t+dNuC1BrPfvN9JtVvJlkpaOYzea6TJkcbQa/sDGzQrZfawckdcxI4WFgD94LLX/kVKQJb5EEe
N8NgBSc7r8elQLrH1ETLnjSzSREv3JjONpXL6zwTrV3JGPZoCMFhkjRthzc7mAvNvh9iHuWtAkgP
5RwAPjd6IcARrEtfXF8sgEGt5kpinks0RVNJEUepCiaHB/1Q4FMJ6GzUoPU+AveASTOQroEyTcVi
X+JHBy5sPeGBsPyW86s/B2mAtw8HROuh94ZZX/cPKfIySRVQEutiXQdfy4Sq3YNyPPqBaMoM9gZ1
4l54Efzq/WmOnt5KDg74jRxzCBJXDXlb1tte5pvpF649OFrAUOuKU8griYIoFdyzZAD6tP4xEvDs
P8zAjUNJ0KVUvEEg99uUHRdfbBjqA5FOUsME7q4nb9NthfkscnDwZruomz0lndmD3ADF/XXxH/XA
zOvlMzsbpcNPSofS3TgkenqlCTKBFx33/i+Ufbw30dKC4Jyb6oyHAcoUo2xekv/IIYWtifv1OIeA
tYgMTSCOHupf5V5htwgatnp+Zaiy0hH5/wKKkw45m/TP983ga2e17aGO7Xb13FGKglYV3xXHe4L1
om/twHd6Goabgyw+K0TqySTbCZ9ESbCdmDA2IIJ7vsWcGBk3qEXX6I6pi672WodaN18t4eoYFGTs
AV9EYu0MJ5n4iAPYapRClNO9XRYGmdeteQWLatcs07AgWfzUyZ0jOBFZrTFaXO12yH/E4JNaMyfS
r4SDj+x1CtPUJBF28JVeFApH4TJYcCoBr6q+Ok/n4AfJcZn16Ng8cN6kmHlXnw7FTY5xfc+2CTpK
dO648pfOirzBU/qLSbC7a0JulnqcZ5zTps3/iunzbtEwF6dDN20j3G0N9vU+JZyNFcpeOFPFyqM0
dWvuKEu2sYXDSrUVw4g1pD/yT7dKRLAJYF4dLrCT1kiLGTC2dh14RXd2TkZ9Xe+w2KJpYzoE2RSS
UcemIj0qyOZHRyWsIDAsVuQuRmxmoF1i0ZqdN5Ae3zrE+nRdWgs/s9pCe9QnW1iexoxZM1HUEJPL
CKuEaCd8W32j4zyte5W8w5XNZ0lGWnhUrJS2rU142esKp/DTJiQmmeSIywU1RbUCRXRnM6cGRAK9
jeztu10XcW8vY+T7fyM74Vr5d0egmH2au3pyQnyb4jNjQKJ4Zk1+tI472PepC0j4OhkveQu5D696
NvSVxP6l+UoExJaB+Cqc7tnvwXYyfzz/Rw3Jx3LkppDZ50VKJUaK775diIEDI//+iUcURGRDSEie
A31REMHzWcp/z6auHjpIDNrXV/txhlzEqchyV5Nj+AWuZhX+Zn2j+wuqNP2IWa+au3G4OcH9LwOp
VXnQihOSfIfuJbWV5a88U+xFr+WQWVjDRYqwPNyc5mD1RtGiAY357AMXPrIrhX2YXzctcTCXOubE
1Agoya0d5o5vsJyo5KbNAi66Xx41U6yc31f2tkCtS8O4FCzwNkPvlYRMwYm6GV7IfWFZ9nP/38zB
FNBaxBwDe5MJOQzjNw5LHVyo+iMjr7/PspA/6OdHcGQIz26WXIjl6KfyKFMKl557XDM9m7l8Xd1G
Pp7MDKF6tTy7KEMwbFtcUSbgyvFPMFKeCRuvLZxbOFzGr1o8UbAJgxC4ZNs/4J32CVTUb/UC6EnK
kYahJ8cue6c7tOiE9VXB20hO51ZqclATS1xB1JbA1CmQvIg6vNCi9W1qfc6SYL1EoYxxnrMVVBm6
HucrAYKXhgBh9EffZRDf2trQR3MmWTkx5pbOmVTNWXT4HgLsJw3GG9VFUlbdG3nTnumkxXN5zNpI
wYY3S3X5GAFXJs7DurgEilQIFnuiHEPS42EKH7lym3GYbZIMiAkN/Pqqgu04ZcA5ttsTjwWtrI4t
8B+9MJys5BGL56tqt3Vc3/jjOohj6LHngOjtgpS9dBnjcDU/6d7SgKu3HUiTQ7ujxknoK0jdPQ+T
VPCrFC4J8MH5YppqSuH3MbH0LAOFJj0awHr/i9zTyFqlBq2nssgvjVUc5EjL6w7c+1OJsyuKbg0m
FRUrj72pMjWcW7lLjg/PNA6KyTVvJdahERhu0equFUJm8L+YM7crT69o5ZzUEnDvKGdNV9UHWHEb
7CIRL2njWDw2AkHODC0k7cg9q+2VY46ujix4wrN4JywIB4Y+wwoviaxTStwUVuz1BWOLxwDbnuZJ
I2fo5nBLLDV8bq6i/jDScrxaW5lRJdosMCDbj+4Qm0D5We0Z7OSZX9yjrMc9rEBJIlabd0CKR2t6
BHNik+Sur7Da9aHsaIVdTlcI8dyubLhbP4dLulVXWPvcjehrF+n5Dhx9UXtexH8PHawgxN0C2GBh
eY3uj6qLsz0m7z9DsniZcKOw/lD7+/W41BrCust2s9KbjYf1EPY+d7AKmEnxAPrnB9coeW5u7ikt
Wm14iYWAAAIqb7hHm5mxR9+hVZM0mWHAltt23P7GeTzzBBXK30ErbTw9K+L+IvWBPhyY7HW3IDuT
ArjIjxO9aGWrjdWVVFaBawHyLs6/ySB5G7FvmmYLabbZT6BNOvSCVciNdUMzgj9D4NIzPI9P8Oyb
DQ6dZbcaKVUKRYDl4GjMAijFQ3Ajn3AwSiNE6fgPGn+LV0VtAHWwbYAZkMEkg21v9KUUVhhaluKC
CSzLFXkmYNcEHbEWnqLyKN7aefA1p5dEt8ZsISFgFvCFNIKb+KhvFQPrFgnWS+RkqBSnTNj2K8Xu
Tm39ISzGavxCiYyNl/0vEEL2vaw7H05uQ91JoV4PHjVYAzRMN0h/InYHIGLrboqStEzYCw0oWkUg
U0ZZET7R3iRkKiipZ8HmHkjRaI70N66rbxVA4RbTGVTxmxQzrRkyv8Z5hrZ/dKHjSIn2VNTKzLCC
Jy7JTN6ydJwXkERvd0KJxLTmNphau/yn+Xirm6y9BsnDqBJ1M+ASAFHCe3HFKAa+YKWG49kxw3zy
9JwsdJXKfi5+PlfDp6qgPEfbDGdq7gzBAW7nUCeDB/31uMDpjV4vk2Tklo18NL7qe9vkcB2wJNKq
f52TzxojmvB9PpK1GiDNtYvQ+djtYH2lV6oQ1Z8mfuUeEhnXnnejKTTy/C9hwXduqXP+n9Krpyw2
EIp7qX0ay4oCVGBkj9fk/JvNaUTIgao9LKW+dy/vT7h9R5hEJz25L+EyENOizCLt8DUMQ+EtvEUK
0OY7VtlVnbVcZCT3yRFWko6+o8DmsCYOKLWf+1D/543RdM1df/g0QrCW4n5iqNJ6kJscqR8DhzDT
zYIx+KI4y5Nx9bgflFqm7Noth4ov46BskXdLBZeC6PF3+OolP2AoqqbfaAmEdAGhI3/CzaIlmuS+
1PpGlM7tSE2MVvHNMUNfRWd0tJlr1ncmJXYPYM3sqAYRNDr3NJHgL6QUfPJnMHxc532BwHrlnX6q
VPprf2H2fDYZJs8Pvp+4dUH8kziEV2D37sXf8n4YTUb9xWTPW1Wg+0qI9cyM25E/P8VApI/SWWqn
+Gz5SasFQsPfc1zs9pa8a1AUDLPQKp3MitL2lHwQF4FrwHpA5SooU9YJBMdMicoi2rBBazmr7edS
XjMWEJ/ZNNrOP6+B2rjMoCMWf2RzAG9OPYUzGhlP7xtFBoOVvwNqsD2f+KE8BpRr7RP87efiH5ct
iZ7dL58jd+KJ1aca9a7s19dezM3aJjWf9cVNWvMP5UO13vaM0jZBXO5JSMBHvucaiQqQqvDiIrK6
93s8A4e0EOohVf9cQnADzrxgzcb6PmM4zN+CTYty6J/xzQBuBO2UKMgT23d91IV2HILECX5JiOhs
39g6wpLpIozF2Sf+v2C3iAH8PQiEnR3d4W1oDon7JPACLI6uRtZE0Grp+m2Ye09SuoZ7yUUCJprk
spXb338n3p6JSFRr2ABsqDDnFTeFXGudHTwdx3TUXm2xf5hyh5v3Z6DqigkfXStggeLBcMeXbSBl
bVmiLu+N0KEppAwzKnO3POPZlYBkr76YtxwjANOPlR+t2tdi5VdTXW469Iw8kyyj7/1puAhRczfN
IQ/Uele3wVg3GP2PSyvhCIas0X2jwOsVbrDSuqTYDBH4ysCf2imZZjJPECo4EBXepDZ9NxWFzDdV
vMiSTjWGECJq1BAFO3ATJ6iTOGdbWVcL+T/Q3K8dcCl89yPpziqno3dKv1MydyM5G6cTomEOiJ1O
prHXV4/pUo4XfpJsvyDy9rq9W+OlWLoZFmpvzzv827qdWVju1+jIm+0kDXWuO+Q9Re4r3X15A/PJ
un1qzqgLT2sLmtkKGYKcOjmIzG+rIfn8o8XKnYSvzvTJnf3ZlfUwbL1xHstyoWOXmSJlVbCqm2Rq
hhAfudOpTD5Sr4+/p5AXynXje9RLCCHbZ14JxRSuahDVXENx0ymGvJC+yz1gCk/4Y0W6mlCnmx8N
RU+3TCr5ZVWKuDuy1P9T0pQ3bGI0cKChmWtWc63f7i6sXS/T3/thJxGyinSnLiDsuX8/WN69AkCQ
azt+X29oPzUwB3yPuCdQj618QmztGvsbXGz5LTRsKaJzukN8YYsxfZfmNl0bY0/lzZ/X5fJkixD+
+FdIaAvVAfXgkZJrwPRmcCefiXqSAl3Bs/LKC7VBFtt9rq1Telhk/JywnpCgtnghxuRm+rivyTOk
4tDWOImu4rsHXbjgRwnuahkKJo1QSlW59Jr1RIV8TH6ryM0mYO2OswVrnRGsW6k+cFQYyR4qG5Z6
ctOCZOq6xcaMyH69Uwxn39ECZ2vI+U8ZJl2ItJEBMkXhJa6TDm0VmtxZVjHqO3Yp2fPt74l4JDLU
wOw2Zacas7x+5aCcgFYGNc5tR0sfn38xCc9c82kz9aG6GvvqWF5cMN8IE82q66vKQ+sgpA8nep4y
BfkDP6HTU6hLBLHxUH8O0MRizZ3QGIcsWYFnQ/MT9fTRElhBtirEuYiU577IpwnRwn9tRG1u6w6o
cLkLq1gAiX7SaECcodSocKDw0b02tJKxsynv8F/fUkJ1EqOpaWlnRjmmDY7kf14IixxpFG1Ns8HU
/QY8KTR9X+GqcLVmZ+ky8UFdTfWaYKktqNCtlhF9b4O1G4BbHy9hxnHYF8jNkdty2O1ZWl5kNYd+
YyhGFwoZGr7LTmsMg3JeBK37nJX+yZ1AmHvD5Q4m+JqTsO8thlwIa5tfZ6NCItvNYF2ifydNR3Kd
5M6KPLOtnB8ojTp3JTzmBa7SMkDCy47e5yY6HI1+XLS2lH13ZAHCQMumO+RnWO+s7sVo43D3WW11
SWsRNdKNhMM2zQ8jowaR6a5y7bLJ5FSyaWQHY8dEeTofTIuYR/1zZtppH3wRPxVXDu+oA+11m2l/
oPr+WVs9c8/FOFIiWTQXmxsEBLKPRGAJbGktethj6bm27Xg1nc2t5d2OTlDZnzv5VXVPe6fdnCip
P6YUNxykup6vNKai/aXZDiESrz0beWjdtYhnCQuKSKiEnSBl9rQjY1pdd4RWYTBrk6HrVgPJyLFI
Ve+JrsG6TAx4SKMnT2bfmX/im4c8bfVjoeA5+p172y0rV4bwNP6qAxny3G7ucAfb6nojXXoYC58A
ivoNEZJEIBtgCMkj8a5JHjvm5kP4OvB/dZ6mIjAi+qgJqwJnMrR10LD0NLYyjOpiYOmhTSLR/qJ4
xM8OBK9KZ6XjBOdOhhlrdSTlrCOSBo3Lya8GCR53wCZ3ASi1O8k86Nhu4C1MVR7yuMtKTeAFaVGm
U8Pl7ge7+iBDwE+mv+EaB+d2DEvjE5obKFliwrO0weLV5APIsRKnPjtrp2QFXWV/ZxRRMG0nuJaG
Sp31xlV/CG2TsCxdW2DFdtlSc4bz29eUYiqsZuXNnJufX6EOx1glIPawK2O7boxB8HCEXo0B36p6
1KEnLSaqlguzO7gRQhfKeZ/ZHHOfR3+QhRGTtEbyNNg71+2qQCIeSjvalJnnOHR+sgRdVepoE/EM
D6kqFAgvT/wJ7m+Ggdi1BUXHZfDN1t0mbJfez0sDzq0ddw8DjGbmiitRCEkqFu9ZT93B/0RBbL7W
Ph0poYUfAn8pmASVVhiorLL439hlb09wfT+cMU7PLSpEubYoT/sb8xJDi4TYnYlxCLTFZtKleFpY
ya4A++7jViAw6R41UeKOqKZBxKZd8p1iOPwl7pqX7s/qbZtYy3pahnGitwfKXafVvAa6/h5SViyV
yV+NGFUelowUpVxhYepu9TroJGRmlORxnpjJkDwaEU0ww4HYe4at/gx178BROuVxuuFqzU/SkNfr
lhJ/lNrZ9hPdFjEnlsrJsXpyPBUoKGghAu+N5wyQ+l1dYuX5UtamebEvMEJLmA0CcL7kVtWqKJm3
c8ES/ZG1E3GYn7k/yTMUpdATZj+Lf6wlwmfLzWVfVPW7b3SSxyWfxKv8WhAsc5zNsV6nYfzjeVec
bO3C13ZU2S6n4/pIkmB0RNwhejf2Ddc8j+JYkn1owz8qzllSgP8X72HEL6nyrbvA3f2HDRcaR1Tk
RzfE0E2tIJV7RzB5mdiorgJZmE/Qwy/tQ4pV32sJaKtas6X7gjpI0yge4Sisty9PIhHiHIHEUSjE
TVyx8DY8abSclgjImqLFYuUWLOxv+artp4WaWW4x7UQzjjGoXhoR/4iXP3hVDPWHEi/bYA5K/OXJ
e5KHd7KpaFUkMHhiOTQD7qwoY4J31jIcTO4KTvKdXCznSBdMbWyeMSm3M0y9rlPWyb717ylV7Iti
a4woK9AW5Gp6IehkkaU4U3vccK1s8K8h1ubjSw/s71jo/Exp46467dMHUKtTdih+Eq1UddqqnI34
jKuVeLS7eoBvTSzUJJykDTHg1TZHp6Gs3PEHWInA3yYY+2U5WNkV6eR3AAeuPf9IOKC0qbklANHz
XlRm0SUAZWeNIl5+UQzMBEFoA75iGGo1L2icsV1X5jjBBB799mEjmqMnUqCQCkbnQcubEj87RNY9
2wO4CPyUmI76u/xwAarji8TMEFMYjR1HphJxEnjfTzp8AaakjXzwbxd2cWibDHwc4NUtNCjcvtxo
JiUhzQhzJs6uOXi0G0TeSDMn2wz/95wL6Q7vjK33eYiPheoz1LVj6IzWjdxsrewt6XctXA74hiqb
NgPWv5qh0ZlirprYVGGdcUDpKvNiu02ljbgg8U9JfoZGLKKW5yqwkr9uoYzcss/XpTd+gNkVum9W
R4RJ67cmAgQxn82M+RPjI5jplevz48YryZ9d03qQSklZxbvUeZuO/SOAcIlcVQo1Jzu0ouv+2vYG
IzU908cdbiCD7aPZmHMq60u+brnRLvjbs0CEDsDsV9Qv7IXj4hERjbGpwLUQ090JhRvq5TiE0fpL
amCOjb5LbDfmSaHx145e6NXHWL0QxkfRWSjpMxAG6nla4a0xG7q2/+/64ILoqlo5rX+eNM3NJ8fq
jTktjIlleRLhYV0AhKbghZr6aHz7KcAlw5Tfj10QlLc7BPsmzNJjwjRrTU7cOdBXlEAgZENURjNB
O+0PUifgNUCG4TPFZJ9Nawa8go1OwxHD9iGRoHM40nODfegfelRywZo9ScgPfJe36GbXglc3dMeZ
jy1a8qjDiBKG24Z8igQc6NW9jG6B6EbfUg6AYp0UhkbL7i/ez4dIvBtrkraBmW01J1eLY4nKzs2m
ssJhPxRHQLGzvuvGMylFDf4a1mxhvZU2zCRG2ZdQdb3aZqCxI91z7m6mUNRQVcoyV6b0PNboswob
2mofq7iAICnQZTJpTYRrsKuVfcwTEGztusrNqdrH0GzkwWTQ7eRNQZ6ORlj19ytVBSxADwpVxO3n
EWb0BdEvuLaio3iR+33OFyWhMby8tN9weEltw0WC+X00lbjoi7e9RSi8l85SsmodmACoFAkZrClS
00iGwztjBbw22XMsUIRltLQFGqLircOLbKqUslFFtEyVy/YaCItKfFvCeqnUW+3Bm3KXtbAMdCbk
h70z4tS1fJ7Neqnh3sKi9yuuSxia4TXFoOtQu3zJA7idnVMPn0QDZbo3l9Wfhgc+LxiWqN7Nnb68
Ub8knFYq7bOVv5O+q2FrzzO5mdYcTxdn9SkVp3D4TiO+Q00E8SIm4iLmqsgomWGMm6oYUte0oqDw
Bo44iguGYQ6vFMkByRldJMh5gD6kbQjn4LaMAkbp78tBgQ2b5WREIM1bkEmA1xD4SNGdhQvoXVJf
jW+BpQ0uvHczLeVMR/mgjmyAs3STdUxPyMZL2fxGae1H0M3t3FfdRXOp8YNRkujzoDQ//zk3/9/Z
1/CgN42VxafUkV0SQOBY4PndtAfgYeaRvpJRH4fXR5s/M9CAt4mXPzTke1YGCcf4iciPSSWxt6QL
HDU7zeANn0Zel1wgTxhf3TDfqrL7yc39oN6ArqhayqpXVux2ELLCqqDh5zeUKkaRnWVulv16bwwf
YeA4kjc16JnHAHQGcgXCXOkBAi1CSLxBGQv1Dq+PVebMwu63erzBwtKp24AnoMwduPe8ySaDIfzQ
54G7kPRDRsNsHEaYJ7zcbOKvupkBth64zf1y/qxirApf+yKSsM66HA6p2QFQHGLrtRAOBCVG1XUM
5chEssl6gotfIR3QfQgacoM4noUuxW4CxMD3EZpRETot+p5MaBMnSqw/PcHwUpYSn/IFJeL8gPeo
6G60rlc6wltwdY5YGsNr8acQAy5rsKYUEz0Upb72R/B4Wotxm0Wb/dg60kWBhp4dlNwNANU6j3s6
7hU0c2xIg2WDIskG+hIJoz4gysF8o5mkMc4JUbqB5zrVUBMTi8GbWurND0spuFM9UyvHUCT/uzr/
cJErlAeb1DpqJjVH6NG2d7et6YWovaWkBs/DdvkcCa1+gSHoo1XH/UEGn+4lgVa+pcmul8kSIJR7
uvk8KwUsDLNFOn/3cnHnM+fcin+PPjT9aYVg4N1Pt25lV8krSxJOmDtqAdfxPa7VoM7G7/jCv9bF
2ZeJaQlKg2vDuDnjuA0F1bjhLYZBZbqq++oW59aSwszxPzgKWwHQgM6gwvuKpT+F3aPeOPy6FIa2
U3Draf7hP+OgnojYGkWHqedOJ8+a8M8za3RTA9KjgAzODUfTCM9dy7I8QB4hvirmc4B0e+VAkKwk
7JH+m0y9DMCyXU74FLlYmp7/yRUt9HzgTX6XFtR6luf/QMDTJoqP9UB7WI4jrPknH3xpTCk2SRpS
LFZ+78i3hb+1kI2Kje/LlLImkVfnE1qsfgcsqkDAQCdfZWGJ7+Y01q3pLLRMNXS6DwlLaRo8YFnI
r0jD5Q9Ejx+uuMCNyhFuIcQus2pjB0nEOU5cl258ju/7Yb/J8cRlJXG9aJbLHRTCYnb2GY+DHiQY
764T7aQb0hM50t2r6PBZXH8Xa0/X30HMc2qpdFTISaok62FToJ40Xa8jGyCzTO0ZdUAwAaRNr202
fecNKkDYBZyJWBotguBAM0wkbbM2nyPDvdrlOIE2T9nRQBoef480wYeq3prmPqYBm+FeLrVz1xOJ
sDWwmOMF3ICZE8jfCGvFHkg+pHYV3uC75ezsT2IRrP5Ydf5hk2Et4x2yxIauu1VXeiMKFpsI+Rqn
mw0NwqwyA9msNSywIlR6gm7k95xaFL5GnmzXAK7BSOue+LNxy0Di5iwSdEWUH+jmHaGR262D9Rfj
PppNsUCDZjwJXUqUiJUGEOqmfIkNzfap8ly/9mgHRbg0j4gF4xNT5SKvqtjDConFRP/32SWp2/ze
TZInv3Nz6G8dEDicDdKZdna4FWmwQWbw3oYZ9tnrjATZ/LQsoHOWqKOoj5IwRQZ3VAdgSJSqhIRC
ORonMJNjZVk12gtW2LO53PQPE6kNm+DteYSVCJkZKwVTUQ4O7EBr/a88ITmcfI+cMPob/XKmHHBi
mUFxuOuTR4iR/eyZeRCPF/Kq3Ro8NbxqVRjth3Vvz/ZMfzDFZBo2NZCK9TKZNCQwKDi5rDgZzaM7
+jeP1tnENuby448cMI7PvwIbC5W6yztPwdiSIZiUBc3+4Yq6E4I6NQF7PaqdiEcCa/2PDIDdYdBZ
/NAxV7M8J5s8qGmSkO3QE8jvoXba1NdTAJNpbTJh7pw2qMewyZ99vpFf+KtWUeRlDWL7FxacW1+G
s0t3G4sA4BYGcRNN0xTK4gPCNh6FIhGSJoF9Cok8MQ91+SN3+rJVhTFHN9ozZd8CdQWVp/NqLjMV
ibF+fy1FUI+Ywyr50urI1ro4bBmkPFICNZeAS0+qQQDqx+80nk7554p8INBCQvfkyS6ycQ7crykW
Tr5laLZgJoAsJAOskKi21PRorSf5P2/vnvu7kZKfNz0XfBzhMKEq561C1YOVH4rws4P7X15itOU0
fgQufRnxHoFaXDOqw13kaU54+cov/dZr8lCczEvLPj5K9qjBgz4/0BR0aRjtFFN9+BcWP30VBb3c
NqGJb10AOm3WXMagPr2YjeasXB/VOW+vtf+/JSukOutOc8QJ/mFSl89E4rkQRnd9MdAdYewCOsTd
BMZyP8E0A7ITI5eSBzfsfCJp/Jc6NF7ECNbc3uy96DPQ1LY1t6IQcGt7Z2bIOTPRBkRPasDuBTjX
QXbzlOwMfkjMaqHlc+Cz9RYWJDTDY1uVORaKx3ChSZgICjxuhsv06gl+Bx/jtJC5cRJ6Xc8ysFtu
lowhAj7ayD+ii0h6w4I0bJUwI94EpDadnEgk9L3MUxmaAZHT0qe8PjIEGGnaVTDWznmeMO7P/ZeI
XwWV8vGRT1d+QAvipAKZf3C2lNAhRFgSpCxN+2uJRYhfJlk1Fy2gs6EULfzi9bbRPQ1l1OLd8XW9
vI+zeIa4uPiZMZb6q26g5S29VTrEo/FUlrhAHq68FfAhv4ZelKhmpDbHIV/8gKRL5d8+UdMtt0y9
NI8S4dYzYN3Eov9Hn7AnTcyfs5E4C9h7lT7hkyZl5ITCX8HhfSUtWfZdxE0slvy9GLSIPLz9D7NF
RnEq/qvnz09TvBAOG+R627RWgDCly1z+/eJDyacpoWF1XABXBDWrPmx61cmr0mEsKFHXuwbG1vW1
rgrK3qjPW4Vu3lLkBD8aEAsHWe5AHdmxv7uWkBCS21afBdxECNynx+TcLWsvim/xbboKbBB3zjKm
Dn79Kw8OJvoTWmJoMF/Jy0dd0hId9+eIwTycJHeHx16mo9LbxhsYnUYsM/IM0BQ49dqxrDO0Hm/a
sr05gYuqg0E7m/mHB9HIAdYUQps/pACmLai/RobktSxFG6fLRKK4BGdmI3sYiJdJVWIKzoLH69eH
0njiWK7ku/s3RmHtprfAWuSb2YOF0AR5fjBE1tUJtLo2Qx26K6Kps/YNTGTMAi7luNIvHPqASln0
r3MROMa38m5VQ1uvlRqkeNgYnnVKyp2Z6y8jX2rQ20WAFht7PoFpsaYQiruIKse3oXe3U1KqHyTN
xVihGSj++sS2Qf8efwmVNHPEBt7nwbxoM8WJdyzP0Pliv+xy4Rp3DRM7gNwQYLsFSAk+10SenLUZ
vCE992nR0+U0dl5zuEEBDtrFXcwg/QAFS+2nSD7z7HegcA3ewkxfctSZtOXIMi1/ahRlH9W562Wd
2GcbVpFW3RdrhPlZE2y0cvG/f5QVWACcUk0jvzMoK8MMPN7t1OTLMxbsQKq8SvRjSENXis4m0b5O
U0NjgQa+9jMSIX5IOZv/qJ+gWUq9PrVFgJP2TD1/8UQ2gITZSzlo272UtYBy3sAtiGv93Fa8IEPc
UQeF4L7pi1gMxqiocZLotyLCN2NNNEyrTkL/sfAOlS8gx7/NfIJ2q8iPlHFFpGIG4WL7mZJE/MKm
qE1QHyPaiSywdBdagSgpBHvgbVtptTWjRI92Y9RoIQJZz9TEuqVeJSu2DACF2fDYlan0W4pQ00vk
zuNUNSWz5BL/TsqjOcpxsXQRXluKjbhWFOU++idG4rm1tm6L5Ua+mMvFEu6VXan+SS0cpgrcd82p
78Oi7Je5QcOau2UeFpwOnG5I7I/6FtiULq0zgh1efs2mSn8VsqHRrBmygWzzSPcGYk22ue5Zw3Ll
QkSyLqgn7z6KYs63Dl0wBysbAD2fmkvMzqOngijvyPZ6eka+FFqhH7xNYh7uDZ6hJgUH4kFta3nC
+BaMpst9FQRr3b6ET9X8JYFkxMCGDiFGAP9WD6m/RbMXq/3JznlkhaATMb7H/8ScOX07wflxgwfe
UyQ72PSnBfY+2SRUVzzZLWlCxHMdxmnNL551BEVYPtcyVqizzzlYH8l2ztdIQ0TXrzVftPgZNde2
6hbgfenbm5BIXs2ay8L/nkoyfDgXa2QNTgL2nct/63X6HB83qbAkWC8PIvdXzI8nKxzXHMwxZy9t
FVWTH20MzIK/GeQRRhyCFdn31kH3su9lbGpwWb+K9jZMunS/1WmIUbsvqF5oXzyc3IAxXWwthT1j
a083eZTJOBSZ78Ki4nuBTIFV02BCTTen0iylHT+y9+N3bnYmdhK6vYwKtGd6DXWbEM/XStB5XPZB
GMADcvQZP3HrnIZw7FdSojXDI7ztPaYsj1RsShgNWRj77OX4XyTPyP/GInyNoLzYX+uENIb+YpMk
oukx5h/JW0RC77D/FoPmHXiFAAb36PZ1u/kt3PHbmcRVY/LCAwEEEEWdsszngJRzu2M5Aq3W688t
iUsLZFAgmYOgOv0USnP5GGDddA1xFgo42WKrhSJWP2n1kGJv8278tOQkAZdGwCZHSa/v/h30Iyaa
g0UwdS/H2h9IF5lW8pwLWiHzb7QLdSQZ46E+qGd1eYKNibl5Xhtf50g4KTXaPYnaCuc7aF+dDtP7
YreyP9rehwsw7uz5Am76fC3f16iakQZL0n+ckqWRL00N5haPOnYpqtX7xKFFYCMLbdR2NDdAb/W3
FXXTEEAJOp/e62x2HquON9DvAuw11+WKxmp228PEq4230G8OxLohZA0uIEML7JBCXXiTNFMrKoxj
ymu9MQpRlfW64Rz8XDwj/PGyNo9f9W8YGo/99U3OYXNWgVBv4vkfaAx9B9+B/FKRM9vvmg2Es4BE
F7BoSpQ/hkRbE1uk+im/UXg8IXIOf9NKoMUB0Hba4e+rJ3LwwpP3CGd6l9qBBd4CtD21FWkxiKiL
QFyhWQKhjMbEGSjxvRwUTr2CN1q0U2x3K1vL9xyXnzDCWXl9qGBbEazBCRJ4jYYdBkPkpAzf/PQY
rD9BzKEN7M/j2bYy9Vz90GhMz9UuIhQS/HE7f++hdlbpHrHQ7qFVDpGz/UrOUftWDKTI7s55QqiK
EW71K6ZFFI6AHBNuhmWJFtebBCfzHrhj2yxxiI+0C/wtmXUW2R6qqgqufsn0d8vWwQtpXILXrJj/
HPyMz3Z6NnRvjVKgsb0/2EIgKGibIH/W3Lj/W/cFOKG21nlJSaSq4QKBWqqMcK1b1VcZe/G0cNxz
l2D9WQonRvYGVAWXVK6znyo+X15WUdVk91WbxLElfx4emrzWq8QDk+B0AAUAqMgRp63kDaOUD3LP
fsiT7HuxfSU7hKZ6/NkrJ+40muw9hdi9y9oJgLiI4HzVPHxeD3VcEN8pCz67VSRTWcmIBywJNKmf
ljTu5zycCWpa32WAplbD1LUiLB2rOolmS7eNFGhRfpfIFewkBOvOwpxs9OFBVNVWA3Z1/h1r0BpQ
CQyM9voWl9fuqrRlGA1pQfkxF2erQo0QDIVXhdWcks780WhevLTqUT73CwtDyONd70eNK9yWRr/r
rapP2BjzqAfRdp8DOuXf6Ap4fMabVlPTWlj+eaOfIg5UYvxnNcrXKqq81t65FDgkEhuHP7QZHifG
lvLuVyriKRKecxy+dBoDVC2kUlqxu+KUKK89X0kN/nv0ZXagr5E8uei/X+veIkT6Ly9zQJWaxeVl
TCr80Ohc9FzK1sT+qTqsPsVNe5dbaRzNd6dd3QrWbuNkhLNs05nNF+kJw5h5EhZI/hN9pn6/tlWQ
P5W5LkGEWJmsyhSLpsTC5fHJA3q84niTtj+Zlt+n+9D3xC4ft4c9vV0G390YbA2Gepfi5Ej/WN+5
9iEOqgh9n4j/X8+Ox1sPhmbzXgsTaPYS9MdE+i/3fpmjeYjQ9wApeaABxJ3jYFtEH4Uu+4BOPZP/
KrZTq7SE05tfZtr4MEs0WscITzM79iA24SsfrAvJZUMfMDIEXhEx02pOoHonWhxQcbiO7j1+aHLA
v0spAWmDMAEiDX/pQgXp15gvSa4l7jzK5g1ZyzmkqYfZS9cqXRbKTaB9BCOa3aXlqcXC9awE66Bp
NKqwi6Rji4cUuIg/lZd/hJt9wniqo6EmxOwkIlUksLps2EVwv/6Z6x9fdjW2KO0l3QiaawYJmuCG
CupFYhYohHhLhngeT+ba3O+aOwszTcyPIHZ8cF52y6jXTtzh1DcvWNoMrH4fzDLayHG6KG/Xe/g2
Jsf6uoVil27DyFOVa4l/d571kEStoax7BlEBJlnxRheQ/uMN11EFRfYGYpm9m+2TBAfNDRzZeBHG
epEKxPs6uT/zapy8pNLyGq1+cBUrriBbjIkwzVGwfwqC3uK7hRWEKD7tBo0X4pKay7hAWWDUPEkx
Hd68LoJSJ8783MEcJP/vA80hmZh0/OE3LIuV3/KIuk4VnH4P6/fMY7jfx0UPXZyZMgNBFHj6woOh
LG2VHQoZubShJ4GUfeiqHcV2V3Gj+XOPgFeDrrjxfJTd4m9Tv5kA1+dd1GeAkEaLC04FMK4Fs0VE
FmuBMdqHLrhFwB7X1hVqtrUbkpVyEcqizDV2wxwYn7kle423SWzsGyLubWLRQvr+LlMmU+Zh6xoV
6GZyx1ZYTQChaHW7nC23FXishq5yuSS8jLPLOzBaim6w/rb50RUfZRNsq0zQA1E52yETyLvjSCmd
1lDtFHryQ5PeJhKS2/8c9aGtCMSICGkqqWMnk8AwVIivBaoDQs4bfNRxre6M1R6KsIciENBXFX24
eF8PYohtBzfJ/ONY0+hNPyMYTMCqk9+uU1nwQzrMnMtX3ucyVnMg4QdeWTRCjRNHD+7Bm/Fjts9u
X6h0A+gr6yNDO21CWeg50Z/Wt1ykQFc0tLGhB3kd4VY1owMi7xFgOiaQ8at1Ejc428kC+p/Tgk23
eZ7z8buipq2/5ub/ZCL2gegRzSHmCEIV8RcJEMNW5BYR+1OX/zlLWUSkNaZHnb967eIr4ka7nytA
TGA/Xya99+jZt4AYupPHRSyFwS+QnPABcD/PlgWH0y7xzCAf9SthDfgvqZekUU+rV+7rCOXCi65i
PLu00ykUlG+wNWCh2bWRSXvh5Ec7AQ7iP4Do4+tFz75kMLiYF85sXm2EC6MKjv2RZnSul2I+b8/2
l4u8wTP5O+K8Bgf+60hPqgIQ+Y6LdxydlYLo3ucm/RB1D14inGXJqhtSNy0Ony+EEajpQXof8/BT
YkkdvtfY3d0wJ219ro7RR3readfugFBrS0MTPvrikqUJppmgkS94WnJ2ULNwpfI2CfcG4ZzeMtwx
kun4QAn9FxK1hKrRPElOGojHD9wVKXt7xDyF7yvvIufLbar0BjzO7iCAMWEScwpSJf3fiiQ5Sayr
wzw00BXnhYnD3fhGg6gpWJLjdG8f4pKi5v4eYqYhOQEeW9TXUcsbuXg4Po4tsfT3dbHWzPKqo/SG
s8soa3KALivo2hxwaG9U7exHQu0M+4EfM3dmxghyJEjTbFubVOKlFW0V9OgItQgah1ZivtPUUVYm
CGuCi/pENCUIu7mjPTza9Bh75RKrBm5G1HzxPEy8gHXJaI8FlvGkLaZw5elz0DIfqOAuaiZcmdLU
7XxfmGdK2Jv70GyfFkOI171kKDX8I2NjCh3LyKJadx0Pg/grw6gMTNXxOeyLiq8NZMkaGJe2IVXE
5jwZt1YUZXqUxVXyFhhSN+0iqp34IlFsmZ4e965MTViEoZzLo8k/o+qUzLaqtae4VM/zddvmB/+E
B85a7rTgdV715Z276uwxftwDpX16VLO/vIj/bHRJw9UGpsEAuFWw8Y4ixVgYAo0mL7qsM84ZI30q
JPZnM1N1GCbDuCgglOB7y/PRiFBScOYZvZh5L00LmvAdZWoIpVYrcWs9iY0+ld+JT5O2Eyth8vK2
I8aS2O3iAxb/2BqVGo98fvTt4RaYKoXwMkyDEbXyFevpM4tPpt6yt5IeYgPSxKnfSDyvavUZU4l0
Bxe96vg9LT4xglQZKD4XDfuvCopO5GWip+Yv5Vd2xZwYBS/00iSFGDpxyJ1UyCBMgrguPkUZS6up
B56YWL7aofHS/5BM0xSADmR77zCPA5pqHwduGD/EwMU6xkjp+BCzQkZbNLAi6csJemfPNOn5KfMV
5g8lKdUShYwqrKJZlXwPBSTaI+ZDR78/HEN7Kcis/o4pklaMCl4H6bopwf9W37NTdIlQw2i1ruTI
Vzy2SOLh593X0yHSeFk7xEDmBhEWv1v4PmsoNWR6SbLWOPv8KvxN/oXEEiqHqxwJDJg7PbNz5Ay0
B2VtVupQfICJhDv1IS3hgl2j7sA6iq6KA9fWFZIl3/cMJIv6LG6PTtqq9TXFs6CX2/euM6VRJ/tv
5BTmNk5dc8+oVFaLI9iVob670Kcrgj/AlORJMR+HlGTnXZsxc9m6GiTk9t/IZxgODIX3W6REcInu
bHGwmpjqcN51+m4YOIuVKfSDmhnc3dt174KKlrR1TZ8KbSMwGQqs1ho/EnrfHz08mabtot4kt+oC
kRSZRjYmBDU2x9ZaV24YFr+JnEKqqWmjrE4cEzBrRGY5ozAvNz+WBD9kjUE9aqUq4N4hI4a6xtEc
dqEjwZm4xt2JsAtZVNjQ7x3l0bLl6qm6WV0gq2GSWOq5e90U2NuEKKHz52v4lai5gmi915v2JS9G
t/Jvg9XpDWOo5mYk0yvmSZyttnC4uBOyu+g2zHBUVvVbg7m0J7JaPiJm0+BHs4XmE6SHEtftsj+U
yZc1x6HNCydoRoV2ZGuuf7rG87r+3lE6RjhAmzipv/Ev71xBoEkNP6wROXg9C0wEQCcErczYYXBE
XOi4i3UiVCRsRb7nWygZsIRVA0Eujphe3Xd68wopMpTCuXLeB+dhYepkbUqiRIJMdf1rG/gIK0oe
I0qP3KIaubNQOqrLcaCxpRSTsIG2cr+sXA29UyA7F1lOwo5QAy7eICVxEJ3evu1fIeVPaHICgqRY
CjAfJDf2rOsalry4PoHU91uaizM4x+kiUs4Rjk59JiKG5xkx/tpvtVSTArexO/Z7EFDqKWNvNli/
SkX0hBN5CSHB39q6Sed+TIJLy5Lyh8+29vGuN9e+466pkRPl/0pt4QRmYCYrlZpNRx5DV9Ec7TM7
2QnVplEDoPfSmYcHvxhS+aMcJ39vsm60u1FVIqukhXyLa8n+YoAPi9iyK40oa59GvV0AyzipbptL
7eJCpRIG/E4q5cImes19SAmjV+GL6bao5MPD3TA1oUL3Shk4mB8+xydqKVzQ29IaYSdGEo+nO5vH
T4oOjSZx4ZvrGzGh0v9Hhcx3L+bRI1aqXsP71Na+erVRe8NKtahS8PgwX34gjLQ9w0kYeapOL/nk
4mC4yMpqlM9eiR1GOpPFWpmyTwugLNAcVXQ9O+77FAaD5WuhezbcOxvzUmROOCfkBAUE0czbJvUO
9kgJExX9Y9VgjqCmXk+wF7Fis0mmrayDZ5dKOE/SMxx/CAbxbqFfQWXiIs6DL2++IMWfZXqHhpQK
NOeDH87pja0RrMge1RD+5K6nujvucXwdPvHFMlgn+TZFkwc3aqXxZJo0nJ00qv0YWqGjDbt8ith3
0Hm9zKcPEw3cnQ06IacITrDkD34Buq1LDgYlHPN6/O0Cj1dPzlWQzrvDix8VDV2jOrxO4dObD6j7
GFM5g+xLW3UANwcy/ZVJDv5Eht4u/zcaW+bqDrDmbCwCgZ4MQkvUdfPbD2W5Ni4Tgpd+TrMDWemh
byp07SIhzsFJyfgT/QFct73FvqL5Cj3Q/fCkKh8ZFn/knB1BlXYSWu01/P9LfWJoR4R7xYk6mAYV
FxSqImS61GjH7KuTf78Icsgoeg7Yqd1E1HQpF9M2OtPzhLqXiNPpmsji7yFMd/rIOl7DD1f51CmN
wwVBEvs1OeN5BwKiju0mV5dB6wnGp7ZN9heP2/YDNPoauiWq5xzsFUq6u5qVFsqN4iHQITIyqMyC
5qZUR+xF7P4YukPoUYGswhfP+61GswoUViRtW/++QwwVINLqhHrp3g4YsC2T3URyXvK9Ov9fj7x9
7BBqurFLzVhJp+aJn5TehtqypHH5gH0tZQ+l3GCdZj8iDdDlmPnzPHmvFeA/7v4kDCvTfyOaWL9m
QAxCrppTEMpr4OTkGviq3Icicyei8+j3oIQg2olCuM8MIykR5jIjaIGtU3XpnkjbwikIb9rdt+j6
D1W4UqRXHGY+WETPb/zMmxUZcVEVu15qH9wcnin1XarQCra75g0V0NQNm4aH0ztgRElg51bYZzJs
sv9Hv9CxNnXir2JweaLUUytsx8dCaI6e5a6dSFruJNR7aXzASJ3pNVF5KOGmRu3DzP/cqlZTk7tC
O7YV5CsxvH4rNS5j1EWBF8O3sgMvqoIFtxvt+jzseZ2BsdzZV8RtiIklV8smiiKRjHUBAOUqHxYi
dck7c71HxlxtWbrDhaHPP8VsECBAUCYkwmweCBadAcvK1VtsSU6VyZcyVO+Hm8gqCHwGmWckawAL
ZQewpad3ikAzpyvOZWKAJuLxglo9qyG6SdEm/7MQpqqDS0rI3m+kuu+iMZXuvSLDFpu6QrBTESWY
cejo5rFM/HtWNEHUChA7TyQLwV6l+pGR3eSJTkU0GtAj1+HDGoFqa1tbqaVyURl8lscw/3ichtBd
fKGfpXeRyb5wu9H2UyxhADMI3pKuMDxX+Pl+gljeNk3Cws6eobjEKyWWIB3D8xcxVXK29ZhZjX9x
l+v7VXYCqL2phKCN85fn4q6zIFfgP+qfDaO6QJfql9lJIG7rFAXTTWeVK7emK8bgFSYfqTrw4V1l
8Gu/hi9SBVZ8wslEPihmcqd2fjhr/0p3FlhJ1cCV6g12bET2hqBoyH60TpxQheTrIL8BuYRIbNkL
ndgHRqE5C09JOvH0YJzuzEd2jDsisCL422KlOWQ3/EpXZiZV1iHV6cFqTCgVWf08gDi+7G7qM99B
O5DKx4RVjrmOKxlJdjHqIFh2pkl0+KVrVuBWDU8+JKWPs1ORAxzKsEQH6icOoUunQhXfS5pb46kJ
eZd8pENdiO1jYM0j6Cd0oKMB3QQYSFyUOxriLiekaEejCb92Hc5fQnA2/kSesrkCnJEcQSUksjGU
u99LDCaBBByj8R8h56IWIeZ0Gi/UVpzgASj55AXTms1uBVnTiIhqa/A2Y5YAeoGRPbJhe0FzaNtH
WsU7uUYHHNN5tLLiGbKfHb7fxL8Ssk/1VTDg6UbrcY+VBG8u4bbO/H4Wvc+GsFfzZWGo1rYZe6w7
pDhDKIf8WKYQFYX/0o3f8GmbLimOZasXgcYx8W/fbyNcmJsgGYR8OKmaer2v4yu1YnmLuSyQYxvn
wWSKy0bhyKTPXKgd4OHgmR4O9qDquUOka1isFa5H4OloelUvr7Kgh6sJl+2YfY+iOBzFPPriwdCz
VlCVIJcS/UiY6L0YviRKJ8CcCveWX3eeR1mxkeVQhLm0OuRVZUvXLAwIoisHh3rd3RzgAHQ5B71S
N8Aa4jgvHj/wDEL+dA8OW+OUDEDgYVa0M+/IKh/Bi/O1UEaSvN7k2JtN7F79drZJ0zXfKV2nz0Ff
MNqWu2SD8c9GZJ6e+6S2q76xUQezW+YofcUCdzxtBisH4C1symxd0qeWrs9Sj7bnsKQvQpnf70pL
gmpxeG7IjapHrwdnQ+5KNgRS9E/pivwRjF0dSe+1dWiTEPaXKAnjz6JiWM2pL38/6FjMWByM/Bwz
P9QWxbn9sVtDfELUWY1miGI7mrulD83DcRkS/ReHM3GyaEsaGXcmu8bMYZBDqS1xAiG9XVnHH2Ve
vQv7FD6UmO4t/VC+me7qxHrNuotP1RbMDST8fxgimV3S2wpQXRo9lKtAiJtvdlWagNchDAvuJD42
+AG8FxeZe1ndAXFah5PS9sc1X2ag5+V1eYoWfh2OV7hAyDon3jRu8f5TGKCqKEldJnlzVvlO5JsW
zHhR3YkWZikEeH6kJJ8lrynhxmbuSOT0h4E3PxzYyHhdpLrtfi8LbzMppQoQ6WYVLVKMCPT0BHz0
q2ESZZceDUkx+rvmNejA0jYAhcfhPTnPcTUqkUUBjic9PPAqWA0WNGzEDoIdkprZe83+S7FPrqek
XfnDAjTUWiQJ84nFa6YNy6i6nUxQmwge8aJX76lk/T9wApBSuvlrGpJVbpL0iLx2ROXaSi4Mo7qK
rFzV7T+Agui7qLpmz4JDyRClkQjA1sUZALUx1Fw6Ewbltfdk5AkzRvfsbwKqxeuJJNtPposeNhm6
j16rIM3AgKGUOFcjIYXDtDc1FT5qXim/pF25sFBo9MMHGS2wq0/wcmaqpk/ZtFHXM0QjPVT3D1Di
t4Z8FX00bhq0+7KH80df7R6+hEHHGn2+vOJumaxqdwFOWF7Pnnll3dA/c81hnuAjnV77BMrIrqp8
kyLCIdfKd7jFXqwU7v/5XRdAV6mtQHJW45Y0ouQFQYfNiJp6S+5/iHST828PJIyKC+n9E8zNp1jI
9MnduR0+35ehyPX2eAyI4JOVmulgk/G9Fh1SUha9YiMNkOnEaTx1e5hhCwLGceAVF53vROzJke2x
cB/B/yN4937nrrC9jJpMEax0vQiZGmbvIzC6JMHL5qrurnDBUbFNcscEHfvLfQB5D1NYCRAc3qb0
ClhQn04uRMSuh8gWeqOXvyrM2rLMYWWLDE/lxORS8IuGH6C1dc7ML1Whp2VHzOLhybZ3LWzvWxJi
PHcL8lumH+2QxTQ1MxUlN2elAO+q10qj0j5fqslnGV2dccmXDHpIQjd+M2NdyFDhwdj+W/GnWt47
AD5gm02524SvUkpggxcfWRRLqAqZtmvgF07SWV3IBu3VAHFI2grMLHjaB0TCYbPZovVnAOMgVm96
7RjU4UdfhwWWsqKvwNANp1vhl+Ki7zgtWbXMfx5uq0N04G+ZnSE9s++wMKRPeHpVpgkRNjKNZg90
MYvMAXepr+Gy2g2bad9OIB0EUhdca8qyXh3xWmBS/urLZro7f3rf2hyMdoLuDOOvHkO1vwWMjCzK
oTlG9iDjzRds9rPRzX3/kMmldePOuuxfhSYygHPXzhGhwEJ1v8pycyCXxbN9Ux7iNBBUfnBBvQfl
tdK0wAIAQypkMCMNwn991UljWoTq8mWXmexZiFwKdLbXZp/fH1ohtIF0GBiPXPk3CERDaywxjGZI
r4i0Ch6QcHIKEpN8E7ehVomg07UlfCelSgfhthQntMpi8S0+2UhIplajgKC3VIYPREO5HVHtBGh7
S0h+ZJcuS3b1jdtGxr1uJhxYP4ep4FaqfRbSU2+VXACToQqte07/71XCU8FmagYqhl8DTyvNUBQa
F2U3D4BiieqQ8dZtLWIDoUf8SGaWqrnJ+jYXiLa7FqJMewE1+yVWu0RuLH+5WfxB9wN8K15w+Tun
W20z16EY9aoqWTB3HKPNU85a8RFq1vgYSOoLWYKFafOgjvJbe8kjwNQvL+teNcC7jgVWCc2ykc+j
R/KIBryvgqcRvVqODyhw3EI6BJzQl50l2S3oMNUig4RJRCEA+3LJlD1uaG5X6P4x3hA04Zaaq5vw
xthss/BaxlnE8Y3XJOEj2t2Jd1lsDseKN0jnVMZ9Qrt7jRFUMXJh2hBsHEMQZBtFlO0EEaiUiCES
pwCyhK/N4SLzZZu/JGszd2MWAHponopwnmZeiB+VGSliQOMHkkHKK1xRIXOPCkfUonKm+485eUqa
WgsaUFLYlpqNqM9h0sVA1JPaAFXaIq50Mgz7wBvX+E5mE/tmXuHiVcZNUPMxEdrojXVHPnSS4UxW
2yU5IRXZZeG/+JQN9/EDPQpUvGZmO66schmZ7gKLesuGcUXw+FbhCUJAnfbCzfY6fRTAyNsaSTi4
fZc3bHsx2RiT4Nuqub9bFoix5LpWCeTPWXueGEduW2T3+nxi1siAt0MKcPgC+xBfuu57t3sXGw8K
wx4WQ8QgH9Amg1PmtVo7BcVrkL4Cf+XM96DnJMeir+u42guTQh2fGcXHTzjQ6tRd5Bnfw9KIy+w+
p2PY0I0/AnDuLYMjYFIR3HGrJ1edVBRcImqujYI0JiXGuvFGGtQn5F/Bnd/whDqLemo+8gM/GNv3
LVto/VHYA7rPrEel8zSM0PhGVj4iEJCB2qBF5oJXSxnbMeliqPUD5wizYd6f5wI9d/RvgZWRMszF
ABX09+XimBkYmHdbcE34Q3hn9bCuHqW0T7G7WaDHKmfPFDlON1GL3Om0NNNBJsWNatShglIxa+w1
4pJDcmcEnJb2U/E2Bwli3ie+vCrcpYaNMH9s4YXUYdBUGH+myg8vFA+7+ptPkDlDheFRQUN/C3li
Ss6WCCJPsCcP7cCnVtfXigZI7+TohI0Qx7LyIFs/qAUp8xX4BHvismrVaTD9wRsmH1s7WsnfjLke
OQFG2XZMyRU+rB86eTkT67QpOgn/YrNNZ+h2JpfEac3j5c6YrAsA8zDWDVgV+WE7Ja5v45u8b8x6
r8/zgHYBLOYCErnOvGFyrUKmfrovw/6R0XQiQjIxHZkDXnzcFbAjF/WNcbTK4GzI/jXo3sJTUwlD
q8CBW/k5FSf0+kXFwTviGLKK4Pt1mvdN4UX0aAf6gFwXhy4qQhrpmUZEjF6tYrlsK1RTAq3zJYPC
94cb84PJ7erPBUuGKd2jeW67ymmQ+oeqsQXTILsHgilxz95Im3sCqASX8ZB9tMdltaMr+/QAsofL
i39G60pr99bHHI/JejRRi1mHUgXjJ+FlRZjxOI8lSTdrFUvCOLadYrrnl1lrWqNTOeIzHOmFraAb
3XOaHWmglhtkG3/FWwZ1XyQCvyDhOkX58PtrRf5gs+1U3teF0jtGiaa5nsB37/UxE4q05h8uS+UX
0MrAdUH2vgN32l/WDJcy1X09SPQ+5dHhDuNlJy1uCuc19v+/69NJn4CiGbCJC7GlFNjkijRcW4fQ
HbrfW8+F9BKs/3Pd007vGQlicnyt4eSm/GNcmn9qSLzLZc2bZIJXmLo94L2McdNagBUB8u2FJTqN
RsRrhxoDFUbPtf+SDUfHNQCTfgV5wU2IlzWIf6laXA4z3cFdis4WRq0pq0A2vLVBdkLp+qiJfg7e
xO6j5r97t24E91Ar42raAfvoj7GP7GLhUUZKdgtGqE9CzEfk2Y/1aHg3GG4zQwZ9VwVULccKKebT
4iRV6r9iye8oG7bNu/AKbbD+npyQMo62mSFEFBDGkIcAnpbU1rD0wQ5vDQrBEuyhH1+Z/b/tqfXv
Ov8Q1mFLYsTwULoQSyT9MMCorUUxBMl40Ai6qQegkc51f76Ni3zOLs6PIzLqGN7T3PxgpL2y0e9b
8JD2vXH3s2nEV6WLvLt3p02/0DrL987mZYo4UkJZxG16sTuS1kbZnBhVa8HLYBhXhMnio9gdaI8Q
mPHsJiQj0QxvrUR0mmEKEflN//SntF/6UO2ZFgiqOIFcAAS/d7fCpzDXQ2k3JDMa+EirPKitCr/M
zUkIh4Ezm3eTWjNQV7QaIl+yGEA0sv7U67n/BgvSM1RT/bUJcqbwftJwDMlhrpd31Y0XufKLNgIv
3ft5FxKzJzk3JtEYVBvumRYdUocGo1ud2fC1zrAw5IPZXk0Fbnq2jWBdSZPFZJrtmGsy3GnTnuQI
VV0kYbEqzSUxlrxcpSz8tsKZxsK5MrU9oK2KWGi6npUfvHWLPp4swmLDQWhDt6QT+rczyG1QX5BC
ENkWj7eytAPVjtvUTl7SrGsH5vzouiJX51+hTLZK6bILZvPcQuZHS9nI76GmTJ3sBFd1s2tl+lNj
cAo80Sui4U00aJyhfVO4jymI+6TF3qQ0b+IYq9zboV/nIh346uNcmh/gpCJ+PVwO8I+Zgs6AcxoH
LN3r9qZOW+Cx2Pfw7xQhFsmLzqKkKgKxfjOqf9SBIR9xNqppNxpCD8Emd7LB4IGdIiT1uzlIs0s9
t2GKBorfZ7iCs8Ah2x6zv4zt04BjzdoMqGKxfEVIBXRXhTU/CE6fsiAXL78A1BfTgnNEkjwV/OyB
xScBtMyN6BrTfyOvNVN+oJhZ+xm0+ve69w520CcIv7wZPY7IzN2IDeEOyw+/rTuqbe7XICjLUkm0
u23mlMIF4SKQoidvzjMpewZOPJLkWl+pzp/livnYF0e6CFzwb2vqK/mYn+IdrmrSRIslTYvmW3Ln
pZ0Lt+S7TOjZoH0tvTVewCufzu/6OlAMlJZw+QlHp/0sgSN8c1VzhFtl4+jGqGgABivreq0E5CCY
lJKt1TJ/R8bvlZMI7OmqtGVA7GrXXDerqi4NClmglwkDY8lL12qrPCKA/FvXzYCtwWZQatXT2zlQ
hzMLD8JmoYW3Qyfgp3MqCZFqb44mkAFRRb71Y5sWmbvcAFBteKaZJR8Vqmt8RgrhYyJ7yg6cHeKN
IYtz+ifViocdUOS4MRSEo/C2o8Hkc0hSdrvLGcczUZS2LgUFOp+vmaaD20+rh5+60oheaIITtGeI
t8NjtyTWA7UYR5gYn7iXMX9KhmvMAyBjfoFaRnzCUw8BVtoEIFQGZqNqQ1psFWlhJQHweSH1eRLV
7FQnToaDY1J4XAZJOGnoiJhkfFcvh5+1s91gyZPtRjiyGl7x9qzNoqE2rCObYJxRdAqm33KMlVv+
eagz5yUMSKbwHElrjsn/wgl1gLrB6CPO1aJcZu4sg9M836BbBLqcd0qKpQpLKelZ6V93RusEpUTT
nUbhZd2RVTsBR9ld0/nxp5+fvqDddD5znPHuYszZnl5HoBtzCe24emSVvFYA/iLuE5tYvJSoY4H5
Z1V/UIotvDYXfoy/DEuF73Q4aLqmMRvvNiFsrk3Gdv1ThCOZBj0gPHlzz6UKGGojcLEgcQ7PwkJn
RsVujU1ILblvrTtm9kyyxKSZ1/y54R56VNcwDVbaloZG0wusxWgNmuvtwV3dOkq/7VWyXfnTavHW
NaHa4EEHMBAMet3sKLnsAT6eTAAA1V/8x+jftJ5kL3a+j9g2x+ueq9jwKze1E6ODyAgeislkaf1Q
JLgSP/GXIy+4SPON6FbhAjjpRKxIH54EDI00nBRgQ+tIvz1J9pYAS5SRDHpc607z9CaBNkHsk9kq
KRbmTlGruPgDGjTYJ1S3yzOVHayUDIGwOxDeve9DuSXVPEfT6X+YTMRZmgsCcAGTIV8w04rzGUXa
yTtxIalKG90T903OtDTY2S4fqXybXZ8CJY21Bhym3ukCtR1xcHLenmAENxiqC3DicfU79CRXcQRd
hb0Z8i7WrNHknJMKdmEbKssoRrc995acCjXavMCT2OgHIKNUbJNZMyHxJXc5Q7110fGRsUIhJVOZ
8jfZCac54o4gcOcEwJkoaiIKGC81IMLmZ7aPxhMM81+TyItGwrUG5gYTnw8/VrETPHzUIsKJ+8TY
5HtF/V6ArJ84wrtYMtd2bxWtcdgtI99xajrK6VvwOMktD+SW4ub9DzkwJ6CYw+Sqw2/hNXVUh6DW
ceUMIbNJHP4J5c1dAldSeMaR8NoQ1EhCUfqEQfTzy9gICa6+xa3xZNYnsaN8/+UO9A4kLPOz8+ea
2xWtlcd8qvm9whV3WlcfbQ1/Zk4XZEBxABZXWtjfpIZWrIjkStPJFrzqDOIU5MxQTV8+dg6+SdMT
rVdDiu4QznvqSRL9nSZy94pBIt4mqQEMx85AbmF+ZbyZjs4B9Dk2uvdO0XaYw9t4GKoqk82P/0mH
bU+a9Gmlk8xA9pZQBbCdJ8asBMJ6xaMlTZGCB9xnwje07GKUYeHYsilVeB9KlomEwwGDsbDPF7Ga
f1lrmwKewWqDm0lamQHnt7T0vQBc3cVoBc2Ckpb6poMzdSeAdhkpdTk9624+x7hzmq52oQ4BwcL0
XEc9iF0PkDHVYiLOTReKlOM5yLfYyNtQQc/W8wG/4qoVBR0QrAlka7g5siPkaMvR1KyobyVem5W/
8Y4nqtVnxYqQJKKUhXaFGVrerAgtFvvV4RXoGdcZarbXDvgRisNnV3XIafZUKJggCNh+9aPDOaTq
Y2wDkEAgdrvOwCLzjESNDQFSr+RiCeqdF6+9i6KO7N4e7QPEKBVJLi4x8SLiHRW2/XMWQFXu7Ajx
9lvJadee3C0SoH7MRGA2utSw81cV5olQGsbSIIllZEd9svwNOeZsEdGb8qcsd7y791D2eXX83vnE
ZNf6I+IG13SUfoV0T+t9g+khRgzBdk3ei01lzUcVz5qQ79ZgKRRk7kwePVYHOTshr2zl1dCAtZo4
bvAMzeephrpVitCu4nJXSFFaocTm6Q5GfdVGv5ljWrg0I21QYfjBvXzaSFSgYY46jBn15Mmsk9o8
QCbVJ3q+wrQETXkVuaHPc88VUJ8rNLRHmJ2haHjMFPfCdwmuYSQi1nFLLHZUdvkZvNqQKiHZXhrT
XbqrRHEFkdkaf1ndP5s06qm8uAw2GcmEeeDlotf3I74nEDpElD+24Ukbng30LdZOR3sXWz/VRccz
jNYUM2vj29uiEkoL91fKKS06XBXInRYfRprfScTcPK+KUnn/JJ/j9n6oFW7ouBFJ/nbohuvKjWfJ
AP8AWWOcIoqUW8F6PiSHI3NeKWWJQArHvqBb1q8QgLl0kUh5pRW9Rh6QJJJIVuHdoLCUc9EHUOQ8
/NaddqgBBpk5mHsE1h4ompMG3JuzNSwEeSAkvZCcRddh5pUY6TxEfWojpQdCyFv5knC8jiW9huas
8fLJDO0y+IB08FAXmFg5nAfcJ4Ed46+jS8ulrFWK6dshwrc+SmnCK8oVToB1TPh/KyEnSLtDTLpo
20uLZXsW9DIE+w0BIpVbvLGh3XwS1QV+Gk8P5imrtZn8cedIa/XosiG1zkyqsrYFpYtphRm7ZduN
eo+7/0di4SR6d+a+OdpIwAquUl60SYrThjwvP9M1phExyFN3QiQzkuniGE3vrlfM5fK01ugND+mN
vDX4DSSNE9bgprbUJ30zzQFfKIxDQ8sOh5humQOURdb6iy6Gt8GiXAhoRRGxV/Fz0PXIjZpMHv9M
gYhESvelrkj+nDnC+y3eDHZaqm5/FTg0KK8y9M/G0hDWIa9/nG0A+q6yKewEl01wjN0hjD9bZPbl
qV0GtU9aWX3tQ7uFe0rc/Jk04dc7trcM62oZLvorY60ZM7KiAAzDTMu44ZKR8Z8gUcAelgylNH5j
F//tAfiYWWC/5fz0R+WOs7zDkwEJ/nMFooXIECQ43IbAyRhd8M9cfOLCht6bEz1SpOJu7D1mhPxL
B+m8U3oYh2M/scvUpZWKCEQi/+M1FVsfM0mKWNu1cLZYWzlynN6ngV/UPeHgH7iPsTmJE1XU7Yq5
AEBKCLcv7CVbfSmk08KCBozxSGQ0SHVSj2hEsCtvbfPWIY7u+LgtdwPgBVeN0n8YGuGv/0wjwSy4
bOpyE7cWHtUj8nXwaBgNOJ483Y/bEvF2OZGMTW/ucYJVMmxWukc6kbbYaFV/Ciz5IOMXOeAsR4nr
kndseRBJc1Y8rTPl2W13dWN/7Q3xnAnAFS7bvNMC/221/pjm+TmbomvnE3hSFLNOdgGV7LXWYiJt
QCCDqXRzGufkql9JePJ15tPc+tSaaO16wrlchPNz3wE1nU7ECsJytC2ARWacUGU4t2kS6kK8TpBb
W8Fpkiyl1UaKZddLmpFnHe38ANA1KdDnFxH82w4waVhoOdLuxkDVycTFGzIgfbHGxkRAqTSN88y0
ztNK4Bnzpx1BECr6dvBjsRTd9byTb5+UlsgcUEskmz5ru3rX3JOirfmdyQxRKiBwNC25PzQPR+nO
4H8cl1TGSyF1tnQvnf4god/iNagmF7hcT3N3zBM1SGZt+JD39xWz9a42oFDV5SJvCHSv1GdgyP9n
zXDH04y9Bbs4HgB0OJYvTkRtRRwJgL/jptKutk3HkS4HTswsQJK4b8J+bdqoDuDfvdnGj1WmNdEA
j7XgoT5E1Bx2yKnCX2SCPTh3dLOrYCh+98lqKFrPYGcA44w/DrK4Uyq/Bzpt2mGab/uhJ2biM7PM
dLtYY5Q8n4WqYbqQgsZ2S1TIA1ziXpJO9fwoGX11Ap1u3gUIDYt9wtT8h52eMEr4uh2UyyFVSr/B
fEE8rIMcL0ZJ22+jnWoRxPcIGG9TzhC6z3duoOC2NZNcxqmiDrs/163OkCDH9YWo/4SuEe4Yl95U
V7puU0FyzI3M9TBNKYmWMUp1bgOssJuX/Qswhf3pSyRwvfGgaBCG4pV7b4Sa6nEKOHW6FFA5hDww
qlgC2FDQcJJT0/K/TJqjjHnqSwFa33mN4mdwjww5qIIbpp+1cYSVznqiNbkEDfFa4b6RY0MUUJEA
EArSsvgFLXvtjI7XMmxfQBaQkB7b485YqgxpeUg4QHWtYYG5QSML9wONCmDV0ewQgcnKQq5q1M6f
ODbUgB4/a5FHfkv8djU8viw3vozDy1poWhScmHnxVF9WfukJa0ItPGJokkO9Y3QlHUTHfrv2LDVL
MwDAnR8QT/8k07g3dfO37zElh5x7Qj/b0XqUjlJX7uTEbTG3hzFKuhvPW8cErOCllmXdZXnX64/E
5DEz/FZjd12+PHZnT1NpdYFE+k2WBcLLXlqNipvcIbRfqK/pPueBzTSvfLeWFyEXsduA7px1Kawo
r/QN3j6s4SRSHDh55S/0Xpt4Mpw6Q7VVqDq7FD8h0QwwKMi0v9poBJWZKwDbN3AjNFu6T++D63Lr
LPpNQn+y/SnqmrrgrEXQPLcgIs+fEMqKuFtlMQ20YBTk1dwnh+ZX1WZq1PKCdU2ydz+t49x6Gft6
osKfi9wqjwfxkwJhR8YOxd+aIBD7uNq+bE3E7PpIX03MKKuyGQRE07JjXedtS2Xz1rXtaT47KMYG
P0oxVuU5d41ZkhNBwaypZGpugk48yKs3Z/6+4NO0U1FKoWLZ8IS4pozGro74M1HQdHnI31hM8B0h
b0xKqFq6PlxboarVxKeuDlYqhQqEoBIfFBKh/hhxLN4Zk15n1bGJyRIY2lW+TL9OgXu3xHJMjYWJ
Ghn+loJ2mMoK/GhoH1KqNntvwxGma74pbZbrABAGPkooaN132aofrsAH7n2Fx+s/5L76+mzIiV0i
95G3edof+bOWq172vDpwOHX2T0p+a4cMGBmwiVB1Ho9VspcAsch3sTWpm8DD0rg3fozzeX1rx7Qx
uQuDr3JNjSJLQ7X0xq4gXQGoUsfTna5O2m/0ewmKPopiWvIGMvZVrqcpYQyEEGZiBVANMqGz8Pmt
mHdZccGBjqKvzf0iRLmnRycWVw9j4DMrCwtfuJGoTF0g8GpiS4FLapJpaZCUslATlL5VeES6M13g
bQP5NYk/ABOiDKT4vYLjSHx8ZIbIahrhi58Iogb73NFfuZMJTISdEnbxQsLfzRfdGCCveiF7tILx
wphInVy7U8CQ9VSsqf4dJV+QeIrCGVcaap/WbtBNa8Nz/8jS9769gapGGoBp075/cmXfm4UWZzHM
+t43nkYoY2Aai8lLQfSbYS0HnkI5kirzm4fHo1FbJTaY2xYPPTo1LchxmOq3aD19GYbTlRjl2cac
5+FDLTi9T0wZedQPm+GLgXLjLGQ0mb+tX0sfEtgV1IAkEr/iIvVfv7POiNsbFb8rrdC41bBhrtE9
OXQChLv/oVhRALLPbPIhjkEBgCnjpJgv1IeUSeie3F4whtv1/opmSvjMUS4C8zI7GGmHvZXeGycq
iES+lVvcvPS51kVFvnWSqjbaEJcyCwimBGfOKZP7847KEnb8nw5K4ZnNCq0rz0StBZ4QiZB6sGGO
zSFJ2OE8zb7K3kOF2wdyWm9Ww641z1hG/esKT2fB5rMaO/ffc66E3luod+R4h4mChgd9KgPV98I4
ldT5mMO2CGlkyOioOfIuKGJD4+WzGMjg2Fw5XxM4uIkyOqZL+SVrFPwgGaWNhaD0Y9pgQTo6V1d6
M3CPPiF+p6Kw1GydEfA6F6VW+JIBWjcfoLJLuWi2/0LjF0+TML5WOO5ixCMjtE0ijt4ioEYv5PuQ
L0/ZrCh2VxXDMCNv+C7xXJM/9Sat9zLMt0EKWMcZ8xpqXdhGss5fxeucpfmbL4eA2hsoNfzhyU7Q
PKbYL8hqMtQawWeUa9QI17/G975XqZflaIHPTDVgCKVUuq3XaFcUXkVMczKbOArfuLeL9hAvpEx2
7FFn27K7Beg82v7OMpU8X7Qz2zk+gZLQ8NDesfIFh02szpKvHcqiJyNywo4AEbQ5ZQhMZd3w/Cs2
4gLyhUkjHVZDZq4DYv3l2KmZV0f2RsUdqDrGOgTfFu4fl7/kz5yNXEMnM0JCtJp2JRFpswXcfcz7
e8BBlgIuJ2XcBvh4rMnxmkux/gs4YGPmxbyeW3WR/kuablJe6TZq8WkdlZtPzfwEQ2QhGhGoVuLI
mksyEq2W7/hG21nAhQJRNduk3Q7T6KyCsmjfzR3woYhqr6kowoeCU/WliaRRuHWVdErT3+m393Q3
iuJI2Z3VrKMy/HdDM0eL0BUJiOPcmDZSeKkWuUjP9vakAp2INhyciPdBc8uF5ftaGff6N8JT7Vt+
E/ELMoMlRiNaeW8sYoBSBeJpka9rKCtyzdB4P2ieIXk+NQizglbLO/Khn1HjuoHFnpGL75fK7Goh
TsIfYUdR0slJVWk8hbfvBnoviotFyHBIQeUT7BJpL/J+lqAsIJx2SjODRzfIYxbkKHts558pBLcL
yz2OS2tBIV25M/PGE5Oy3rWb4f+/JaPDVv3P71ApMhiecTfcBVD4z4KhRJ8vVEDMOT0tQlmRhNzg
Mdj6FPXqk/C8o9QDN0M/BQWX7tEXlwGIqDzI3NDi+wLKEIpEBGixcE9bo7qZAq2R5E2IYB6czV/H
61NXogRLRpWJr5VLJEI9Gja/K6vpV/P+v3QsJcBBTLHRca/cuJ+V7LAI2/2pboFVGcbVzZCiCTHa
yUR8IHUMur26lm0EePKnHrz6QM7wHyoetfGHeIWCEnOY+tUtD93ib7OTp8deAKL9uXl5n8KM6d95
j7szpaVm89+WK28OmWhkM9K5QiUZ1rnA/r4yVFEabGe0P1GstJoxzRwqkL+iAsyBaUmDrsk3khJE
35XOb3JNfi/p1mlkDr5/tlgdhcrfrkY4QkCpRoLng0EXUtY0hbjNyP3g/vy4XefiyPJ6ubao6Imw
kflwP+k8d76+qQDQ3KkSPKpB58Ec/tklh5fXwzSxMHTxKgJ4BZguHU660kc9Uw2ezAKP1ViAjF1j
4xgxSkz/lE3dVL15r1tWSzeku/izR3OcPr5lMQrV4ZVJltmR3G3pKlkm2CIAW9JS1P14XYS6gpd+
D8LqVPEXX1lf1b8/xMgjagSE6labo8GqwYWrnbcqtqcbybCWANxcoE3pozp/xZnwvgD+lR+a3/vp
5SJaUyHXx3jBIJrjYZQbiMREIK0heZSROiwn7/ierpPL8nHuS+qHIkpaHFrHX2mweg45fkBY+gTg
DqOoHhnUKX+fLIlsZhfGvnnK5V0SJX3Or+f73rTO2xfztn2k+EPNqGWq3K+6zCpyn+qx2jo/T9Sg
wdBMTfnM4hdkUwSz0ELEmFik6FW1v7HQR4ORpsEXkhVeK7aIU6zoeng9wLeC6qb+9oqe8ks9Buv9
ZLtsVthny7+JIXPka6iyuWaxwNjD0cz3vY9sz2DSlsV2uq5ZJj3QfweGbieSAYpSTPyMBvxikNh5
GUT/pqT6FfF8fhXPNs2PEE7DHc9hN65Fr6CT6lroo4qLfMb8A91w9A5T7OLFrA27JNR2w3g9+NSG
d+ZmIq8MmGkTh6q0MIxsXZO9NCSPTIONsBRuaat/8d1U7OqZ2dRfG9wg6PBkmB9PmfGAMdwh8ssn
ZbTiGfyiI2YusSUpFkzZhv5Uog9aMwjnIp3lbqoLJ4iBMxRSZ3f4JMuwLKhWc+Y4wtiufbZQc2YZ
SmV49uRix2PeYb3hKb7WUHZjlrnG+Oqos3GfcrCTlOffCNsikiTyaQMcK/1w4V3wEkJZanoUgzuk
JUoQPO8Dr6EXWXBww95v8DszPGHzBEvZIHlKtJe0xMet5PQ3XCKGf3bZfBNnq1bJqzx04vgIbJMh
5jY33H7gF2xVlu2viW/oksSZY4g6sZR/2IXfr7wAl5OQOSzVKksSxfKqDlFQza7vBPEZ3C1090h8
o/GPO8ZVNwfI7snGcy5+/aqbbb9P3YSw1tsD9Tz3kpbG0EoFBTvs17D6L7k51hHG+v4a5X0RK4/W
Ab140uPsgsx5h/L9zquo+OdgFBQZX1vnk5+DX4Bm4yjRSJmYqo1WX2wm9ysOIrGNFhpKJ/XYSwOT
08J2MJzBzKsOe5+5wwetcPgD6XFmCf3GSGl91THwU2cjNkAz6uRG/xnt2lKg0XXFcE5lx3xZJnFt
c4hs/wQLjUZnX7iuJf7s1+x0e/ppCjxS3HEJ5d6HRKxZPlAR89SedmvPXlrFOL+AdhJjx/Oiiecz
aS+L84aA6Twi/BTsOOUzck61t8GuyQUfNfLqdDo0nCKiEWnn/qQN2pUzuKonPP9EcmVuLAwiViJs
IgjxiMKUgHdI7oWTXy6wZbUoBC5wlyCTRaWdrztuaGOU7wyn6Q2AzXMeOSCiTHZbwWgsnLSxM0OG
tUOgiaOr7uwHiTtfem8QvVbUPCSav5T0WVDthiN6mbAzxZf5bI+vgkXRQDD0OKwgHvR3bJA0y6IE
UZIJtgK5+80wZ2Qb6dh3QRwBpNgCJGwvRehKW6QF1XGMlg3wRZz6hugp7S5iDC9Mtrag4XMmTK6I
4FMDnx2KNBPCerZ9gYfxx6G6uTN3QOebTUbsI5JXFkYbYewq5essqyuTwjf0jLJ25dlE9YLtECqX
h+qlR4d8rLkcYWo4WRXBIh8pP4k5AmBWyV3+ZHbG+pE+72m5cs1H1+ku/TS5dNHaGW/e9kx1kIbo
Q7fKor3N1200RnBsfzlTeCyUQkZHyD1tqD6LiTQp6itbZr+QOQ5tvPMiPRkzm7kGeQb1BChRtWIB
qOZe8tEaZAd2Nf5y8GRGqtQKf+yhQpwkw0WH1IZDAjCl7vsbNTwXwnirGEuS7N2sPkzQ5+hu5JNU
3MBbMfWWQ6EqAmsD4sX/9tND0TAozwCfEIuUj/DbckXrQoUKsTRbhlLTc/ps/p+U3tyGFdQHWGG1
lj6ceHcxgMixMpnvJ61QlGEiSxH2hFQquew15f77Gumi73x5hT7PwoDLCIPDs1HU1t+NqupVnLCs
vv3rJ0Ep9av35sVJ1DtIGn9cyIUTDdKzfNnygatAgrDOT45VIcI5W9eigiA0TJRA6m+WT5R+BbvG
kT7Rw8mHUcf+AEuqvfIZuI6Rga9BDyMWv/xbbhQzhqBRlHVyOHa60RzwRH5h4jflWW63wyeALqX0
IE+PHw3IjFpcngxk5DYea3bQIMG+zPx9S+zgzaH+wMGa/7uwht/+Qbd+RkVXC66CkmApLvrskZom
C+RvBBbcX3kaYvsJv7T1IJ4vf3WLo0uaCRdgWvb6stb5LUlQOrr4yAmjSNevwndmQNZV2zBuVrcC
TZzk82YshMH9TbN9cRVTemuYKJmthBJAqiVNPwS364Oo2AuL080aVRgXoS4wRVJ7Aqvstl2239fU
Q2Gxlrdfali/Tb3mV9PANTueNwFzMKkHfB+5PcQp65GbdhMWqE/5ff9KValOLQvtgcsVLijNTWpI
Ld8leNZq+0KC1H67lH8qcqN4BCtKAQwhoJWYUFWkrioBQGs20mPikIJjun24JN4yQdIHEFGF3R80
VEmlCdABP12ra5HvRej0sTKY/yjIdpMgP+OFL+picqZvRuGDL29qMDq5T0YDBwoIBRyTwJscpSmm
VY6rNjv+u0hBvtxIIZIubtEgUWokRezIsbvb1k4l6PjDFroRn5mRc5GNBKZ7OU0g66QIiq6k6V3r
SK3kEh7qYyc+nVVCcrDBXiX0uyOlXFOv2rOinUAgdW0hjqFB+ksjfCWns7tpUtQE97Q02NGbHnLB
/NaRWrQUfyAjp6/rxFGif5R4EO7eiy6bTNPvtgepANQTu8osszPLpa4+GCiqwMbz65CovEMvyItp
mnS6BM6eljbc0bn0N3BWdw0FYZMrMcYlbehiIdOeStVFLwAGfezknMWq1cYjj4hN626OIlh91MiK
0iVvo4bwCD47n/329R/+hIlj28NXkX0pNtYLA0BoixgDQmajTlOTeNFM3zSTQltkGVKB1v7PLtkj
6MxbD2tiWeXhMDYSKeJihpDvTQQfWwN1tEKutSdk95t3lQi0vllma3MvyoJEBTaot27CLB+SqJc6
FYeEXZ4PMdPJB9X6Bct1WIlczlRuJPBO/oCcOc0aCvw5ApzNKQr9D7XgMQ5+2L9AVYSZkg0HlNlB
eaO0U/0T4RdH88dWiqwZ3NRKcjpmTbkwQSZ+9PJCjcJGj9TQ18mOeok893Ms7jUeSo/d0or9M2zA
+jxceHyZeNGzQq8qMYd2xNj/6Brt6jH3Rn1Q6m70hx0Z8Tz8HZHYH44nizh+EoJiJkZHNby/BiwE
M/Upi1dAeE2XMlm0fMEPTSubeLDTppW78wwQc+SUoqLrePIPNPLvuleuSONvGULi4BEk7PAljKlm
4w1JvH2jGtRrDyUSAqWn3dF8y6vSTFbRucmTWvf+wTENJTxGuczCS4WQO9W0dmRb/GSUlTR//BHY
RxKvYBRslsokD3Avl5xbemR58Awu882fOGvQNLqUUGiBKgp0CywL37Niu2x4QHCwxcnQNMtvfOkd
TNMRJo03SvzoWp/ni0ytP2XNRa0x3QiO3DA2P3Wg1NB4HNUTcr8mnfx8a4sI4VQ7l1gkjf8Fo1PI
+F5pEHAA2EBvayKRWKmpBfqd2HXjWpDV/mBk2QYx9J7CT69a0kzWZrPak6Z8LTcuSibpkPZE5I2p
u2iE/KoW/1nhPtiF/VEqksWi+dDaxSVQzX5BBbau4a6uSoVEDa75bILS7lnnbv7jETUUaYOc0rk0
jXhFDNGBMIpVTCJU7P457vW8usuP4wz1BIL9diGdx9fMDtlnDr2Mr8FQbhahVS/+wEYQqQ3ivB3F
m7ZJ4fWfip4Mc0+v+igZayijnyPrZsG0jRpPvoCY7Wn7sHsSGYmpL5ACMaEIX7UvtefsU6/Z7Ns+
WPMjFJ2ssOqnokqlMG9tAPrneP5Jh+Z+EWsbzWPWZEsZP5dXJHq2iJwEsP9db7qIXvKmB/hsb1km
m+Uqe+V0RWslKZV0XEuDtcoTLxGNppsDtUMz8bCaHbjHPgYhheop2RS8Rfc9MY8nWq6eOX2eruBW
O/0LOXQTaV1JwzUyrulKcyC78OT4eZTG4vcj0qMm0atTN3A06QLF4BQq6g3qRxbA2JtfSngjWLBE
ieSWXvUmtQXEpBk58JuEcCEnGVtL4hZRGL6WkREqyMxD+zwVbV3+Ble3mA+5LNR++7uTW4rLYUE3
C92+HTkvc4X4430qZ9edz69HiY064cXPoLpbOcjy9wRKs5Zg1wr1Gqul79Km7AgMjJHu7EqsrPcB
BbTwDWDVvjN7Y8KilhRIYgYyKwJDKG5TVfkuwnUxLcwaKmFZ9hul9jSsyJKM8MpQ2dkUeVUtX/AH
0KU54Xyv5Tmm6988C0mJXQV64cmtrJGgz2WRTR/97wJdAp9GJpJ50/P7Jyh8usVIwG1MiDDwCsPm
FSymM+R8tpWzF9Vin6YH3TEJ1+gGUh/XPB+W9UFELYpGhlKylbbhY1ZeDesDMTChyIOJzfFQE1FW
WhXo/2cOEmROI3JssZap+2k3goDG9442L4sFD1lmho4zHmuiPZrTe8OxwvkRB563dAlpummouh9S
Q/yfwXOToAMLDiaJ7OcUBOU5uZSDqdV3JITrDlj+YMNFczprfb5JzOp+FZuACKLHt0K1i+9Am407
ZrsV7RdiEGgb1Ct9ZQfO5wWRYm/my+NL2Sw4oSn/NSaRO2j/v/qX/BULGocrF+tv4KJIpeOmPyaK
7YFFpLqw6KJ8MiECoUKmmi767I7/VHDu9m1odIJ0MpDmEVR3e/DGBSWIwr+rt2sNnWDs7dgzJcuE
ufIa0xFMq5OtXa4KLqQl7RMpDDN0tOm73gagXre4+GYY9EOheVNYwI2UrHw/OAEga/1nJ4l40xld
5NYprjBojBPZAqcxdLaeZlNX+IX/aE4/rDYDXQaGSb4/zudgjOWn+32osOGHRvxCoX2wkmozRXmf
XG/pmL9oQUCxwIyT8vJcjvLOvPZNtpsRmI2PjXlZ4x92xPd7KdRheUwsAW2+qXrxCo1n4/j1kMPt
YfZqTUC5NCWJLuq4nnZMS5bz6Zp72rKgl1Bs+oVefeZFL5BU6LX9Yt7pg1hkwu3jmLQqrKnLrb4x
Blm05H2u22FXhICpSUm25Cuq2H3IaIUKx8dXU2bI4vXqAGTfdNgqN8Qqb0IL9VRjRJMx26GSJZij
ki1yiKkf6HmP3/uafjnwEt6WfVpByJxg0m0ojAFB68TJoBagRY/sXyoM7mgbFcQjCPHcXz3N66my
jqViyXtqzkzS1tanKxnoYrxXzSigaTccmCAQrqz46MgaU0cQSEMvG+gz8d+7YKrn317iubsiE9dE
Zb9W7rF1iPmPagvbjNSRVW4KivzTtsogsA1T5UwidjgeXxiGhg5g6t5AbqOp6ctGyz+DrJJ3BrTH
YgQ4HkSk7TdVJBjVU+ummXpfeaPQ4v26Em6naVyROJJ9J4tw8NZfjcWhyeqBb+yAlUFzlJ8uDFT2
iF5x20ubg7qQEhSGV9Y7g4WDQjv1CwnLXbttHEPuUzfbntD/2+iDqdVXirkFSnDa/UOjzUWSSZCx
fxaP9n9vWD61hVTLnx+7UFHwiHk7YvenmzYDrqDuRqk9Gba7cCxc+hQtLEK6Z8PewDD+/FsOatmW
G1fXKcoKqkuweYEkWDX42lIwsPDj7ICgBonCRgpjFihxQM94TQFl0bH/DsG66sUxQ7mkg9QlZ9d9
dd/HimLXhmnb7abtlJ7F4wW613mFsmPWTOCdxYJ9FNMelMaz0zTImYsyG33GUcfEYLte9nnrhTGt
NoVeiiPTSlp3/XkBt7YdRQgQfjr4SCbePnzfEkUYQ60MNZb3RGbAyer3TovZQx/GLnsSTpCn85lB
BfAzeKM0eyuCl18g8LeM74QBEDTzMj4F3GwfGOCsJThM90wNyJNL9iU0xckLenpIZ1cpB5hpU7pI
0or7KyOM9pUv/YIyjozVFrM/kHKuTYBEnFe6hKRNXXV1nxxVXkPdd4ylSz+c5xO9XsHbcnLUeV7r
YxjEoNw6adiQCFo37T5QwEzXzrpj4dP7IfcC5o3bmYwjq3PZZoAXnJGb8cscxGvIRh3c3Id25Ryd
GZqISld8munLueQuYa3CbmpwtPyYeaofo801dhKvTlnSkLnF5OCWTfiA2wOaFEgLp77EoeiVP6Mg
wS70ELHsip0zJIWqg66QeYx52LY0RXQPyO8TfElYUsB0m0NOEapbl1vV3nXwO/wBrDO7fsq5YO1d
udkyy5lFCBU9WLmxuKwDb9F5gi3aEjLC5hPQU/i1aEQaDERmTi1yYppXvy+lW2u/82/7fDl/Y6V6
BZAEA/OzniJMdX/XKMofRGZu2HTGt2MX1Fb0Xg2k0Qv88FhBI2eSN6lXvh1IRvIfR9t+q6bZX+B3
6E4ot/VVsRKTajFtlb8/vIJ5gy6Q0Lo2QeDoOJ6H/rY9yBEvLZGRmrxgM/O7R8mkcNMkNBZs8qLS
WHrQN5tZQ3647bkToPlg41VWnLSrT4UfmjTfNcQn2S29XPWe7TsjiInfGIBB4Dhab+hoTY3Bb2ei
62v7slGHowfCFTeBdt4lDfZf7O/XXIiyGKa1/Isy/TfQt4PeB8cKWIE31xkcRIWEs0SzAYVEKido
mxOtLjJKGA9UqHT9nTEP8zMHcgmbiGFF4aCqjrYjgRqaMoM+suA8uPVBNpyL6uFdvT2JyLp4vfo9
SCt75ZUzaHoVJyygruKlNJUoHMM1NKLEGjONfnuTtty/Kp9KjHDG3L5IpTdGdqvHVlD9vaqv93W1
UrjjhMK8EsInJh4JD+/lC6iSB+ilueoinbw5b41jSZtuYLcG1vsty5p/wqy/i6e2BUHw+G5QrqS0
Sc5+09Mi7Wx5nEQvvAB4p9i4raWOEYuPjgYYnafEbBiHyCBXWpCktJ/DGzig8KG6ZMK/Q6tbl4KI
D3kRmMGf5WUhkBr5IV/sTBoImstiqKDOYRsHnrOHVScPmcvfAmAC71e6l+kFHYYu0sanlaqf6oiR
AFAXEt2t2g9AGmo5SzIIF9DhbOcIpfXP6aymWb2kK7RvGKeqeX/K2BQ7DHXLbzhbKA7iG7ktj0MZ
EXwGhec2bmuR+Lw8Z8fU8yrjlLEFBKzMOzb6Cfws2LKOr9k8AK75FyJxyBsdNBExjRDSYRE3QQkW
WP+hPtv8v4GsnXTwfI8AmFuGAhwMnImrobl+LJrmmls8hbdE+Le1FGJu/Ok/EKLXFYOB9BXaqRoF
w9yfa4toVTMNew8dtpoGgPuOSb/HpCD3AMjJiFvbUOaUzzlddtb0HBxoz8zBRm59NJ+yIE9Z7dyt
Wg5pf8/gI5/hKBfHrq42o93/l5irAkTWBHDrcaskvl9Stid+LFxW8Lklilly4yZityRxopnY5dBV
WnoUQYEDzI+jTzJ8XkslxgvGB1U/a0Py4EF5G23KGOsiwZzNQfo0DFnLWeZinS21y/N/zFz1WRTB
sCKok7D14SplxpYKry43EfHp+Y86e++AVZ/pAYjgKlgDM+1WANl3IW/c6oCMBrf8DAlvcjXtuQrk
MvvCYP/2CpHtl14UqVIkP5fSMSAf6nI/XXE4IRUVFOGh93ne/rD/K6jc7+CUilBj+eaalQHJymTL
Cl/pWfB0EB2/F0XO58uXo0H340CsL9mO66o2cZ9PD58hwSgvSz1YodAzEDTgQx43nD1c3fnOEdDC
6raDpnz2yTNzKeQACTjLUV580gMkKF06iMAk5OPs78vxrP4NdqCUyTSR7wvVccK8+XthFROiUPa2
P0KqvslOVGwZj4o5rtYHGG1ykpkNFpU1RxKgxl97E36r142OeuOZThxvdrniVEuprXYKPe2JNpET
ffSExxLiuEKf5F2HFcYl1Aua+Ut7SseBU1wRpGM0oZr7ks9AzYAZGB2vI8yGTN/gJsDSgJlcKXXZ
G+vvDBa9FWaLBKabZK01T/Djxjawi4N2db0xNypuee6nTYTGBJIpOtLmwXOloM8hGM/R8l4/heXo
lJPed45O+ka1l84TwXwu5gFmX9Xxe+dmYPm6aPgJK9N7FjBTpMyZDAOp5xpWN97G0qekxk+0kY+k
ZN5PiFfOc9W7HUjXpeWvEw23jH5eReAGEkfINQNfyDaWO58P+UL5kHMb7RZKM5ejBmNg5prN+vk8
hTDNvN63Ny6W+y3gEMNvoMllRz8sUOsV33rPkH/HkrdJLrUG/iSH7gLhuC9f5wJsDcgGVYFBp0mV
Kkr/ocv6LtGwhMb053Z32hVWwN+v9Y+g4L+6CvIZwPe2Ft8QDNcF2GSoKqBtfoRPVahpptlJL+S6
3ZAW0HJ5Bd2R2/OXHCY+FWjvju48OW3AUZROyJyl/iuxRZ62RFW5mMDYcPfd4nhXqwrsWA+8EPIA
4ChEBzvYOt1mjsBJA8J3dIkd4fcx1WCrb7IdU7vrYZuwYY3UNchwPB77/U+VNMKmLmOXKkjSnYqb
/94+18SVhrhmVd6ixDwZFmxWoQpvzhhMbSCbxnVTCGbDtijbwykA4qsSXpi0Sf686/gNGcMrrjCw
urDJqHtqRAWPNNUG0hk+PL53T9Kb0D+vGnOPbOqqPOEy7wRRnMU/DR9EMkH8wGNb8ItQuZlNyYl6
XTjGPrlwHeGfqNqT4a2nIUUNEovtTLyC4te17RkqDokZ59Kv0f7MwL00sB9BzMPpLdvry6L8w9Sq
60QMspfzVdzdcdTOfOYLmvmlna4j3HMBRQS9BuG0kytfCNP7I1TzVOvdT6nV3Ux+M2Ixdefu7I5m
13+eeVXDrgQG1fDfK0ANg8TRpMK9noTShZzo0emoJ29nCWTxyc1Byl28IaM1MBjpEJNgIsjfFLv4
xDF3V5m+CnBf/vl75vPYUWb5hyZMicpnAN1d+K3SIW1n7b0ybgnbJSCQ84uhOTbphPiw7yQtvzwO
62PNHd9tMYx+c3QrnKDQys5BEuRR7CVYMoDlv/nX+ZOKtZgVoaETmEHuwaApbPSwPSA5vDlNGCVc
fW7v4PIFkQI/tqosVpvGGy/ayJTj1rxeVrsmibZ9uGOjb5FR8H8mhfyKd4mNUcqZJYo0BxUvCInW
V+mSKjLpp6CXKv7lCvS1laNjsLTSYzqONq0jUgj0DWl2hWKnKu/mrG79Rny64y3hWqB2fLUasSZL
3qok54KBXBOvuCXjJbcsR3BlXWP+JBrHiUCl5xkm8gDPgg8gUekhNS+7gPn8/GxxWo4NvKBMD1nq
mFBOEl3Q3Xf692ovDyhxSqwPu06NI9N1xWc1hIhXK7a4CD8+Gq3MI2/A85BlP6CTr44M4ntoZ2j8
Q7zzHo4wSZr4so+QI/vA+cUVQ/BX24RBAO34xd2T+8097W+pjoCHYEkNTDQLlDnf/Yrj/D8JNKxp
pNlSSTJusABIMRFGXQEOh2L5ZMFlsiBlSs/vx4lyTArigL6bNeRqpEl4XwHUZqB9mnBWLgbYyUYd
Fc6rFkZVrJDSfH+8f0bkoKLt9BwICWbnfnKlcmthZgC15fCeGbiIaCJ3Ck6/qiDUc0SfRICO2LSQ
LKaQIXZHIwpYrwOJdY7VFaf5VzOZ5gEZ+FWSVD6WehssR/PQgaNYZfuAj7P4xo9tvHmSsBKCURlR
TICmd2LEenhZwntxo1p1JQY5VcEFGducCXCAcQcUGSpZXuPkLCnTVX9tkS6BKtLWH1gbB3u9i54L
ft87q2ccOvIUO46iqXOG8cOfrue9F/KzJasO7dOX9VsQI5ef6zYj3CKI6aGRswVhUALgQqb2N2k8
qy2RJ2D6SkfJowf/qbHwpqMMuEmIjGD10Hv9jdsS8DqIAJUVmCM14KCVEDJk/yEVr4qm1Hm/9mDa
alSG+MfxjFEO2ZIxTFb9ZlqUspaZNfmdkOplMCXyAB4HeGXGQ580TeZM2t/WgqE67TSlqngftRZ5
0DuwAX1SBwQKcJsqu8xq38w2BWfzf0PqDXN0bFw+0+c7EEA07K3L6+YurjCReK2Ywkwi8vD0FO9E
tYCQSWhWIURQs7UUamfstnXGlgBZSr2+3F8WqLRQiSClJJul82drEXkst0Lz6Z136KArsnF5iXls
OH6Z7P4q4LK3EDyk4lI6yRGHOFDaEEzUz3NQc99rjzjYaRf67rA5AcGPikXCtWJHVOOR/KxFO/k2
IjgauVkGf23v5wlY/GujgwOONxgaFog6+tqrZg7CohToh1wQ2lhxUaqdcbeB+/oev4FqBjsAPQom
AxVj2Il+cBR+oGAQp24UE4W5zwqPvowtaZEUU4oj+sL7Vf8Db+WnIf7U5lI9Z+B33LV4V5AjJdQP
q3yqF8a7JLBFqaRaCESgIMf+NlzZau6BOSl71gGfravr69Dvz2ef4clZtEr6AA59yTrin2hPhCU9
S7HqlgCFQQbULZqnCqeltiXWJs1o9nmc7Ij5A6/0pccw+BOLZH1DCpavMLxw6UPK1Q1Ntb4Z5TYQ
ZEwKeETyL6hMKIuxWQzoQwzSLGkVzV0Y0CQxxELPSuDAGl8iFFK9GB6TsRiVdfHa3eLpVyRXj/Uk
Q7pNmi41BIWDpdqvv0kLve7b7Vsm9rZtoo16n3N7cr1obia4ZBQU5mrKhQXWn6ze59fHdv2Y6G2s
4FE5T2uJogquI5scZ8m2abRuU4Yl75PIL4+NvozCxPpj3LQKKfDSyfJTTcZfFptYpq4TWe7vBJ3C
6vVkvwOB7Agbo+jAlMhCCeS7v06EHM7X+Rq/xU+x8idj+xDwb5Umw/Vz6mbLB+0RWij2DT6scYl+
ZZfWZ4PP4sltS4nlIuKGXqJopI9M1M8BfM54tU8/AQfZuWsuutYzFqYPLXFq/N+YJSZ/JlRJC6fO
3kgrNhaQpLn3kcVykOjNFJfWNd+ggiTVxPyyXq9npdu0sE1eriDRmS8Bt1D0fsx6x6DkWXJvJTIM
oavn+YbQ15je9iM5BJ9YLClopTTAx9G3N7w+P+Gh4EGAObT7aSCUDZEh2pjxgvzdaq7Yyz7U0VIz
9623WYlcbWzYZ/DjfqocjCGg6bwwZloEgjmut0/7n2pjZ54Ka+axSLXhnAeqRQ2aYgmz+mF5ovKi
Tf+65g8bb/lIMj3W2PO2ZLjt8K1Pho26Kqd2+s9pWa0qmL6JUgwxiyqUk5G7ihKCa5X+Ib/WR+J/
I8LK1emGmGjerbscUyskoRnmugVyo9lsAmq4KYhvekv4CoZwZms8S0UKAPweQDbVqHOoJRpy7QFl
t6HLy6sLqPTxLtSyFJIL4UiDfCLj5nG8AeodIwUtbeBBqhDuNSJheetXMb10OWeV5Z9asTDK+1sy
0i7TFssTIrL4Q+gp7VrgWb5VuiQytP8t4kUiWHu/qmfpC30QFfL4/Uw5rHTtu4Tp3yCsTnbb4AXD
hQruyhJ7sIw47HuXhD5fGfAK8LHhxEleEWTaevIF0X46TyHWYstLbjNAZYjpVVbSavO2KDgOkIoJ
bQLQu0K4fP+B73uKg0lw7tkSfWcIatAGBqeDonhnYbydXfeu0Hd90GNe5SdTXescC/Ro+3RvT83Y
FgHIai/PIP84QYNKCWtaBYqOqffZ1Hc4Gd6TqGn3CEI0kjojdSAt0h4yLa0iNzofhRBol4ev5167
/j4svfA3y055TbmzaH9P5AbAAYjwct3QafLV5tGWTG5qqTMkyXFX67hoV/dIZR6PqIImQn5pnMJR
UyXqVTSKT2JjYQcUrTe08JTcS0cAecn65wGdUFEtD6I5ZWS65MQUgYncML60aOUQ5PtW+1WzfKw3
iUynWqZgrZ1gfY9SlXg29jCJ5evWQqWtfwRkhBmzpQeHuSIOJDV/EU9DeFA6P9ObEQOvP7u3cuEF
BuPphY54bDqHC5VdMz3BBCFRY1WptTaz4yc2jOoIsmqQtpy210RX3RQbQa+MW38QboRpD8laX9/S
x9O7q/gO1Vx/vf+i59wnFb3AF4WT3wUVjpYMM47opdIG4FXoLxhiLpgUXVQJSZCBwfVuSRCBNVjK
Pt5J/kGY7T16XwObheA3UxKFgIvEoERn0UGBI6AmAtmtH1EAYmDyiqB4Py5T+BgCw18umvh2U2Vf
e1bVemO2q0onpy8J+lbwn74zOtAFPXxB8Ib9RTgzHDW+b+f/wSeEVXL8GVdErQxrqSLH6aBbRhGW
/ooBfxtUE3w1ngH5pbTQa1Hi+Mb8BjAtPjFi/BsRQBdtJO6aYuEqvZtEcbgocjRUcY2wjcy0gVLs
6H+EYgJIYbRgJDuoYHVXmgIknBOgBkN8crFK9eSqoR+DIm+IgKaqoAfxXxpOFgtMz0hItQIUNFB8
302YePhDOHCC1npZGIxwgaLB54+TM0Wu/YOy0HdAlpuzAWpVifweUWYRe6O/wzckI0Ld2ZGJkq+E
9x3QAXz18leGTEn5P4Ivhz6+ZvOQAB1tQ2KMML29SAqYKqTfvRfGco0x5aA7752ugyVsNl2sDzEE
6dV85FVOgvDSdcygZt4d5HxSoEKyV0A6RjcB8Zbv6baAN7/hLDZdCIQO63bhJ8ianB90Rrijp5kG
Dctfbke3+aJslRSXzuMWEe82Epm6y1iXUu2eNsw9vUPTDUiW1LYb2mdaz+i/NXh6f1VCxyQna/nk
TBAHulihGRWLAlTeA8x+0MUa463s0Yblnb2ZtpNWLbFJPpDKsAoCUQqWIho7sJ8Q6NpP/H6OtXl6
ykCUaFCn0qfcHAzYm5fCKP66P10HlyEGLkwMAqkKtDbJIKeiRwR71sJOpu58HQZiUB5vBmjL2w5G
UeZMGyx2ncZlxjiB5SvEmAgEvh9mfFXC8hUCgf+p455ZDLrEH0xJHT/wNXp4aLPjD16bpJ2vBVn2
s218rNl2hZ0tPRACY23dRP992VInc66xHR7g1ytUsQm1boib1CaHs8hwa1W3XuUVyWc2/dJYNV6V
OUDxI/gQTVefR+oQnYMz7Jia5EzrYbBJcBNHSLiyE/vmKW+N3jSZFrNeIQwiuhzwdYOp0CbAPvdq
mSr4guyReA2cpF1aEHijKoZA9ZwqKyP0LKR+KUEG0x/6ybdm4xjYz7iQZpTuo8nZ1KQ4UugxFwBr
sER33gX1zbST5tfURaGH8PA+mhU0QH+kVwKq9/BWmgpOd35ZO4XSE09/lboQB4/NG4p1icEZK4sD
V8qox8IHty83oOYaiODyXMtgkADupohyBoqJdbiX0c10NAqDt6/neWGxIRS7YwBz/jShgxI5icHT
28kBdPHmhBEN9QZkEyCTmo2ls2CE/N0OEgWb3ChSd20xxbwflrI8fTeDf93LmL0hkElENsap55Cz
cde/gMfMMilmUNQGUy3Q2RGOsj6RZ4KvjhbCp6AErjmMWh8OsxMS0G64EzqDtL4g0P2UE83AYbb+
ku8LdPkozGV0fogHelK2TQkEpE8LSCKtKQ5l1V8+pffNeGA2DTRjr3otOhPPIo+M/R5sGvS1OiyL
xskhYGkAG/W41YkX2kugjLrbkr1UNR4Vr/p6P++louHfgIb6kTa5cRdCtfgEKJvEqCKukiYwHIfA
ovU694Xg9MXumEioB6Gkc7fgF5t72ltpCVfRWYeUm0Lrq/4JUrY2YUJtL2VIX9nJQeOfTQUaKfCC
r3rpR8U7uO2Z5EviTPkCrR+J5w9WSZbEzOYewyu0KWDkbksytXZCOFlmZ6ZrErBHIHnvYZczxNnJ
5Ywjo4vk80bHehcMJPPAZXD2prt48XjSbRLpNHnkVaNINR8eOqCrzK2NvkipMc/1Iw8OHGSxE5I4
ln89z/++vfccQU2ATxYLKj3Q8gYfdpUjGOOSHmlLbT0AUjkZ3fFP0pPzYWgyGDOcrmjddIvhGY9u
mY5F1iSDBEglhq9DHlR/3U0+/AwcISjyh8qjfiZVK1I9IalXW3VSkSv6FAjuxMkRuPuKnZOl4W9t
yVag/E2kPpFxu9HjKeYwm2kGrCDExUOmqaHZsakMqMFwqa8UGyRblIMTu5Vbn5eq9KMkeP1eAC5J
AybfeGHzpgqHV2ZHpReVD2PWZp90s4ztgK1QV93PDKn4dNJ59X46ygalFchLn++TWogZ+c87rqMK
aNki1PZPTxXoBsfZHOIQrMXOVlqeCpDWXTGfyZdO7EtNgSbdj2ppCeaA3ByQMNHVIrpepPABPI5i
Cz3X9ZWLSmo//gFU0yGsGN9AtywwnUAlovXHFDo/9p8sUx5Tr55z0W2QITV4rW61NSAWJySc6oEu
eRTQ2IRzAs1/p6v1RJVbF7s7D6FV2v6ppPJCuqzQnoUzI+qlRiiscol+YH8L2Y8UJAHQ6TZSEKWf
5Q2+l5ou4xW5vviWVYTmZrckY1qZ2qrbX5DE3g5mgxUWfPoyIwvPsvqjGb9VypETeJtsmlvrBA4I
EAPo02PuoqMAnFjbmfz/jsRsczb/yjlFUHKnmH9BdkeV/8+QmKWys/ZWGDsl1l/vLHr5J6HniDG0
C7F2Vni+lkTISjK5z8T5dc9xtmSLhKMPS4BJzfZKSth9/Vl/y5oQwl947KgzpOg1ZCJMwj84tDUJ
xKfw2O5p2zDVly3CsJDOYa5pBEMKO88vacWcgjaulfhcJFmp4eIVPFffSEfcHDuQfC+bm9q7E8e0
bh3bdBwK8ZzUjk7Y78HuOl2cH7i+OOPiv5QMFxCpXEX6eUOGVgiLJRMgvkizT7R+Xbf8bNhAn6Af
rKVCYExqTIBXqo5J21HRb5KUEYwCrCj4KrfYuiK12ZlgFk0tD/VlVgol7mUUwyQY6jjdYjcwT2Ko
FO+Ii5WJgRa5MTkJh8WqVmi+Gko/NPDf4ZQRboycvQd0TciLgg+0dvGnO5muTGuyC7J+kSK8jNrY
StTUePw60pgguUI4tpTC131T2Y5042GYIJ73b9WR4myKjkaQwHRAZNqwUC+RtsDd7CjsM5vo/dRp
lPulqa1MBvFU/UjGOd1ntuP/OO8tlamDydZ1BLzPCH6Q8EWrCy38ENrR1rkiEQjAbw1X774VWPYa
2aMS8ciFCX/17gOPmBAsGOtCcpdL3AFcVMrK3R6lBOK8oJnU36psgFqpJjtjqlnT3yT2hguK1dpn
3qxKKcA3N5g38AvSjP7JddVHU+X/4aL8jgV5cb+ClJpXlTtMj9FH6YAqBIGsy/zKRnMM9UwdSJMZ
PrWy8Q7HPwG/ddN98a3RAoX5qvRlVImDkfh1xEpN3d/ggfuAdoZM6Iv4AqPvmWyP93MetXNWaQf2
FdrGBRZCvMAVy37Ru289d27oz0/7VWym+p54hRjxZB0B/rdexEdtF1KivNSDheaGtky4Xn/UIW5H
+fDvN9Q//2PAbNe/j1MTbvGtslR5X3Wzp7XEwOgHpP2tdjNQRkVYB6hqEfr9fpyoSDyYDqSaGYnM
73qqAz+sXC6v8xF6GQLuIM8HbgXRpUg+jtioBWxujaDtrXRmW4vTJPUvtwh9eB49Jhrnf45eh4mp
E1sAjjnxbe44HYPqi5fTRiYr9aGE+ZBSqv6X7dHh1T5QBpndBbjnRtRIf8/lQBgHvto3qEj6ABX9
5k6KeZaKm0rJWF1vi4Ub8btj4WHF+b8kAu7V31EOawAH7qeJOOp+xR/7AI5kx+HOrglpPk2r0w3N
KxWwraNMRlKrM0sQbTORJQNPCDLs+dsYqjQUkSXDJ2lqgmtULSJWE73t+9CUY5YFnaJFMeqmZOh8
blDY/REUWs5n8VAxyw3EwHuLDeg0ZAimjKOasRjtD6wq+ELfdLgDAG9MHqGUrJwsGB79QH9Ljz2h
jiD4hJTpQjEGkXaw1y4qLVGo4QkzPYW5YNPA6P7zisXZqcKzL8uMlfcyPXqodkavqDdNLopdc9ZL
ycgbCjIRr0zmP618eO6kKKbmGEwRVdIXZe/nibIME99hChYx/Jcl7ZuBVfyU6c/SHzRFn+1OxfNf
TCLT8lv+bocuceE/A5fsYIO4xJXN62EhRWojjqOaDuqaHvWjYI0PwIT2x8xyNHZbcLwNw0AmIpSx
5V+fTUcCH7uTYBMJ/g+5XHvwvSB6UmZ+NnaXN1LBqHvTQGuIZqT+5VAV8m4RgNuLq5BuyCVmdjs1
geev29Cweb7iumiEtpCj6KwnEkeEoaScEa5btrFUAx7u4YO9QxG1Qe6qo1Oy8Rln2p5H30cByjxU
d+ImkTwtpmxRoFfw3SZoQHc7ulyaf2HpskqcEfNYn32IP4q4HKAUouskfB+UIgG8gYTlfgPNFAGQ
KQt5UQtPy/PHDwF7peaFZr1i+fxrGzxcg/gOJ9EnY0gkCuWV5kROe8nLupvw3af6tH4Zza6rOWcT
WfmAtF/gzGdwRH5cWc6zrRJlxXs7wN4KSjjxyQX0m6TmFgu5eGtd4HFAA4ieKgYqDc7rEmHS/gI8
DHvPosEDVCHaZaPtklcW8j3/uJGWycL9kOb8WjJ40G4nAD8z87wXMMDDWTR8jbksPDPBbLdGdZM4
TSED3eG+d2uEUq4ityh6Lx+Z+LsZ38fSbDPOKWg8hvoHUgKmRqNRH2pD4+duBhGkOWnH1Kpa0SDN
UQOtcMLceMDzUFezluboA/CQDzZQz+/YPODKE14qALRlN0BnozECneFaZ8Xg5dXxF4l5G71MPrlQ
/PPmwQ5VaMqB1zvGCa1e6To7ZPhXkj4ugg3UqC4UhZGXCQYfcLc+jdKSUU/fI1jvI4XqrYlsDTwE
Lm36+AmynVy273j42BcCbtOmv/hZSW5/+B+gJ/kxq10jA6ed3GcCG607BSBYo8X4fe8dxAXWttw5
84RXMO1xou75Scq02D33vkPbROKo+Tx6Xc7piKvS0xqEZu6ClyK3aNwRyBaYGyON7m2hz3Hj0HKR
yxG5i7zCU+A3Ud8BB5OSBu5wct0erlkwiVdHvDObdcY49rHfSa26QWAyIytmjaSPs0uLheyfp5FZ
NTYgY3Ab8hzseXXjqlxTXY4BWQrQdivPoKEiRGXTpTG4flL6Uu2MpZS/9V70nwzAEqfYPcnTuczR
XIlrB7zYB+Gtt4tJiOOg1zWlhlOLYjBuhAyrqHwBM68KwCwYL9NjOkfTbHjhrJ0z/HLdSHtyn8sR
t80J8/HAz/SMDMG7+1QnI1a2vNoLd1j7RUtRUtNmep35rh5EYRiZDei88XoSa0hiikD5GfM7n1ra
obTbf1o2ttjw27Ec70hstR082vmXyom9zZZZwz9rNYtLljBVWiZafduOOdlawySTdrhAjCwn1BqN
nEx51feLoci2sF5jTVYh0cMiEIeWmvSPVFkmemysY2MXvT6UI1Dw3yemQXp2kJEgGkIK/QiB3f+f
DkVmG6Il1W6qQ2S4rEGcOX2J6UsGAKaj3nzNlQqw0GAxJFFneXGCo5ZMXBQkUTdU1V7mFENKSBvd
Ul5j6+8Ugl0AHfmkIgcDGRQpFTfUPuO/zj1DWW/TfzIlLPjQmr6RknQyYVp4b3hXbP0VUoSQFbwq
+k+L3UXwZUoN9vu8LtF414L63MqxMyvaE0LPazndgsFOZrEk8sz/FnWgFCvPC183baQ1tECoUZdK
umxmXoeVic1ccIn6Qknoiu8oWr6V3PqkNzp3KkPVA1x+OM9NqFPQYaAY9SIF825HvrzJiHJHWgZb
hSBApuVIrKvk6/1Qx3ZSTI563Twf38hIycRsiKJFbGw3nITSL7EJC53EzGf+0xXMZjgjGZKVtpIh
FZ2Vfn1MBYqlo109xRylt829R/28c6UxdhVMfhtmWS2/smFYFTMOLKX8R4SNtwbTnZbPrXcvNOPC
9jAg2dwH/abg8s88kI6pvGp56rYBjCOavbMCTDPkrsxsR+MQo+s+GNsVbgxnTCf04FREeRY0ncgF
yP5694xL6A1HdAJY7k5uvaonk2J8wmlhZMYY+8gfCfJdvrGkrXDjmGuxwhLUEVgOTq44Jr74sHSb
s4yYNQNbuYER3EQUIHOzYlG19gGni04sG5yGBb4C86jhw/VbQXx1vL3nvr0gDl/0uYLg24TWuIdl
9lksXso+qN9J+39+8eTU8xliTUCxX4X7L1IlIcAc2t4LrtxbykCFSzedegX/dho2m+tN24ZFshO7
e8joau3cGm5qogEsb9n8dD68HP53wrrpQFUVCTvQQzHBLM06VzrB9TfHHZzV7Kt/vGiI9LyoWtHX
Yv4W2GAJa0Q3z8fb9d3BmXPQ9VhL+ub6V3CPJOt0IsCyMp3CxG21ugUZLvvjMLq8QilHAJpJ26tJ
6dbFPf21Jzurb3JrQNsX5Oj4gve8wMGnAsqhA5tGUsDGBIUdY7xMrqowWZEp8oudLg0E5VLexfD6
t6y7mhbAysLuZJRF0JvxmK70GjE3JjoPy6fsFzUmslfcwZXXbKakFMPnR9f+Rb0QDz1e5SXJcZqW
nsvTai+bf/6bOx39QGseozZgNT1eGitXOO83BeeZFpsbBttX+NLJuheohMinS81boTLmHsnBnw3N
rW5BGbSkjZaDFZwMYwM6eUlNoap1kkz7QPOdM41JgvqIGHTd95+rmaWQa2D6VbUzgVrLNekX1ubq
QxYaFpQs+IgEs7B2uXcdyDs6I9h5YLoLwxnZp7NPTaII3nNUm72alcoAoceUK37I+0b8pW0SA/b2
AddqzNBQP6PKamPWebzgnkyEtRvlL54RXAcsOvk3v+3AuDm9whaHaizeQDZdJtH6fhA6OC6nTw2q
l85BDv9yyqW/wFdh40WlUoIJlCOl7J+wjZwmK7G2wL/sbEUQyN3OAdY4Kpz6hZGf3oEUklK5dTg0
NWbXwOkwIpJ0k+//O8cuCFZm2DDdgRssops6DIasq0akPXEiE/mxHl9kiSNu6b4evo3e9uKrXC4L
8tgFhrhyYhmxfbD4J50E7YmdRpfi/sOkM8WKvzYsI7t4YM4iBd5BMX0hEpBtAwzn8QfdQgWlI3+C
velRzItuYPihF1tMzEtTdFwPMmfNcW3oYUBnxCHDFOFn5KIkyBtn2bkKfgA6OChxbc9MGVN7jSJV
8MnzEr6AkiHhp493Tyj9dTThtA2Ekrd66DBy56gpSkbMG3stRQENj062EEswfwnIaOs0eg1G1z5T
haolceYBf263cg6FmWogJZ9v4/W7v7U8hrdwstRkFsxN0Lb9ATOo5oHt8kmabJRFXYTnHDNODe4l
MZz6SNvnab1hsaH9cVIBUqi4kHgcFcFGC9KSVu13qkEfniAoew2U3iarO10aO2AjH7z52TRwQGTL
NK1M7Kss9hBUtkHqcne/wljmtJXnOCypw4FfReYXxEnu/FgtrxpbszkrkExddwX3Q6rizK4TF0gD
FclYnTdhUKoSIVgXycqmv/zJmqEITtr5EqE+hmjo2FKnFP/mVA3Y4t40IxIQ5XgMIw85T4Wbl39N
VBnvIaVZH6F/Hw+4gagAdagy/Cjucf2W37CUXE9YZ2CbFDgz1AcDRNQmlNv7/SOWkqCg0nmaDl7N
07DMOzoGsdC+rvXZX9kTGupJWcdViil4KXNuzk9YvSZBRn5DybQ7vkZXLQTS4KNT0vlB1fJyvVvE
qgllLLtxVEALbtSlvLyYftyZuxdli2WzzGncwSNoYVSPXhoSkqbIPYR0hhP5iLjLt+0qX5RcEQI+
ql6U1/NwIzqabQxvtGd5rDj6r+iSNVWZuMLLdeCw1eGnE3/iNTCwhKAT4mNqbvVGvD3pr1MOBZ7g
HRY0UAVoseIyZohbBxiJioeAV0QqMAVRchXklgnIEZgf2YllM0ZUkKAPFAGOSWGzt1j09hkICUHv
GVDOe2FleM6BnqcmpyKOYqmTqqBBWwcAIqBP/61JyAwAtRSKXk9Bg8zSdhRLJNLzpqw82nx9aLPA
XAHBGk/jl38RopyZdFAU5k2v5guY5LAhwdJKoU615XIxfawU/QIinQGD15V3ISIQxjbSbFsWdZtw
xxVRhelEQ5YP0wy+AZF97Lje26a/3FB90TA9uoiqRdgLM7TDXuaNTA2fpXlWJeY09Totj5Xs/AS8
MJLXA1E+vUGCj8AV8OB2xelWNr5Oi8Tcp9Jz5GEXxi37lRaKUzWjeTOBSWrwlhVcCgE+bCASl0Xz
nKhh4tbHOj8ev/eh453Sz1AEq1rviey1l1mTNZkPb8arHakvwTMn4ybWy6sq4rhdhYrf++7GpujZ
x6+u1ea2/DDydfDLy6zO1hD6txSoreWV337WMIZ3coRAvBm+mPYQtjkdNpjwb7pzj9AMZSzN3w2i
/w0lantjEZ1sU+6fHb5b7g/r956CiuQDLOhMmPSB0NMc36bJGhm1PEytkJz1czDVaI/s7Xjvhjnu
KYfPvakBv5ziwjBFVcdebu32xNNKD1ORpuHICUFS9zzgaIS1SzlnvevDmJDqVKKSpi5BZNmRuH5M
oygqq5KqPZGR0GHi5JEKW6VdhaY60g5PT+aCQ7/om1nUORcQZc3DTfDoWEbsKZsI+ubSbYMZFA5a
RLc3060Y26xbleJgcuDOfsEBBUqIhyb15bK4tb7glA9pMmru/yxHEzwyJxYn2ooOH2fBA5wHIPJt
ThlccsEf7PAZYj7KdV3HMvMYVpfb2sQroedgNXc21x1t16KOYdDnyvBcLPznCcblDPI6jR5OwwQG
pnMRXGd5kXIx4VuqHdOtY5G9BGTNCiKTtOu3pMucVec8alIUPvEWFyOhLJIhi0Kt2Z02yGO/HHnF
y5g1xCbDGk9ONqs6dfzKPgyrK2ZrYb4peLTXprgBQhD9cEfEmZtouk+zH4qefcYw1qrScFXyGsxv
9ae9mI+fV1oMkUH6TEm5fjUVwGSAKAMEKUVwfMkcYWzhn+u1MaqAqEjeteQuQA1XmogkNvFS6lNQ
QPdk6M4UipvFekPAKy4nTtHv09VbQWd5EBk24zr6jsqtGrVBA4AW6Im+zAEoaly5D/vvoKOVpPu5
tNv8saDTJpdZEpqaBNlJT0QP6T9o9ucSN7cP2aZl6XdQU7495kxp/UIvjbmBMiGKpAMT4Lt+bbxL
2cuI1yep0NY9L9Wa3tSHdNK341buO6Is4r2+JETlaJWBrNgFvpVqg7kkc6MZ+bNd1yPNA5wWtaol
sfchQt6Q1Kfqh9S/JCIZBThX7UZxNEinXV4IEng6b3G3LOijiO1ParGmfFxl7uI3qZZBEnqcG7Tr
RURG0FLk6WXuIULYqgyWXW856B//RyzOysEtLk+hnFjjHQu5DaNiwdqTaQkCJ1UdTBAZX/IKkQvl
lBt5SgMd1VMw1yEBQlWkY6UEemc5hL+ncy9Vj9xGZXjObIvIEWjU3vv2Q1UZKVCOIhtB2EmwpPsw
skO/DZIJm0KlPCezqY7h4704gk0HNjXI7XLc+pTK0DWDgjvyZ+ikCCd9bPcUyFLpVyS+ym7JLaLl
U7IxLhV/PauJX3OwQsvxMRPoXY/8Ysl5h8Jx8WxJzhKhINgHbIJmRpQAkVilO3JByuMDiRp0nnDE
7uUijBAgZYFWmZ/RNcn8pmTPIjaQ3wWvV7x3s8DX2DClJ2s6YGAxnbdvczNwxb6npqvkvJ9hBcvQ
8aWglwiFNSIVMk4+huc2hYfyodQPQ2WcJJ2FpFQMPikDF6Chgr0L+RGsmOY6MYbvvSUV2cC0SvmQ
9cMz7Gzh/r7upKdCec6DnazlOzjfjvMFPRe25JHfx0U9gzopetVUzrrZ9cg4dcF4gqxW+bVvZn8x
zODnTag1JuO+ZMWZUFagOmHTI2bqSwwR56/CqoqSuD/UaBJXUwmUbTk05NS82n28Nsfu+vw+eqNg
VGyjazelIwlBxIgo4o6O5UcNOWg4rm2PrMUHf4h/w0p9H1ERtuL+ncZXv8BjJ3AGjAKm4eTIRfjJ
FPTgPqpEJ6QtCHwKkk+3nojjNiEeD4961SeS4Q6PcqSWrPCXz94r2Yd7vM+2TNGDTUsFfMj6w5ac
x10978YHbRu7PNODJnizCGHVym+mFG4pmeWFBZBwv7QZh65Sp6SmQpsvldj0WjMfbk8Z5spPILnd
kE94BJENKuwjL5b/RhEuwa/60LUS7d5s1xeUDtRRaF89MDVioEILLDpyFadwfmAfdNAxOLrhADvh
mNwhH/ghqirhd6v6GsBB5YmWNYyBX5VRsZyXFXNuajSq21d8P3m0QKaFeXNhoGjwFhGwXJDAQE2A
KvDiSN2Yy/dWCyA36NH1zFNRILh76n8kJn5RU4QFneteeVoYLdnLaGRi0LOPbwQdPWXQSWjov6Cs
vp85ooP6uOK7W02bQa8LBgRl5u1lPeUNMvpNeZnbn9Y6V/ztdwpIL3fkreTfG8ghgAb+3gV5JXDq
gaWPCEAS5OLoiW/w6Jct8qOjQ/mhjioz7GwzeTN8VZPu4Ts/diQKoPjeqjVO6VgtPciBojzkCrl/
awaNydc1cwtht4PYvU5lsfDU8RuwPecppG3dK3x5s+EQlpOXYKagcjc7P1JjOzBxbFOS0pTGaMPm
RxtZeEuNDPKCO83QVPYeofbgnCSnc3JfPDA34D4JfNRxT+VR7gYFO0MX98BgcH4nUK3XMkx3NpoP
blzo1+etDVppngR1hkHQ2c4IbXD0QufJH6fmkGLRGSlC9DkT3ICzeaBep3IshbzXWLKflbUOLN6J
nn0VD98/jhieEUgbLdDSuiqACYgr4kf/W+sazjAePJZ+gPHeNET5KWSRYSEqvgJ+bzzNo8OtM7aM
7AZT3KVknuwbp3CEVTYq33zDIVIASlI1HoPRmfjEeMWeLHqICzg17NELqmsgAcsTQzmJ+rolfbOy
COjwdIXt2Vs3iCy41dkB3dUaM5/+3Sr1gD854/TWTc+FCWdgBEdUyzcv6ld4zGszvhX2upZWqTDe
Xy9/vkszQGW9XnLEX4iQc4dhpjrjtiQgIhFwT8oby2g1uEGSpM+KBXxVrJvm/6PlStub5d5OarF6
UATKQ3L7SaAzO9nvq3tBWzdFuUNTAKv+ZUCL8GvilIE2AaEQGsIvGSNYIekS+CVYZyTvCdE4yKh2
YSoHXPu0MY9SCH5z84G0FxH3vc1hx1r5E1tBHtSouxNVOu9bzNSe4EvWq0ZBT19eSNSJTqs/jFLQ
tpUmfE5acK/8xZqltV99McNAC9JPgHZqfRSyvnoRjkOY8kLDKEOICvC3+qdV5k5cUFndmcpxj8ul
hXzp62DKkHOFSggxa4Z6ghYr+HdfeHMAzWB4FWKR2y1nNQS+IZuFUtQFfL2X9tGgvREQUxwHeb8g
NyIJ9HUx3DFHgoKAAJqEMufBIZWMjQnERNgCcWBecL0CtSvK0qz6T3I0f+2FDKWPEXBUfhVNPEC5
i89bstv387KrcCI9uxLch0ULkwxIFdg+uwV6OnsLwo01MlBWtBkVFaa97XZf6oeaqu/P1EFrOrie
/Ic5Sp1nt6O2ZZY46hr6ExUyE9kJo3gcDxuI/3OH25W4XVkSJBXpGjbWJcZvPMvvn96DW1RAQvPX
DsX07IMuHEFAymkC5QGvlQl1YWJf5JR/aeie8bv5b31Ll7OB9k6L2+AZEe/OGasQBmx9G+sbkG2p
mzJb+bG+hMg1RJACa5rptGVSNESfIwhym9m23gig3sIZBBp6tBo/iJzY0t/TkJ2MY6349RKA3diL
M8JmNl+FblIjJdRIE8irvr3eldTvjx5MqX5i37S4Stm9UoflxwkmVgpQY1lbVOVDslvVaKRp453t
DHkPJVp190OcP6TH7cRxGmRKRW5kuMiUVuPpWfK3BDtntUAwusOFdjRJFO0mIvtZpgO3Fr/8W5Zl
Yz+jLixAct0pDcFh9KpAIVrLRGihGntgh7OReK8vXX12BCkAOme9YvAk4pmnTbQwY6IZz+HfxKJd
1ty9qXhJ5o/taI3weebZgcUklaj1BkPdLR3jtUhLRkpglRbKQ0ZbxpA8UJLjS1PrGQlAmaLu/EJ7
vvLrZ8F5qpdksMo7JDuInsZxvPFlUoOnRTmUxooxp+85WauiJakdwAbTS+zF/NttUUwPpPKV4m+q
a0Uit24vlFSO1dl9bZCHMqEeghok5C1JjCBuQg/PhvPXEmAJ1dyr5u/K9KX1IMvvhcm6TVenhtAx
pzuFPcFGrtHlBylZ7uhY2G+1ZMIgiO3J4DjsAYqVqWQmYWytmzWS6Qfn32qarSXZ0LAY8lqCukVb
iIJ7gCI7m8tJUSpXA/w9e8fY5U09VUiWA5gOIefit4oK0FtYwwxOJK9qjxGygG88I7EB7MjFpxVo
0c3bykbUr2rozJwOQbqDWfLceD9cuwx2AZI3sTucwvmgYyl9Mc8hq7EKC9eYcy7lAMoqu0c8zRRl
8bKbhUHfx7Qpd7R4VGten13oiLZIOViLgTRAOge/urfWECqyrDqHIFgPVSI2Jks+Cu2uW4WwiXrI
xT0GpZzXLJ9Y+BZSbdG1jmQyHCRyXg4zjUSn3YZEofBLwZKAtcDVNtSeGPkDwEn8CG3Zbvc0vyOl
2t9acC60YKW4rArLv0Qw6v7Wr71hLJlNEBy6aZZl0xDfy86N+Sb512z3vrAr1Z/ymzzeW+k8mojT
9ZQFXEA8hBTNN5ciIMEHr/fL/yZy3t+sJc/7EtEI+sJiEd6qfHkdEWYChVMviEypbyUqeviBTH5a
+Veq7sDTT7jYwii4QAyk3GCXfDn/HQjSbh3RoRGOb+ScBeXRqY2xN1Z9omzt5ynNEvt7VhyI9ydf
zVNxHWnQTY3oPulcpUYmW8umVFmE3J47zM6OVRZAj3UWfKEzxjiXstcfbkMi2A2rHi1atHjOcOZj
HcJMNRO5WX3OS9GsBHnGBQwb6jwmFEJriHkYNMfhGX1BaKar8r02QCH8HGzU+a9BbhSfIl0nIhYr
Mv50BFOlYhawhqnYzO/vl7UYg7Y4ywBpybNnDPLbC9s9wq5xbdJ0vjS+6AdYFGLBJXHGscWnWXmS
gybnTZCohTRIt9eYFuMLF2Mm7Yx9zfzzXryXWXN5js9x8OroH7jpDeJU5L9GZckvu2BbXpP41+qq
pG78X8qLMgM8vRicgpOXVFte3uX1lzwYibSBw/16e0NQBlIwRuuJPoyjvt0483Zw2pePWs7x1nKT
BGGbxb1fmA/+CmmAWvTqHc5Q9NEZKbRszf+pUgiAauzAPCrl8TV7Ds9Z9IrJ6DqfXrokAonWOcuC
4vcwZrsTbLkRFQweIpJYK1rtV3HEuAMkDnd46udsTUqJkAfFbx9MdIKMQvTiEMsHYpV3PzkQbr8s
84YitVqfDyeYVNUebQiqmPyE7/FmAZWaP+GCvLOzVBuWLtjR++oOLRo8RCNC9Dw3NFyr24F2TVdI
EndiZtz1HSmMJ2dbn1J4nKtCjlpntX9HFnHJGAIn/VlRU/8+6RtDJu0agP9rKROw/FadjmQC6BqC
1BMa70bz2tqQ9pdoKHv0xzN7ylThlIIBrDn1TIf6Wn6DPfSaMK16IocFlUZFpFajtKXUEVp6PCGR
olN9GjUYUfRBIw9PxixOaciu/yvVIOw76Xxy8RGyqOO2BRxQGnHIvlzUuLsAQA+UOX+TMD+UOfrj
r4GXR7Dk8uUJm6CQL7jXG42FeLAF3+7ZgNaM/VfFj56YjMpyQd3Psg0DC40Bm5pta4hga3dIKf9x
1tCHFmNtEOZfoDenn5tEcFpCdduWryv7hdrVx67gQSZhT7cm2yiE2bg2qdFReq/0nk0aNEqC7P+9
Plg3E3oyKphpJGoAMlP42jkQzILJvwOPQuM49yTKKUcCP4iReUOEjZgabfvuPSC4btEnbBxg5ITk
+1QgEevJ8+2/MvKvLhm1/tUmug7qnp8jj1jGzDat/TA8pU1bcwUZvY9qmi1W9DsQgsHqo4WxdDKl
CfQOfah5p3MUruIcVqwKN6uPU66H90JfWl89I+My6kHNSpE1V+nTzUIOuAi28tq+VtGwmxgDZwt3
LXxXbnpkr3wQrKlcOzdGeJZ3H3ZJ2FTKT+tECvA0OSPeWJAiybMB/5O5IJehcKJ8koCQWFc8nWtC
ssNydijZmyZcgj9G/nTprYXbSnnxxqjJ0nyRFQt8SjjqgNmj7JQcWHAAPESyUI9AUxAwhSPspkxX
AFy8YPIzTV3InTV8b1o7l8Y0mRhCwGovEHvjP/utoEfHFbXy1WiU7dNIyA/gpuYrzPb9gOwU4O1q
rXNwhkWO8HnHs0wmPAkQNcdzfo7cVB920vbVEL9TfXjDn0kRVA7WuvQeQh0JiBtznReGjkRz47Vt
GkLJnEzHOIHlaAaKKeF8JOMNNVJ6e12gpz2PU9L+Pi1xrNwdb97iquV6tmDXXxsEYoCBVgdbDw+w
2iUcE874knf6krx2rTDGbi0Q/S4V3sDqIdD7UhEhPfDC2HuxhUMazD0byLDBmEcDPdLhCX7XOiiZ
IEdZn913PnaRFXe5K3J+l2lHnnzCHEKySVfy6JZlfFgGVwvHJ+qi506s8mhR0ijWFbfU1kPOTO9t
bBmL6E6fTVBEY6v4iQsFruG23EDLzmSjN3r6zFcyGv5V0NvHztTFU9MBFnW6uBmvJomwQ/2NGs/o
imH0/ngfY7ZeTl9ukzvYhfQdIh/+i98ANRyTOAIz6FcOMZU3mxRVNmaRUgQ4FevpqHS0JsVjGCWI
y6I4qzAORWt+bBDO1b2hN7I4J880DGuhjwXNMcpYZUCkVUNvpYqewT1cYMuqU/KCxnR9kYMBr3za
teHFcC2r3ZpFDbb5VpoIgLsYf/oQLSvUr4oKXu5hU2VgTt/GKL8k1WBQB1w/qA0OP9P/ExcOuWvY
3Cglapd26JVJSGys6fxSF4got4FHJwzzoRlUzr8jDDHfThWo0tPcv50myglvu4qPdwyVR4SVronl
p92N8qscxNC8x6Te+mIko9gRHbBQSja8aijb9FAUTASpLX+KgdVpZIKmKVwYGoXJTrCnKCgqtumw
G1Yihtl+JUQ3gYkQzyNOJGrFUO7iBnQcx5D1ur4Qru/nQ7tL39WpFekFtnrkrlY7GFET6PSCq023
WtcIxaSZuXX9OxwciMfG9JWpcQrfNxGc8Cd9dPvYGbDCl22+tqE/OKWBisnPyZ3FudDii4sGR//p
rhpNrr5eOaUo7vlo9kRQamhfAf5xCBJIbeSFff17+ShCKzVBClJylSD7LKpQaVBYtLggRNoXxVSh
Q3CXo2I1dif4gsIHBdgyPFCt8xwFiH0qLkRF1kjc5fT63dVruFweFFwDfRn/utDi2+2DJZlxyxfa
WhY8c4XB1evXedplg0t+T0s+f3XW+0I1oInnPaxzbq75YGtXUTFOWIpSeekYj742ZoXFTzOql+80
d4gC7VK5LtX/Ytx9BSJ0Du0qfD+b9NhhI8zAkqUgAMJvBVAVETtuP0WoEjSv5bM3jOukPoTCL+a/
ie1LjBEsDICRbE5lNKuIdFooItcCWE5c9GCKHGUxcszNhHB/QFumZO8uivFjFh1OYNAPk90vguMW
4M0qmweL6XZjvkaXW+gChQufQemDxIjNWed+QCQe4/x1gXfrUMvec9ZH16BVvgTRg8HN0t4M1xCL
nxic0X3LTBsCBPZSVv+F/ZoKWL2Ul300WNy1fRiO/I1io0P5LgO3MdEu+9NWoh7QXZHwwfofb57p
zTfRsF7u/+cnrlxENDl+TozPwE0xVVEdm8XIDIAOEGRu9V9Cvdj4yb1CdkFVLXWnl0icMF3ui/Gg
bhvfmur/iUCTjjKYsmczm7Ycvn2lXRYT8qQP2R3gzoEdt8yVYW47W+IEuweKnC7BnFLWGIoN9HJP
DJIhsGYnSxxVyS5nognjH6bfwzYhKgAqw47MWCNX5WnB86kyTpuRCR+E/F6Eq3p7eGFP8JGlykoy
PzXjfAiolUFHA3HU6QWllo/F2JIjDcl+unxHg95Bu8cQ4w8YYV9q7c+VPmMguQtozmZEJzuqDOVC
bFGud1MoohM3xx/4UhtgrDmcjfac0sxU+oCXwu3cWxoRQMD8q0Zu0xCS75e7caDCorNHdLb3x2rE
wUXDjZ3lhz0wavdUgklRAzA18qK3Bj0Qz57oftHvmb4lqUX2Xt1QAk5RvMQYpa/0zsDvVGMtsA/T
+ZiSGXAyYwlzyoCh8afc+VDxYIDXmivCUK5Bcpn0RvHt1RxiIRw9X71sSkuYO9YDlw/0252vXpVc
xjRFooZqLq12M5+g3oImY5wjnC5llG+tRM650hC14aohimH+KMET8TO58e2HDspUcnFNwasL0N+Z
2i7aTu1oKOp7kgnqp/phIMnYJ8ryEYcwN0hASroYFgCfKhz6e3Vxi3NWaS1lTT4ACQVsaIMC+Fe4
LQ7B1SCVxs0X9A/iANwaHL2lPDjDtUcGECXQmoQvroh+tPWJ3DjVGIahn8mf3o7TanWffeRuRp1Y
ZhjwNn7AiGAQ3xb8rhiDG1xaKjTvVVGOtRig3PWOBvYpGOX9ds0IA4qk0g2Fc8/pN40c/17c9Rec
gp4/t0jR78nDIlnkiletJuAHTmI49v1O5RC2Amj/1tv4B6qERnDcKlUigfseBWz+S02jz48JbIpu
1EStZrf6M9LsFelmaqy4baUXvU/9t0M3ftfvRC8BCYpr6xB5P4xycSTrUHPynmwKkbFFK7wFz20s
A4E+favbvn5uZWHub/lyvhWScJ9JOzz+xpPuuo6SVgFbdL0+zzDPEErjCefVtyJ/zl+3EDSwrXP0
5UwP8IgCeP3b/HHNH8OtQwLs+cVfN3P1N7XyF2YzEtOIHVh1v2I2GZbFTZqQWob/Z0Aa+tM+IwwN
ci1YCywYnvV4puWFrJM9ZGzA+AP/0m3efyXqcVwRBB/o/a4ZClTDkqmw2GWyTkDwEYkpX2NPsfwu
Iz+nBaUt1wBSm/uTDYDcKnN9jLOCIcv96bA2nHo/1lDvGlvcrmE0S+vu5+kW+zJPY8b5bb6Iec9j
q2LgDMoWgbXyP0G9p0082oUai/nEn3Ru9BmcSp3/3aD8pyJGQpG9eLcu0nu2Vw7R1P1kQrlVWcGp
MJ2WPH6HaFKRvgwnHuR5XRr4JyrpTX8xZaG3vFijklAB0dusW6NCNXvYHKPao9mtA+IAHs/zKJ+E
AsmWkl2eBPhQmBsGQJ5wiiwUy9HeGvp47R34Sv1G4uY9Uo7w3RkuxMxFyGNMy7dEcWaSTBQSgFNJ
TgZUe2ki14yIVd5V+YtVSxlwjEPXqFryTapF5SySBLzFGZP4KFbzT7cqjkAnyIZSB0lMYvqdIFfC
yhnjUtrdl2DhIfFhhOjTb4HQ7f4n4TZDfdH0wpqclWr+Qjr9p+XMtII4t6cx6SkwxSqWAsoqzCMu
dP/7ZIn2eUfokTuKOoyPv6KSCVth1J1hN/9xM/5JxrdTUEggxTcyPTRyB/5oA24WLvJcsgU943Dk
CSg3nA75Do57FZa8RkiInIu2E191OhQykjdMFmpdbS9M1B7nZ6X+0zQiMuUsPQ95m2fAGyi6XrgI
uOIJFbWnQLbq1VtpvW/uPe1Qg7N1mH15p2UbmnVnbZvLqtP5uyexq7FgD4hopryyEzN9LNW78DNF
R2cUCRFLt92ZbBrw/P8TjqporHdYG2GrrIeBWxAMYiBByXJF2Kv2LdWfAUKDEubMKs9mHf3Gp19K
O0QD7NkdFNCN9RPabtXr2RMQ+FoAyXGLm5iapw5RZvtdLI1qXep7SpNkZxRRZuBKjgUBW++GZoV9
giNH7I0IUZtEL2FN2JQVHMmHrCBJ353ZBEmCbXvYee5sWEEtMmdOpHrVcnF9sQMybqnIxmkuWK5t
yd5tJEiq9Wi2AMfyVbdg81t9QseyHVOyOEQbTi/ads9rIqwjeA1Ee/iflKhnVqpTUpcg4r6lZeRf
cmNoom4pUtkrJEHxS7UyJyMgSFiiCmEU9KnrBu4qORyo0ulZMtkErnnPEEJCx+qBm8KhFPlLGsSc
VKrvJYukihpHoH53j0q2x9uT9WuQUIJSYYoTDRYQ6yIrQAo5oix1dBfktXNwKp2d8LRsxNzRPr1h
zE5yrObdXGPNKjI+GJginCo0WzVdPtTq7cNqokjmC3FEJqx3+oZEqWyaDVIHO5ChsL4nA9JEfszy
svsp913v0+FbB2N6U765SBHmnBIjacEsFR92A8eK/gceuKPaDs5OKULiRCNdbvsmyiv7ZPKe4iE2
TpKgdJQDe6Ybfjpt39fsk7FLFvpidySWSE8XEpFUCoYEnyFJ8ryso1xZvZYRTF21O+GhG8qu/DM8
FvFQPx7l50GUOlIUtJ1JNSggks4+ProKUmaJp1/QJ70j5+Ga9uoTVXZzlKQWWZZZ0TFgi4TawQTN
vLbiYjxjtSt0Ndp7y3twFAGc7upCPB7bBJ40DeWeToQ80BNY7Xq4wmtktA3/1VroiCnn9wyalu9o
LBBwLpqYB/v3RXKH3v0fus3C+wVZawgSFbdcSV6iKSJ+AJkZhQiIbEhjD0p+xxzmYxjIcVq3j7T1
w8gdF4TOAj8mOuUREiuBdAz1aZOZhcrAZsTcsksWK+XGj154LMs6atHj+xXL5Uz5ZKq7pNe7bKFw
jXA3CI1Q4vrM6iT8nC9Ds8HghK2ZZrzxs/Oybv7hiqB0KxjX96PiQJNVvUPcKI9NpRDuna3Ck7Ki
nDK6l3bcr2ArifYapev1f9L7L+Hp8nTQQBi5W/y0zZW94zKBNvyL5p8HVzG0cYN/PkksI0nXdiVD
RNeOZVthEi/zbGI5gMuFU0AhWQPCUQawLRtf8WcVb4Jw5Nx74EogIZrnJHOQOu6cUeu3J95jrcfo
x3fuxEf2xwThisVyr3Ffg7Q02I0MfiZ51vD2p0J4pyrFperMX5PJS9yhrHqW2P5Tyjncy0eQ7+dV
uyWT/znfVBffsbffN9x6+r1Re4njx4Ok6VIeNP23HPZwu5ZtYN+58qNWU3Fk5LOOhjiN/ezcKTBO
FQBIoWyfB5nX8cGoHVfBeHd8OIpOkmdyeoF/Kei/G1M98JLIa+aXExYxqg+MIVFTH7/zongCuL8R
EOAoZyg1wDFvq51VzImsX098fawdl6pN7YV5bX1BaoPIksVNBqeOxd81B/ZHfn63uocHtlr8Mmvd
BQsUYbIO97QipYZnb+edZuGeNG2yWSKCBSKjg33YvxCpR8p0Kn8VI4ypZ37EbuLA3JwAaoFH+hdC
neaHOyR85Rgs+KZUONotA9BDl3NOEFoKvJJRZOs1hIbDDCv6kux+WXFatY5EbfhEyLTS2zz35puI
0nT5Qup7aq/4fEGycNVm6trcJMAaamIWf9/+FpzMMOOabYm/F5nxogmBfWPZoybPJbZo6mediH7p
OUUGv+2ITicA1TH1RWQPzf+kmdavGV8vC+4e9AmnNB3jw1NG1XEZ4JBYl+8uG9Yh2nW4fpjv/HuZ
8cgIcEv1TNDYzuHrsQT+zpeWdViDFrPlT32ReShwS7hlWjaphMB6RY9ELlF8ViHlga2ndzYPCahH
jNo9KqS6gqhXOY+RyBoLrNoR+l4LXwowaYehkYGlhNyTknwsIk+A9GV+NDWg53AOscN1t3A/gBz1
3/KNv46Z26ypcuDmpE72PKc4m0OGlH6DR6wlT+gT3NSv6zaLfpBFTgNJj8lZ2QF1Wr//32dmy1Z3
6ZrPRQ5qfa0IW0Hkk3IcvksOm4Bdkc/NTeBLANjwLVaqcQqLGGdal5FyYJJiguSCWPdjf7OjMo9r
YH8opcVVSwE2h+DcXhhoS7rSxuDrL+r7cznmgoW36nqWweqL9zgbtgLkCy9y9Rd/GF0NromUDE9I
0Sy1jivXMksNB77Qterkx1GsWPJprj8Vqmgmt9LtGAO6qKh+LcI71cwHzehozuwNbJf7mJiNXctS
m4KTmxT5J48p08LrGXZs96zkStis1jdeFmNJsgRhp7wHjWoCa3ejz/Km+OTjy9f9F0MjWMG8t8tO
OLw3iDh3D16tLuuVD5Wx88e8BUkhZ4/NGGjfRgBvaDxpMpgpy0wp+iyJie+cOTUpKA0PCiDxm1BA
WK7KMlxmsSYej16jqA7BxBF/fWQoVd2XWj+o3kpAo9im0rKARK9MXCSJhlHO1nTfzKusH7ySJxe/
NYTBcldqkBURf3dBZ6NF+x9YPz6EEoo7xKFw5mJ9WhOI4mEXD7KjCpe4MjFTpBevHaHxVmXouKXa
tRViv5woySUsTWKoMLhr2SNIHmTe0f07/0aJBVtiI5urOS3FKGy7MLv3CfXj8wGtAsjSyouwNI4z
fw+9g8d4uAgGJS0G9ZWBmvqNwv0keII3nD3ZytBlznLT9u789UgnrlkhJiR4JQXJq9IwQGVWIZyv
4A80mkBrznpmkYTsdElF03ULeaODnnMpuJK5xohxqEDqRDpF4k+xkU6/mUXFGfa0a6PY3YrOn6Vp
JU/jVq9/Zgkw1fsIZ8Tw09zrswB2lSmEwx2lTsCeHYHzwBDfH2X2tw0Vp6z3KSRKLfSqndvwenOj
/OEaov6Q4S2r4Jxln+0tyL7sRiXTpO9nEANr//w0KZONgB6mck8ufhocMLleLSwYHs8zNbgCq6fU
ye/F9Z2VpOKoraP3VEnW2kXo9Gm2sbpDJiuQ7tWlvg1XY9K3FQhC0k/1WwxNvcUGSkE/oT03gjw3
GvL6zTb0k7A5qclhoB8gP+dc7kXCuLwZ3KZDquiY83raqbko37Aggzmqc8lc/aRnG0iQFSurwHMx
2pl5YV6KJaJFfeszIx3utaw83se8NWK0PsN3cccjcj9mfx/lf8RXF2geHN38rFcn3g+l0g9gu5oI
PgTIZfS7t8SPIqdERp/RW32UXXKi02EUvCw3bGSOCDAd8ZuKoj7EPDRbYqq2K5Qpa2I42UWpMVhi
mUZnGUak1j9XATKyZ3c3nhWyP8FBL9l8ssFcYyKwZYgVKu7aKB1lEQsnpGOo9FUitk2RoA0VH5/T
Vga12hqo3VbwNfeOrBYbWbID6k5dFiWxiXhbn5zrBwwxGhWtC6/FA+OALh6m05y4HapOW2PWK9HH
1X7q2OaqHEbJv4rAy4LCRsZrmvOnM3GeOddswvn38MjhD+CKfwjwNHfg97YmNmUKxZuEtxg6uIey
NwTDl1KqNhDwrIAL3YP9lFjAyr7ZbGIpLjNeD9kagVIPx9/7f20DwwkMfzrL52/C439qY29uc/k1
yknQzTCqf47beztyVihgcWInEhbu0KxtoAj5lKt/4DudzumXPah661zhMcjw8vQCk6u5dh5wC0Xz
KdtIgjl0BkYUlGhkRvH588km6COviUVrtLZEPE1aqr+p6dRJsEA/d4vzQqyX0wllyqDWflxlG/CU
JHC1SEvVmG4uKTrrMbSelNdR+YgAoZVqB7WEwyt3EmqebJ89StPk4uqFRfEpWEYk8QaIwqwovPJO
9BzA8m+KonWrTN0XATypRIZ9kXFhHmKuL2UkRJk40okvPXb6zHOvGpxAPbvv042GZRJPewdJwRzA
GlaPEnfQS+fRCTQnyicmWy5xfhAlURqy7XpWIxiryaS7pVALQX1uwESHhEXAGl0vIfKOOxbYgZbe
7ySy6k8yVru0f10pmOeJIP7h+WnRcEiMwVMBEvPEepRoUsuyGN9+2hFmrQWDgwIsxveUcJTGglUh
sZfG+hP8BeNhOZLkNYgcrpoXiJ3FM5iKLU1SKoS+Z2vCyGGL9usZsHckfYGNE5nC5s9RElGrP+cy
QDdivN9VEGpL+L/rm2QeFqFfy7auqgzm25140lXllgAhpnXkP5yiwQCA5GmxyXiCq61m/FXjS6GA
RYN1u487ScbQQ6Xz0m3uzZ8FUt+J+fFlCZLa68YauDp2NTejFA7Tbm82R+QihCtaph6MCA1I2Jse
bIBi1I/D4vla9R1IIJkZMZo6l6b5lxJ/GjTN7/h2ARP8iKYd1y7vtFxb/6kXwiiWbtj1GAuyxeT7
fOxNVayxpxcLShxmwu4KpB2wg2w1VQm9CO2MHzTgVQO/Wq4Vl9nXSv4tpb6rj7plY8/KvyFZPnvy
ha23ajs887SBCt9j3spGCFsP7PjchVc4s5kr8W4c+HqqVjK3ZEywccit32QvLxbCAuIgBIUKUXE+
MRcHSp5hFbaTdlSq6wyOcbU549Ukz4IdQbMtet9OHr7ONcx+dJWXwFXhVg6sSFfNhUTv6VtFhU2+
bZX7bFFy9MMAywfXH9BxyB8QqPQ/ITB7GLubk1JFEJMtfntcRGRCpzgiIplV1zTtoKYAMzgEWuf6
zLdKjyiWXRIrrNnGgP2cI05BGPazxUhlFDegfAh6ROG0xveqHrns7ux03FkZJwRL0lrbxItcVIfX
UbTGoP+pszQ5u3mECIJD+WNmSCrK0MsVCtCPMy9id1U9D/JPjLx4oahRrMUjGjCantjGjV14qWVM
hOaI4qB1EbSrueUdDNXxJw6PRCS7j7tHxNCCf+Hp3XxSZxRPh9obNTBCxS/pmZ7OrBzHRqoCHy6H
4XKvTFwx4DGtPqgjZkAJZokKd4LOo6xL9C84elMNRMJTWo/tzzCBAmzjGGtC40ZfJ3kbYavrcvMR
kKloXVFv7PBfpLA5/ERIUBuWb8011L2lOtu/AJYfWE6W7XCnRe+w1kACx4iyZZ3TzILj4lRlsXym
QLrp6BqjMb6k+3ZtLNJzWZkQUWmCUl0PypEw87FUtNnisyFeOYAVFe3CS0v5j3SF1yY/Xt8MaBgO
YbUHHbUbyJ1c0RPMD2vTUhGcs2XNON1iQdHzMkn48dyLEnDFwpZlUCN7j8sJgVjZ0W0+gARt0jq8
CElpt7h6RB3xmAi19KL05UDqfMuV+0W/T/UORn3W6RpDbmrQeO/jD/kJhS/bbZaFY27dATQAHknA
vJ9TKs6fhC+Bb3uITwLx3Xi1CX6JmefW00nXxMcun9fH234m6+Ll+oDfbYB/kDvndEvYoKyGb2/a
Pn9QyJG4xs/3AaPiKSuae8C3ye5LfkZ8FVwu79nISgAGz5zVH143hG18uvvB7pr9V953bCcNCtry
dwi6x1/AbzqyEiyuzvnFZj2ucoR6bMNVYAX4Hrd4H60UtuU6oeNxXbT1LtnazaYTkoCbYtqzlbSq
ZDET9CUKg4jrbjCpnpeUpxf3xKy7ELaJmDEM8YCG4K82hK135uag/O4SuEIZLGjGBehkXHTVtVm7
iNNItgOfnHKf6qPqh5yteRew9mNS6t10iaafHmAohAnhmoMgu+72SoZncj49QhOoNL1yBm46ax2t
Qe42c5zAQuTJYSTYQGOD/dNbw0qPHNKVkhYksQyCkmK/A8sg55afwujF4ACTdBhQoE1IMrh7bYsM
oqRtrDdy2e49FVAKY8RF2QTivzDekkznHjsooDYITj9jFkaqsjNHT+p222ZNHV/kKJ8aFUJbFj8Z
H6lrwxXR3DJ75h5CpwPlC0atuKuh+op6gIXHQ62d/oRQo8li/SF+NimLhT8MK1T2LDJha5RO+N/W
OgPYFz0FnTPdKk5cL4IVdqcM6+rY2aGsg3aHcMQ67QI752zOAqrllHvEDrjPH7g6hzCkzf+Cb+hI
pA7R4JdD9WoWCDl6NVoHPtW6L69V4ECgZAEGs+mQo5MRj9STxNEhtMvr1ieSJdvnPv6v9A8sQhAQ
qMp12b2jXUs1tk1hzS1a/eGM12vncw5bAelLv12rK1uVBk4iysusZsG7H3LJHtJTydIbIBt3h613
EN9cIp3FgEk07hFskEO4UKKtjpIejnF6xQ3hm884/WOGV+RnCPKUciMcrQs4/F7u5l6fGsI/nGHM
2q0J8UBYyHcNYvyKAwBqVYp7krc0Pb2mdWd4Hd7SVyHc6g4m/q2o/7RTh7e0FZZW9PedqnDoSVVb
RcUMfaZqzv9+31Fq/6TxV/sgf0Pbg1CO347hST04kJ3cMdCwb92uDPXrvB3kaS8r7tA32nzB/XKN
+RFMZiGLjQYnkIN4LACexMDqUUGZwhIwXYC2MbVZ1BXezGywVS1oLtFJZo8IF2ow7QYnXnxL+iEa
mUe8m+1RFAMn7R5xjfJ8Zl0fCil3VwIf6CqWL3F+zDHQIQqenrX127qG50JAUQb67ABROub0dioq
eyK6PjBvpp4bdOPbr17/oB4bwsldLauxYhhV0kduJUkgKN+u5QsRwN89F5kvytpSDTDLY+XMaraD
aK2Kynbinhqr5r+nJ9csqIq63DVAdsOg45IHaffT40gANWqFgM9RURj7R01NL75inlgi8CJLy7Up
QGfsx0wTHwSp8oUrg1oMHcmKr8TjKQymyp2gZaBk5ufCoBxQE3MVLYOxg9mtk++PramCeo9tcVOy
7sPnaZUWQvssbQc2nZ9ESg+rtcVikYrqTZ5J4sUuU78BzcxinXr1ZmQYfa1+lf3tWpdgO/g0SmId
miYk4kQQaN8n/xMEiVu0if2iwsqn18fD52DNCW090i8O1jShWCP0egm7Rsl2+vaOoNGV7tGg3yxI
EtjE4jCuTuZ9wQltxo/xjwqK2SXi/4eV3ZVEkDeG4QfzkBLmfs97Z/1rJ7BgzBtL2riKL/63QGRt
q5FwtUOrPJ04Ej6Gckemxccw+7lhOU9+7dY/yEQq/EP4Oth85iBI5XKOgdA4sBeMYzpHGDWG/Swy
90tv72A5WlwVQTh6zFaqfLctQFPJ90UKab833+TdPOJSCJsQTgFXHG37JgLYEdGH6kg72JmtaKVB
k/WJiQLZ5gWIMgpDnEwQdy8CfmK533NUE74Q/iSockkZ3QcB7HZ8pL8GVAgpzamT6MV8rDgCiLtM
lxdoXFgng3n4gjduhvOizGNUwqcDPeeiMCy3cVYe4If5NjAGJPsa43SUe/fs7kJ04GMZid5bf8bC
Wk+dBKpg7zY6Xzx7topGL36KK1fC8PN3jGt83DC2ntbdIysO9OBtkNzs0z+8rXtRRZwGE4s0G+w7
L68xuAjUEQgPmyleEC2h4x7t6iX9VZRrB09ZkYA4VNMjRlPakN7iM+YAv/uE3YkkHwo2HyPtoJ2f
JGlSPoDY03Qg8FiUiQds1Cn2lZ47m1gttEiwlOFCBVz4arV14QRw/CdXSai2wVRvfjTAT59hpAmg
EkPNOzyYHIpffV63+AenFtRQkQHO3VL6GMspQU2tfz1HwVOh8b0OpSCYUfLITsjh5dhLvWOLwSU9
R9QMBoXiMHOsXlJhNLQqB6HI1FgNRgAzMtEkXH0gwJF6wsezH7mdYv2GfgdOchiiNNPRrgrMftKE
cGy4YbNciqjfJau1r7MbGY201REmB25HnkKVTUh6pdmshYQUe+3M0Xc6UmaZIUh0ok8hPW7MckIz
IfO1+I6fi+viQ5p65X4/crd7Ohu+QTsIiNOcEjQF3w1ur41NZVa7fWoQC/0HAteRM11VFCMGd1bJ
q5r2kSEfBh3Vs9OGn3w8I+bUOSs3irFL4INodDnOtpFoLPs50lXjIMV8ruGed74EqeZ+HOZCQukq
HvbG9acPwvMJAcVWsZaVGGPQbnkqlgYSO6Fw2amDt8By3UVta4OPE1hL/uqbr/8rlBpZWYJGniOY
YIKoppIGyvVhwFvQp63UasWj2DA8vlMeSPSN/M+35gtqR9Qf6iNSlTi3yiP1Oc9QunFU8pqF0xbb
hoDZa4HrnCoT2Iza5PYN0JHFnlJ9WCYGF7Z1OtAeJxO0t7hVSgJHAl2iZUFCMjmq0ah/zuA6CUSB
Y3497jMV+AxaNajz9feq5OAT+JsijpXRMXru2scOcai6CdD3zZN+SlI7ZHBxWhQ1JUfOVJBgqIdn
USgBXfOS43gTg5SSa8DwkSRVlJn2IVMCKOxVq32rrmLPTwg46SSmCo1a/QErTpyskHKL8omfkQKB
Wk7hoKhrMyHWQ72QPhj7QxkOVI/bPMqUJuzOWj0/nvKQJk3Bs7a+gxcfceKI6h/TR90U2do+6AGR
e9u67Y6s0sQ8Dx9xwoJgu+S1XB1FjBZjAAnvSSBmTflwUN40iOIESgHNLFXoTKFF9uRdruwjqDUY
StohrPrN5BLwhM20ZbuyvdawJxza+JvwGrxr+/UZPWY8VwPnIMTEbofU2U7uUO+fBJCO6DQusmn/
1vj5MW/ORR0ZNbs9zHYF53eqn+ZyIg/DeWEyJHY96sC9wJO4cVoFf1QYck0n+mgYEDshE5WjRYlT
dm5PU4IW4fgInQaGY2Q+5rwNw6HjJ/FkZS//b6+rZmdwtjQRajSaYTb4KLKm8PjhntCHSwUoBt7O
9/LtVVGObbK8vIbaHdUQ8rs2G/cS0W39kbiCwhonYJ4MRK+jaJ6SNNuSD4d9LJi0HthCvN/V7xad
s8pl2Knp3lZXmsU9lvcK9ClAWnnEeFZRB87LB2fEdGhQoX86rWyVZuAzZFT5NTamFYECVpOkR/9h
ePN/TaXHewE6J0/epCOV9xIzPo9zYPPMU6ba5EYR2b+QuxnnshmxrR7uMMgFv0cbpSdSBWLImi54
T2ZUUVZJTH6UvG01zHUv+aOj5kmGkH/q2cH8pXD1yswumBbzG+oVq6q/AWtd8URLtmtW+FCZwCdd
4gyn3o57LWxZT2usSSKDSTrGnu6d8AoCMjt1aXUKanudxqNvA13U6qy4xO7FZ1AgbAHIJU1a6nYe
0z5zGlmOlFBVDBKewcVq9KD0JIdVTivf5Js72os8FIn4ZS23aRwVYc16t61wezaku0R/qv9CNRto
cvX7yMxjCLjUKDrGKbeWOYJmMFMnAfGfoHw9Q7cgKaY+v028VXBGZASpldP0gkFA+8d5IurHe3h4
QzECJIRw/kBirMzGdpLIETskmvkagfdQC9LHSBpwNNR+5s4hUeky7DPF5HwSH9lcTCZyc0a2i0u2
cJMcP6OGjW8TTeoNrnto22m6Qy0vEGw27VTfNb0g1MGhAe/r7Cn0X2xW5cbALXJbFtuVveuyG0ry
pDQaYmJ0Y7DxSLcZ49rghjz+S5pTHQvVoBU0orLzYJgBovxsjibhMCFjI0fUTJw334PSGEcGrXLh
T68/wkAcEI20hNYib6T7wtAYY3nWvKsngvEuHrozovO2ZdIW7o7OAf27SkcaMY09Ai+HWrhn6+YZ
0eumfzgASXgrGqoxOqW0XePXG3lOFI6GdWerO7U+xNyb3uPihhl2Ne1NZfh9YTjv31flkMsepOwA
SFqicA77jBkTnyoLgCREe89U+XHGJ4EbaV+UUEKUXoG1d23o6IbrXqItlsUySutzmgLrvfgEDio5
G6ggaR0trzNRGImawfuoFzrWEVs3mvsfbjnXnQmzMBITZ2QnFSrIqtpdwAGNaOQl1S9QLwROrmGI
rBTb+k/JJPrh6MjrZmD8oR0BTuWNynWrO3eNo7uM8pj/bqjNXNaCXUrIIq2MYB6wlWc/g4+vGWOV
UcBiw5EKKKADBj75S9O/+hZBzzhfTh9KhtM3y+4Bm4vFrDpYSsXSP6m/qRTXTQ76rNOxrh8D13JB
Gg36L13xPEA7UwFPuYy3OJo4yfFwCfIrSnLaNkx4uv4qazvgSLRPS5ZLtQM2Xt0z/cl3Rb3ckIMR
NSOBoAkprwe/O9rleHvEisTPmgmvymED4RyjcJNjOpBqKOvUmlTCxp2ZiokzhEXbegV8yCaCd6i0
0HX3ARCzkVi8u4J+N3DZThNNpHebfWQE+Y0U7xF+xTLpclx/N/DpTp4sc+Fk7gnLEtizmlNdSRSe
pWJJOScmzCA98i5jQt7iTKkqu9K9KYbn/0VpUJDXQQvZJosP+SLf8AXi6WfEV/WDwed8sborWjSM
SvpP4MceEH1CwhHzG3xOcg20mCGKOUqoeSYZKMeBgZlZ9J2wNJ8L2mhVaxWiOsMC4hj0kUzpi4KP
+7YEYXsWtgiC8R9fC+/sgxiJ0QTDVx2b2ZVQNINhINwkc6iVa20OomQNRsY+SeNtP1mVD9yiod3Q
gDeNlUs3J40zWVF2PG9xmdOKtaxOlfNo8rT3an5QuxJL1bB5IkOhMiJoUwCM5ndEb8d45mi2mmM2
Ufz24yvydn00f9wdsso63lB7nWDvAc5WYP3DpwqDwOTnTCI2GVE1c/IPZ+L/ltCnRvgjjoTxu60S
4iuI+VQFvZ69S6WuxJZcBsPXb1Xf54NyAEQnfvI3Aak03s+ZIu7CfugP+Cym5bj53mK1j6P2rZSq
CWvk0Tf4CwUhYLXscq45wtcdhg8w7VHu+/bux4GRn7Bx4MbIXYXTYsp10i8NfBFLyQskAuDp9PkX
aYi+NH7eQ32Bb5a8JIpulErTvKkGcwnAIDRZ0JtXJk/J4J2PFvBH5dFf72G7pRq8G7J4BnjrXdoN
GvOHyrrarOVmye1aq62X2/OeHKHHaToaofQcOHiAu6r5bGjewdeLOIPO9f47eKkVLMe6OL4ikKwD
LmlqpOL94XK5tHXQVxAbRHyeJATTQE+8rshLlsgglU/LZtgfMw7xrwEBH7xi1Ex4eWMXJssOmY9c
XnQ6FIOJoDHuKBGFoIIzJcKvjyG/yZBOEK2aBBk5Hzz7tR6afsR+vxoUDY4mvlcqOhya7ulQpU9K
jTWhAskxsZzHaet16YKZGoMTSXkXZR5To0ogK7z0Gmc/B69Nw0fmpSXuXRT1c2BCF/kNlEs46P/h
9DYJuuatOpEjL1oJFoVtPEMGU4z9qTw5N8I9hnV2pkK71s8kwVb+G9TmkOJeQmnIEolgaqvpvwTz
BQV+gUpLQPVCyC2wYb00wHexnmrTcYE+zsGfgMmpN4FGEgyYAOicLlD6HaJk8xqev8v7GmDC8IZZ
S2VoNZslquANaRq4bWz42yJAFpchqE1SGng5iG0albwEzv+UYWpiPZDriDt4uhmOXqSMX+8L5+ZV
rx6yJ1yfzHpWkxTqAicrNHbTtotq1kaMd9b0hdjzxv8g/T4wUU+KF8zLm8qSE5tzJR5xgFEI6WpH
293TDaaGGydnEl0kgZmeDz6C4JCKqK8xYpYoMcxBpHf9+ofg5sgUVL7k1rgMSW7kpPLTQ/cO/5mH
W4MuVqhtZ/1egnDGCZoOe4cbOV8JxKL55affjafj90UDw1MSOWV9+C+MAWkTlhAFlQojiBzMoikJ
k34B3Cf7sLu/LtoP8QgwIM4tY+2lk9NfwW1jWhf0aqfBToEbbZZNylO4qpuCJQFoZwpiuOShdMb8
l568tPdmOY6hm9Q1zXMwc3j3VLq+83QoXb7FBoasnu7FXrtd267l+Qy+wo9gJj38LlwpxNHUhS2y
yXdPJ9swkHsVLZtoCdIgfdVFe6MzWw+VDKslTicKEXDW7Scv0oRpBfIWlkhalvxGLjHXCdAVyqlB
L0w9zODwEjL8GRzL/hcFD0tQPDYDGpvovx2C+PyB5oEcRu+xsR4OfPl0+0cj3CcyQOn68197RclD
7Mrlzwfj/44KYSU2NHTyBC6UST2PYAPwzhPfgbN3DL4KjRGAJL4E+b2oi96X0YmYKzXbwF00D2uM
5CeQOgtRhudS5WCTPHeaPjjx+78L0529MTlNw5XFiGikoFuM1tZ18FhtWrN8O1bb0LyrV9h7fRi/
ZajmcrvfEjTnhC0rfQZcwDO/gIaokD6Xl4FsU6Z9XlWwcPXF4sGgevCwYZXblJ9PF0eAtlefjed5
sMmzGVmPTgyaZ4NNdFTIsm0v2s8Zo6Z0Z9uVIPkzuStqABqp6c8CtsWpG3S23g3X7ETw2mpolF2C
aB9Xs/GICKANyQ07x3y7mU9QavDTU43FXOHcsUpN7YU76QhkfEoL6W2OeizP8dDCOHqcksIksdKl
ah0RytN1bKWPqitkCApeawx/2nchBtySYcTs/tqluXLsQG6TC4x3+J18/XjkPM06DbWz8cjAO3DS
Hi/cefAExbtSq/vBEqW+NzUWdtshCu9fuMjeBNuxJ4Cl6/WdUQCyQ3OscwoLFrCcuN1B7oEyo+/v
euF9oO1wSRYa8BcuDcBteuREKMDrLR4MOyHvyIGM/0gN6di3joJdfX9ABsD2/ATLwOEDBzbeDXdi
2Rdj+6BcmifPr0TOpzWITGjN2ZUgy5SK9SpkrF8Rdwl344eXaxC/VLf1+7J9g8IDXGU8PDj6a8pq
PZ3o1hOhoeS0XN6maI+EGU48nzm+SKJAJE5FFJvlsEbRlOLJhhtBfrlI+PFQ+fqQkBv5ltkrKiB/
+9fLSWM8UZ5w0jGLkbPeLmd3Z1fiIfjtNeydKsLhME1r81DU2QDzyncfjXjJV1IO6+PhBY+0oR0T
8wB1MGF2nbHCyPm7yA6GQBzBNhLnpVuTSDTFcj/ED1CXamEZUkjyhXTLrs9V5cmLg0PP5CQ+yPaK
DgPTX1/PZDlCHZtUlTHpBKFSL2Hpo1sxN4+25lSFc4zXTHgTHntErEzo76fRaSACMZwNmuoAXmI+
Iisi/oaPGplWP8abZxLzQFu1mXJ6lcEftNN/uVcqdOebXgghO3PD79d5rkB8Jru2FA1/q6ud1ztn
4hsvxxe3cPR5fo5IrE8N0l3y+0YQjc9N5Jlos7hjzjATlmwmZr0yQK9N5aSeMTYo7141F7+s3TyX
Gp4X80vHJJIPqq+cvTZkf7zZmUoEZ02DxzwwoEz+3kiY0X7jO7NKhPlR/IQo1iEirnyu4xOcV1BN
aCzIPz/4MNSWxZ+UVDpwnk2kHvIXf+hvK/QEA1UrxKyTZKUqJzdsLsMkqmJKoFD3Ez1qPSH8qybf
4hSqlbDS0GPVnLn2Vv2bPw0SSOhbjc2hGvH/TRjyhuzKcX5VZg67zgeXM9aqgxwgBsCQhBflWt7A
c1QdTKOdQh0EujXXTr6OLpE5sVcRzbpXJrEVYyb2JQk6bx966MxzvDOf/Y0kbQ6N3dEy1TBnTwdL
jKbeCzaloymbyNpDVAb6d8NM38IMNzwNHPUJEfMKpqC4UKyfVzh9Pq+gsAWHm+bfiT35kSY580CP
9uDQjpQ3uLbhQmRfBdhJe6B14gaJwmoJPkkSTdXWTaUgMN98kXxLBf7OTaoYfrAd8/MYrRkaO4Zj
weRUyEA5nJAhqpkv/0WZF9JRFvsydvig/paFOMlQZggWkLoQvCSNg1XBxJBpehYsMTFIY/EMlZ94
lMrtSy7xmUGUnFJZWCa8xyRJMQFHI0mXAhrHIGPWOTVR7In0ExX8N77XBUrzfzfGFHff59AFvPU+
29BBBA2Uc791mBjnGZwMCS5ZmLJOVKtsS+bJJZrnuCwy2TzKrIEz7n1lShAFOJDpSJaMkK5OCX9s
5dkxvWSAwEog7Njk3ROMxc1QaOYovg1LO9o3nvCzUPyvp5uJwyYZz/ThmYpMRH2XQ8hF2lq/FAnx
Dos9DhGf6g3Q4JPpAtgR/8pYUN9gF4E5UQg5hPq+J/f4jUFg+Wgm8TviwEagQUUrhEnB9g0lIZwB
dcAVb9rFEDW/XQ+X+ghi5BGK623VECQ0F2GhCqaZqMd89zAwur04YV1wzJzwZdq+BhL4Gk0Yej8W
gTWaDJeNciMmyLju+6O4ERZ+ss4AQMya1aXZLFUE4UmgxFWsecMAnuMyw3CD6piPsab8Qin+mTxf
m8iaqrDywTc99duvKpq3hs3psetHdpqaLHX2k6t0F8lQXOeQdHeOreiYs96TLEWbrJrEfgN1t3BK
7xPrGYdYbuTBSsNCaEVr1E016vnzfugTVcPiGLqT0EgJQ56jlU053MTNmeTzqrdUA2x3BoFzDbW8
k2cyprGuQdat8cFcw74ghkOrz8WLQvui4i51fPtzjQiYkN/05yKgu7fhjpvu/3L4igxaanwEZowf
rTUB5OTAOLVrHWczjbdTORBMqAtX6Bmqo4ySRe2NVElBEekBqnsJRDeEU5i56/CQm+ONvlInrWy0
6ci8RhBcV3EHSrB0jyYUmgPffA0rWkW8jzw++Y8rmfOaWnNJ0nJWz2R+pbzyP4dLcJw2WTOJ0vyz
VRuYN4ETT49md+rocSjuoQVMTF1vGlD1p84icluk95FoYxo5J6rsVZ/Vwome7NBvCKumk3lbKDTX
BQBRzUP6226WkdbTvoriFwkPGtUaXGF2KJIshSvGg2G6q8L/zxKvnjhizjbYKOghMl6buv5ylYEV
XRO7OzYuUZwlek1G8KVMCe0vcGBWgx3yOg+5GiZ5gEG0t9MzLer+fE6Qx31QJfAaV25x9iYXZ44Z
M+AGs2z0fVVc+ycrm0mAX64OV9KED5nECb9ZcKCJNy0feUSozM86LqmhPT9GUYUJ28c+L0ahQRuJ
2zpYOmwZxIvDqSb+xm/lhWuoUlrs2pxNtcPx5xc9UbmDeLTbN7Ln05VOKFhVX05oQewZM8QZMOBK
QJhxSdFjwOXUcyMZgCcSpxSXUt+pKfYTvkMtwvDyfSTTPVtNO9kPbPDR8Y2D/ZjLq8NZx4zZf1uZ
NejyU0I5TRASRLyctMv3yoFVToCEDso64M1Eti2bLeBsPmG54C5g5diujlLwPkd1y2djufMo5lsf
X+eadVX8mMLZyq2PgE68cybRu9kq+hL6VXi8CuZp2l+R+TXveUzRs9xbGejggGNz4nE3L5aMzBf9
U7wJV63lrRNIAN4tttqiB95623oaOgDmCO01+wL3Nc/vtB0uzKvRi0n0wNiJs2gf3TnvFGHpIPAZ
y6kplOVkfEjnB5JKXHk5vgmUlvQWz4gG/diqqeAab+5o3n1ZZUfEoJrkIoz863VgV1y/EqbtK5Yt
nlrLe97mBzgOSM/b6b5x+jPSP/EbuLDtfneRsj7oFPmNAg6b/fxfgkyZ0t4SrhUjsW17qzVYt7CM
JEp3yiWGjY1gMJ0UdC1sHyon//pS0C1KbTt3TlllkqUtrlEgUtyNPxOAKvssB/tfb95sY4lAvEyS
hJlhut3nFKJSaYwyUQ79dFTj2NU3cNdF/syUtdf3hZuG//2BRcSwLc48Yw9ekLaIuZL1oQ6LEomz
ElTOD5pkm4K/+xsWEaop0igUQgDuQ+ZloP7uQwogMUa1dJxTiGxs4cI3X9huUuJbvL7HatHZya36
ePSgop3iWwUf9T6cHCAhDgnyvmwP+ArsYrbirwKvMes0my5iRuxjSUXVyNbQcYUwrISJDcDh5Cch
b2R91NCKWLLl2b3fsNzuz7aWD3TnVqqpVKW1r9ImOBWs5WCT/lImoPGfLteCRgcbT7LXUaRCH6Fh
jGfrJ3xiQe1T8QDH9H62yBo5hH56svD5mv9aqU3oqI5A4UKB3dRHA+CThFOmTG0KzyKRu2BzjMsk
zMdDTgEqppuUW2LNymzcpoDB8AiR/mlykk7DirMUoqzc2m2Y45ohV1beh5/+UdSUtEhWE1X39PbD
eO6M0RNvVMtsnX1UcmG/jVkUgS/SB9O1ljzZqWKXL9uyf77+327jRjz1SXyCwCajXEJr2pudfFmm
Wugir6vK3R/eigya7RgTs8J95BDNWgULQn4L/Hxk8wudRxcSuwWasl10yPEaMc1F/Dg+Dg0oK7u/
pp5HC0swt8/e+o1NWyFdjSMZzscLdLNM31wm1Yuj+b1N2whb00COyLAncpMxh7BeJKcQjfNl18lG
LxKcNC4cXdC3OdjyjlTa14UtTSFmkA1xctcfZmwDUaVcCWNxxX8YbuEBq5SHRUMixkKV/oqR4afC
IYLZhK1M7shDF5b9JBbmo2FaiUD6LKzrv3fIfIWuq6owAD1hCmhRU26XufpT70hOjfAS1TcP84sm
z+zfIOwAAFfK2HMZxv11N3Rz612mdGfxaFO4R4XKrLx8LIxZSoIAMRCf/ighckRV6lKmGEJNnpZQ
d01WNEVDFG1S3niFpCPm1Odya/DX8XojiHLNjvaqYvInVbf+pB6X/e+uWCM9kJfdjKJnP/90e4tJ
wipywrQy1AJ4XuC3PtquzoWb49uOUgUXNzU6kLM0ThARQEjVdBu7kBaqHesdQXrFN9YCUXfbtlJa
ATmZFRpKQGFNQYMp1WBsW4ArPwWGn9xZNH0vur1kYukahWQnRSwhxOnU3ow0Oh1Gu97O6FZtdjKL
AgDXrH0MgNSZsqUqcWzmSywZWw0uNC7UgUJd5v7FWSMOik9/LqMG/YfRAU/jYobGOGmAomZcRgCE
nKExRHrdiRLf9sf0hV9nn4IVWhHL0ZDxY2S9X6vUGlGCqILhGFBL2R4ii/XH2JGARPY9cp6jl6GN
3OFl3U0NIrkcZftsU6mzxCiepZ3NJmZGZuqwuNzQ9sRAXP9Qjw7L/aS7SuhqysFXmNXKk4rSgb8/
gt632yWJKCNHYFECXlOaMuAggTY6WgK1fux4Oc7YH75Fl4Ahhd3W9YxVWU0Tug7PeTbG6LYZfXzM
RYXSGqBZVT++JFGDjMaQwkApAXXnVjUfZj3DhxZvasi2nQ5PthDOXBP6F773IKxFDVyw/2n/x8RJ
Ce1LIJTPSR4h3QvFV5GP7/ShB1NJJIGo6weqb9gu15m8upUMyru37M2F/VGILXlcKwJ2cC5Eugmb
Bnb1TErvc/Of9WndWvBW8AP7YMOS5eNyH0Tv+eJVVLn1q+y/oOoqnp8sJVeQaKjzu8ffGH8pm5ul
1ES8F261/VlPQbWVq4UMcmek6aami/hBgzL/HQmC21dL8pglefRT6lfrVPLJp2qxzb+PQisLsmrt
S5eCPFS5CIHvCpfhkpIa5Gy1V2M6u0yKfH2NqW1ti30h3dczIbJv5ycnhDMzqF3zZ4osKsU3uHtq
Vw75wxeQC9WgyVe7M3wprKkeS2rmK1SBDUuez4/ttJwmwMrv5AmEkA+kB2NZb0FpN+DZeZgZNK4u
FsqZxEze91fqWgo6jDUlTkztzdUhmoYAN4faIRI9eb7ZD4fj/Kcx4pXlPtp+cr/mKP+4HLSHNBLH
wf07sVP9BwepRsHI3FlcsTIl6J/QCUzHuovgbGnrsImlcRyZXzy3Fahr6nqnqz0FHJDGSxsIEjHj
L8QKQDY7PleIm/3kxIFoVT8F7MvQorWyeYZedYKEdHZTDcBlAQ3JvEbTQlc3ue/ajT0C3BDyOGzQ
cvxmmSKz4NLI5RoXMJMCklK5xxISFZ9ccmysbtoKQcY0GbZkTJJ1vWtLMq1kLMY4oMBiyeRvdizH
AzbdSNLqCyblWRweTilxjnr7Cj8boKQ5sHI2A4QBfB69CT4pWJFT6c4sJ1WO8MXQ+GXRNLlaaLXK
iNc4h4dyHOprR5GpOwZQPVPWDXnrwbczc9z6wdM/xaLem17Czo3u1su0MewwOStuu7gt4x+jPYrx
KeCgkruzEllZsgv1gv99BvG/+18vmDa+O4X59L1o0/5viRw7KBuAzy1RXJtLO0/195ZVhl3b/BaV
eWea753pk4H31/xjdr3gIwp9a6JipZL8R318J7c30vz2WBTapHw45XhZXSp6k6vJQw/Yqk4Nn3pX
TnW0Q6M3l6m6rCsi3NSKeGA4dCGAzhAEaBcsM6wpCZYtPpZSfrTAhZX4JRext4NkQ1vDW2lxLzzQ
hN5ldhOQICQGgNyNu6cEEbUKnlI9Eaqb+csVAhKXZMfUp/7hpJxtunyL0M6kj/sIzXD1Ayy1+RR7
AXShBbU1tEMs+QSFE2msVLGJKB2htgw81UEG4fVBUzKJ/GOMBjy/PA1brjxgpo8hbSKdaQH+7FT8
3hyGlTvVE2+cZmm+RnSLzVV3stnPoxqOyBuc9wmlBQDiX4qg7yuRJ8q4/LykfMzAQjDddxEsL5B/
KVsdjX1Mfv2Kh/1mYoRh5ZCSNc2RApR+TW855YjPFkTh53cHpRweupM+MngOOkrkdAVyDifFpnkS
eRndUc0GNMdS8aNdvpvt/f2g1W4jW8aeLBbnI+Dn1QO3lKaLf3XSzpPNXbWB4wHc9Zqlu0NXW6Hd
i8sSe7Fg8+A6XkiEk8+fOJeIcsmqqeZ3SEGBK0is6zrThWGCtGDFNQvwHh0TeFm6wfI8t5KBUknx
XEhjSMaRcIAiOIIFzcgjY9HEzcA73hWLXewP7dl8aNedBZS9ydZsSuNFbjGUUW3munFjDWqctsD3
9FuCpd3CvZ1jRf8utIW/3VxBhf0iFao7kkH2ZvXwUTYzUZNP+weWcvMIEJygO6V5JOczbINJ5EIs
91kW42FMxwOWF4OqBXYA1SMbaCf5xBl140h53Lu5OsNm6DPWT4tJxHZY2UKoW6Lg6xtUyvc2vhGG
MhAzMo9GEQxd6E5z4WWBZWIcHM7sEyCYKTAn2vl2D0FMhmoNQhy8rw1+EbQfhh/1r0QpmFj/Gpu6
XEn6OEW9xwXC87laaU4VLsWQRxp5zb0TvZfwjUuRySiWsZ6ILVA4yd26PW1JtyQqdKlY3oEzust9
0M4gYSEV3hBlnW06lTP5XtqkjZJV50Hv4USkMf0jVzN+OX4d0qz3wlihYRrkEI1GNRmY/jCQ3IRb
0QXmcZqqdPaRAJlAZCcznD5HFMcvcHgc9vSNxum2W2Kjp46Xb2bAO0NWJQk+ORS2pHOLnms4LVBJ
qyg/Davo1+225v/sw04pjCiY09MwskEMh88ohufUte6LGsMNDbIyrFo9tqGoP61nBJKZ39+CppmJ
eBToi6HN9npBxx1XT2qwUPPqF5MmI81PaahiUsGNRwiA2XU7vOUaSoSEOlAEcWH42OO7awbeHEc1
xkc5GKhD7haHKu+wYEXq9cWCuGo0YiZcKaAzHgK2WQHQIF1rshR/B3G01K0ybAFmhJUySrkKgsEc
U0gQ44unbil6wNflZs+AhdTLMNK0yprtPKLN7SI6pbLNFZBnuHlf5TGEG3kJUss5YZn9C5/rg386
r0JORghW1IttbUnHEFwXRmc3+bQgxDL0Bx3aQ07wQ1tBdR0e8iQxSWR46qnALrnGwCyJpK7U9T1e
cPaeJkRAAEcp8bXCFVxEOYncnnhvndK5ddpnGzNyUEMOVjtu71Hx9wMFXLLIscGbD86kpoI+W2fW
hMd3VCODwuXl0IaxYHPkT4aLG5eib0HAGq4Jhnxa9Aejuuafy50phuqFGqOVMrd80UhhQDHcr0pj
aVSma4Z1AdfNXwKhNRlSCEiQuZ15UUVnzskkhXDSXW6WolGb/oOodwK5JykgDJvhtFk2BphS0IxM
UH03tTfD2Xeu4h8EuFZnbwh0x/vKyNfV/hScCAGPdAgNJHwXgGgl83Gkjwmcvc9xi5nH4x74LU3a
BDSlTmnsklGLuCj4eNgbEVvI368LhrIUd9g6ONuhjiH5jNe88+LPfEjVfqIKYKHmEMH9sOMDqZy7
8r5ET56FaJNAkKFEspX8gHgyxZQJg1bUVqATnXDkbAHFHy/tSJ+X5yoWolJ+BVlNp3qod92JSLMq
zK/E/Hdz/lVAhs4tueBJJ4+13MEsfo9pi6ISvKfJ3wqxE/eafeHKSznYmZ4T11DH9PSbXXBU2Z2U
GgOLNlwjfrQiZtXzh6vQxCjq7orTUtH5II5FmkVYbMFsfVtroZgx07C3QB/zanCJ0PHlFoi1WoCP
LlK5TjnQSS9hXV59jMQU04Xf2UbftfBQQjtZohoj4Xy7KQWpQrkX6AIQV/dhOOmyE0IvL4fbk/sV
6hCJQHseumqc4k44giVv5LmFmz2pT9mFqiNnmp7P6SBJGcJR+G4kAihCq/psJMzBRNaxStYEjKhn
wU6V6uOWxl/+NowLCpip5zPZXczcgUjicPYLpEUCEa8uFy+X60xZ8qjzF0JvP8iQzvAE/GKk834c
fgcQM4FRhbm6awkIGNB3sni7Si0I2W+AmC9Ba8wtJRY6RpCE64Q6MDIxlJ4XjRZ9q9xNnzINN7cV
PBVXihMywDkUHRpvDIbqtf2nIVVKylYZ0ssn8orsdJzOQOuBHw6moOXs4P2ew+ptJJrGHaAHXSDg
rb+brLcMqnlCmfnDkGQ4RpdEruMpvTnbYxG/dar+26OC1ZMTMsWpzkFJTCviHm14I3tveoYROvCY
o5QcMtEPtTBsEQjSbKbJJwOGOUzOXoqEscTHK3bIdTDcx+rwmtVoZSbguRObZw82UsBQUyU5fz5h
oL+T6RchptQPnW6LWvkdKZUFhJmT2WVQr/NwZ0uOWtLGHzJyvqpLQ01OQiQzqhvQ6OD7N6Z6SqR1
0OZtSCo0pY0VbYrzdZWEPzDkOyy4Yu2a8oLnC7CLl4RQbvJYQrzKh3v6rTZFd2+zDrOjPjZiVzNn
rOFVjortFWX0HtCapj2TTXeNLKmlkKYn5mb7XpxYTrIltCrDTe20casibosXSvcV6FI+PGSXweoB
X1aoxZrFjwiXmSwRdL0oTvYhnGUvvpfT2/xWRd0Iv1HTQCFPdyqeIxiazGnzLNCL2TvE2+624Lng
j40eQ7acuDH4wvOBu8Xf9pmlBjHw3YRNGqxpgvjEFNulXWKoo9aDgmdD4c0GFp5GsU0L/VGW02V9
dGw+qYKzcrKxTXdUz4osBzbUGSU1FyEGIMshch6x/4R1QcfWypnAruZFgyzNe3nGgGexSp1QWK12
FJ8IS4Zuy5Afqt01NAJYfaXXVQjcqdKnq9KJLG3tXzNTZ0CsC1kJEjC1ZtiRIRJg3LlWkgjI8NoS
RbMg/ZD8KzFsNehdz5N1+xM3H7MNShMYiclxJwFktW+cSqi0v2T5zy6OhYAh6EapUeKBQ/U0TxD9
MKkpH05xlH/2K+FutFdvwgBNItjiR47hGjCQ7AqbAM1yR5VDMPdzq7FJXu7DRvu6Sc4bvVjPeD88
UcJeDoIl2F+Y0YbOjZmhZP3+WpCA56u6YLT1RjbE6HrTgQgCAEICB3N9H8lX238a4BcRz6nQrdsj
B/4dHVWitGbRmLr8b0A+0WkroThhk8c07xBgH33l/ZRoBQLOyK12PIO0mLqE8UO9pkD5cdnGTYmi
7r1mdROVD5zYoqPNURDVGXNN/MeLSzmr9MdtmN0qc9K+5++Khwn5SlA7gyY3x4B7RYFtwkcQ0LTV
gXA+T2U9abGgsAoldv1izq6ksfAL3hvNNwD4pZiM2fUqBdl5BEeg9RgyuqjTnrQ5/ztAIE44GdEe
7dbVQupKPpDmBaYCCIdkq7GX7sbjx77M7RngpbXbbNdUUUQudv0RYCxvcSixEmb4HMnZX/bAXcfd
Fq1//WN3foSLinRMSRIv1q5ULMWgGvzOiN8FtXaHzDEiQbQp/jqxvq4BBUBLpoooYR5e7GsvUwy+
dv82euVGoDoqpqEHuK2x2OJMag3JbJ3toMz3tBLrAM+KvM8NVWRvXLErxmnU5NbG0jBpdC7s33C5
mcnzuu8sZm+BeAICzNIo0hw+oMRH7hVbWpeUDysq+fUHDQ5fOnRA3UfZwG0eMcNdM0sLMFqvuLCO
DZQ3lzKsv5mQJWXfNl3/lqPAMO00TcyBND7V4f7ToTZ+YELz7qHX4DBKwrdIzXOfMFeWp2D3Fm0D
nW9XBE0t4fRNR9rg/ZV0Q102S9O5dhITpkKSA0/AbFcTtLYTepY2prfV/PPsBvhwR/g6a3ddY8jB
Rbh+41GF5PdQw05jhKF9A5iVaMMBQqHaL3odR7MYyhNdNJ+tYc0ixB7bHVvgGhRdyWleqpXzGWv9
jcM7Ri9XKTbH3O0P75G9yFbVew0ZL2X6QilkPWwghzSwicvFw0C1wQ4PxuseHTCqIhNGGcY4T9u0
1yutIT9inz2x8qkkgcYE+e13x+Vx1MQfM+wpfgpVy4I5SAUgo858BQQDu7Ezx4JfChNUkztC0RyH
VZuBlKPwPMAW6zxju/AE7WxczAvqt3gC9WHpibZSDJpWUUbRRKMtuunxPjAwZmkYRkLt/bp4PHDx
gEsUndEJtLuSBOPm+ZxT6BqTDfQ3r6ZCGDqlPEZloRl+o54UigbKEp6/iHCpZOILHgulo5UQTKgi
mw8Qrgg0UhnEN4I+eTRkjPIqNjObhEgJYgduysD7A/ZGcLToulQrAMlYxi7PWa4SWWJOVunJJ3Se
VWCGsbnxypmKs2k2MIbHrzdA9KmLEHLaMAekCLCwioRc7PQx2UcKMuaYPFBQEk4KvaqD39QNrEzS
6UIMB9RqKjHdJRePJ5up/FT4J+YvcRTULtymPaT2kew9jRAOF3+mzY80GQehsNDyRA0oXt6zsUoe
lyXkhr2L3J5qBzU8QbHKtKihm7W8OjhDy0InQxksx5aBlENMKYZ1njpa29Pu8YMvdk6JRiCIKZ0e
x+BVVrv0w1RGGhuoWYqMAL+RZbdm0xSzRbZ6+RKi8dHk94iYC1+KwU0XG3wz828wJkXVpMVsQKez
XHot8bLu+t4f4pANGF4LCs6TlnY0f/KATk5W53I+SE6oMuYHO9S1kvPbaOpWU/f8ZruJD4jVq+si
yPiYnB+MEQ6vBMQxGWRGza9a8HDZG7+EY73N55lizHEHabP4313LNx1lxRqnADmAGUXPRpkdDDdx
sawr76tsX3aKLQPzKsyBriuRPkgEKMZbGlliCyh4lDuXMvaq6pDD4CbCEwY070Ep/Po5JncV+hN7
ZKIRnpiY5obkO7Jd3sLXU/5y02MJirZlPE+Lcd94EIDXbJYhCqQ9f5HZHxmC1llR1b3gGItpBuSE
nsnNDokKDFFPFO/LaO1gsmTbXw21R5ZpnuaUuBgHZ2ASbokFIJukBazQ7MnhsW6c+vXnrpEngOGl
6WbFXW51EeW1lY7Ylez62p9uQMWs6+r1jGd5rxbbhO5IxHqv+Rzia8c4r8/1JSYe2OalvHtoaSY6
JIShRK6HYKsKiDk9Knr91q04iLDd/KxkSiLR/M5x2Z/IvdMJe0MpEtqxo7FyCouR0Vf7IsvkkeKB
wRG49S68Rtop8p77S73BZ56he4XmRfHV5NL32gm14cDkT55fWLSZa0Lcf7NIhfCo0isf7ECn/Nhm
ACx1HkGL6Pwc05Tx+EwP4UzjrsBvKoozrRdNEhk2P4aTagHgZ/haRNt/Jld0D73/M31U7LTP8zet
YAQR3fzHMgibyxK5mojijJWBMs+0KhlcHf0EiVILiONgNs7NHbvRzhb3m9veISYdkKyNVTxoykTB
3f1dM0cVJm8ISVsIn82Rhkx4P6gG5WLD0SXYmWNYOtV5sgYFlHtu/eObRLefPP1jaG5bhgV/M+QL
TjzhevgmhCQpfdDxOrDyO+KdntiGLwU8MgrYudQU093f2mjlu99QSnmrWwcD/CWuj8Z8V0R07SqD
UjUmfi2XFUc36AOdPPIdkQRNtUG849iN42GaQbLbpdoLfmYKZD/KBNnNz+GKCBH224QRx0EqQ4N1
AurlrVxn3CgWInJxEO02O3N9ST1ucR3Wlc3Vl9iAltqQUFAIFigI2rjh1/3J/lz60kd0/KAaFvNe
YVQrqpbcAW+Ej07mYipSt9A+vJlOxmJkCOa2oHBfwp594BFcpWBh8o82ragMtgbBMKr38CLJgfLG
gVxpUk3xc1EmY6f01L8Ie1Ue+4kh007df7qBcyV4OFX1J42okVMR8HLiL6/MAZdD4e0TbIIYk2vu
ZXXnqxeE61WLcAeFoQqESHTudKdDRkp/y8H9lxOKaFIwABaqzKvhoS2Z4FC23+nv3OnAyHoUk7ha
M3AgrkTscOEOrUH8si0l7XnBDBa5xtweGbOOTHF4TIck/GWvoczXlEGc+yL9DIxaXXfWZICXzJ5F
9jQGwKJ7Wk//oi4fJe0TujPJUY8w3yJPNQe61CAUJJK7+ZEJT+Ejz5LWZRFQCQa0Q7zg5Dhkb6/1
uzOSzps5yk11EmZ0SFxqCKvAbm1OBQWdzLUORRxkZDnHiPVzHwVaVuEmlwhI++FdMaimcYg2ofyy
6e7Wxg51uElKem+AGfRUmiG+D6zZcLZRn9fue45AfzQcVE934+jVr1EkfvCyrvvt/BEDw6WCzyVN
Tc99xn9oHMOnUXR3t1eZLDO7s675uqHG5T8DCHB7IZanCdwSfYUfU3AY05hICHYDtaX0uWvaBQSp
aHDmlcotcueqy/IeQALPFjLlFcftm0QNp52+zhPca9iCLR6dPQb7tSkJkgUDB7kVcPkwIWg49xvx
ZSeDzaX8lbAwoKsc0gtHBYllacTcf7v9ft0MeIrBYHA2CDA5F+1ilfVuVC9cvQ3o/+iUcEWMhwZZ
BVQt0jLiEaEOoSLuyX7+0JFO0AG6k5tiwWUfJwEh4o1Gqqg6wkLI9oYBFCfxZVAbap83rbCoE96E
YpK5W85GSS8fAe01LE9nBRzsLIipYIVhvXSVV4cvihl5QiF5Dy3U05HMAP0L7LLNCVYBljbkgBzw
BprBs0iQuLMECzV6q/u8RefZZ6W+AhkA0nVitC8VYUvvTipNa54k65L3Xg5ndbQhJNc61vIRZl+N
fTHmZd80n0AEzbWL+O1PSpf6AN0rMLDChR/nOmY2V0KYEGKxH4YtpUgkXIdkmnuO8Sx8IbCk0YLL
EbqZ330hds7HaGd99uynmVeKzkaUUG1lr6x/7TbLUe7yrb8cEDu/t7iGscGb6w4NaYhoBABNfJi3
Vr+Lm0NN2bALBbZNZvf1k1GkLcQpAJYy4NByzIauutuFfDiFm4qQJzsf0pQQAu8kv/AkZEpC9CIm
bAgMfOBVjafKSL+nitUxMHW3uQbZI5f3YIU/dWK8oO0IVtgy9j5OkyoqBkj8ZiTt/o1fHprH/rEU
ckGkSOOUMBXruFekui87rt5m08mSnB81ZOKmNw1z1hxUyxQFb18fGbkOItMtpEfCNoc7McYJBlQn
dhuajlVok6v6Op56rMTR+y2OnGNIz6Qag/KqwTesXexrXNYgkRM61LINQ4f/tfPIvH7ZLbkIdSC/
dzEWvv0NG7N/+o3XLB/DAxVsL3khMky1tx4nv1rI4igZvabItM53NqilFFiOO8Rbg1na/qIrUfMb
zADLAPyBKp5k/QbaiAe8N9gwGVrlZVMQwx3HSrY64ezZKE0GB5mEtl1hf6snuzmDSQvowO0hqhCe
SeBuevp26y+fFm5KI/Lo7Vp3Zguqeb9he/HaT7C//g7I+5s0TpR0ayGAY/+0zEj/O+JWf7/F3EKH
8lBKgYLIemkV2+v5+nUwr4rLxq2qIG5lDTE8YcdDarwTGNm0FFicl+BFhUdLCrIEFqCieghtXAPs
Qjn+06xBP6M8JhhRW8Z+Geo/ghmeX/yeC0NJEnyTUUICWShWbZzUvy3bug/PF2GtcwAXfuKK+mMk
OMdGzfiTJW8MDMuZ8yW+129XY9hxS+zI4O2/WGLyocETIPlpi4Xz890l1K/WsDkAnN/ziZhp7oCI
MXZXA/opPPuJXx7vhVw8Bb6n6gfbgPgfYK6NkHY/JoHcYeR1nqiTjo18qEw+0drE8DAu5Z5oQXm3
p1m+PiBcVzjaMhXVCu+0qw7VqaGbn5TfTXp4Y4Bwmp+mrmji4PR1kilJiSHhrUefNRAK2m9KBHei
efzJZXxh9wareY04SdX03IbqrhMv8OyeL/scKP/H5xNr0iXM8pw38T4CBQARlEXlO9aD5eJNGshc
HlFge78kS/G2VH5JGJJGqwlfPq8s6ZIbuTUwA/JW8/xDyRh4KGQqstbfzkBUBqx6zFFMQ5kI1Qah
4VAeJNHUMrxL8RRZqrtY5iIqIqIT9eqmIv4kmQO7roVSVjtfnuLw0nyQYhYCgbY+0N1iNGoi8KVd
8nqS4O+xA5e9yx3O1CaTArfTe8jQE1IsKCNCCVXftK8GJbYhuK27rcBPX5NwwC7ROBA2+r/LMYlC
uNCoy+7VvcQrofBj51orY+Z3B/4V71WHGoPNxwAwWi8XhGjOS6RPhinzzpjk+uqe8T/zwK8Q/Etx
oD2KrD/f1VBh4cVe4N7lKekuv45EX96zw1RPZwNNbplGHd8+3uY9FUdORNDh9k7nO/HpnPpb5jZT
Ah8wLPPu/bFyMgsUpRn2lCYkY1ritO2ueDgS2+pAYie19xzCU0OUJPOQ4C7U0tlPZlhDExF2TuKs
PRBYaFVu2mRT95Nc46uJXgDhua1MobrPy80yc7sNVS1YaxTrjsCj2GYJH/Z5o+nuuC3wiQ9qDQbG
aaYdWREDkc+sQ2UnXRhqXGVs8eiHrSjQXXm4Y4yyaJJRexd89f6yNg3H+mHi9+OpC13ttziz5R3W
hfdw7qCxvSc8botQqWU2UmSNc7cMSYLBIsNDKPdh6DcHdzFp/f+V88pO0+GAqS7EeZ3wRPsHL/mw
4IPPbKvy1xHPKgvrAFD3jVH6FKdj86Ndtls5umauc8t1/RjagQUTSK30hOSspTIMARc7qgOmNynx
FKlLWiHSLNwFF/8EQ7H6wozODczM9ifQ4xbLJzxB4COybp7uqPRdtVZrQuNcwsxP+Yy1TgywPS22
y5QfGMbePM8C0aqYRP5Sc1pmhIZE5KWImZs9vLwMjdpewGw6ymj1ZUqrzWmrLGaX7MeCu6om56GX
fyaMwOGWfAch66mB4t3NERmRq6eXIpoLiUZ/Iv3l5bM6puTrfGPUJzKmtN3mW7CyeAzxWhS5esjZ
cilACrMwv4fB934dfikC3+8s2KuGZn373vFkmNoSIVFyqMmsLML0Tj2eZWEbS1llwaUDy9xUOWg4
oIBi+52rmTzj7t+twv22KtqolhweQA9m31bRydT9o09WDrbm71lLNsKCVxq20fUDrpz8VwmfSuC7
YtoS6u1EMaWSyqhN2Tj7/DsRfvvHu5HR/Y49Ch7rhIBwNuqNToFiAJEyjqmXaJlNBLq3AIavcDH6
1ctyzFNZuhp7iH2UKeS5TRxVMSh+ijSltKMtayVSRyTLlQ2qbxbxiiyZEI/DX1tTzEZAhU6PTsD2
ua2KtRu/FgOHy33SFHHOoVIAAPkqo40cindfAugflKRuzuH/HUqxLytK3hO3WwUW/H72EpNrwXZP
i7RhoFMjvhH+xyqDZ74ZY9A1LcOJWvVs9qygSiL8xsvsNMmfFDcP+zWuuas1u7SoA1uqtHELcxZe
O/PMQ40xbcAaXCDcxTXiBQX4aN3EF53lTKva89tUFfdvBqaWiGzEkrZojFAEhVI2pPtVMYbkroix
0UjMreCJQ05mkPelw6EJQ7SwlaWvCN2AsrYDPMvkZez5OS0Z5vlCo1fHRyWY3fzF88ohiATSGsI4
7CNCTcKhS0fc5v1btmZ+bC1gexhLM6aik3pyiw07E3LK3gKgi2OAQn1fp0uoywmaoRKh03B1jcK6
PT4SDrk6PTJMxTmddoKrQN32gV+79PG5qktGXnHEhm3WRbEgtNnp9H79ZBwa5pOmTHnBn7t8VrzN
SF35VV5eOvYfVD+znqElUbtoh+vf5eInZWvnvvKzBnMpeTg237FxBmcqAfnIZaXIFuNT913Fsh4o
4q1yU2XCIewyTEsCwcgmDSkGH8eNpptpiAmmIc6vW3vis2pFUoTUABK/PXfzmPftqClofGt9nacN
WRLXJ3M0g8pIgyqc/4CxvFKbuRa/YPznPOJsm0v+Vrm2esT7oGX3AocJr5JyACgqyi7D9NoD7MKk
cBB2GoXqGhGhoHXr0eUNZnYZr2rgFWwejzb3xtRerIBRX4CpcuCE5kR2gbIm3aLYNlnUS+ictttz
Z49uLzt/e4jzq42F1gzgonOX0gCnPFmCS/3BcWAUe4dQGO2wO42leB7ns1V60sIpczH/cPUMJhA9
+ieoQl6viy00tjrAOjPIqL9cbDolA1bQnD3YsIN/oco4u8xAPyZld3CvzoH3UeE5bwa2auI3F8vE
4dWfPLQRu8KkV7pgkLr28PKTUijxCtH0VLr1XbXyzrLKrcBcOX7pBSlTPU2Yt2x3tgOqKRIHsnKJ
ADkh9XYgledPO3SCDqcn+QIu73ouYI+nYYcIn/8Zyyky6enV/7P2Kr1tYanejg7nCCvkXmDawp3+
xTCLyxcavFXAtTN31Zm+7nnfVcKA2AJtDBuc4HaEtM03Zu3gxTTqSHZ/0r+OYhPfODURuXnp3b/F
6RoKIeQy+yVYJ8VifEzxBv0lxap20b44EPx7ZAZ7kGeJV+zra6wnVqDz1ILQEEB10qudCJtF5QCb
dfPo/ox2xQn5j2NAjjMsAoGia+hqhNicFbEI5P9v+XGgqxrPGfTb3/qMQ3CFGEgI8+pe+OGeVUlg
R8JGz/yam2tDMqQcQNxKezOFFua9IWjVeQ2H30I4E+bXO253d7koBLjrnJVE1M3EFXQ5HZ8fsTXx
UZ713SUCsQ1kWSyf5BBiQRn9jls6896VG1axiz2KoL+t+clkmijarsTN6mBexWHNeLombNgc5xOv
uUbk44F0D5qGXLQO+CLSm8fjtlS7N3m1OWUs/0yIt+7TvhdN2/KF0f+KOpp07aBlR2yAY97ZHTiN
jYRtk1OzY4coH9ilwv8BLYfs+w0uHF0FHfjekLTpxr4p5OFjDqwFxcFEKcRbs3jGmD4XGEAO0dK4
StDL8aDMP+vAawrbFJV/acvDPxbaGVLoKbOCdUYFcK7vw29lZJTdJoiqvtI6ngImSv6CWUmni/Sa
E4JFg1WRcx/yqZIlCymwaSesR+DKQIS5u41vKPEYRmn7iI7qy1HSNo0dw+My/AYaik3X7Kv1uG+5
jLnfbI7MpvHiz8kbrnVfZ1eDv4SPxy8ambr85JRW37mffwyZPTWZAI6qms9ha0xM4eNuvZarnKUG
GuW7Tja9IjA7pvcRiHgdmAo2tCgsxIG9VllZbFMMnBAXeIyadiNEWysSS7GeKa2LgrMO9GS6dkBQ
Zs+xPiYbFpDQSlZJA91eGPl3kkmdA26NpIHB6QsuciN/kG4rarnbM1K9abQUK8nRut4umrfQ9R7O
TC2EOmFh/X46cNJxZoxFfxk2IQHoBEFpxcvmj9ruJkJVY2JegqGSRY/dv2JIGHj/9hBLVC0XhKzT
6cSZTs3dl9S35svzUmgiK04wOcL4liL+DbiLenC4lU2/MG/9E87b77W8DZbHUbeGlR0ZwyUPaWRM
uxu0ugqJYDdMlS4OQhII8X2nb20jR1srmdMBQCBT0ajeaFwoJiIv0yzTG1Rupd9Mncc0A1MFbyXQ
cUKo4miIsT3FvXqyhB3VM3LTB5AD06okn67CK5eWIdT4F5Oj+F9rt4zy2jTs5mrLRm8LzzojvAEB
+XuWEPnLnHGhPKfeu4GxW0jO7xCnjfsOhTOCAXxggFZVwDEevDF8ZfCfYzqYYHUJNmBtaDMm4hT+
0/UCuk8arEqyZyaMmuJVTbUh8DXhRQb9KAX+HBHypCNiPdz0RWjEzGDn0dCaW2E9euw9Wjp67Lpo
Ali4EiqF3ruNTKHrV9nI5bA98m/Zu6jMzibyYYUqnQUFFfjiynQmln78VHmfpMNai0Yw8G44N6z6
ddGnddJ6ucLIWMmEvY44wFWNGKP/5R53HBhA/pc54vLWXZlHlfgIAsMkfwq4zWu+CS1QTFJx9Oc2
GLVm8tEyauNJgDaFYXh1s2INa9rDQKzjExZrdAnajudY3fLbq2L8vv4h0SfHB/FLqf03AkFMyaIK
4w+7zMX4r4sqM8wSriSWkRibaG6wAbVjL0cqI9Gw7hSDHSy9rVIQnG5bAedRdNCHTTthlX1YuSCc
ZHKT+fFPyplDmBXQPOIO3R4bk++Qg0xbjLd+79TAeAMS0O3tfFpRYedjolJUZbAwauWWEMOWL7HP
Z9p+n5rEA8WAwj3Ylja3UUvQZcKcx4zVib/mG4ER6zxRugVQL4SKPQ/elxWlQX1BwoXcXS35GzUb
tzcaTKzftDOIlsxqSk3Bl5tfoATRSlNcLnCJFCFq1X7CfZEwCxykTezbvX0sGaK0T2Rr6OnvOxiw
pWQLI6+M/TENdl3+kDPeVxyEuMMdZ+aYPb2xNUza+Y42BaXzuSeNeEWrywcmxoRUuzamyP3rfxQ7
gDdP4eIhjx0e8IqHxiKKYb/5U/gV46lxWCnAYt00EmwqQz6anp0GepuNkUM+TLUGRBCWHbcJolXi
3pm0Br1xNV/VINGMVRAlw8ubDfNo9ZiOtHkLJ6Hw6NBCLFvMEp4Nt588kWJaLyIltwnxJLen1CNZ
Nf8Lx/6tdeWw8yt0f/lhgDFObbVXyE+8Cjn9QF7XOHAv5wesST2txFFBMfjDsIQv2RqTWf5ckBeq
+/C6hJiYg1a/ATT5ZmMsnBO2l3yTQ2Y6FCuThHjgODjcYZ5wDhodro1r8/+A3+HXrxR6J3sp/RaL
5SiTIl+e84TPDUeMNE9xPs0SHH8H4CHb3wmsRijPHDS2Kf2EdyG1S04GiVyKt0dd09mZxEMLSyO2
0H+QbBZDFNvtMErzOxR6dpGkE2I/xdWKJ9u/z/IXqoPD+DD4lJQ1MEWk8RDLaLiOUBooH42vMZ6y
WSdhYsO9GFOlnHEMr69OrUJ9j4DjA8kBpZdIgU1u5MmJmUN2788wNa2QWi7nom/DDCvJ4XaMV2ZB
a+Dey0JLpmZo9b859aW/OMRSPc5dhbcmMgLtnQZ4ytiWN/q9hSiVRWLqo6v48Nbl/fIYQuK6/gCQ
haStNF2wJqAdlhU4cnpPA3Wbp5ERAwHi/clEAF+TotldI/6igpQByKXnz78vsskiTWn9FQwCCg3k
yGKrUz84dz+3KUyLaN/jSFHUOHXHnuhBPN4fYOi6LuU9H79oga45Dx5hE+c3HZ37/izFX/XhQWTf
24wuHyoEG3D6d1yWm2ScMnf1JeHTx82NFnYpixUpzO3NeDmQsfdMECLF0yXVKGyd/loxUWBAegWD
xO5TdQl2g48xL9CYurTn3v109DPhFOhysVveqYbNw9/2BGmsyZwAFNUCQF1okuY+/lo4ovToViwG
2r8KTYaKghiDJkbdAIEtA4H+GBtIgvxavEeYI5lKk/jB57LrwuMWdGFHNSez/BveDB8Fes+gUMvQ
1zj7fHqy/4Y8ocvKrIPnV5irxF2pbyFvnR/77WFlueAsD2LkG424Tnh/uKvkY1X/Niuc545ImBJ5
gHMblLgnffBBiDqOqWACOZtrLHFch0Qcaqqz3e2PIuQXKqHO8xBb6fQ3wEw+3AW6RkcSAtJJsg08
2BrWj8gJcvIzyV2AVLNEWvgU3xFnfAzXk7b+0T4IO3o4wipRLYeiI//hN2/8xQByIUCdcn/2GXZl
maYQ0DEoGK4IMAKBOcbi5gh+FSgTvzm6ExwSjxnziM/YfZnyfjAG2W3gyG1dOqbVBRSWrvKmgb0Y
Hw2mPvG6zq6FFCqSBipugkZKokoBjAbZH8DBBhFPtZ2a9KDSMNsoclTsWPA+ZHVn24lC3REf1qSp
Mh5vWPGU/oJ3LfetTsIJsojOj2cwnSGCnLOPEhZ7WnRch6aI9o37JQmSaAvVYPgXnfBRWXQcCHrk
PzQhlK7oTROqCLOsl5P8WRawqwz0LwvH+NVjrtMV2mr5BPaq386aoUw3EYqGcwikoYMwbtUirzDw
4tEfZGTaoB89NhtZMKM5YuH5IynMVZjV0lUd0cN2d4sQlSwlvlSd/wtpIEjkm01UDk89LA4hQF6d
iD6kXiGatdxv7FGy78WOj3a7IgrNrDbbzKPkT+qRnpCdKbl8gchNK5chCMXNdOdYvVYRDoKI425v
Rhg7/Nva/p3XMoKgx1J/LzxCr463MMzwek0i8yAnb+8UH30Y/qeuGSvsbG7mWk/DfNasijyIn9O2
YgXPqMP1UIqfJPE2Gvw5+KpDkVkIsLZnz6ti2ZA7pbrENMb7l5RXPpd5Eg5QYxdR/KZWSDpxaG3m
cm25SFXdd+zLvRjrRTcp3kz2iqKJeFXwdvZJyXJdr6LUzwbFSeFznYWN3MQBJB8yYCxM+mTe+5t2
0MbGKkJ6qma/l47kB67QWl1TG+2jOb0Lg9tdWcjYLtuJJ4oRwHNnXBHnlBnMEQu4vS57KvX4ALgU
N6YZMtM8uZHdtpueaV1I44AB3q1MeTBI9oBt9KArsmVhZ/6QoKXw17mqxQ4OaAh+OajXdEbz4xZS
ku1uoaMvdwZPXJmd2j3R6spafb0RZf7ewqO5gEayTRt6Ysdz3fUUCq2K8o0rjPrWOyZz+lRErMUU
nmcG7jJ4nZf52Qn8o9MwnIdwlsT0WcIhoUj/jCH3z0WgJLeNxoTd+d+cT6MFVSJNTYnmgitj/bFO
INaVXWP2u4tAlUSQJTEecvjZHkBsKPHPwzXoiuMDiSlUmeOL6hPxzC9Bn++iLMeAwViagZCa3voy
FqRRi4lSZBsSIn8tx4K5YTc4ECE3ZdqzGVYotY53UhfmFwQyJDocR8FbjmuzdSOj/0pbnwxIClu4
KpjWpuYdNk4jinYGIaVLhysmptA2XgPgpByoo6MQD09ca8NNWF19pRyDwSUVumukexZrhIR4oEBS
ZDKWH/yGvMQ95hWqgcmUMKgzfIYMW66mrztOCwHTc0XGws9ozBPCh4HC9yhxXlVT/btC4aVQFpz+
KynSe4A9oPPE007rQMryivN3GYvRXQAAWFH6+paKcC6wIQvX/BBpVrgE3TDvV1JfAlCpTiWXkNC1
m/T/DYHd4f+2gelaIvbu/ibC97+fj35IXUX8j5zfMx/B6MDp/htflvmIlupZJ3qs1tQx/jQMKDhT
analARdQRRpPN2UktFrtYYVSvYz7+3nayGdWbKjjVIhlWVGUa9sphs9QdX76FHs981JAGh83WvGZ
1ejuU4Ey2L6IKMfU1kdtg2X+EdR2N0/geo0zk9zhNjARY3pUKyNhR2eKsT34Woj/MGynnvjBHNg8
ktlT2/p0D2xtYgjGdZEKXnaD/QB4laPMZRAHEoZ1GGipGz8OT3nkN8KyUGGOO2N240wOaqMTAwfU
g70DNLv4x/j8vzbBvu6gD3bTu8mN06QuGg5CCGbyQhI4xVvrbdatOKjWfGGoFhgrRidR0czWunU6
iOdqmH368/QwbNmFa/wwdBnSZ8IZ4vFJVv+be3SdIxmw+aTZJy5Kg4ovxbp2yhPPOa7HtddyD/wX
pctiW+sMIpe17ymD/8vYAGuoHuM3l2aIb8gjMJEuSSuHqBKQOResFNTUT56bviUqEQHbTe4D9+42
D33yimABwkkDfbGGmWhM4Ti6yEZBRlrWJDATuwFFg9Iy9/tE2Y6d+Gr1dPfmcCElI3q2hjUg0g62
37wK52i6Hou7U0ZcTEV7G+mJ97dBlqSFC0Pl6EHTZJKC9gnYg3lWPNA9HZO6G/gywAsqu309LeMO
AJdpulJ3VYq5RgGfOyhI00e5wKW3oNNaCDVFvvSTKVo9ivHV+LOy8LddkeqB0ooUcPWUF9i9AISV
4CE3/kN0X3hIhmzKBzlcPhUlAIe41bIiMHOPW8EsyjTRRItKWZJXKB0iMUu3spl6KKK71eQctY3Z
tuzxE5Zm/KO6mAJnR6+MepAmiiZuAtaxn4ICMYoocLV8x3ITSbC4MrepuqQO9JVQCL/p+1gRR2f+
U18zxR3WtHu10pJxfIlLPZbK5ZG0HNpfRqWyHE+dCCh/0cdGZaXjgm4F3MjrX3XUsXbDlnTJ16FQ
iCVCulkM7Q5sWUPl75ljdcTJWEZbZa/v1d98VXe0z8RC5DfCWIAtMqTnCdVZ0HCVQJ1+xmFFlJ94
VAHj/BcB+d7k6zr6yQ7swLbzXLdGM8mAeZuSvEi9iTlxptcqvorA0kiWvFF4cetsMUYsZ6murwXt
8asgSrxx8nVqRM61JEYV6DDmOUmxWkiO4xkpJWcTfUch+QzRXFjw2hTZJ3LKuBApqJZqM9dBoqfl
2al0eRXmf8riBJi55M+/d5pfDUlUtLJWxHrokkttGhj5NtTvWuTQOJ9T8ePSBrb7rM70MmSdJvHz
sA7d514icUSkeB2H7JBtzTTc+oxAOyq09zXv8H0cecTi6wk/0U5XJLhMgpdYeK+3xyzPZIzPRlTT
tAAFqNFGtHciHbRuEvuABQ5uZ/jp3Q7PUbpiNJXioToc5TuWD7Oh8ryq+ufOcBn160XHWTGvdXNX
gTyox3bWKkOauMUXMOf0OVBPXSCD/r3uyemioJK6grEF4jJkd27cL4NIbPtQqAUndKxgEy+sHGXE
XsrzqD6T7xVn5CiCpFWnyznXJqU9bhhaemEGc1h35RaIiqwVdlWQ8/q+lNOD1Jl5yd0K0BjZcOhr
JtmasBHvBpLwM263I4NYl0N9DP3vGdseOeLEBazQJkggE5wS9QfV+sSCI9eRE0Tv2SOuOexsR/WF
y86uGUNF4aQPOk1IJGIh6C/IQ+OZPJXp3uKvWXkLq4Ca9UV0qrixt05Idjl2h05KpI4SfvojNcVK
04bbZSc1samyqrgvYbQZuPQ16Is3YCQECAOpOJ9x8ix/vMChZ0/e+9ec3xnfmH8A9KDVSwChPhzy
z2Qr5Eb8Pf7gaZVgTqhsOUmm1WeysnN8AiC1awyp2cw/4/JQrdJjpYODCmSA6t22Fmcq/iLhv2Ro
24zabLDIR8rZPXeNyN7pOEbpYqhd3ONjHNVkza251/gjuXC+8J2Ehm26hCNr5wdN8oyfhuR6zK2s
0+O8O1YAiKRVfM3mhMtnrPh/cZUMhjbRCECV8ZgIsiIcpIQoHT0iQbYxyR4MHbc2FfbP49KQqjcZ
/mHofSs1PgCjfw0u1xD1fiA7eoiTFR7c22+nHfXNAU3tsxE67nddKfkgKXqEGjyctBEzXmT7qswF
vXUmWmeVEfo5NQuJBKDJpPyvOWobBoj2tbz0n3JYFqgdkK42ufxwfLKeTMoNVjQ9HR0ISjc5xwex
bnuWbWMT5wkEAnH5DTEe6hhZT/6LwXTZRxCJLLh2eZyQ2BrSRrDe24RUfO0EqeIl7sdIdQxmZExb
mMIAgy8vld6GX5vPaCglyoJctRsHSnC+eA9NsE0XY66o16Zi1qOlRDCkYJdhVJgwnujvWHjEwaTr
635Vgf8XDD2fPUP3jr6PRLgwEyWy1d/r3axSvqL4pBMwNZYwVLeWQURhpeTNYp5Cga+04BCyr0kn
GANMUk3G+MzYvDQoV0eKa2YSGasqfz7UX6/Z1gudkOFcbORud1zCgiZSy4WQJE9oxF040sgl2SD6
8gAA52Y6FbvZiCa0ZZedOaL1fJNcWVU0daZCXkkDmq0tGD+LSZJDWZE4DLoURo6swb7rT8izZ1Km
BTpzuaoO1BQbKHZ0IorGjbZGBruiQXwdfEdlsJHyeHaYC88dnmH2NUeV8dRXImIY47fTX82nkfEL
K9hUviU0V+U42WM79iiUHaNo/KJZrv9HdORJ0dmRprlvAcSmC4lato28qT8mMeznm19rAGxtzd7z
vxz8uZeErLCF1JAfj36TPvqxakt3qWk/1Gre/iQcYhX+49lo5HqDfQdHiIaOkb8hIkz6nGu7wNsO
bOGPktIqgqcVmoCoLA4LvkjH7IPiaeUG+bFGtcmMgyjX++6YDvcMVVGwNHQ9cUiA3UxlKG7BKcpN
suYrdk9DR9poA+aS6Af65TDaf/MSamG+co/P/6cmRNAuXZnPNbfsDANuaHtdpOV+XddWVZkybP5p
8Qm1UQlIZbp8cnB7sQXfH5f2Q6sX7N8fcbBaYB6OhpnI8GpdJFf+ggyrQUrv2y9JQbGJ8eh84tC/
tW1g3bpp9HC+W2AhAGzzgxSL8EBLmSF4yEEUFGo7qGXlIdTeD83F9pPEsiRV3/NfRps1N2htSFk5
QkX/HcHw9aXyHlLp/+nqJH456NL/aXBfJzX2kvu9xSRJ3m7L5YHRrWEq/LEU9WQcRZY4bjxAAeDA
0mz2lbROlbp9k5IzHwxeiSKZ+iGjRkw0XPEoWBbXPE6uF1DZYq0ZdLYFq9s8CpfKlkPoco4BYJr6
BlEz6z170hGsBnc34se05DFXDxbbF8SRPEp9bbYQq5DKg5vykriBKSUXLm2ej6V7jezZKLR++hgj
VfqASY+OWqbF0Zo1Xe4IcbR/CIGPDXhXSsKZIUoMdG2aSwWpvLnBu8fyRqtq6DQW8uxPybPNqh4i
8fo7027JDheENNKXeor/5XDPLNfZnCyg+1O9mMq7h+oQq+ntOkWPBrWz75YbUTeox+E6nccUW3RQ
ucgP0vV9LesaZhfRSZg19tgGgtdfdwLdKSU56mjcn69I2j2LJ3qDoux9tlHujXTrjbn/2HaD6Stf
RmDuy8Ydwk5l9vmf4EF8D6MtYe8wOUM5Fp+FF049dfi76BeWSab1UMX9MOCpuwMjIV+SuysWcu34
F1IOfT1FlRq3csgYZ99tkh295EV5PIIVpv5W5n04ykHj4TcUgS1GAvAyVenv4wuu+v81xTuL/DBZ
WI0cw6uSCirxIB/P0ygW+0Ms6R0oXVYFUBx4F8KVg/WhZu+pVeKLVZvz7RPCZ2s10LZpr8ZiGao/
NAng2dXyTFt3Pe6jbKwGaqVfo3xuNcQlm4pHICniZ170KLmUrRhUnIGhWrETme1B4YS9nDZc0wAD
PSd5SrNDrp5GDdhkCtYs9DCNFE4iKX2SnTuuJMrUXhWfZxxLYZnnWHXb6YjodmCyQIAsfj6Rr6X1
CqybeeH9j4a2S31xY7327s5o1wJnmcXV6hj8UVaEVPW2JvIOODcv2GPjuX+5aTleoMiHohmy9jT4
wmm9iQXs8ONsTdwUyvg5ANvvAbvujaci63iujmSekbiRIhSeG7ucyocAkwbeXQRsOujluBYADg4t
TqplbGY2UuctXc2JbESem7e8XXMD7Y3QgFrAxWGLbge7l2MQh32YFEPITMLznbumz09/Ub3rhoMI
0vrnbK3cuOpF30Gc0UjUeLR3kclpjCNFqp+IEHewz3mJBNrAF1GVAovPK7/UblYYe9VEHgwQh7Su
+jvSKEClLSc4NMG+JUWxaHiDFUB0l/lzozr2aopqnq9HFBZTGPF69vFLPstsyr2DgincaXl1Q1U4
se7UmfqOQqDX2x1BLqbO52gEYDJa4N2dfFwnAX+wIO4bfwfjCgnjZkAs7nqHR4+ipWbnewLhLaya
Zos8cCb9OyhQwGoHL8M0FG0V9NSVJ19C/2ao4aYe+zW89lRy+22TnATN4bVmnRIM4cbytxmLU10T
Jw7AoerTRzbEpu+/xw88sqCJr0ItGvnC4CtUHQSA/V3yiNCo960qfX/1KQ9UuUA1Eg0pm+LIIo9o
R/VoYXv4GxtE/XiN0CXIBwClAuJujCRCNSLoFiFQ7xkLUl9kPVpkNO9bVFGZR5YfrH3uk/Z23qE0
Q8zKIwH1EI2yH8Mdix3mtIx1grRbIbF+YfMWTyHwyIqBs0JP2RIWdRkwMbSqWF14sB40+x4bHwEg
uLcho/U6p8cyfULCz0Yajz1oZ4fh81gDrwOByLld+cvknn3zXLBrm30PFCrBYKqKwxgmV1gSp2wr
RZzR3sGshTxWaNqYAOXk1AM2Y7AgadQtnLd7hwDvmdh3ociHv0LUJpSRGtUZAos91qTlLX8upyw4
DLJh12VCvqnZhWrwLcOWhVCa5Y8siEWh330OIK6YAs+wLm2yti43+UEWtcKYHWcu7CcWOpx81Rvg
FTzqclZpndFljQjk0Dxmw+3MlTOw0wYX/eRex7UjAocGxYahJWfgSa6KQFEL5HwgouUc+Rxzf3HO
9m330Nk2vDWMCD3GYAi4m8k55HiyGP/y2xXgxgOYVOn0KigslTaL8Hm2jnmXP+a0nFALAGrLfwzD
lqIzqRcUJP/I3Fq4tYORwsrOjsO2DKnY1JsZd2fmBtzlOIV/s3eRfFY/N/84vEsRJ8YPZkD+efoI
2aWpFrvhGCjgSXe1uUGYUkNM5kC9hCLPti6C2jAz+KEte2gAMBtHSZiV601pU8nOYT1URQhQlN3b
T7Jf/5+y4fLGqhqKk3Nd8DU2J2xf/9rLF+2Lmg8Iw0hjyDZbJ5naRZ5h4KfSPlscvPlFJ6a5hnri
q+FAr5onld5/ThEls8w6ComIhHf0zVfOpw5OZRm46h2nyPq2tzdPAG1zSV+hl2L/mY6RuUdPsuKo
LzwZevnczh5Sx+hBNxUge0b8Naiy0KriAwboAdMMXNx2B1t+8Nt482lERW5dw5EyUyOuPYzm83YA
2wrwT/62f/w3LHGa+unoDvy0jXFshkfMI8BNXbExzXacNt60TtOtUcDo1MF65Ox0kSSe8x6a7/qB
LPQo1Ubt6aJFw9XgosnTV/7fmPipnTCxW9a7j3Rxz1BXBCEA3oaCpVSeuvNpeDkBxs91TF0WmoSd
iedo5py4fklza5q4hP6eIE8mczTHBIBQlNqJlCtCphv+YvMTSkAO+S+hHNnLsspsBWUMuElCa8tr
kwSKEuUYVE5/kJLBwcqx6WU02LmU7CH06ZPyJ1JJFL2KkqoF+LRpor+eubWrqvhAAD0/LQiinFm6
xy1yWNbR89SM6158iPbRe5mAfb4V5nNlEX0T6tCnkBZb1UI8HCIk117w1q9WQXHOAwmEaO8GhqHN
bjMYylrva0fb2kekL2BP9zXRDtLz21c////xoJiYVIMPK3VGb08zh2iQAhnnV0Bk/2C+nzG0nHyu
oiRIb7E32nO7pJrJvU/AqBFRx3HR2qethuQZQtcDe1g33V9SnyeUZCIGfnD/6tmchZh8HwEneTDN
8aJO0vmJCMhMDID5fRFi2Zyg3/9xTrMmnhX3is/QZjKBuEU+vYm0YVfOFgHpYSaJ9Uv1Kiz3cIsl
BAFdGBTJReCjNSA68+zgDXolk7mgjg/1p8XUIt95dwReoJcGEz31hpuGN4smlGnfbLuyL0P2V6gf
lfgkQUt7Gr1XSoGdAhVQHEKla6LiEGnoDBEtqe+XlYZ8srrsr6tCKDOBQC3UCN1y20i/kCNp/Gk5
6Q6BHTSVNhSOqK0MyToFYvQWnasIMCP9ylWU6SYL9v9JC+CJeD11wc0cteK85uAMsNBEVJaLwzVU
ttH5W7/W++AWn0aRGlHeXoeo3IX7rNkrjFwk68ItDU09kJdhtD+RvJ80efIbfiOV13e6GVfDwAlR
NyO24hZRUAdy6tIZtVz5b0r8ZDjhT876pQdhiN58jb6FYiJ58QhJGrz2hwsp3ndk4gL+UmnMinj8
TWi7WvRhBAgo/gtW9EKjfj0U2YslnEY1LkBZIVnoZvjwNFsIv2uaYnLGdCJ1dOh4KsySUpKAi2Hy
zXVTLIuR5GlbG1Ca1KbzHbeOCqtDjM8QGFS8r7Cisv5Iw5NtVfQRSvcBNXJRtDPfxWhwqf3oN622
ZQt8mjW9UWMZzUYa8VB3QppI57YmOBQNFrd0vXZL5q3FtsaCYPGLLtvZkdU0MTS4vmci7pXlfuIq
yoLwB+Sn78VLI/slGcDFKG4CBNYOy7XxZ9Xc40FFgEWm77EHybgWVGfZymLnQL/W4rTLRFY+6wuF
WxM8bIMCk9T4zYXAAe12+2DzamsHzhqax7i/sBmShtJrb9x8xJXH4CnwIMAt02bEhhCJawn2xIQe
+yXy2sbz7bEh9Mvj6J140qJuj8i52nf+/EXJOUt+RHg96clC+umEi0rGedkLxJawGQzqdfdqT1p1
KVjeVsZE0M1y9JOhy9gjbcWbxlswQYRRzKq9BEvVEJWnAA/Yl8nNOExS+rHr49C7Ll1XnTFBKZ2Y
6nS8rOi6Yl3OQyhtS+4EmA55h5025+U60QMJaaSD3dcz3QAzaRIrF46o7JsE5I9+k1SDaprurIVQ
0Q9PuoBQxxYthNC5jI5evV9b7dxd/Iasw8XyKw3Aa9LcyoSNlWs8pSSFpmhCHsfSMZMgCSUvGnHc
LdoKkNDcM1xOcw24OwxrMHEm89/VPRTiQjoQ8Xgsdw2kQDN3PFp0BYnDSl5WSRt1yP1DYrFGAKxk
rQx+L4PCRkcLuP55/EHn+yDI0QvbWr+bF8vouX/TiN8u7DwEb48ujiy21g+rEQw8GfMvXBH8eYX7
P7FJkuZN0QCv3HoHRvyuKiIjPiZNKWKTI4ROkwwpySfyq9wSRvDGOPIcy3yNN+qJ9KXlllmCnglN
xS69jCm0AjSKiXqM1tncP4YQP5SA7xXFjKGzVB5/msL/SPch6psB2QYbQaxS/GQEA6P7Z2XkG9nL
9goBbryh1D0Sgb8dEgEPBnJdQWWf3YyUNeaLdDQ4b9wRn8+D6OdZjcQo3KHKbD1++wm2FraBBCCq
ln8ssit3yMBm1ti0x4oq2EYL1kMMmovGvAI+5X1zNUUTgVSF/mvsSpshj6Vu5mfQsTVY3c7HYIyO
SB0hHq0vYew74Eegjv7tQK9CClKfwFlrslflC0Va5EMq50DDmDELVH3v/CcJyEuNSh3CaMLdURZX
y8OO+aQ3sxv8LLWNaai1ndEBzBT6BEeD6OEvqfeTZeMPveozeheAl0k4f91eppq3hxNAz9/9M15t
CjRAGNAFJPmRZIGt/6Pl76r8sZn4IM1biSW6ObCYvaoteuOEPa78iuz15iV9fvymJ4BSln0Ps7Z7
KfL2LrGGje0XT4lAEXDhdv+KUfz3ieDUjeYQ32ATumLOQUeRikmG2W1Gwk1iqBI2LEc9ZomkD4zk
SBgRzRdlUhiNkTkU4iueTTS+ZIE1MCOxkQcSlrNLON6FZlEEEQqlcdIvT38ENGnzGlgUazxBb/mT
h7/mCM17S2A9SefsgDMoTxReFHv0DdzYEFqkUSnwyvWkRUi+ZGCg7LKAJ19AdCg74bdZbZDBx2Ah
w6r49bmsRzARgUB9i70CJFO5SJpJ/z0itCdiovhbWJxz4d6XRjKSqI3WCZ7y3XsHnoGCsigDLNLj
puut1O7KOmYV/dle7xcq52Zrv5J8mOI6WTv+GZrtvAAMC5zRnrMnzFrIpNGUdxa16+XDSNUeA9FV
E3BoGk6ZgG0K/HXmLkmXQkEwHBi2hRsbOVA4ZAbwTGM5pAA+fOe9l56UDBGnQILmQdTeNJQGtR7O
2fkZfr3k29ZIp9gbIO72w6YfuXdql4hcoyfvq0wJHY2vMcOIFHtIJ9XdA4X5h4B7QEIpirp7EOoj
7co4t3X8/U6GpTYbH6cezGTgKyRllcOxtf8+I48CeJ+4FDwrqEsRn2BF1biUQVbBtJ54jUL2IGfs
uyp/W+07nrFLV9K5KzcbfJg+bll6+tXkDMiP7aYiMT8hPXXSGFz8cFiqO0GrAZO6yV9MIlDlCgR4
OYShR4AtFWctokJdymie3/mYeLg2nCHU3YdwrFhVLvVCafYAoCHCu18Ji/02d8I87p6fyWRvcTNl
X5G1ihqWT1NNxXvetcATcX3I7wNBA29L13af2GoHBEvxRRqww2SfTvQkoPKX8D9UQ+Y4Z9P4SFKC
M4wEjrOhA8rQxxiFPYSB6VmJl7olqqq9/cOE5+rAF0iYLHDvH/XsSkb9Xyl34Pg3JrKgPNgRkP9p
+CbXypqlQxSqwiQgCnKPptN4/MeQ5yGnVaNVn+8bLDs3LvIoJnVGMxZKfy0vaDZ0W9DgsDB2DNRJ
uksbK26tawILANBNcvGAO2zRHQZ26YqpV14B6YSCWpLSfjd9De+z1/dUxhabX8E4Nv8lwpIqwRqy
qUilxO2GDKZ5cgXBl465lAFqVAoSljxdLmascyJAmhJ34rCACBXj/yxWAslOJVnr2gbaNrgIbMFd
9CakznS85Pn+wZB+dzpxcld5KQRFgxoZSUJMvak6eObnJuWaBZWQpRju/A6bQT74qKzxY7MQig5K
dAuhqgdK2YOJ+MgpFiV9XRbJjHCC8TDdb0aGgXDAVKfFVgPWWbqDPri5ktuS6Yv95q4EU4CvHoQW
Gkrst0aaHf78ye9ZXOMwWoH7qxAwZ2AlEF4zBIyq5yKoe8FqlOuMmisy5grVYrOeB9od+d2RoykD
7tbgAoB8XawJnifXTW5LhBkDAQFsFczIV7NihifnqlOzpB3gZi7NkV82t5GO3Vh/eeaBBSa9QBFI
2hOc+xS/WPf/a0PegDX/t5qzrupETsKlMIz977gx9HuPpOBYtQYr9xVs9uIrsPveY/gaVjlsyrmS
PhpxSR+bxN/RW4xqXBhyt8owqfyDYJgXN32rdLc1M+LEtYhu5T6mEfRJ544/E0YQH6CwiUUZaTzu
2uobyZ1TL3VbajXOhk54x/UzdtUmOl8PaxbQRZPkEYC++NxK5+dF/rraNyqsHLl86ftW3aPmDhCA
7mCRYk92b/uw64+FF48VpFpEnSQ0RJw2J8Q/wne4fx4jdnF0O3IjkIuTSCEQ1moNtxNg8J/QpoxM
yZMHExJY/BoIwQcF0OYE8TjgFeds0pYoJe9W8gGh5wzcYlBFC88vpsIiOL5fMjVEEqdYPBr76P5v
3MC74oNzwbQ3nXFeqpc0B0h9enxHHWQ+dhSsm6TYPb7RpokFbaLuqkQqpbDx49Gvua5l1+GZpDVx
7fOPOWUbkVEpG3TfRAuwyb2vdnIe6wFTaCiCRUKwf0sKdEk2XIv/GO994Cfy1zgNe6E6nOXB7snj
jXize7efn3o9hwg2YZ2dXvu7Bzfxzh5l1VKsyy9gTeCqrGilMvzvw6MuRp8YNcT4qgoCnqwgPs5a
QRyEhWKBqWFi/ve48xSUxKqf6j/DyIQkMcmXYhtV+DfPWvAZ8eMlsEDKq8S8Dgkuy3xNaaajZzhg
JHlpJRxNgzkarKemY8/aYOaUTc/xyr67GfOST8BRRb++MS49Se9UgSaieiisI1sipdpypRenBRGc
e41dhw03ida9M7lLUn4ydB/mOSBu6PXPUegbqBZmLNZxA6eh6JR7TthcWCkn43DR0oIheIDxIqjm
q37C4h/LY2VQG5JAqJQspwGzML70LlDzauPV3KKBa68mQ/Q438cH8Iix7YWrWqAvub2Hx7pXYPD3
v/01y4mMEu9muoGoiQGcskm1q8cfrw+aebBQqOyS1dYdMrYt5ClctAjv2E/ucGBmZMB1O//aHPn6
irW5Hvi2uJen+VaftiVh7tG9wz+ijsIn7oqJyQRXtD7YFnJ4OqmC1F1NKeGBe4Uk6fSMI1ZWGqRb
NXcUsWfsBgp75kclsZH8G7exaqZRlfsiTtfjys92IhTWINBBO6pA09H/48TcYKu0jzqiV4L5r1pI
IIjt0bv8zS8ocMm0TQrJq1H6TJFwGgPGxYU7xXwvhjhSM0E+/+jBjlqRf8BS4A+BGQIUGJubC5sb
zyiLyg5vhNiZ+lshp4MlX19qHPqSgNmIbGkAomFCGQWeYbqPQ+E5l53fHZoJpBmAbncf4TXhNn8r
m6F8ZrEuYpQz5wnu+of0Q4ZfoYGab33F64lCGWL0FFKZfl50fw9U0S/abAFMSM3hQYhoFOfW2Quz
mEEe2OQn8qHoQjK3Dl2GBksLEolNhFSuykL4E6p61z6Hch4ZcEbdg5qLNV2J/8WR1k0Y3FKMvj3k
o2OX6P9p/OtqzijORxDi/cgKT/oVo4M3/REGoQilrN0bLjir5KjkD7He9pShSoXgoKi9k6TF95XO
k91ClqqTmzw4flKbp/ikp22GLwdX07SgoGNm6nm0GEkgX3sSKUCa9G/C0Sz6pX8RYtF/Cdwwh+VM
mmMV00XJ1KhrhXLYVDQo6TJ3CRLS23tz/ybI8hSjyxfoSHSTsqNtQfa7dpiOw0gWsY3u6uG1EnOM
VrpugQKogpizuwji4P3Nr1br9yuc8J1dr1gFDUaD3RqkAjmDxHGie0YN5bD8GDEKMm+UmItT8/qp
ooNQCpMm4wff+zrOfcCvdxQLltoy1QRUzxcHY+Hwp8SHhjpPwNioum1tOr958taSOzBf0cj8QdrX
Sopwudc2kBU2BTkL8GN6+Kl4aIt194kH44F8N+nDl/vPys/zuy10Xk/IFb614ugAnrU1HwKfeGqc
58Er2K2ATBLCsJM5l2G/eRt3nHAzQ/h/FPD9oi98bueMe6gv0dRe/QATYK02kRrjLnxLCn3kZgBQ
LMjkIvavj9UNn+Rw4o9sz7F90NbLaQuj/Z7t/Wf/ODhyxe+xqewWaUEqsbPYaJZXOw0/QocAQrDx
yjHfADBZWFJxLe2/pU9h2IwQBHOEefrzMvn7gk7jbZ//qMfUXm0MS7mKVnn+5skY2Q/dYtPHz6cb
t4rhmY6ZHBYIP+ASk2P+NQ9srxYr0JPyKXPZECUJ3f0SrKVPI5T5XV6AdpaiFnlQF+HGEf6XR7HX
c0BvZGIM/qOcGB8ZLZhewo5QQbPRRRh+nNllnVXMUdxlRTJW4vRg9ReVaophfzAWU/YvgbqOvuuh
enP3hwuaShzHw1982Uxc8BS3fJ4w22gFu7J6n4Je4SXaHrn8QnKtYdvIkcdHyuQwPMgDCxj97W3V
/djf7t3Zr5dJ2bolKZAHgZjw8mFcCl+AFWSkxDZMMiGhGkhVdk8YV/b1Z3deeiMdA48hxqHLGvM6
P8Y4U6r8HgVvMC3/dLKbJqohZvr71Ha2SLf6TewCcCaEqaZTOJuICljypSRjO8DAxY6/Wt+BhenM
L7nMbvnjbSD7BkoFOBH/Z1LKjbsZpAmgshjzFrGMJwV51HGbZr13ZbBP3LY2G9zj5trLpx3lyuM8
rzM/x+s2uNhh3IImo/Rla5sZgOi5XIz91yUDd0hGc/SIL0pYeWoRFrwX2EAK9Aa6nGAbLmoVaQLL
VSNjxNou986dD5lZXU5w6qXmAo6CGyt1tZuZ9RaodE01KdBRdVxumXviARX5eFfiQUAwrcPuoWk6
/Z/nKrEhxiRrlEZz2owNnPkZB18jAj4TXQTziRx6xVk1UcMScSKI6Tt+nNuLLGzimIcvykGVOHBL
TX8DJ4KuwVkYJr7zKchqab3bfvH19DnEfywNkh82a33VNBPT4MrfHpD8UzvotD6vYJEAMBdqJS09
1SPye49Z3O+8XfWMBYP/vDiH/zbzEwFPePrnSi8QcxSe9Uo9w2KKsrMvVznUa2giQ9jY7sm/vgmI
O9xUHBwfenVwvMuOVukGlIfvhivFFmD4RdEolULNOxLhYUaIec4hJPEUMsex7ypzC+jwsVnto2cQ
mF3XAGrbF8Cr4Uxevz4+KKIMvJVeWBdM9y/atk+w+yGMbq+hiPppXi0mA3purFBvJNebh7FFme40
Q22CtT1boJBGvDOFjS+xE4Eti7+0d4mG3LTGTtTe9Ay1VYCd+YuV/9xJ0bXceh5xwpI5KIZlWg/2
FqYP+WMIcDiA13IfKwUw4+cuVHrS8CqnwfeIaPVdalELgnGlgyWBbFzMYLXPvz86GLCZgjtq6BUY
0ItEeop5nIY7yOKxjqeIMT/XxNcVTqTHGR8BtPLXF8+/TBs9klMyeX7eeCW1dF6EfPEpdzK+aNli
JJwcHfJ31JyR1/HZ9TdAKOfrhVu7eoRw6/3yKjh9j1eDhLX+IAKHb78RodD9MGRlS6qL9Omj0wNQ
eK9xLwsqrgK1ihoHoHMoEKzQ7/sQf2WhwjyH5dZBh988RpqBH9YLgpbiqwfmkJgI6ygAvrOSIQb1
5P+KkGMO4QoMkKh+nz4qGXunrAqbyfKGj4Ml8jMHXE5xzZJkNCPjH8nB+jtYF8cUTsr9+1cc3ZMa
WKHi/Mrip37YuqczpYJL7BnEBwR0VEUz7JeJrc7sv4rEraP5AlsV/KNxuB191nVjKMPUBosT4YdN
WV60fd/rWaenbg/hetjhrPMXn9xrsNPivIAXKer16mMMk1Dy9S0YcAA+BgRtou0BdS6BnF2XnKoR
xihGpcYECjZf/ciEumsrLWGJGnc45gxKAi+PeuQXNWN5g0NoeEx7cf3z6lK/W9W1Nm3GG0ga9lfi
rdEr8B7ebb3oOpigofydMX6RoNTKoHJtKpBQIXhZvn6M3NW83V4QimxlYNz6QbLhh0OPYYb7yHVI
xCffT3VtLJ9jAwfLcvlSFbga9V3PGt+j+IPzq+Sqxpe9l7/POl2s19kUe3aj6A+PkEUyIsNeCgmM
/EQrecIz3WKEvgOa+WhVQXl1k2c5GX8mlG2DIz6OCBDnh3emKuFcfFuTVVr+0t4bSIiUJdJeFDAi
cwWmQF6ROLwoB1Sq3IFkTuX2r+OufSEm28omB537DYZXfZ0x8BNUHp0YZnK7uWkeJRdnU0g8w655
hex15LSw26RvVb/RJeSZOJOJDVHPKib9EXXtaEZfxJjsUb5n9XnMkUWpdgYxQubBFqXVjC745xtq
vAjm+8PVzzdUqZy6ZarAkHU9JieDQhgQdXaDHHOlfht5RfYtkhwmWdPjZ42dyK7fanfXbaNqbu9G
qtsh/A1+RlQanhh83QdIoMdeU6xLALx2XbkrllI7sL2Ei4IqYbxFYGSsunnRgqpGK76V8li1m+k3
KFGiOXdF9Ns8LLjD91nY5VqZbH/P1N7AAjXRu9GiL6E00tC9SFKVmUH/W79pEUW9rNw8wHuf5JS6
lsITa3pC4WMEAZpMFXInoYwWexXE7XG8jZ78tLx/KByTFn6HClgnSaiYbGNk/kK/1n5JTgaiK1YK
fWeuQLi6b9RF+uzncAFfTxugTBtq58phCbVznexbYuZvpTMx5dI/99cO3uKXKaneeC7eo6zE3LEO
lW1QwcNBc6wEQAChRG6XJ+Qg5VQ+qHQQP7JgqjLbpUsKIvMGQYg29Z2zmZTUNZH1+En8Mujrf+Tf
tPhRvPMAV7VYq0Lnw/c/wkbs7/b7umTdyQMV3y8zP/FWs6Gqko4sIdOxOq/aqF4cHY2/vQh28NNB
lvyt37iU9aG1zeUv1Ck7sbu06r3f3CGiMqLjv9qzxDAzjt5shjT5ehbMbsfxzqH2ZwDvVpttFs6b
G8351V2ismOOpB7Ntq12cHhvj9/w9K7p1pqJKcyCs09pQ0ApLB08s4BfmSLi5PNI22Q8S/ArWAw0
wgpJJMuJyPzj8+uOyUXgiEwP0KBx2MS2+UlNcJyx2EV3JzaVc3gYaqLMgAC4KZFdZ2PoiGeJVMGk
wD9psIZf7WPpEjiIA+P9YcJ7zbIb6g8UknpOCcejen/5ntYrRB7JpOmrxHizvpZkabdF+rH/dFIW
I3nJmtaDmPHzWudTDXRIRbcBnR2RZhA7U5XW+jcxd5NCBRxy76Wb1QoIAFY72cwcNsAFzruW6jzJ
4zdN8NyKPI6Xxhx8D68IVw3nFKJ+jx8pKndOdxbYZoxTNcGr/0YYlSwQOBbEbGNEXMm8FDZVloAQ
mZJPyfF8iNHr1DWroWBXAQ37fLACQFUQZVbpBXI0Gv8ukzk2SGSDgsUBOsm5DgcndDMIBhYhY7Nw
d7c4S3PnukRhs9l/av3DGZ+wnplVLWvvq/+Up7G51YQnjj4XLJlyCZn6ns05wTagIEy8MICSThLl
ftMIHI+IG1/OjM/CKmo+tP2nBlnVYXIoVg1o6aDmGMxCTifdUDMMD4WthpYGEiIYxkfB+q8mtAEd
eyn+FYx92eq9bbDUGFIY5YiN/0M9X1aVKdow2M/+tnk/d9EuVa+gsyT/sNHFx19fAtPdyiyMFq7R
Bns7m/v/HamfTlBvnaPoH3OsoDSbTZ9WWKj970dFqBjrMsxbp2U4OGVSbMW2oimU3Jmx6t/35OQ/
/tgVfH8NaMVHFI9UMRjyjMJg4XsVCi7Eyey15uEzle1Huq3A1O5zA+zLW78W/NdrDAw/g0Ih9+xw
JjoXYeiNjmrbsPOYr+RfRJUcu/vkMLjJvPSABLBjypt1JrHzw9WYbuBbcLuQsSaIMvAlFexnhs1w
EI/tU3LpL7FYrHVdd3IrdgcETxJleHCMIsE1ay9l43gw+gQ+CYx/CCDFF2UW87ZTo76KLNujdqs/
WMSEIXr2vf8/i0GqP+1hn/6cr4R30HYQPD5V45gNtSpT9zivomCsYPs/p0ZE0otNFfy49TboqgLj
kwdSSODXgZ3z6ZY5Zp5clB30VIb4HUCjBQds1Kah8+kpoP8U0Mm0q0bPLtKYskjxX5O7E36XTWsY
T0l7nHwHFl9isJtA5qYy/QfdUQ4NgOiyE6z2+mVBA13OeMqUJt4BQFnsyLlfkdzzBreRmfOPlbBK
XiUANxECitLkKCesiFRpai2+ri+SzQ9qw6ld0FArtkgbXiRJk4Fxs1j0mnEBEL+FBPtP9APrU4Nv
Zl7mB3MoJL/oQsqEYZWTdZzOGegfT/PfjtdeQam7R1NN91Y5VBME/zl5CPWUXPjLJXSQPYilsBXJ
i7BPTd6KjYv3vNhHPDb78Y9S0ckeBQWtlEvwtkUHz/ZpmsOMdfLpJR/LwO/5z2lsImeN7g2wqe13
lQp0XqBQ8XL/vlIRHVpFo6+0NZUgGpkJ/lJWHFl1oIu55tIbeHFl06PcCGHNOqzsU17XMMhDSWkp
FqYGpqmj+OMlzC/707pxeeosQZN5RPgzcmdW6odKD3NgNn12MQjdZG+VNaUXDDXhHuWnAdw6l3Yp
wVB9nn2l+X+3jeTAYP8mslZnk6Ii2P1pXbw7bEkPDXeqGbtdHkpanmXl8Ks8Gx136rs0hvVZGA6P
cpnUScBpwDu3rqGYSuwZpaQ+NYYXarB0XsVYW5MPjSgaRhNSvsHIFzOg+iPGzhoyrcUeXW/chwVX
xM1M5r7mzLJ42IQzKmtdUDA+jI9jQjVLpV7bnHZnCwNPx5XBRUh7J8fxcylygJ86DfGGBVfnPVkb
hjhdpQOMbDcnhUd2Ns7jmmkbdetKK8PI/fiQomTcEyrhS7y+PTxtiZvsSqIfCq8b6LfXhUOO5E20
3JO21FhZ3VgCUvyPRYdpJbnAlWo3eYzetPOJt/f+VOSOrlNEdypZQTrvLZRDWO638RtCA3QnWIu0
hjjkx+yWoXcQ4S/AA07GqpL4idHL/OJRVwARLi7TQzgne5orM0DlatIfeYHZqqyCNcmzVPkPL1nx
5DHu0IV7Dm/oE9h09BaI0WC2gX4QZXGA90Xw3vxqovs+DSnbUEaHSELjP0SZTBeq1jzXtwE+Wj5a
6UrMIGoWh4GTWJ51JUFIR+GcmU++hnaTtoxNDOx4zra2qKjuk9Sd3tUCyna/Ado8Sl970qkaCSMO
Mv2HmoTDFKIRIYmCZnLK0wGMuHWz84e81gbW67/y4edvH986Eh65WbO2OcNHPjICxbl95DwitNYI
tJa9WXf5LimwNpYIW6w/CUk54+utLSiILyF68Y4EzaeJ7UPDn5YzfwKNlZlBGH0ucRBbfyWOo+Wj
8dIlAoTKar+Ak32kG3Sm6jk5c/GCboFmzTovRdoamsgd17uHPNnsVXCCvDnXrJMg+SyEn0AVG2bF
gJouCHf0NfqM4gZD/mQe32fAtgEkhpBpeFquAl/3DbWx2QIjpGDHbIf4pNHJAwaZ6bvNfZ4gCE2A
kuN8NN8fg1KrqeYNGrmPLAI+kbMYFjVbhQO99+wUMyeFSl+aZOf3M9JuMLROoCMJ31yT255E4Jt/
AAS9cqa2y5PSRtNv3Syq/xnZzB/ekRFiYZr0+H4Cs9AMhg3Kdb4cRO6MKi32f0EVQXeK9E7nOvvj
J7/jAlNZdJut2PnIr/SCw3hZ9BcnwwNEgo23rNsMHuewrlMcWviv9y75JgsGxoEREz6zNVsaP4bK
lQR6jRmf3xe+UUokCdfTmV78XC5l4q/v4ndOXwVX4EPM9Cc+TWGDP1Bo+4iRtAD3evk8mAqCJntM
cC3dOFH+MgyQOSMELA39YedqVtH8rHufuIwepT0JdFr7gNTNWjN9tx1zQrknBRs5YADh7AVRduMy
xwGkIFIy+9IpLun612ooILqnZqZcZlxA8URxgFJzk+ohmn8CGXNbby4FJlFr6Dp46c4GKddvel4c
ilQBNjZ1eVC9a50xZiQCnWVFCI5/hV8YL5AsaF3LjlFozsNjQ9BJPU6dzLnUZ0y/NyJ0v+S1CjDp
C+tufRYlnH+YKn6TK5ymLGTO6p2mkNK8dQCvNBCDEFNBU9/cYYe5jbKxr6Yp2Bbtxlx+Ym5mggBw
8c8PFP3butwusFahTpAQaLkSWt1ZWsliXv8y3gWPA9paZsWIN7KEquEaSvlXgNddyG//YcP7i2rI
jrUiXcXz8rnbqS4MLm1THmYPpBViWIS2g17L9lnQj5Q0p6v1X5B0kClM4FofAZXQIzhJQrgZ0yut
JfpRpf+br88Izz100pTpmfSsZke/bFfjEf/ME0H9o/TKSlfms0kMhmfQE9GryIsDT6qgx0G6HtCb
SDj1Qvl6o6DIA6/82M/Rzb67ZjT7H6064QkYTWMCySUBPRruzVcK3nDOVQxPv2FdhTRg63Z/jl+L
+mBJjLqdxjygJVuRZ64tTsDTgWV/vFXqu29q9Gu8k9t0SJK29ujSrpZFfCf6RUtDAeAQhJSSUAEK
CUKzFKIBRRsYv9kkslyebXL0EQYWFcsMp+fRwOHMxZ7NC9kMXwvYIjG4GgDN3dPN+pXY0GncrtW8
LX21QgqJriOttOcKPfAYkK5mtmwGnNYFTBApp1Hv0ZbvKihkNAtP2wgkXgPtqme3pYiBOH0ne7E7
qnIYEH1Zr4KfznIaM1ej46br4csu7gKIdFqt+TZ767pUEbgONDYC45adKbo2Au7445pHwlA9vVi1
BoGuhgFukyVvC4MTqKs0A3TX4PBxfKJyiE7RNmf+9yCZSc3Msi+w4LSMPORjkS8DWvQEQU3snC3/
yifQ8RVGYhFbPZSVLGOZXHEyItbDIjujsuKE3OaNlfIVYYIerYG3fdJp62bw74uB5PS0il5b3SxE
91e+5XslUZADLsRXW3CMg9sSLldnDUefDxUNHzJxhtz78mHSi4OXiOlgahFpdLJHv339+QsttI1w
0VB8HYA3TTXI8j6kvudlxhvdiOpMBfpneNyz4Bko5Qz9NhIWjvItTUlzMY/rmfEsdTQ7OTEihhzJ
dgCq1jXIbKc9FlAOi3GWTsMVONUuromzOcCt/uxrRp/YwlJPCO8/3ZVMVJVQI6qnbCc/pgZIKfhP
utMMyNkAxhte5B6MHCAnZ5QxCM3k4Jdn9YdeH01IXNHq7kHA+akDsBfrn7IdAR0LmizGfzSneacT
9dLBDYMOOiyeGzqylAYgZCHYr+jtfPCiHUe+bP6FYoyBOQQ4TNWp0Gfo+6A+JZ/1pSZInje4oHYv
L7bLhhGugpSHr9AoJPubgIC7G7IQBf852Jsb4mHPpzLk01uSKnzADih44EcoDe9CdxKoi+jT0HFL
ayYeLrlNVeTBgSmX4XeTpQAuBoC48ZhLCO/jh3aOZbrz1rDywozc5lrrTYhO92TV5Agjc6Ojs0sV
k9+2vRoiCm13w/pk6EPVYukoS9KyBiEFMz1NaQVB7l3u5+HWKF89vkzZ6MNIgap/YvivTpcXfXiC
0eSiWM53sxmJBk0shgzmy+Y5a0Qj6jZ98pzsV14t6SQ/dOKtXgF4EDYcUBvMYvaEPEHDQEtSU2Yf
bXuQVOrgMkbNoLeYMQ7HjxE6TNFuhpmQrQlAfsIAGyeksTSVRyr7Z+PhpPq2giwwQsRUf1GB0cMV
siCa5X9rVy6iz62b1PvOHorPqgJUDBc1b8QTjRz69rhrQm1eWXp3KZ3N1STWkMoOAUXgUgbE6hSs
K2xghKO0625woX9oB7LhM/xgzED0KsoAx/Ym8bfMTZEP7JV/gABB66j8vYW0Yj8dpnjHNfSYD1Lm
gnyU1cPcOQvc5m0o7QxsbS9CTI9EVOthsp+6AB+Entgb3r4fzU8oJ5NM2x4GMmpXx6NAwIzUNCvT
UgKP1M8agErTsuA72bib8PWf2BrS91jK//Q1Os0iWjVN4XMxjh9Bm+jADKtd4XMwsFJEWrOXnuUS
egIzDDEm9Hkil0SXc+mN+RKD8bOCgeRfpwENpYm9MsMabxl57mrjw1SKBKK7Xt1R2ekTBeA1oVBm
WflJ6KZogGHNjLiLHkhiWRscmLJAAzmUflIasdgRUYoKYOFzg+gbb/IRNG5Qg8jgGupoudDQdWwS
RlEbmmzJ262fd32quzxEC5K7PV/WUYufna+FOfAWpne3RMhRacNfKDGyEt6qFWWJZSlG75A5Tz4W
ae4+qHMZLh8y0WnIjTO+EOTjYZ2AGOQ2wzJPMPJpoWDDYhSUjhdr9rnNdxJVwy42Sw1dvE0Jix0w
PkVs2SkZXvdWoc6Z0GGiYqDbZCHXGu1tG0G+Vlugj5YgQT+vAj5fDm65GnjBN01+FoBTAe97JnPi
6UgoTNv59sh7U0cDBfUelYk+zk44BUD0w+f2TTDXARh2C+C7lCMZCdGt18pSnkfoFtwc/4LKZyIM
c2osCHx4NO0rHMZGg2T39PAgERCxHOgt+5C5creuF+eKtnJuMOvM8eTdUhE3ww0UcFcVhgcnGjo3
nKkl4YffKtXmpKAfUwivMfA6lgVj5f+PbOh36JHVdSrED3ZFuPqx3fH1f11EGuZydtPjEcXzusJf
SZGsQmiyaClIeCJGUvb8mlxiMquq77HUt/5jdttWYoTaSmWUIITcV2o6RWh0FcAxHDGP+ebbOf0f
s/GJugI7BjLMHtsGlByLrtbm1uDwgVM2//1WHGkbrwUZbpuTL0MwmWxcgalwmOIQFLWns3AUlHWt
ZnbcM3CHev1gJtJfMCgxHNSY5xCYL8PiGXg7GEZcQSpy99te9GeZLklr+NgnlqtWIVe6XXkn1GwJ
gsD7eJCpxXd+qnrhpUr4rEb5702vjMwNVTfUUAN6ix6/SsRV6c+uoidX5OLeQYS8KMA3GDZdIG7D
O57O0+KB6HNV3CkS0toY1sjvQVocw3iEza6fRbnoL6AjJpOMKQJfXvM85lH761ciBNTo8B6xwVcE
bde7oVLpZW5qAHKjgm4m1EDhPBm1ck0N5P83H4mrTXnksRVGxdFBVulGK+jlVoi47EqOGGxTXZRT
fgWOH3yFmJyzMHfGZM9GdEiCSuQZ2WrJofi7fyRNeqzYDSHhYyQe/HA8DsaiSjoXoC+g9tK3tDzz
P8kem6i7wEULLd+1yRsfnpCl0btyrz5GHDBfzyJK7RuAt6WRC1gkg3CB+T+eJKt0rocPDql0AUhd
24EK40wjTfGZGQLyM1PsGDZM4ku+EuMwFpGdlGKmkVj9zuMMi/cb0mexzQUYeBlkJuLRffNhjEtT
ukv4+wmW8QdOFviIxFhUsa1Eds83CCM7vBOyRM3y+PymorMl20mmSXI+lmikennaej5MxziCieck
Sc9RvrRf3vHiNeoebx0mlzMbe4orCA75qnKloUtgprkx9Z7SBhcqb/b4kvxwHbue7GvUbQeBus9l
Z7ar47/nJIDvbblEoiSL4JehljdbisL1/c0h5D9PrOIws4NLf1gpgZ83Lf9DdHYbpGfOimnBgj4y
6WfMC+lvcLQ1K+bbEpXg/2L+cC05f94TQMGGu0W45NvneUQHj3Rs5VRSC78ylFrjrZBuyR4DOEUR
ZTi9pwFMfq2aXgT1Od1cpjY5mXYwZLbbJ7E5vsmFhMjqJHQji2ycwlISkBZ1FP32VHR4wJixA+8o
NtiyghBA+6FoUMaMwLIYIKFNKJmetSYTIOq8Q5jTGyb3pAMDNbeg6iabaCdIBYUsJbT8q6slVY/n
NcU0EIrSTOVJohUtYAf+LzQC4pl2KsZ0tduyxxzBqWi+2JHz3YVo/pWTNODEh/zHz7MzR+qPrYFk
xz+h0XjC/CZlzdNvZOHzoAdHJJbyQFZfCjlE4OSLhNpjZhUzd+sQFaT6Z6GNlZlA9L+JV092Op9q
7ApR4YMEkFprOOP5HK01S52FSQCLhX+AU8CQkCn5JF4RgCLRPr3p69IdRvxxGx3Qh27FxOeoZPzw
1q/W1CI9NqC29Oku8CHSp6sLqT/G7LF8+9mG18KIs6WYcJJ29Eb+w0zo4fPzbbGQ555IWtoq22lh
RQ1VIC/Fkqbi7o/96QrQVgRtOPFffF/otYHddf4kXc4S6QYx5/wLBgwYGPFbQZ17URBc1NT1Eg8H
BmYWeFIy9Gl5Jg8pNAkXs6y6V8AYAz1k8fhSMms6LqD6xMapSJ/XiDKur3ppuBEfQeXBuWEg/HgV
dxXQfThzvHKcpZIwfMCU8wJg6t+Vde8+0TwAvzoNuwTteb689vgiy+EJwr11t0ysGyl8fBwQf3wb
I+bKVM4tsepgzdOjg7FBY7+458wTQlmTWCyGxX7wXeui1qTJrQbO+W4iIbk9LrFRBIKyLp6I7nNR
JfP6dWTcRGG0OOVGDQc0XNMNg8TAkRsKnXrYNQXb/xrqOZCa6K3MSNcJtRwcpzdGXW81B9fns6+z
BrpnxbriS8fItFeuWGuEYBFbSNMgR6/BLdFus9ahZH/tz4EMG5dXcMD5DZJI0JdlVSbR9YsTDuXr
TzWqenj2FN9bNZ5Ku+7FTUbMYBzpsPOHyrSn7A91Ip4HEbDURMQ3iRZ/2LAU9eKn+I+vD/IBc+en
i97VDtcQBBPJcWzq1lUSkKFpEsSujEZGWNykKSBYMYHHGY02rUzqKjn/QoYz7JulWHSeDC80rFsI
Fm2fVYMcRUavejTspEv95ffMjx55b/3y6Q+9BHeC+rq0PJlIcol5IA7LugPwjs0LiSoRvRM/ZGy0
9CAYqhWUMf6gY5wiGkqaW8dryeifp/nXdR+c4Kdei6g49htiGb6M8v+7zeKmAcMS+rTqe4B1eie4
gZY5Qp42oxK/W30l15f2z7jOe772Bxc8vyAC1jlmPWb6ler+HVIlPp9hqMPYqdf+hHSDoSFB0U/Y
qFQzq6Dc2yfV2ry/5OjXQUMLMQS1mxCuJn77HacUH0hVxlk6gJ7HE105CJyFzUGIlw1MgzJJgn5c
17wpRtRZy76OiCIRTkHg7FSUetrGP9WEPVtMw1UcfrKBVCSnCBHhjUwAZaZF1ks33u/qJpahmr8Q
EQJ6RIh5r1fu6SIYGbqLZI/wKXL+a9CqeWPWCZcpTXwfA7Aru6DrJM/WRgf78bjkh9PVvAJpopi9
DObhQ7xc3SW/cUX7GYa8zaf5I88GXOTPAYUufwtGwFBtLUxjRrwNUi8n/hou/amBafMfrVGt6ln0
t/ZYUacxJxUL/eW6fRXxbOHS2UMPDfPwpWEtpzs9ctskL3z3aAk080Dj2/WJTVEZf9DeaRpDAD/l
9jcOWevRK5CQjTlvcMLE825LfEdZhRdeixnGtPW6DuWPc6cQAYyNqszTp6hIk7ESUEFP3hnpytb+
58IsPAEYJvtUIK8LTEPodOIM4v+6mNDieW55qA711CB42wRQLF+HvrYYpXd80e/yyenV0v+GRCmR
nXrPNeAUj54+55f9C523UhjoqmuZ0lh4W0ABVDc6dPMMGUvoey1TanTwXyLE0ZULpxDrULrsyx0Z
2F9u0qRDo1zd+aeWcq+8LYvdbxRS4qKrI5d/t4+ccWxQrhCJoVALg/ybfGAdEwl9KmXpeprjiBmK
w+TU6sAKra3K0UAd09qE0kLIoKtH+oHWhpAbvCH8Nn1CucOUcJZq+mJRE3qdImbHudAcOx0KusAn
RNVTMajxnDhuEAHioEcSyq6q6mnLepo/RNKYNhRGCIOp9VyWoTO41bj0cs8USDbsPyHvmtEGncA5
9UGmnr3Nwv6q1aQqhZKAA+aKouavHgQ0/4/rzBdm/6l8k/7mt9cvSTjhD4xJMX0qn3NFl/kuaq7y
VTbKCAOsGGPT94oAv6cUMYtD/f5JOATwR9cWaMrL88j8XZQcisdw0Vl5iynEu7VH5iBeKC07g44c
czFwedf3WhlqtL4+JqXNgssP1n1YLanFLmDkZCbtoSyvz8VtqkPlFw3B9LjZ3UdBog/w/832T7aU
wdfzGgZQQlLcnsx2itOeuBRd0nQ46K6WqPYhECg49nc3n4/vEotZFKD6Yv0KQBJEP+pB65ugj3+c
CuAWUHrj8tPbeGVbncBOeWHTXpaxdKiIPp+/5ei8C0JC1RkKaL2t+1xg3lH0hxaE6IKW+pZxyhNr
j1JgkgNFLhKbq6MDOh+ZBjPh7Qv+7K0+thTlCJe0AqBrUzk70gOazgD1ky5TS+fOsrAptbNXdrNm
jOBX7Htv5komUcv4K7uPKu0PBJrTWNhf+Tg/znecIA/OVRJ5tmc7T3FFcgRjL4tEgrY9Ghz5cd5S
uCyROBIKR0DWlYeGPAAhcRL3+PA4oAphEu2u1RF3qGkwJQlMcQrI+g7Nr1183zrDU1zlJqojC18/
xsYEGAn+Ygjpv1swAReG3X8DV2N0NTxixft16kW7NtEQiV+UYvsi9htIHYjWBt+FhxzI0+pKBGgg
ju5MHd7+RTChWFxtoUIQOsUa+wRtMhqQznibxiLPUGWh5m6EKoAD5E1uWJIi0YjwomLgrsz+rE53
N1x7YNBj/2NEBqkrWTDHV/7sIdid8JTuz6kFO80cb9V352onvJry6zQ0c3aMihvhSB6kQgFmp/zj
/yashs5ZGj4C1C3XaXhN7SgqVzBE53UaibhTVbLk93uZqXIxIZuLoYWLn/MnSdYbXGxzwQMiPYyo
ixPNf9Z+9iY+QgVNo3AN19TbKPpLIb/hCqkI3UXdZbFSSrKAmUTQgm3s7wPbC9c31TjBw6GsTSPb
l2ebCaxdRQbcXzFE5DKeYN9eho7Y0/gfz9YLHf9/WL4VeYv1J7zes07+CFf5DUa0lBAfOXc6l/Up
43MR0FOAI96zNCVVm3S2CdLWkXwQoyG858Q+QVbTLmR5ChGnXODShpWxLegIDlVG9pUcDlzI4s1g
LJZdQlx8UVEAyW4fe209pfcb+fgsgEplpQPGhe49l+I0vPEA0z5KtGze6OY4Wd7Lmu84NsU6tuMz
NV3b1aUeAjJQP5mKGXnfRMv2tuPoy45C1QDqF6TvUhy1ZW/2ksoe2RPtjlbNKtO9tNL0KnPRbW4q
ucXqobIBcqtuAXTIJRLEDB4cwgug350ngm3HfS34f2ASC4m3xt+FySIlEFJL6F55XTAIGKyVkAtj
oSxDGeRZOOhDk77qKQstCHLKjfo+ifUgeU2OLPFwR8h6r4aq0lV8ZsI8lWsWs5WoCa85KMzmcElF
4Xg8SbA5xTIfWqrGtBXezaQSx/fMohIqgVRpiUa0nkzMZGTZc/+P4kROCE8zsowDdSst9w7ZEIBp
o9P69c/mOtX3+Mv7wsidGjeloqNrqnSZ3tZKRO5Cymeyu1hjkyLX35IoymOJPLIxN6Mxzlo3F9nl
GgWz4gZ2fBwsJh/+I2FVQJEjC0Zv+fzNiLPvIHuIRfpkiCqOaWWWWTaYRM22EvUL2mOHwjKCHgO0
f7cGni09Mlj193H93toZFz4IR8w5dqv7cAZEJGVMD4pcihlzAjRB87miTIUtbkDwY5kqswl5kU2v
TcnVOhHKezFNRIh7HjT1Xl9ofKidQCJ61/mrHAt58seKpOqmUVWR8Ga/lTEN1rsnTTimLIDiSTsz
YfkP7yZmD5VfJanl6a82QTQFTqaQZ7MRr1T05qKM32XmXbNzInPPXoMBAhPGHsCLpJZxS6lwZ8IS
hlle63Zm++RqML0+aEvGsIZXVULRamXikc2uRb2ix8oO2V9cmBbQe6KnUYKug+vYHiuK4hVMVP1s
+BJjvNer+pr2P9920jq827QtyngTBLIHB06QlJ6/fFvlKchc/74GKqmlBnU5pR6M3BJyuq8b9Kdw
ea8hnjE3dxtLtuQfJCHbsoBPR1aUhpkj4pdZUyNBO/mmRqhQW5mbhLyZCMcnJ5t0hgvdT0ODt2vV
gSdPHpHkSq0ouzjtwTbkYoHaxxdW7D2vgQk6Q1nFc/QJVTgFZIh2BDgRa4RtE0UOWc+G3Z4Gqkrt
HQenKR47rujG/EK8AE5hHA/z1v6lvlJ5ZLDiG1/NhQuA1EKGJMSr+IDcuO0/fBHbtps/PrrlGjCR
jt1LWftcHOryUWpGl1eD1HgXcDrLmRaR7OIcXDuGvG+KkrRxJ33X4J6788p1pWe2WQ+b1otLk7JS
N/zfRl9pscIGSNGydhTUMKwo9P52CUuz78VfRi/e0mo3sJN3eqcGVGiER6dHWEn7kUPJRsUUVazx
GJn0X3KmF9kt5brPXSMp91rPx3Ho0EFPXSY+90Vr1tOCMk2Ry9nHtECzlmCBgpbBWiWSXCJvVc4K
STFHANZgMTRGwfMjTsV9xIEtPovzWkL7tE32fYMT8vdYUYABY0nk4/V/qU6mlBHsnvSHkkGQbMOd
wo9HHX59wxvU+1D7B4dFO9CPq32w/Ze2lwvv43JxzVMyR7xVgO2a+FI7UJuHH/JrlCSymoVcCQjb
yMIRMldY2z/ixD822AFCcJx9JmMZrNa+MZra2eDM35kQ8eEi8DRp0cjbz5vc474w/9EVaN3Dpu2z
yfZhllywcOZzA1JIFkA0ZlHY7xoif8Fqm9LO8aSbrfMczQEEcx9EJdmjjJJ0zKdrhMcCLNcKyzyj
Btp/2oOpjyfDcpQXkusOlcwS1Yn3GDZaXvFqWHcCa3uNmDJKYKGDnw5jt5ENiMia73GOb10N2A1v
M5Eynrwe8xV6tzRJ1BQXT4oLXrAr4oM6Qo2WPG8EWeZfnFmakgLiyIgcwk0ngFH27fugquNS6IJg
NMq9AN9F+3BEwYaf6ghhPspGj1hhPPpLgEPJQiH5vNRlPuLJAkuQS57lKq5FbXjqf15H4d7CJAFO
MI6c16QeDJ2+76yNgw9m41nM7S85Nflis9kqs8Ye6eZMBCw5GnbsJIfHUxcICEg3l0JxJEAccXE1
mUvWuecO+RPKFAgVF1erMDNiq4/2B8t2/oiITE3qe+9iqrdgN29zru3US4SNb4wjGqtH72aNSAsF
zCMtelQ0EVuN/9BbiRzJ1O6owW92Xhzsy65c/DxPZZrA4Ws2+afMez9JSsm+3UXz0Sq7B+VdJh7i
3CewX3OH2nrWM1vqmTs2Bdm7rPDfW76mJQaeppuDnOxwEH97pgUCW0N2HqgOry5JliXKB06/OvAD
FAIEy5RhYXKTc0nDwcm7kHuhp+n/WHRH7pZxcG6NJvTk03DRCZTFaUt9vZv26BfP7b1UZEQ9Sndl
bqant065dsUE358RW4/ivcOt4LSQ5F36NiS7PCbmQAQDKwGM0V75U3F3tA7iFeXY2EoBLYdHtDzo
jiHPuUrIrMpTFu2VU/SIhRyhMG7wVyg1LYopwVZdrAS+vQ4J0E27Sl+dq5U5sG7rH3t8dsq0Ofx9
eVY8Lwqnt61wzbS5eZHnnpj+FAhweDDaLyeep8rbeWnjgGzOP+fVdN4EvZRECqC0fu41IFXcIVDG
7qLcKUNbEk7P5c4T5A9bcSBzh0GbH4QA7AwV8W+zoV5f77JuOizayGit6vnNZ8f4CRauMJdm8JSh
1mUMDO6xfuGeDykNJUKnBJyiYz3gWa/wh/MQZFJ3YSlzTmuSZsYUcAoYtVr28qTGf8u+EURc4Lcz
owVMMjBWiNfoSqeU9vbnw5U44W07dMBYB+QdqeEo1cdnsDnwcDAX+osm1xsfqSffL49gDitCI19N
DAR8iTZNv40JjoL4qpysFJgAWG4gY7YVv+k21cVSV/nnHj4FztCR8geK78swj/+lZ0LPID+zMt+y
/aWkMCc133BEcxYDDg9ui1kLHqy+UqEqB7H8DEfvLNkvUvFR+ootN1ooxAPLwbRgLkbaKAcWxbe9
AEWUCDlKpLYYqOkscXJ9VbJef5alSAyvZuPtgGGaR9Iah28zOOUQi828enSP2ZRh2vO9twQcgt/5
xGYazQPkv9aiPDz2bvsz2UHOed0sGOh+5MSo13q7q0+iUOMHeMlocqcmg3L1bC3FP4MfswXF9eq0
LlNoGKALTgyBFELeGEXp89ussl6azqybNxOQLwX8QoreEXri1aVWWMfmyJXHSVWGaIRnGSP4/USM
HwElk++Dxjzpc98nEpI+xhy/quwNI4Nss/6GXjM9Hmvgw8WPSG0uOrpPriiDRugw1NGh5ojpqH9L
+1mvuU7NncwXVlaHFqlH2MlpkB/t4eaImxb7MQ7qBwa+JW5pdImOLs+orEHB4ikC7G5T894Qb4bS
v8DrQXjU8AppTDnd15cU9ok6Aak0J/AJKSThGiUDU0DrusGfc8mpzz+xNsw/0F4W9qkcubMSD3rd
iXNH6Phm69Qpe/MDL5xrltBt8kgEJ7c6FfgB9N2MjqsW/2/5rVd3uscS83c7piCGpjZ1wcVGjm0F
Qr89sNqRpKC2Ww4q/B4X0t0qIFqQgiO9xAOYc2Y4uodEGp4nmFQ1oABF9hBSqZEepL3rwzMJTtyh
blZUx649D7uKPtCqKrmAVBwTBjfdH+KyiCcFLyQKvrrHYLUeKPpEiNQoY0ATw7IN9OQCVwXSXSqr
/yM58g/Ss7+O1DetoGC9g1kCZTuRGTG4NDBxjeUu/3e3njrCchr3Ao/wO3NYMWTISr/BcXyRV1q2
DfO8z+GoF2vNoDjp0n74RTm9/LfMROgF92j07BNxJZGvq01mTEoowOij3JFrRX9QUh41y7/3rgTH
FxS2j8aOEcbJhZGTkeRqkBmMuiE/dqUreLGT8N+F9uhUnZVRXy7qkLxlEll0vmt6+Wy43+kmbPAi
jq85dNOo49tgjFRNBK6gEs1AOXMQD+KPF1YIvBBJvvviwhrC9oCk5AiEsl4Pq0iGGHeoGyClZuif
kpFBB54illYTpZqK/7bYsAU3j5L7KswtynjKspFMGJpNvSv0zRAGnnPb2AiA1G76df9tfT7JOkGs
0+nan6YyGxV5GW8ZrT2zjibo9gyojhL+lD54gV5r/hniui2nsmSNbD3jPTNo4oxgTLnWxIl96XdY
f5L5kpFYHko/eeAqFO6q1ITV2Ms4EONAvG5/0LQ4yYbEBhaX2DoBAcqhtgYDgHhALpGdIn3cdMEg
3KXPxtqFItMTbVZm/lrHLffU/Rg5OZQQYRxJIzrGxPbO5ba7i6cg+Zdx23XJjmtV0086K1CxgYGe
ULZetRi4sXP2duS+YrrXwZlKvEKI1KrjyPLxOXXLTaU99HHLDLea/308qYhBWHmEXLB2Hs7VBq8e
v8ylZGW9DLP0pLDcOUiPD0bySZLlGSv3AWMUqRWErEhH87Oe9MCC63gFpsGwwb0IT6twEu++vdP7
mDf1simHvrz72zWPCQ/b424srF7+yB4K+RNnh1aUYqRuFlq0+0dXUMFL7Q64+M9zg9875NR8zC4x
3/dJ1RcGMuXIKI65aEVEADQqXGbenTpj8Qgjro/wUq2oHBqvbUwYf2+wvte/M3yIlU/3+gqGmUtJ
sRtJVKSyHkJ6o1H1zJuoGaEcr/UCdyGYfWafPVgRji7mkuGB4VXg/j6K9RqgmiTbG8UWsMBHkhxX
YfnHIUnW9tLvYTUY+RY4rcRsDsx3rSKZQHQ2ygg3uYMEsDfO9M05o+OgkrvZIB64k5sVpYBmL3ZF
0Wsqpb0m28DkbPATYE3ER95rLn5h28Qqp9yStn7xyFFADXmLC9FR/WQdnjRwWRYYQWLxnHYaf77h
EdgEyEbqnzqSeAmtSPygA7n9Er2znzwV8wupvym+1CKzFIssCd5e7QZOS2eG79um+ElBKLFXsWXU
JRYYTz+8To6pP5f2KBgYZPHJ2UgND6spmL5KUwhvtGrT9gzCVXbdATmms2LoJLxWF1szEbLdxBA3
ifKhgIcUZYGjn07ReivwXP/GuYgl7S6rhL5lHawdHuCZJ+WiCl02/NP84ZKWC6cqQVpriPh7XnRC
u7pBvhL964QQJgIDTSMPcx+p/1PIZR12GZzN3L69sRYpWKWtcKAQEkvWKFRbkE8MGCCXpua3u/xm
j3bAolPtgxzmkKfVJ6wvK5vV/nf1+s4FanLWe4kCaGAfUk8MN3jr/26VQ7ZXIcWtg7SY8CHr6GaL
zzV25wfJPx/Yll+/V9WbUpBD+Qq7G4nf/E+x5Vhenr71Eu3g8Ue6WNwh859InOUgm/iyd+wep2OR
ihHKZdEAlROfhBi29+t0KyPPxdqGMq2ZE4pTaURmd9mEfJjiguBFikD0chBA3tlE8/txHvRL1JfH
QLRtM2jpBUbrz1KvGNn1JN/y0L7DvHSyc7W7Ecj/BwT+YuXTjEAcSa9wROVaKWb1l/iuO3IVRDCe
yWSxdNdZc5JQxfOuEU/B28vEqwkVNdX0lLiOKGDhsUuXGpA+aywG1jpUsXPS/ZEZOh0xmrjEau6l
yL2VH1Bt06CNzhZXYAIoGZzGSLdUXe/akD/bWW4SYjeKolp0vSTCNxd0oSql2cf9nt2GWn8qNE86
UTaVcRvYluk/LqGaX1V+tgqAF902vMkt8a5Z7kLNxeobDlVZgBXjZZceJG97234M3axDjCJLTXvJ
xoWrHiMCXu2uOcM5yiX12lmsBwDvEHT5xgffW+/B79Dus7HYPv6cN/D9uY5ajzMk1w8zScaxkkhE
6qDN7xj7BdYz2VQdAuJh01wNt22zR22PuW36o1WZlFgGjNuo2D3+ZNNssWskuHuu8KOkDY0O9xb5
qmEzIu9aT5/XAgl/ZTUQ4zAH3o14cg79cDIzMEoCkPHaM3p3wJm9AOR0yZjkLFHUdwcav8rn2Yf0
vZmPBFeqwduCMFmfcAN+l/xsGmPTatLiKVltnbuTyLC6Sa0Z4efweOe/dwJh5va3zDwvBqgLv8gl
1Hjstxiq5qqdz2dVIgSJOxWkPzE4twxRuNTqLqZQwwna2nc8jebBui1GNPnA/ZHuKVQvF2EsIF9K
Qp0wg0ELBVPsHwTISzAVPVWTGrX4u5vwa3XQeQEI03KCIqGqkDwOc9eE5gJbE1sScn//2aGSz9qk
s0WwdiPgOuEDiIXP77WkAFo3zrcRBqU6hQjWyShKc3+gMR4CB1eLdL+vaPnSrT4b6KqdsCtvnv7g
+/qHuiw5Py+GuneVBLOREzEc8WLOMCNfhQmHnUM5u0LyTVwG2j/5bcSTcBqiHbeAiXBUqp1nTgho
lNpfLW0oHo767eDWKEaR8s8qUnA7eOUBc/4eHO8Pi30YGQk8AnwpUTDG9V1a37UOmYxODs6G1Gii
l3sxBs0CB7bopE6ewoMIqoKCXTcb3VWZcP78zjaxZLzAbvOnGEvtLPvO8ns1KYcyKsBIZQui76Ir
FCNMgVBitJfkV8dPll4kPyyASkZtuU2UQi9wSs4+mlaThaP/ijfOfijk+rI0sPC1B5Z5uPkI+Qu2
mIYtrNiN5N9ElpMaR+j/644kJGHURtFo/6BYdrcMf9Ss8vvjPTdPLkeW0UaOrDaOQ2DVGGKfr/dC
GF2Ml+1j1jXrLHe7cVjunJZD/+8E8PlxWZKEAgAU1Mrs+gaTYbccAA+sVCiLueIzUq9WcGw/d17K
PKAh/djDsgiGyTrzZDQyltlWfHV+Ggbdfa7ekC/2phnP6hvppILJiSewIq+ZsCJIgPZvqhSAq4lx
dYMgHSfL8jSeW/q0issNs8wj0Q6+4aC9yWYkmjKhkcKM+w7TrTwnBoExNqEK7PRvnKf7R1i/sRgF
wBcTt36MdFqWKsNo81vv69kL/sHfx7CBJEF51YsdQKv92sgTufvhwZ/ynxQ5JfrD0tagLLn9Fqit
YiLYkJCdOY+a8ByqqKLwj5x9+P2dUrKvPGEOgHdUv57Cmsuji4jymOC382yOYMLVnHBQyrg2hLXy
5CM/f98JoBP6VREtAAPdxn8QEc8ACuRWrUNZib3KSPItVulbnp5tM1qW/8cUqaLwdPdjS8ixoLjl
qtZTMzFgh5CvBk3d9y1qj3uosxKPSFxCAezaNKQ5PqDV1vK9YX8p5wOLlByYV7DtVpMGaOZpjcrI
Qr/dzHaPOAOTMrDEsfp6UbN+Xrdzvn3tXcIQl5nWxl9+vZ0i75uoywAtVVdT0AE6uS2atw+s0XTH
Mv6i1xIdijtRlmdQLY4mwdYyBfaK/zkMQJo4dDsuJxFYKITs0otvh1Fv+Yna0dsVYJQZGDcVJXJY
XRZmvZ/4r5LqqvloLbomEj+M18Kqtu4+0k7R7DS+RgMA8/vmjOZOyMeHtepDtGyQ5LSb90aWs48Q
37z1ZpLhr8EXRfgHT3YN3OZYqyNQxrI8x7TO4Qmh4dlAFz7/8gXoZNz25YPor/nAxnkbkopHk8x2
YoSu47CFz173PIEETfPbm6PQJpRcXrrVqZR/mL42uiS7eKPwtmcmR+jXug77R5BeaVmnX6bW8hXU
S/rBg9y+Avl2Bpa22cfJkthWm4KcEXTwnnAXxHHdGTfztLPxcL4GjanxMwuKTkJzIrG3PVf5z4NP
BNvStRY8urJ6d7pxobyhIESDjGd7smHAtc6wfzuBOemedXVExPENRyZxEBRLHoo0t1JyFPaBJem1
CW7Xx9fFvdZOfuUhWgumeVS1r2O6ALL6vAgQ3tne5YstSB6ZaOLV7FfcsDUNdfitkwxTsKh/j3sT
nn+EXC0tUcJuBNJEXmdRtuZSgME+cNvsyVGO/7vvN6SnWrvT2ulY+w/FcQN6erPK6wZZKB8B0VmX
daVUBcM8+DOoP7O5n9m41RIbGN26hgJplN+a+He+OE9G6+vDWcosBqH59q85XbryEKD3xbZG4KKQ
MLILiK+r1KAvAoV9Qy5571BX/Zc9HSUfTlkzoaMh0xyqWGjwGGZHG6ylWbaM1uJjAiwLVDi309G6
/QIkj3TUuYdeIsQXrZNf2kp/oyI6nmqAKbtcMdT3PDHw1PROTrcLPXswVn4zUjoh10gY2pSeyQmj
emu0CluCffxihJEGNKfHQuOJIOH8TBbN4GmKd+/Y+f5FrKuPIKQUnVyC7hvGP/PYhCxIlnS99TS3
1VAj/fSmM1dHDsowNCFuxARWUseCHONWYKBwKXdqWHS6R+UUQHw+YGeEC0VhRfEDWsX4P/uyp1Cd
DudzSqwROKHxSw2nzL1nvyrciv/CISTwPG2qTnksb20qKM97QnxL89LXcgrba/hWiUGEU6a/P9pD
feALXZeaOtEe7l0xt8FaXcELjLaEb4TmgwX/8Y+tX7qRnzodjInySaQxz2KcwoBMwAkZE4uAlN2B
OQbjwSJS8ADBYYjO9m+uN0M+ZhsNOusPflnV0brDsybFySFLThSLqsqXO+pxUQovP+DFH+nmxt1K
bVp7e7XlFNA6rkxCd/ZJJULNyHKJePJ7G4Qaa37gxOYgOBf9+fXgUAmS+IqxNDen6LWTOKw2WeNm
pZ5HrS+12WxCf87lMLM6L/eED6dJiPxy8i5HaS/zfz7szcWr1MGe2xOUUS5BtqOforV7sMNI3ldb
KvwMT2qKBb0gizDFAe6BRIpzO8lAPeMDfpPP6keIAOxw7gd/gCek5+iYitb5annWb+6Kr+BWBUe1
onmmzawcAM0hzC5AR+3aEl52ZTUQ3pW33PjcWJiAX/6oDEtA5VfKUrXMWAftcfEiEJ50aC8gv9l4
86MjTXzp8tICv0YHLtphFdgRoYMTh5UOMBE7HIW3w1WB5qIiz2s3A8DYXfrv9YaB0FbNEIsm6ob5
N01dj0cIsqT7IeKlm9Fzy5MJIMaXT1HBV2IE/PnWUbUGQvRCLjFohQzAowTk2yaGWOCvSRnO2bBJ
tFdM7IZj6/H+bjEntPq+2LOFrs2SRkxOgwK0RV/Q5kbcXacADI+I1fHLQJXyL7/1mIa736qEv1F9
iAJPDSvH+1LMPAd7D9/hHooh+P8Ppn+kqT2Rm3gRzvldhQBvyBk4P4Oyg5nnWND17sqRZGBDeP1/
o43L/rqxTXaDLfEtEHLCCjtnUtIKCX0sAMQpGPW5ZgA4v1WK5LDoFlI0ohmY+Enw36+6GZQtudS3
jlLDPrtlr27kY5778sSWempF391nqJzIXBOalwjZ7fkgwcFOCjYHaOoILyAkOEouQhRiy9vdMC4Z
ceUDxlDzLBCIIT0WtpC/S4VO9AQrHmwatjtipP1WkubipXwA0Ei6QZExtfMkD/jpKhqHzSM+jRp1
RL0icEWlb2ulbEYqtVtiyHVuzYZyPZDG2iYEr129s6TQ94ZNNv/5GQXr9volFF8giPPst4NCMTcU
9ejmHzTfJQ7Gc+mFxFQZ/S888uwNzrZV2oTX/yGji9Pf9tSFSNN3MAqF/ur+Sy5B19QLn+o61otS
+IrPkFQXTH6Ng3sK0Z416Jc8257BZN6tSmATejBhvEb8cxlP5F93WzK1FfeKsKtQqiDj9nrtgt4+
WdvuidSn4NmK0J+9mwiM1pXtp2Xv07p3judEBjJDyTnDW3A6IM9fd8nWC47jiHDotn+oHYpjdYBW
GHOiVsuIbikm+ZPSwYY5PjhA2KnNCx4uEgyo3GTDWa3tjwHXFIoz3vFBmtjosGK9ZO9XRASvw9cD
MNz3zGbXQmCwj+dej/QelJQ58U3jLrGgVur7Ip+ShAwC329IEFJV15KzkceT5aLTBu93PGjafynS
kjBpEIuj0i/SyihgZzBZddwFVb3JYQDVLvzGlIKFk4wz6o2b8PotTHiwhZh9SKHWOuDSge+UfCF2
dI51WUfw5Wn36B82hswEoPFiHQAbn/V3xnfqbQ/XRgGcig+Myuw0LOXWILFdz2WrU2pLc7FfA0vV
0W5tdNhDy6UmUL5T324pyPUsNbuHVUoOnOpNCb/Y8MtOCZMiKB8Mb16PqgT0KoVSFfUcMogoc9MT
Q4nydcc0xOe0q9XdW3ZvRS/IqmM8p0EKu4526EiyBuDs/YDAcS9nPKh0yGRzkMiNCSX8k8UinPVK
B1tAt2uD4F6MhJUTGRzfVgiF0RwheIN3A7E+arNgAZmn/G/B1QIpbHgyxzrqKBosFFDaX+kxdwJp
YhplC26UUmNW8YqkM4NCY0c/VANixyhWz9hFrTpRhXnNoLKRSipX/TXWIN8HmHwA3YohqUIFgV7h
hp41YbK4ZtS2ytpCa8cnR6UkEIOhH0KmqagV0EoIbhlM/Ha/+BK6KHHLF0StUYcJrp6di0rRrKwv
JNNhEit3XlfuzvP4scIVpS6DLEBhVz8+Atskn1nWFrhZPg5goOyoWUATEPEQc3ThB2XH3Mcpwpd0
Zz+sqcWOURUpnhK+0Oml1jcaGFSQjcGX/GHqT6mmHXsu1DtUa15yYlnddUjsqNazkAqNW2cagUrO
ItPdOSrXUvr3PG6RJp9oYn+cXZZ4n/OFNcN3thBpvXDZ1dPirqliK9CcmLCzEtI5oVizGJ0H0UVt
2MPt1a7UdztK63CvjFj7SGtatJcMNQB5O1eMOBY43t3YHJIcO9D/duqw02WRRlqOS3M1pL+rESZR
o6zrfzOJRIxZ08brBa5Y8HLRb7XM9+jLjcj0Dz48tPtMXjEP7smIe1JR6vsoe45PXxPeKxUMuHPj
52hS0GqQGq2F42kcOmKU1dId+3aHU4aJ/UQ5fCj7xHmygbnn7LXqvv2yi7iCX5uMgz6SZZDYBAvd
hT7X+sI0XLcJ7k4Lfv/Y3dCEGnButWrpFG1LCD04eXnbiVJDOA1RXijGTc5zOGolJOu3q3Drq345
yjFitKTLcSN4CuiduMskUnhzwNP4DAlbfUUrACBii9b1Un54tnV0VNhJK4mpEmxD0RzCHj7Pv8WE
q17iikKBnWIU0pJDljq78LpkFGJfOulNHElEsnBq3zbBV3JFQhQUoDOUkxBe4RfWu67RUPzJmAog
lNhL+iev/iuk25S4xe/NYrNbTYCnOiXPPqG15pQ8t8/WKpWw4nMCrUXbccx7w2OlEGneWSRdNYND
23W62NjaEdQW8omsqj8NaytjQ1mfk3H42WzQeOzJxIRKL/BRb23bAnZLjs4CJ8LQILCEZPML3IJM
7cNM/Z48uiOAyk+9oX4RVbVrGNAHlxJawpDARf1slGLC5G3m9DR0Kit02lGmxZBv8W68Lg9u+dl2
a9JUSGo9f+QacwW9jlPZKXGiei8ME9tgKo1WnStVjItQQRbZ8WbL5JKm7WIQ99dr2HaqGwxp5BUy
GcUtxomXckWeORkvY7YwQEi7WGxNwbWYKicbG6iQZwqJFhixyBM2Mur2PYCsrjc3LqHFwgKFgCoU
8nLX4dg3lvrFpltPTBiMSsRKU7oG2WTVMXyWcNAHqYJW/bmhlHVn43shCh/kzQ7GYw/uz5//OuyM
k/Zmk9IAuUN/BSK+jYMTaQXOQrFQEUCbw/nocM9ypq3Yo0AOkya/ILW5AX7oAeFkU5n5sG27fgER
RWy2VuKMg968dXAsBURrlt90wxfAqBYwQ9hu3jIHW94qRZAEhB3NrWThR7+qCgMSTc0Vpe8tcxIt
YcmX6aKiaVNw7qAYN1qiXgTGeY1apHEvdKKt76WqxNTw7MCqXpzEcflfKx0OAvqE4Kg4mHKOjVEX
s3DIGaFqbJdtzv7aLwgY4FNOa7GoiJWHYLQS7mJWfRht6fC1dNiHCqOEQZuiSAo1lFLS9DIMz9s+
pSI/b+DIRNsn4mHjM24B1mRBCzapAc9CRL7G8PnSMpIEbJb4plnzha2/1ib7vKABhtlEHekF3Vi6
Gef2Df9KZPACFkvQxZYlyg4wMLVyk6xTEt7ZW2OStJpe9HOYHt9dBh+bMyy3wmUcvlg7jDa9+e8O
6ZWXfjIqmua2kxThtsXoDFjoutN+Yzxa751qU7SSNliU0LGbx/lerzhumGZnMhg1ukW7rwEH2/CE
RcFsxmi8jEb4DrtDVyWCE35hzzMgaYXgiB4GySVwUkoyJ0mdkVxDo2QGAXQj8yaYCpB0Yvbv47/o
mmBlZEiRjqVKkdLbEkvtEPqV45aG05lFDgzmmZtDOH/1V1T/HB1ygUIjSkivL009E4AAEAMwLns+
4cFYIKgafhazJe6O8SJriTQXkTWoWC+G8ijG9BHSWDRitTr89NSgirsFTXkKTyb2YbeOAbkgx8bR
lTQhjcnr/z6rrQKHzHE2g8vbeK/vMdivYk7qJlcnAJb9q2FjTQCZN9B4cw0lXXv17RLgnAKFM9Uw
ymkUyFnCuEvVyLtCYqB/VfhY1Hw2xt6jt99tSBsK2i3qlTqaPYUyqQ2w/929UiU62AO9dZa8RBdB
Gcty/3KmhP/B/8K5TbBo77WqV3l6XEt2E0Ojo1SnQF1nyw5YsfW5vmEzeXqJ0KmUzs4y5Dr1dQnJ
8HaG/QZBdkPoU9q01gPjjoxDWUr8qWCKPq5XDhg7qYlXl5PvvhIM5/yL7PXopQk6RkyDqp3zFogm
644TzdmTQcU2UMsv2OFHEijK9YXDGVxD/hLQ4WygAx81DbzILYa3mVpgsegHQvBvE0KJmDBd7bez
IVs9AClYErcDNfKiEbu9bldqPvAYZDH4qZa9bj7v9MzAttioJ7Owaa2Xvrftdt5j2zITqUjQ4/f+
wnTFzVysRJa+LuH7O7mQsixQgIXXfPZzT/Y6/t4y8K+xvxy+mkqU1KcGR0JGKSNwVdOO6PQPTlAN
/mu9xdx23X2XbuQqxdvBWUP+XnCZ+WPo0qBw7o5JKvWK5xBTfnz7pWkZr6QIjMtAy714Cki78/8L
hKX84TMIydghK5ycMrjywJ5xFqc+TmSxbkWiwkUsynyFtxqOm8rHUnrTkWq4iEbmu9ccJumOKhN3
Joqqgce/SvqejY2y/WYhjKnqR8fJWqlUMbUlugX7gxJu8X3Gp2zi2nqPyDaPz4pPIOwTN/clH8jN
GtJHv0qSNwkZPh/Z5xNGlCYaYG4kLCkMh7RyRk9jotnIlAnmGtg2WLhuEMXGn++NdKLL8qLg6VqG
/S2f9jx9R6IFgfEXsN2BZTvMH7ABCtd2hiUFUEJYjSHRMKzwgo1DzbI9Z1rsp8RZXH6WlFCa5smN
Wc1viIyCv1mi4wUGYYkVDVxJ+4bq0ngRC/6rikOcXvRYaR9Ew567gbw05bxijeNdgfbjMoEJMpv6
z7DiNw2Jjkk2KVSgc7veqjdJloVZWZiwGIEnjxHodFUMoymc8trG+ms4T1jITY7lofqW47N0+sVn
8HjAjuVoY+G962B/l+ajK0kORQQAzm+nqynvE2pCEZ9DVKHLSMQhabLi1GfQhUXMr8B1E21EKpAk
p7slNX91lgZqVyUt2mxCTITpaSo9eyNBGtgBRSqEiWJnia/bUPuw71OlUV4yi8gwzfTdR/wf7/72
GuULaEkG9RkdP+/iAvRed+U99t8H80VRU60/E/6Of0Tgfc5MgQHZTCXGhBaajFi+E75ve2VecyRt
eCxaURQBbRqKcVXPeFxbqK3pJg5sQHaFARhuWWYgeFRIyVvstOSrK2y+VZeFsKeCwjArsMA58rDq
A9yTGIYVPbt4eNbVFN+z9U61gqYRE9HNeyk/SzKHX+hz0wdDPPvMM9Cvexotel4NeiXYNcfr1zrG
mZvkwnTmc4zPWqTmGMLY93dOH8gXGauF8jro74nPsa9lm1un0hUDOT1LGZQ5iwRWBbNpEv7wWBcD
rygV46KBNA7Hb5fASA8AZ8N5YCryG/LS0ZioD21zsifJgbMr3uslkN6dHTLjQDy5kp8dQ2ceUcFh
E0xoDRXR+uns4IhDWwQQu8qKiG9GE5roJCMWEva9xMUNAdRSFV3anIBXDSPWxmlYoBc5R/PuVypf
2jx/7MFg3/F/RatSz6cH/1Gtaw1UDeVS4kQlANGxO6uSvVaFdKtLwDZFC0QrKPjiqpqtX8pMO9EB
QnkcgoAIBeGxEe8cD6OrMfj648C2NYWFezUQz21tFF6KLgaRgm6irznf9K7ty37hB9yGbSJx63yu
W6kYQCc1ypqF1OciMrK/VbPIyK1jghmPXgxkZ2wLu6P2rvoCnZLtcHh/guiTjeDebUz8Ujqf7Du1
f6+5x8An0NzOW92o9ARqOtRWMxwDSTyVR+9Efvl9OSni7B2RxSrjg7FGasWf/tHGuT6OE+1lIUOO
+s7OaWwLuwEI2jAlOGxjjivu2nQecIeo7Xg5MlCLixYm4+3Y26pEe6bUv2wWf/rgd0tpv2+TDATC
7VlGQuYQFGR+Y/Rg0um/Ek6U3RpkY5xohsJSfe1O1gFamn4+fHnGiSMwlNR0foooB2L7BnAgdAtv
mrFV5FgdJzdXXM54c00VxZIwiCqC9NRLzBqeKaasTgJOaBsjoQMrTI9AXUlvtjab4WHblnFfvzpj
iyzVTZLilnRmtPjdOk1Up9cwBx6AMhGnRIUwU0HDstNAEmozsLIg0n4T5L2+7pQC/uOQIYt1lSfF
XZ8pX5cdGsijTUffFy5Pu4Ie19V9bJog+4Eyn6kqbMO7SfaZ7v6aKcZ3OpbqAL5yKiXK+K4m1flf
veIeW5DulbipoxsC97yO0wuVyrr7MenkKVTNMjQubhRRKlYWVS6crCg3y2cOJTLU/oklD7uJ84Vk
A03oCopcAFxLvF373WeJva71ao5RxUI8lPbeFyE2w0VOgOOoI85YuUGDfng08ssIMzvzapMrBhsO
Z0Ez0nRkmeAJ9F3X5UWjKOGVuqJjWmgCPkP6qKywVrWuDPogomEJNZk6Ky8weUw1GCsLTd3WWJFO
rrt+rwKLVoCGH+KFBoT2ygE+6Eny3vZTzNQOpuTMhdQ0pRlZuNmkGfoMK1pkehkCNZGS4HQfdsed
xvjRuSUXVADumWzeos7kwjp5Kes3Wk5DP/Gak1V5JHns6L34nRrXev2cP2gXtXSugKJF83VW+v5B
/8NPzvA21d09puNE6hylFO9OVSko4E6Sv3uAjKhTYB4oet4EB4v9nS2ilZtnNerknFbW27ykT47H
kJ4df76bFkDbjHw/08dVx82d2wogCt2+tkb5rzjfQ+QYmZfV9XI/ncx4oZq0qS4u7LXxBs1RB4Fj
Ze72JLL5Y3OJzzoIWenks9w95n4jFqzp6bOByX13mz6IKBhJvNx3OSPdPZ7L+xoDLUBm07biOAVJ
gKAX44d9OmD1xF8r3WO2lSPhZWkaATImSC18IN5Quw1GUX4h7VPum67uEzJKfQNACTFX8e1gGtCM
ctPp7s6j/eywYCv2KxRfBm99+sWWjDAuW85pqZJ7/QkWmPb2e3tmc/VJiej+itt9VCP6ZHNIiqIp
k+X/JOF2KsJAt9ZAvWMYnrPz7clFi4dCrcJ85yDJI3i4oBd2U2Dniezva/J8togck5T2S8oHlKv9
qwr12fDRIye2zUc6+Asc+UWnHRO0gdgPel2smPaHNRgK3td1naT48mGjG7PnB4yOp1NEQqGyN9fw
XbqGQB7oYI7W5uMMfn//hjLHecnT68pm2XX8yLVPROIstFirKmqHN2b61Bk5MzIzeSojFEi2r6tT
6S5Bh6AKYjOqMGbVnDuF9NEuSg5HoN2v4uIpUOfZOHHyJuaH9htQWx1KYEWjuyQ5pnh7HXUK5AmO
eHdxXxdxh8CFVbXOtWKWqFis1EptzglPyy1NbikQF4D4amSvh7YZ6lt3MAsQq5A3XqUJ9r/tGaf4
YOaZ3NULb/fLtQSCsC+wIq1aRgXooQDNi5TveA46bgjfeI5oz59sgy3VNieJGa2ArtyZGHFQdGqW
b64Wk8OcI2Q+fQymIqK8zcqLoYSV1CIB4bTwGZQ4IfMdq2RdqM6TRFEeUVGEStS30RK7WxoUDPJa
+92a20rl6EsSGeQwc0z11tCC0hvnRIJGvvNZJjohbvq1PubyfHTEkWYSD9sPl13JL/KkKchvhzGn
9XoNYqPBVss62gvD0uanx/9QjRpV5Kt2PjyqXz3MDqgKg/Naxzvgi9GfsCXBJ2j893yIYXI5QpyE
TntPo/Olkz54/o1QbGsS5dhHeKvfXmmrr8nXX8kZ8lGQIT0O0VnXx63qi7Pv5JPo4NuZnyJpQrlR
+cdl7mFYwdKQY/2TFDB4RCw8+0cfV7g89Cd8qC4D9hJwgOmGP6Zf2ECnPQlroMJNJr6McB9XmT4Z
dIAVBrducTzChKDlY417OxakLBzOFldQhptsvDkQsZKUT9DbykhOQBnVsxC3rZoO7OMfYPt46Ex/
nItYmWVttgzJAHZJhDVce0c/oVevVwM2Nvf6Azt8FThXFihzOOqFvasLp0xB8NeJiDqQa6D/VCno
rfN/p+SJstVg641zls3qAZvGFXqEQ9y6XHo5XuzkwRHySBS7UxsyDXCT285YaxtJaXzoyHcRT7Xr
pxD1qHk+rnuHSRKcTnhUSBEf5gkYO5FPgSX+Zr+M9UYS37I0TNpszeEtrNN5QeolIkp7TAHxt6SS
BkeHtg9+vAIHbK/I2onI1riMBjKkk91XoMxVUKQD1BLXpGz9dy/+0TAz3Ky2EXx3YknLq6Ec5ISJ
Ryzvpjsu310ap2QOTZlmDED3aOq8kyQtIW56YYYbFGJZtTzQmqJ0T/tPAFnqRTBOhLuoQaelvUZ1
ze1jMsD3scta2GAVA7BiNO0pbbvwv8yGfS9RBESdGwC0OwBPA3a5EVZQKU1cBpQGLMGQOxJsMhgH
XTzKNMn8zW3nplgw48jddacK1P4S/kBOtb36Y3tVfU7WlWxiLzrgYUVeWal0iw4n3lMGawhtH/rs
2Wq3JGHQnvT2+riwsv3u0isx4MD72SzkXMZG865P8HG3QmpKfu/g3DWakwvyOqTLFWQSKtaU0bFD
QqzLGKlY+pZV/yVxDH33toVMDyMQ5dFW/zvFoVru8jvPDoOBB7+A1xHjHhQn64ueth0lUSoPZMSe
QmdO8uF18c8mn/L/kDawcNOVeWahjK1Z8D+XmJlUmyIRc3nLrUjOp0BgHjeWHpnivKqDxLfJ6x4c
WMDGLMt0AmDah+Tisy7JJxsCIcWfR/nqaC5/am2dwgvVAuAi3EsYn8i8CfO3/nhadWtgMz8XunFo
ll9xW4TuGZ1z8xqFlwhk21pAaoLYdLC3TkojXRCpCwcRC7ZFJfH+rdCulj47SRpsmtIAUtBpnasy
N9OOq/j+lSGVwq6CuyYJ/jXJTAR5KUPivhL8JtnnWnpVsdu+nf3+/qGHB26BraumkzO0QPlQCriX
t+/1fKj9v8aMpeu30XGThzXWMUrJSQrSvkFln+R5rhRiGavOcCXnE+m0RGBUnPvphXqgbnnGRGtK
8vSMF4XeSlYZ6mWM0YFQ1I5Rci+Eqa55C9Ep0TU4lx76M35CXWdGlOKAQmbQONuAKPRelKry6voN
STx0zH03XDolMckMMRF9vwyZxiq5AVsHU/aBpGsWilxTQmOVgRV8MBDNPSoSCDx+itxeniQ7Ba0J
9Sj4o9azNuQtnObttnqxwRd+QN5R03myXJ0QiRfUGFTGrReDDl2tjLAD4DruPnfv3g2JZNjvlATw
k2nwufTqJkGKJWo2MAEOE+uRv1x32obtS6MMzoajk8uEUyhqXVB4gCbkDGm55wNajlG7ikUfnYpf
3XCHluD20oVC2jvYeoEs8avnFj0msg8cvWjjkEy2UhPzXYGIHckaETJHBw2Cjn6RppTq6KWDtTCS
aa4zGdzr17PeVxSHKBOkIIGumCPbov6/WdfaJZMSdlRgbtJnGtJGLIHOSIl8Zakcyzh3+9oaQdNH
g75nh29ap92ZMnyNzy/vwXXSmG/9C0LseTG+jbTCbJTlAEparN1pP095PFyKVRGTTGaIP/Z2lU1g
oXxR3FvuMpX3a8oMmYG+rt9ymEI1kGLPOPHF7bf35LvtBVV9H1NUjpcyFVu/0fDL6XebsrGbtA++
oxiONLUwesUru9b3ef7TGND2JsVJQDj0XDJhRWto6nc+9jX00VlFQskF7Wl71zqG8iOwfx6iMyH3
r+pJuSK4c5g6fpGFwN+ilVJ0P9HSXbo/iIOdk9mSIM6sxHz5U2b754xLbx0z1V7sYB8Gc9BF1szA
iiHrYUadnI9YeQ6XS5dhH5lmFRgYItzM4BRX10o7RftWY+Bn1hUukvYuC9oWymIxZcloyswMYWqN
JZ0Y7wPQU6B7DO+Wp4R/GetvlhkwaLzRaqP+1T3rIdwIAvsIQaVTIlN0zcJJk+/2KLSQgqonc0Ol
FKS3cmmJb7xVvpW76FNqekOIXVK/LOmVEOgDmTo8KAObXOeNhVEAEjZcgYjcnTet04k/8n+/D+U4
ZPZMHKxHFd5OfNcAtXXf1Jbb1JUYwrnCJNiQg3cyaGeO4i/HcqRjblVOfQSLh4RkywfNi3NYa1HM
yF3pdnjl7ySNfuLsnOlLL9aa0/7mN9yXbkHQSLtFLAZsWcBdIV95GKVhc1kNLm7vMk6dG96CEqO8
OvwfNnUKz6g/skDSkW65hvVxLZNHxbBnksZvpB42CiPM2cv0fXkUjmpmAfxWwj0QV/GSXW2rJUnl
oGtYKqCWranI8/zrsuxsIf9X0j0+RF9ZZpskEs4GS79ye85cVvYEi+b4YWyfZ/XPtqsTsiVWj19R
J4Q3HYpbo3QHU3vKVvp1MvOoyFu5C6g0A+mA7j0AjdnUpJ/+FpTSqcTJ8Pr/bm3zPeXIxvSI0T91
VPt0W33bwFdeRy0MzXzsnIQinSmkxTgxVuntSnmmdWLMGmHQq7pAFNiqOiFubO6AS1nyGbffa1lP
D6nyE8iYHEa+0DU6MlWYdHSbZELYw8DRfQlXardR7F9F1B/gMYQApShpkObVy4eNy+6iolMmMJtD
OCSIDCSuBvrtVFvNY75SiD/bToxuJYwti+LnR8AxT7Kite70eQDskV2xGXC3MC2bMEfypaCoHMXu
CStbeLbmOZxo0J40GzsYZbZ48BCgaj/Q0mnXqy0cOT0lKCQC2ppVFMoxdek++vtq97lKobqo/65s
wRUQjwpjNQ4+nvgYO1WYXZ2dajKUsVdOPwDo9uwM1iDyBI5a1Lx33BnaPyR1tuLHXjj54yBO1dCm
osBCUijjinNPt5rtfSq6F69LuvNN7yi3/MFr0rl82DIIkSeGtRnLAIybGHaT3UIid1QuTxTs3NZy
rGcdvnIp2OPFQ6v5K/2w4CKtLn4BbOEzk8ZrBcp0Sv0RzZ2QKl7RyCVXlNh+IR9Q3clTFtf2/DRC
uI8e8/INBlEKA9BYUgo3SjYP0ZlcozXrI5Hf2hx2nfQPMfi9nsGT77GTTKSB2APS7wyd7SgTDlyb
QtB7WYg5JBCmQnHOj5fzTSsr46G3ZQaON9ti0/9u3QaqeddT1RppiBLVQ1r5dg/wv9rUQJmhY+GN
7KYeQ/oZZDZvpBPVdYJFGfK5pzsXbQds5onJFWWQSju2VNYNDlG5yUryB5G+UeiIMieW16aFN7fI
Zc7KbGnQ1z1WXhaoNoSbxxQAivi6QD1URoBzLkI+tynmbZPOOQP0G9aj1Eu3jzoA95TVjipBcAFx
y9qeJDzLsGb0fXUZuQhbNQPq7al9aT5JHdmXdBTrzV5rWHfmIKaY7zpuENH5OQoVu1odC53ofxwC
M64bsmAVFlMJ8aaxWkfAPk6UkrhMVcdCOfbo2nlRQV7TyYTGozdam9Y+rpXTbOu8eSr/YWQxPIxv
QIZfARrT2btH9NXqmuf7MxAOiHgXr5v7QN0aOsp+TW6j/T4w4A3LMT0zCZUfY7YlT2JAmVrmX/2f
Y1/pzgZG2Gr7OPR9XN1to3sWWRXz9dMI7d+LKE/tEB+rxcGbRFu9/lhvn15KoQojZdRW7tVpWptw
b/xemFWLqwVx6valH6MMuuB5thdUCNSXyIuLb6Nl6gzEbq/ThHl/nBfKe+PCUASmWgyZwp8mlypf
7hJdjvk9FXpdNvTl7E1hP72zFwIDyhW8H/b5xfEyBvW6wQIUZtGIrIPmJ6RBsda0xGg4HyIuZK8K
xa/dsjYL7toSdsaJ4Vq0K7jAump0htwYD6TCc+cT4RsJ5HcK0uE18NO0daEHROSPVAQyUdecf71t
wQ3vxOJBGR3b5hGTQxr+cS6M0AH8bC6Lc+fM4/cP1T0N08+eJbG2L4mOwJ1xGBY7RJao56qwnsyx
2sPJAGX9t8kDmCfGR2p3TqGCgruwbr/HnewLA/GuC85U99srlEMopquiUCJNOfua04n1DSrbw2V+
E35f/Bllt3YwrI1e6kSz0z/jv/0vAeztjsXMrfHYvadbdUZb6FmHBAnnbTtxeBQknepK1vcgybxw
2Mxj1/LDkAytV3LnuMZWOrWD79D1JSFu1TDFaO5nfAPR2EmKbzcJi9KMHeySUjofiVfPErDyIzma
ZU1xnAErvNfIqXgGscmzR9tbuoIqieKbz/pDABXmt01o4y8fIaKQ4RarxLADZUtzoBKnOpUsudS4
Y5KLTNqJYzQHmGv6NPh8dtkPvJkHaMyzxzx8wS40Q4SUGpoC8lPBPmFuc6PRaouM0m+IHBzXzLP9
xByiO+F4z6aU5iK/qQv1Y+/xqTjHcqbgoC7G/TTv3X9+XqIfLq7/tDCWXp7bwCmz2bURx153cVK6
wpTSi414ML8lI0P1WDAlnWdKBm+uqWVNhjrerUb8hWpE8Cs57ev7iKSmN8/1A0ooz6rEFXV2aPPq
lqkcUXbKR0MRmt/QRQ29cIIoeO0mEZiw59oumwaNdvnfTUld9HPnZadqF4t7w/FpN+v5KXcHbnnJ
H7RW+BzRH1iGM0Cb2KETQ1+QKJqXbTfCQX4oQzbC2ByyoHFGkEqLTAa95cvR0e++6BjofDR5d0O9
80pirOB6xjjkS8PlyneYb6ZH+6BwtjP5/kVxTreLV5qH0DUnm1FZZZ1/m0JSqiyHa8UcUjI0gMf1
dqd/72PO1zcFn5BMRQTv0V0fKWYAgLtsbRI3+K3ADSANS4ALpowp5J2b+VtQdL+Doxhh713TzO5n
Q55zUg+TiveQoausUEv3qKLzj/qtkpe9Aai6azar1YD8xl+ilsZdTY8Ml1UH5UAKROV162SDMDnD
ZO6BnvCMZSqszA5n8io47E1z1RVQEbiA7uR7r7ja3+htc9IIrQVSGH/qyK8jyOWsDKtvUk0ynioV
OJve9gLpRQMA4puEJCsE0uoSVq/p+ACyMZiwEdT480CHsPG30CJhO+dmvTLBcGUJwAE92wRWpFlJ
raROoyisosAH8BtJAi1knxv8VYVOzL+wS19U2KHml6Rvqtub8hpvF8fFrDe3Kq2ir3i17PNAkJR6
JqLLpaWNMDhC3FcHluNH6yf5itxtQRaj9k+NS50YYIxYpi1buv8nPMtDg9lwtzzsDVS1LflYUZgT
liUHZNFcgRcpmtDdMCTAZdz8pYZth7sDvco4x77LqwpxX0KQhcY40SS7GeVtTfELnHEKfB4vVM7e
9ljiDe5fSeJ0Sa1lJyXPu/OpBLtERoePdNh46Dj6406SHwtNbNy1AG7L3f6MbWgpzYkxwcNY9FtY
3HsKDF3y1Vz7rr1XAXdqqzjtqOaVELrPsK4Y/L8F5gwUxIpZ4vAYGiws6oGQcP++f35BFTsmbOsd
Bf9fdm1J+pwAWsiWuIwr5oOQ6kMTnz1eXNwF3X0JLe2fjrPzsJ7oiArFF5VNwZp2hfGYzglZPYPm
0D4x+D0rajiZEJdgfESgxf4cq1tRfnWbtNkvSjw8eWQsp4ca44qG7YkQ750DOmhR5XT8B5FoU6gR
K4M0lZogZllyKQYD6P3Kpfv0f9+oPEmk1EZunF9JLclHvccRy4V3d1BDYx32yXCqNe0QHTbQor3P
cccMzylBabmjUn2FahbbwcfCZPnbBREgnW3KTSeCqk/0gjBa/uaNY7N4zlrbEcIbASMVPzKucX+K
tGX9KukdfmQnu7AodHP70svz0vQ/M5Lzs3fs5V+W3FetasKQdLSc2iQ9KyEehL8JxCRbg4HQR8r5
v2BzD9Jgwdd2IgtrDTsawm3+j+hTGmuRA7d/bk0b6tcKwto6ROhUtJurOjSVjrH+UY7vac4y6z/g
GVU/ejrY7h9y3XMdByu9ooqB7X8Jjr9TtLK49NgzhykB/DNnBHOi+VjWTvmD8IgsLUddCgmUHyzN
3ip0ZIsTbjwJWxOZVGmBQ1pRk+lBGzOdF+rPSAjIHrXBEZS/anDTpjwS2W9JjSocOUiK3ydy12PQ
MXWXiAKh0VDjQrmN+ma1O/Z/Yy+qBHQ/DFse9LIvvCwI+SslOQvWKblxHIGwEwyeNzHerOXv9HAw
bjBY82S+YGJFCXzKMpT1AXoL6U8EMVtgXeNG9MfHueePNCTRfSQoD3Kqz5vM5ARScG/zkcPKeUlr
1u/T0ZYRK1LmnDWOqqPwgY9HVT/p6rqhmnOTYiF5G93fkGQa6ageZt9AG/NY761zCUXbsKtfxxbr
2wuYldFr2rXAjFlRVpGnJitfkWwIyAYVtI4DCeJe7LZoM/AQrDbxjMm0npGsIszII76YbuIMnICQ
qR9Ptyw59M6jOsMQy3YENRxZy8F20sfoBgLc1SqnDiLPwVRkA5P47JL4kqw0aeGUupRVtNXDgsq+
ROJPy5TGYyj9JpGc/oXGp6MZMi/WJr/VZ06HBarN4+jLU786vJ/sfUCgwMh/nZ3jbndCkpEwEdyX
o/lcs4S2HhKPjXOo1KDnUemwKTqrjGNt5WM0aySPk7WsBB6VIQYZMfXz0FHqm1ctD4l4e+6sTkaz
xS6j+UaBjfMYs+k1RUC8Wt3AEmAERhwV3zlkvU2aCzUQEqUYCCtoJN8hBbxbNFnMWGTk9Mnx5MBF
EoIItlFvfi7leGk7t4Riru7ZOyFsNla/DG8vOrMOn8ddhQhjfpomuENuuSSURwp1b+heMTgrzlNB
KlIZIb0gFOKT/kAC3ZlfDJwcBeWd86Oe2NwjORQOwczXykLTAPaSRx0/x3DtRTmnw/CnR7X0z/zQ
7U3C8uFaJZH/CQmmwyWcrMHe2IZclCqUsNhrEr833zmggI0rU2pnw1W/uh4mNlg+pgxYbBk=
`protect end_protected

