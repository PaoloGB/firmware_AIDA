

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
j1+IbdCEjp9rON6GmpeUO5JwtCtNnN1RpPJWXPb8z1VONUriYeHT6geUliT2kj3j3ruQooz0qaip
cnDlo0luIQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EPib3HSaO2+CArAeOvemjeGUyGUgxzMbveLbA3orGi9nJ0JEazCwIPCLYN3/Fp6jpmXKleoSy+Yt
8aVlSldbRVUL0JefBQZLZTD12wkF8wfBQE4Sp2pdDWcEHIgUNVWl9DbkyIQLwYHP0oTW+0GVZwrJ
ZCU1E6Yxf164GIujPQo=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xK5iaFQJoJv0kMguY5xUiPaUTDqZRMOZH8/ZB1Yxq06eRqsbzZHKmtGE08xScCZRlnVLo07S7cyH
RIMH/BqEnGQvUmVbCRTGjeUl4o7tWcHHIPT7lNNmhMmPxgEJyobC71LV2fyJ4dW6SuDHvP1vvVE4
7qTX+iIzcBALjrVcJ7M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GvBFNkACpZSDf6d3aojglxv5RKUE+B8RRKiNrm7zUWZctVRoUgnqpA4jFrIulgs/o7tDqWN9mBDb
/q1cNTL8pn+ZdOCA6HTziWecOxCYCUCd05u/Vxp4e14C7m5co1IethhXVIP4JtgXmF/SDla3WE5q
uIJzYn6zdwgJSw/7iNz9Pd/+0vi8THHdMW1+mm0kUSsYmtTwhVGpXHiiWb03ht65+nT+gwGM5iFJ
nzfjybmQSbF6G5HKZ3PlbQAsYUk5eFkKJRqVLf/0XMyHdJK+9ZBUCOsM8Ktyd5syTAA5chBzULB9
lQi8iw9dNvGUbFA5FS3SHWwwSTZPZuVVkVWOPA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rgmQKXOffXLszxMSUgYbFQZ+rONPKKXl/cfmAu8056ONyDKGiUoXTrjW8PjooSi/Ud4/7i3j8v35
RjkT0tmK8Pvf46x0y7TIS1SoKTUOKDZdb2rt3k8TO3qZgW5nKyaHrn/4xAlTJYKpUChEczmgzwjp
Sz7118D3XAR7XuB33NPGnKLWNF6XTiXPysTIYvAUfhtKqXqNmvE7P39ewWO1Xk2jXBqJCYgyxHJp
ExtLkmuxpjAWsYV2ruEjfK29oWd6rRX3RhNtzQOuAuuf5qOSJbf8elnfzSQYOi2u+kcawpUMxDXR
5JWF88ZQFKexPoKVVSRVZzZXo1KKEbKFBqsECA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YkiJ9jZYjxcmbtSRgqPcdSlRRBRe3AGVv150/BYf+XDcHuK+xaSmOYiW9EOeIYH/CxXSZdUt7CQO
67odBlUa1pIQdO33H8JDlfyt1d4rhnZyqpb9+ZIE/VSi3Sb6SC1Uy1TbW39KvEafDFBCkKBaRyIY
QU4sWxqbXLS2y8GktCt/6wHpRzcW9/8DE9uFzDA5AaYzLqMMgFHGihcIrG3g93C1JExTkj6GUN3O
aWtzydUOoE3laYAcY7AbZzdQHUjaATzo9ki73FwBuauXCOi6aak7/MhOI5f5RMOx0Xmdt5lc6+Ai
jK1AxS/deBa9TULzkyostDgQ4eAdNJ+Bn49b3w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
uBIxygOUKTacvV9Xmn4qE7CPGF5QA5CIrYjzC8SPQpMe32OH7NUCawkcvj5VLC9Ft0A1BVqz5gub
0C2DUavDJNde63H4yuivd7OONa0C2aULDdInslecLjmV5hkzyJNsHtkjHO50vgMcEBtltqjIz47C
Wdry6RbNXl8P8LqoEMkrEQO/xy1rwz/HlJQ3G5w9WIKc2fkdg06vEvQx5zs6oalwwYSab4WZH/39
pd0qgK/SpvOP6sLL4q4FxhZSkTBFQVuBoVR1WT9ibHb8ob7E20s9LPttzaXlXsROtekgPsV6ws/y
3JXmcdaNHkox+GqMiT5Eu6XV7xFjSLypzDTWwysYVdgklajCJmgQa7OY9tM7QNx6ogEj++d/Ib01
14Z7+PrWyJkJHgkRz5P55hE+XiZmPceV6ZHn+4J6rSrBnW8lJ7xh+dQZIe+yeTn+AkoytEP4hEsO
Juq9wAgWoFrdO0tY2TzIOmEwJiXXNqTfPBkfooyDlMmMOTCjstpSnaoOCywIrLbMMm6wd5Sz4rzy
JA7NXc2wY7Kj/G2x7g3srmpx+taApEcaBbkn6grFQs0TtEgghRI//+nfUzy8IpWEvMijcNekLZt9
/tClnWvkczpx7EkZ6m+4cHZZVsJuUca5bkM0XQIp+BsWAzNoUWCCvzx0dDQFWAuIW0MYPM6WejDT
bttKpk7VHzxa38IrQT4qA9lzMXzBO6o5yb5Ncu4OKQCrcwYPIru7myKbhgWwWS6rrVrrZaYSRCGL
gGa0LZS6Ha1BlL9Nhi9qCjwDg1IbNeHm5W0hmDfc3KnZ1x+MC2haxI3MhgETwSBK3/nqqScHBQb9
iyoIaHCh/qL4XCdqJ5Vm72GIXJd815J50hUN74TjC7SZKknq4NMveT5foX0jYaYqFhPjZgbD1HwU
4hKieYtVNLUqKeXDog1//R9iudvFw0CRr9pyHHj6fydsx8MM3ZjCneWZwV2k68RQSbuI0xT/CyIx
ItobxchEasxYlMtWvjDrkGepgGDV9U6Vx6yxaHUxg6VcrnwvaSO5UgFZREWZgzyW3x5OmBddomDm
326DX/OIiMNTXLnm4E52nCQurbhBwFcdS9iISGCgYKhB3hhawZB+Fcr7Pas+LIAeYZAZK4QPeUWN
d02P2MY7vTTSt8zVlN3L1GzWj0tdO2PrdnZoLsT9tKxygDjyuWl2clPa5v9sFakKI9cunLPg7DnK
y7nhLYNTN0lsMBSUFLmLYc4U2Kz3ZH9+ObnNf4WxqJ8m0MjeVjmSJqqqXZP6pRlowXzWmzYW8fAI
X/26govLUePehCCOUs0mKI5Jf0z6tVFUwhYP6nncd34xqkrE1H4EaualyLd0Rf92vEdN+o8N56be
hJ1JH7rB8OcEfmwh2R5U6F7vYuV48pFUWF0KvYL16s7eR+bNYa7APVSgv3Ca2g+1lh3os/sGGMPm
cRO3UYx+cAedCcCYIiLv+wa87KA4kT602zx6I9JqJtZu+EROchzoVLa6ByDvrZRtgXfPaPcpHlag
enfkZFfBTG961+m1GeCNXQv5xnvonZ4oHcSmY8/5SmjutSvs9TvGuP743N7FBPtO3nbmePOH8S7t
uwjKd/mOJaJlHM/4EDpMhvQ7tb3/ZbKyi3m+gv+9RXaB1zX96a6DaakpDvGUuaS6sYA7j8Fz8b5t
szKO+/eRKZKWWYrZi66rXUUHYdaS5xnXJzg8hsrUZ2mqWScZXKumKmDuRtj1BWARx1FfvoclLKS/
gyKkOcMTMCVXhr6VjtscFADNVfx/6o+1Pd8cKgrc/GF/RQbibhUT2DgjJfnJwoKktWOAn+/RZ25I
Dtj3BmEjStVNqjxd9stySBifxAI4mCcH+ChFZ0QoyLgXfKYRh3D31aCZvm/240CJFVm6h4LaeP1/
eoNGMuyLwgON8WhCXky80Sd4BsEj95aAyv3kihdBbQlhvs2SZT/OgoXVcg3YVs+t5cBKB9lJbeFO
dJbUA6V6pflLB4MlcH2oNTtgr3qLK7sOI/CQnJwjVFZbQe8cvfL+hQw1bEx7/RNQ97qAR95rJtgR
xa0YahAgeYryFLRu/zZ/YrH05K4G35NVv72j0l8YYrT93gP8yv+iK+azxvTe+scS1543E0j0t10H
kesZlT3gIedLpSGPQc6tMgEihpzk/lKeep5tCKRNtf9FOhKANTtN3oGN1HLEBu8GwhiDcquCgGsx
5FsYOF8K+zp9/9rIglljN6iSa1fNBQnyG8LfF20Os0NJdrFPwuFGw0Jvdcv0FYpCboE7doczMj3W
St+YoVbS4UkBgwUUFkw/IotRti3R0E1KOZ4WWNgjGtzuuzrltOD/DNIsqjhCmOMlKrNGs52TG3ny
xcKsYoZ28bf5fJMO0n0bB2anwD1JvjACWWfT8hOvRslIau05ZJh2Q/fHSLebIsrSGxOYw3qm+/WL
ZTvEIuuDhYVUtYHtWSJQ1Y6Fs2ATlbDBt1KBEgM5VxlB7ODinbOyQaTC6znBAz1uNb7akDTTEpxa
Mj4sZogj1zOahv2q+IiI+/y8EA2emy7l/ZjL4HoVHagam8mzzbCcNOFuShLkNIU5FibAi08wKSoA
DcSTnS+SetY1c0Z5meWgwP748HGYDj4ZwmPGqf+xv8mGOGnDnSk3MYGsaVjhVdd1slJk3wyKOb6R
mZL1qzEEXawFsmAmvTcBPpo7VQ4ixACLh9/5LmwD71FgOerWLWa9EAygxLANCHnUFYSD5zR1fgdf
0yoap7KgemlkGFHzofZJjJ3vGLNRrR3PJMtZ0eyGBKeVmU8epo/jPRWM2G5Jgnqm/zrw3uMbn7IG
/LjKcnYzdIOhlfi0FvxDgjndhYEqA6QTOpfpB5s7ImY1iLQi/BXvloL4Zy61KdourXCrtZVMRsas
f5rzEcrGZzu0zW7LHbYynnDD+QLgep9HhYuRp9gjOZdouf2P/HH9qsaUdYyNRzTYZitom87HXAbM
VWks7JEqNUIkN2Om7brvc1gkzA5iVyEr3imtrmYSsQKTiPaUFWw/EsthUl9uFW/7z6cwuPQg4P4N
2Adx30ZU35kVXfz1DQjnnDCraMJ0cLVk6ij7cdrpFj9jYrrVWXCFvCzr0b1KeaPXDurnRacC+Btz
oYGQfbEkxH42eFAO9x8ROZ5N+Vg01eZpHlu9mIKlFLF2qINYq3StmflssFzKEg6rXPjEdKEM3JYs
Fb8iJBivqrTZTnu+LrNewYDL4UC+qKn4t3FWJG2n+OK1RWejdpdjtvVz70H51KcXBLYiQAt+xgS+
xkS1PB0dktVUzsMFEhsvoo0I/qFJBguISKsw0Rps2QDKNx4zWoQ829+vAZrXh3xPv04j0Jk5gHeJ
HKhF4FGPjKVwPigkWxOXYvBP1RpbvpAsFkVPxHsmFQZNY8QOQ2ll15RkgLflNYf2XDn/kfM40m37
lHVop/dHC5BcfzjG32jnD0bEEE+GxwsNr9gvfZptyaytqmWT7p7lExyRjPSy7rpBxBwvesLl8SdP
B6z1l4oI7gbsj1/48uRjY9Z6xKU/H6plXineOcZ1vViMJFqBeXB+SvyXvlXej/OU3EyHEO0ANSeG
PZ27aLrFpk+3ndwDaRSuVV9P9Svv/MQ1NAfQT063CRCoeiPUfq+E7BVgqqmwfw5PhAbYx7oYSnQI
GmgVjD2Rm3zujnv3gIFpA+rYuWAp1z05WBFD1WDoAj+MbENj4+XGHf2qsAP0wlsndaq8g5P+P1E0
u/eXNUAOT+xbG6BThFHIcMrGJtC4EVJa/2VySG9cmY8v8cCJFhUhzcMwZ523oz3mCbXiHKSwAFYz
Urell7wIIsYZGxOmcwWLM9IfpE2tmlLeUGkD8a3YGzb1IplHwOi0UKPIQ/6rnQ+hkPBOJJcLrW8Q
xFO19kO9Yh5JVbmg+WRdH5GxI7AJvX7muL4wgrMp6DjJz5S35XcyGUN+M465hCU/8MjNqUiIuWT5
AzKz6i5b4wGN6oEHkDHZdJkx4xrr9zVupiA0oqP3xgVO1ZonAZ33YKJK/UxT3GY8R4vHQ7rJa/J9
cSuy77PIykzhqsMXppYxG6NJsDQZusW2JBFhLYWrzswk6mu6moPSz+xp2JwpsjJoqJmrZ/FKzcP5
udFi5W+B/x71RSLY4BoawJ6t86yvkFyWj6Co0sE64nx5jRooSRnSYjyX3TPFQS7njDbP+rxQoxDT
9l3w8FqTUxlB7WJ9mp99TagLmgRNznjEu5F0t1ubJksMQZ9273nhBgTX5lA3dnuaiokUgfoQ8MuA
QF+JURhTUq5/BOWEUhvHiYt8E0wIAvEmorCC0wzxjF0Rh3L46P/C8SnOljtnfq2sAMJpRBmz/nHi
8a4utqwK1s799AdjHIqdvk+ILk1DfrQaaxt2WiQ7lfduEX4+bQpv5xL1Eke05SAGUa5RA1EpTzcH
VU+wHX5EYVZ6Eqp8O3bJYg2K97M2+uneeNzqZQ+mozUJoaHrzMS+SWXg0prYYI661sP0kLNmkrXQ
cIGIgbMfl+13FT8T01d7HkOgKbHGjUm3/norOW/KfqmdB6K0UA3i7QKNJfvGCbTm+iLOkd7Q6RmM
ikmQX3l2nxoO8eqAo1qcIWbwCK4zIfc1kNVl06wiRCVY4UN5DMGJtYln2LgVKo5jBdxniVw8Y9eQ
J/rmBdvEDTmbCyZiafWGNU0tpgANlGNk4KDokreyjV65Unv8Uu+zzrRY7Gc4pPSsnbUFX/KeS+YU
nTyghwpEuG+PePmjcGfDMpHRcEnRjgy44kGRVEDaVadiHaAzFcZq9hSq36cS2hTsJkqRkmBWh0/U
FjQb9hilj92TMuvrBZg9f4CNksJAzuzMtQ9LE068V0jKWjkdsiuPmpAJB4Gjw1I/ZBXhRe2uTS9r
Ss/WpVX1tYVxuZnzQwtSlyngqjXRi5MnQ7keINgD34+fDxIENDhd6YwQRJpBRgObneAnWDMFxouL
6mpkPYhIe5pQDzCQrsvEsrk6bSDcGuO40m7HN0MhcdRUzJGf8qvejPFTDGBoAMyuOGcLsOdSXXq+
FKgCMT5LYL/qywtXrwD0BZ9VAbKmUV0IFvtkInEHQoeN0jgCA62PxHOB2Otc8ZDxJBsbXHoZMK/2
9N1pks6f+3sj1vz/vqDzAz8i2lBOXy/Yn+7x8A3i3toXO2TDtvCJsgCuHhCzTsC2YU2jX3RT6g5T
xLVSQSFjaKYCjDyM8iFsqimXGusOHPSrjc65i9oe+30SjAJT5Md20AHsWJU30503my2gnFCwTG18
Perpbfq2mlcY3j6GsH57dIg+KucSkEXdbJJMltcdy3kWoDPxnDmuQT5ZEScXrkzaAimfFFdPciCq
22Ovjp9DEeEUp1laPI3VXQ6hpRZKLTquJXMj3C6GmIHjLdVH9Si/zy6AOj0ToWjvBmA+epGTxFOh
l7dQhcpWCjtp2mADlrSqMGNs1xmIxaueaMgolw3nC/ZFVjT6BqJGMp8BxMHkKWTjeV0UGmNWg+Ki
1YDjkOINa2o+vuFAGQPIAVv4Fq3AebPfcA5DT5VFglg3xYXdHwG9HIHuwtqyuM1YzKu0gdlmBeS4
mbNdEpCwQLIaNTllKxzf8m1aluJ1CuJ7iXYg7xZ5E0fWi3C+/sXuZQIUpzbJX87hnRTkkQsMOdq+
pEyKr88T4XqDW0uXINPe3NNTyRwHZEwW33UF17lO9Kxs01Y67igOde0NtKmD95f08BvV3Uba49d3
59Bft9TLZanxD59yfnKE+ej9Vtftcpx5tfkXyd8lOSkphI8lvgxFUgcXu/47iKb1LY9ZNHZRnk7Z
h7J9DsAnclEE9cs8x4ASxpzzeiqoyux7LOhx1CDp0PrFJnw6lqIKsLclT10s/yWNYL/eAs1663Tg
kngM40qTv7a0rvwrzZCsaQ3+dYf4xvgh7xPpXGmS71nMLUz96mdf4bSIxuzkRmouF8OStnZoZbll
ZLsbxj546y5+XY4LRXm14rAFC2Te5Unfv7UVk0S+Lm8k+U6yT06sPOCs2ltc/gMLdZXF5bPCVPdH
T1YhaALsLWE/7zyAZyIqDMt75/5BeCUpeGbsrfjTnsqWDhXbO/p24BjlD/wQtIwOKhLEcEcbmld/
2qT/9DmhInTQGycfju3JbVwR6mrr80LbFCoQ7rT8IIzzDBvGrVYJeWblNt4KvxSl7mbSWS1qQq3h
TwM2yR8KHZb5GMvOV0DuX4bPxIc93cmjd8XiStq34w72vUkGEg1JTERtp/D5dcMOQ/Fg2yse92Mn
eKDBtnAxxpmV0UU7cvrHLCDIiCNgZBz4THxFZ1GEYzs5SquUBnpIXsoF2hJwu9K3sNG5Fu1tfvnc
9WSviZwVh4fKgXrBpGD2zXK58OIVA5Zmg6mnstkzSo0i0J9hnU3vZHZPWFeFSiIJBHfyTHva68hJ
jRi1bRqMqont2mygAEWC3WaIQMDGiaJYMvmN+iOcCrUl075baTtudGWrxV333H5mmPIMyq9xGOtA
mB82sleFdoYuJHSjN1Eia3WJoZe7IzDUPfz5GJ+EVC4mamD6TNCFc6ig1J5Eni4jGa3NmjoKuRHi
wmkwB/P1imc5jhKsl8jVcwfEVKLVu5z1TWTWQbTYAXByVGkPfMwAiX1AcZjPukZZuvdaxSXHJPEV
MEpRHhxzWtw+zIyu71LWfp2ur7DHw5f1tsM99LgkAdaM6/aKGr3Hu7mzgxSLRim5lUc2Qo4uiBgW
5bH9XhtjB5+IAX5h7A5sTWg5JQzxm/mOMQIwREfh3W18YTWhYa7tqa2yrVSfdpFC1wRr0l2+bbRc
Q1645ltKKmLiFgLWXqvv7PlinBotRY9GoZ+Cm/5CLwLNzMQT9+vh91NrBcX+28yj/jdOg0YaZOh4
6wd6Kv8WwBI/yPBi7dNPKN4cRgI9wXXZQYTYnp0PYfYZIs4lktFDO4ITZH1hjMRjdAfHbLFGD39C
YDt3ApVezuxXyUk4HqRANrepisCdVEihIRXuBb+9+5Fi65Pl6K78oKfQpTPRz3IJXnqqY8YKTnQH
Rbt74RxtuksXSecfjbj9vBdjUwvZH+MF/a8iLxVcAXbHlf/RxerJz4AozJkKmv8B3vnL5eUuRGKY
NSBvdVvL0hsNGHEk2ChMmpOmvFFMU8slFyD5CMGiXLVj6h3DwBxjgishtCyYWAdekn4GyHHVSgMN
pUv8kX6vS14aysaEIfOSng0/04vrMrryaL/jXTA7bGwcBFSSHLacknLPP32qdz/2/K9R12MzB1F8
hdQwhC2wmqhsqqPg+BfIhNkRcqFKkTcWi66wvS5jxOQDMNmVDQyR7sh09/Tpa6SIGBROjcpGMtkv
Lv3mKm4FQ8K7se9fG8VdRMZQs1IHzK/raLrSJ63bSdBPXhPR/Uh3Sv5CQam7k7CFJrfmX5vGGhKn
9ocoGTs9KWrUsCwemLAE9p8/RQ+pOyKRE1/12gPe8kHE9d/Kh5dvNyfTZdOXTRJVKbVYB+a0JLWM
+CcqXw4tKnydop8PBgXvfwTGf42BqAOricPNW0h32bmlLzflTBAv/IR0vlJ7AYRbV6BEQ/mB4QEZ
f1fHy0Z15COgXtKBz0gRFlzab+J9tLjky/V50d3BBCto1yz5ZacutvtNEG2yIDCWOrHo4S24lSwE
yuo5XdSz5zh1VKz5lqvx6G7zkMz2ruujyi1VVLa/+mxbKiviUlG5MRN3rz8jcAasesMMUjp3sbuP
EprzzfGcHKcwcYaFF3QJ4m3PVwsFj4ifA0wOKM4/juKOwtzkPGgueCl1bG9gW1h5RAe7kJYwl7S5
vRWw7P6oeL4MbH7/QlGU3z63QJF1SatV1jxD7+fZKk0KYb6YCRHVM69tYs9CshkPZvVYPrloZlFS
iBZsU6LFhcCFAPT4IeWH7UBN/mwhVf4rARzebqbVnltzNmluJNOMOp4+Txd9zk1WLyEfKHeO5G32
EDN4J1AIOltUProM8tCd7DT12s/Hqfw68Pdpro5kfRtS9/Ooq6sPKdyBSiEHHLcw4KJCaaXIa5D6
D/phQ4ZH2ymdlMIMs+jSgFFYWSMxXLMAHGNehkN2/vhyHE8KMdo0LZ7Hz4FO9qbSqXxcWg0EdbkS
5eU2L87/QtVtH0d92jtFQ+ET9oy7coCDDOFbKgvz4BPGfzDuy4cIMHIEy+S10DBxLu4xGb6LW3nm
cQJarUoWhVGSW0/ew80St52axDl7iIiYYzErF6mxr/uqdzFCXz5iwECXRNcOjOrRJ6/DpeoMTZSS
NoEdiHBHik3LWflQcqQZQzEq6rOu3gBfXBmmpBj99KVYL8mQ9Oink/3wJb5PDkjXpJamuMNvZnM0
9H3G1hhZw6AVhj9w6vbLx1fzuIVBoAfcMTUgyLXfKGCLMcXnVX4JlIZDIDFZuvBP+1DRuhRj+3nI
O8e1NchPSNOIIEYMC1pcf7m3HPkTr5MP9JynzoYtdbQq8pVqcHzWMD3d8+OLISMkaYGDtbzhI7N7
qxCfH91e+qVMFt3+YT8nLafNLy+rfLOzLqcFelGLzUctNMq9ew5KYUWnHPaWX7d9LYcUKuqjzKue
q2sou9q8iluisTQteMd6HeUgALujmkSepXA1UcLKSpbK9BxEDqBJtlkXoW9Wf42EfKN6JCUn5IGn
51Qe6/YD4HRZy8fSRhBZGykavBev3O6m9kma1p8WyD8xn1VZ96tj8TuvzUH7kyHWhxQNqa6MnHOp
GcTryJubArZliwn1CJcGFOLn0nQsISf4TnOBQ+7Dg/LnvWRT4gbH5K+WJDaYlCdEOXsvEKB9h3w2
5PK8ERbwZduNZzOe1mmk1lmLuYHnT9tMb2j+9O4bDQSyrXi0JoTlncShz13RFL30mDNksz3EXk5J
a9iLdZYPL6S6BlqgZYeKlbaV+njeyHq5+J3UN53VvwBbYdGCKbKJQKNF+E/TpTmfUpBQExlNOEUv
BOH8+b/ir1Mf0yM2D3EIe3d/2CvquByYTUJukFSLmSOQ3nxZZelrym3tD/ngPFYrTNZldg3pjArk
OEQkQ5fCFnjMtF8Ml81UeMmb2CJUgLgteljBMQEfNtbe3XBUom5oZxrSAKQKhjFGTA11xz6XjPiM
9R0K4XlsOUkLm0yO5169wP0uH8wcsD6ZygcS7Alj2CRF5va+OIslbovk7vHoNSFIHTGBBP7hHB8Z
dK/4YK2F/QBO7ECWcRDAT/qkqHX6HUhssYllinrOSawPuTRJ8sl1XYYRncqwObyxikGCohLn+cNi
ml5GNlYmdCkVggkoWLQF2dkknbV0CrHh/pmRPBThRCNl96N3KYn3Mw+IfAe6PwWiSWLEaM/XH0qG
NM68zQy69BLFMfjoPh61XrFW+wCpwcXLcurgi9CexQWhoU5jGRdb/B7Efr3va443MuXPm+AvXfoG
DvrEgxi9VrjePEI+Nz0jRAAPlXJBxy0NvZmC+5y0m4hDG2YjoLTMDPnwCk2jNS7V+cg8wI8NTZ7c
e14coSs4obEqpBM4sXoGDDvI3JGLquX6N1CYuY/ULQm0tFgLjO7jxbVFadxPakkXbkEMyAoIuTk1
jX7LvC7EoO8Xql7pQ4/s/klRc4xsz7T64q7CMlbIyIRByOOdwXBtdTtrzDUdWCxEg3F4j+44J86Y
uSqjOY3xYCISb2tLSq96X9zvkLfs2LrPr1/ckTKMwFPbq5z+qmGMFXX1FGenGslqWICP8Gmry4zk
tp3svwA3RxplZirIyFRifOt2RrD/7o9HOMev0AAffRY74dsuWWdSTvfE82KMNr2Y7OPvySZWSl/h
Rt/+0ozDqRV+4VI6D9M7EyPIhCtrKjFqxD6gOhaDU72IgOn7GKkBNW9KsTk9Kj+laO+skmjS+dUP
XzEHKxK5I7+x/sskf9QSmCyaQXdiWYKAfCOMuQ+4okTyemgXFfkIhcGsOEAGARheeJwXjJPIXvEP
Cf0NmLaik2K0P1tjy+vHEVy5SDwoIImGKcGUDTNZQyR03BIdm9KQi/LLpiCcxS9jABs83DsQ5UMP
2oGIbPQM8wbaPWhtUwXNQQx+iT/x8UMdprugdsIV4sX5QRkhojcd9xbblK8t9g2FEZxN/V81HeK1
aZhW1zbMOVHIRbRlQw0T1MO7DXxYvnm5Fss33vGmJn54UYr7k8SkM950YhwUqV2za5TLgMoJ/AbX
S+6OmiXxx4wFi2WD8LtRUHAaAMWcd2J9tHEzHj2CYMuN1Qk1J7/Fc5h9VNyTd17W/TNkgHHZd89m
kVZoZKYljFjLC6K9MW6NZ9aUIIW/AkBF5FM9JWAtB2NYmft9izeq8f0p3NNAYyefj3hPtxOmUULJ
EMcbpBF77pYx11c9i6h2/6Elwyhqoaf/fdfsl2ZcnrOpl47vHixKb2k5BwXb4SREYY7H/zjyYfgB
6wrbv+9/aojVwiEdMW3fLLfxtynz7kN/60CazVRPMbDuVFU06z60CjPzEyMomnM7zPgioptWf62x
HoKrzOiN7Vfab2W5bVB+dBBkUu/n0N9fZuZdklSpPZ2TVkY2UY/cO88NW16fYWQpD96tV30+5fVH
kGmLVYxPJEg+/rPSyyFnVhjTuL9hhsjCAJEqNsm0E+o++kSXnf38DFMvkeCNCaLKDLfBZ8+d1YoT
+n+eR69pbZd5SdqRSCG0EuMyvnxw7GsLrQDYFV99jLCaUaPUOAgISAl7afsFLyYq8FwS+HmFU16U
GJDuTioi4ZQmHaxQqLEu1id9v2oON2N4mr0AATRtxpqx2Bax46kJsrEwIpLZyyFhDUVpeIGLTk22
RRXWgxzw5eBgG4Y/+8yVLC3OHGNt0E/JbByibj+iitcf90K7jN5AOaQSYh8+og2mNeLo5uHnVmnp
MmzFwt4oaxy7R1LjX9yPfQUklGNVy4FvIJvjgq+O8BRD7J59+VRxlqSEmETtdJp56HqkrjNkJabL
XPqkfn0wyX9lbk6FfFNImZ4RSSHFuzhI917SzWGS0nm6EuHaFGNA1E1CBJw2+PkRi0s683yZ9pya
AD43aV9IgR5MD8jSzrc4n2CxbR+G9fJ+ZZfp57mJUARRmwGyKzZY30qeuoPjW6Kw2zKlb4ORxNH0
ZdFYiFY1KaYQ2G28p/Rxz5rj7JwjLiosI4CUwnSyOk6x8nvjoxgoEbAlTtYEnnYWXcHdLBp2VNee
zD9DpEn21pxI9JgQj+x1lTpYWQkUXYlVE+4STT23De5iUc52t1SGJ6A+xg9WFFQ3o10TqjCxLAUC
QoI1iolP5Ld+zg4mJ4DULeOYaFg5Y/LXVgsPZQa27+jjiL9IqGM1cv1ZvstIcjUk9WQU5I54d51X
dHzVhGVuy/uollqpr34IFlCB6tbRlJ44QoKnx/ogZHhkaiGmEwXmxgg424sV7fqpmpK9foOI9fFY
9oKGGUhIEZ/ip1tn9dZh+Z766t8X2bhv2utqZ58Usi66myEkQsStdRJ+DtC4+5bFfKaxqWAIhgbn
ABM9VSISvmRk1yQzZFsvT9IVaDO1trR5CsEcBjSKwoOLzA8nE0w38RnLuw0rOrCdHrAwIJrPalD5
i64tvRT2AVJgRlaw+RSA+orgS9CrB7C9G5myCl3UY8mAmp0hcU1uBgijQFBFmbt6LihnNYLxr3ag
ibAZibP1gKAeqTDIrmXyLcU/mVOk+PaCDSDRyi2Vd9PhpJldzwhQKUysfiRzypo6O8p7R2yb4FtR
krP8SDHdMe8sgwhhyVyktxMtlvT43GLq+2hqEF+aJzaPIGtMwQCtqdjOIXRYsyDua3j8ttxhTMXN
/owFEWcp7nfL50VEJTMT4XmL3+i0QSGmu78AVe46m3DS966Ihq9sihc6RgDe3zdGRfY7jWEXBt4r
FjLNR5SU+oVw3jyHLJQiZYPYdCOz4D3sovpcu3OA6baHOeuWvfZFB9UpR//C9z7DNJaXo+aYUkTF
QWk4+VReU9U55zcO90ZuA/Vmn4ETUYpk3Ggy0Xy87iC+afcx31bfE830RZ8eDjCPgrxJHLzd6D5T
IKXFi7rDjhAQddGYLh3p2GI56XejxGPfRhGUyYnI9Lxt0pbbaXC+tDy46h130mnBUYov4+SqTNSL
Hiw6QTBFeecWlHf41PY0IiwJnsKdJItdz1eGG0qVRVrT8qz/1m39TzbxmR4UE2gv7Qqh/c0HeSAd
jy2FnfIp23oe+mo25wJC/FMonVI1X2HqtZ1gToOvj4Qv9AhINo3SmDJNW4cshm+u69sr5zenIN9K
FUq6RQJFe7MMHYzpfsueEBg/czKumPyDogD0AmZohVQTqDOzBQgMwC/8H0dKMHJ3juoZ1s34c1v8
k9NvOVf/tQARVi8AFe/9U22/uZD3pROFaJfigzVnUKZNItz0S2mo0r3L3K7FYbuDOcJbNAC0Aary
ddGV4LACKn4XQPDZ5nk0aaQD0ykjvtco0JPn7BTMi7/CylMAEI7RVEQfkdc/dMKF1ZF9A39Q0V8k
MBn/G8jlSACa8cjG3BQB1yEsqdALev1rUA/wjjlfLEuKM3tuIppIAMu6Z+a2oNPrgEeeVBZKwPFe
I1B7qVhHsbEqzKAfZo7egltR+GCuDnE+SeBjTblueXOcGIPL3nSfM1dXMl3jI/DV1xZTwcaRmg/3
PQzRiQCuBzhaTW88lk0KaOMjnkyZuoVZn40lNCbWh/byOZIifBElzjTs8Mqg7fPtKUGQgbCrE7p7
HhhaMortZyMlPzYRmNLFy0ba47Bv+qe//fcUmYxSk8EJhmY+eG7wCZl8ZkJo2d/gjUWpVSbT9gFn
JKtCLJxnbtjj834fFdCg/yNcWpGIOUWIXN4igyrx46OmH0fFq1QIQDZIRJdCudv5gCFxmL79PHhm
kZ3HWd+5vt1FFHm3C6vaoT0kzVWT+u0ZENxcN4uXqZmW6EuywNmp2jC3Kz+aKuH/TuBqsL8sBg1V
QNaJNUIIf45EY/+KxytGEzrWbv6bKIqhOANECN9+Cg5pucdw2yvvsJMIaYrGHY8NcjnyZeBs8V8c
jgenotry+sF34xF8cBqkrs2rDzXSpTc2F05Vc//Yj+48TLHY7bjBEyCerbYw+VgUSvS5jEKP0Coo
DjVeqoswafqVrJ+b1SqTg+8t4srzrghYHW4lw82uzxqTXuWp/fbnGXbx5htoSiGfGJlLpfd11MV6
49KrV4Npoe6ao2HXCE84am9L5m/tU40hln0U3YDs497i5xOP2EtRb+mu0HQUm8Kqvm21Rk0e4Vou
3HuwdPVPVG3f3HaQACplKbD2VUH1NVwmahO/9SnAud0yXWGPCb7g9YASyYPXLcn8CApKRZa1zlCX
exRUmIZa3rBC12AKIe28BHR1FRHhXYDgKU25WuKGQ3NyR54pLsdoJQUgKSixcfUbtfJKm/fvNBoz
OYTYM6fRV1Inut6326GfWCXmzP0O8vQmPObls435wjowfKYWtoHDVyuMSzEV137mwDlhl3X924Fu
PlfyPb4FwaAHvKRRE8J9xUF1+jyLK7ug2cYq0R+JjX4Cb/7z2C51FNWnZYFCazmtFkXEDwPDPOD0
ik928Fmgl0Z59AiVkkEmwgFTYY9z6LDvOqmXouHuRJSG3scwgiPAPzQKnwCsRTU2hgk91B+HCagw
5fcHthwV5YxBgYUTtj5233IipqYbJIyhd4A5VMebHHPO0JQYgKBjwZpKtGR+tHEccl/Ff3vDGQD0
dfy9XNm2xOz1k9TOblfLh0Fe91K8KNIeh5CjSOr+Kn8VPe6yVDx7p5CWcdhMQ9CCjULaqRms0qkf
7NB4OWVxXrQqTifxH4kXswB1xCpD3f+05DGHC6foLMHc4i4ZF1iwyRfFZhxY/hYn0WHIYC08Hpim
azEXNOcugqEh0oiBBwbD+c4lyTjopZkDidCop+g4aVHVUARtfrpPwniyU6InzPR46RRVye3EreUv
C+ZxNzwhDApvLbEkcuKtxHOtxm4dhIDzmnQ6iR2W0CVB8ZetHKqnd6T4gDtHkKSAXaE6U6QSWmI3
UQehtilZz7R8GVgrYqH0NoDJVmLXNDn8nyl42SXl5YUXEzfdUdmCXqIYIRq1QyL1lkdEmeEMRwRl
KWyd/2swIbXr0wmnva4ZwjXPYKtNRl/0UWMz3r2dVi511G+t34vvykTo5VIGaWXsVjt8sNz7q2nM
7z9gDK7CxxBTeg08sKrE4twfXRz0GdTOa3ds1tp6hO4TfZUDacP5IJ6S+7qigSgmY7xPUXHDD+rV
AinWAiNcnbnqtsr8fyjCq6WN5OAwswE0NdEqJ+XMpz/FkhIZmN9XEloN+NVet8Ydqbw1dNiQS+8x
yYdakx6FFQcL7/FwdP+Jzj4xlnmEzF1cvLl4L7SG7b6bEOeLC3vh1hOgTyAPUJnNb/vJtU7mPkd8
BReJyqV9jWkJlRyAR6DfkXW1byEmY2v/Z8RWtKbj7czHgxyoWAdvWfOCWppBkK5AFNjUqaLM92ej
s7HfV+3/ih8QRt4vj+7uy8zm6USFoP3W37hH7Qf9uE0P77EXHbzjWebBWmMmbIP6kNOr+6hvH0rG
n11MLvpXp6AmDS0TAjZPuI9WAZ3CLxCbaz3QrTHDUpjP2B+aeNWwGWHBoTZ+6O/Og4z3wAftCPrX
aspQ0tRkT/HSEFlird0+SKJPtabREsFOQ1U3zUWLnrV5INZFBtoCE8VYHk3qdXhf1cQarnvAv97C
ZIA8kmPDABKOsxLtRb5BLT4zsaUovxlTLgvG4ifCJI+GHsDiwyA+luIPeZ6z+Y9CCc75taN8yMTA
TmQcONb07zfZhCUr9s3N7vVV1YoWrKs9Z+QUeDcqDGZch6vQx1nnHAw2AW1jImPxxzLhIBdZ2bYU
0S3tDFJBLWlk5RLn6hpeD0gM1GB1sqP++2uT5IxDO/JqNhEkmJIZIc7vyujewhml/DDqv74qXREa
xxqArWdA7xle/XhUz5ZtQ+TxS7AotTchM+1UcoRkcm6nWAiBs1Ku/74akz+R/+G84GZkmXh7Il1Q
AZN86fIcfmAN+EH7noC84cPK6kTRfLuI3BqWFlJixHaGZGG36P6o1rNavo5XRFo641Sc4qdaiW6Y
NgNUG4YUYU5qiaq0L5J2tT0zYMxUqbqugWApRVcqid0on4hKz5NKoKpcMSyQPveoHp9dMwf1flt6
2uuw/oO1fFbuRoIZfwQu7iNWSC5n1BmhXvgOXk4ZMWpyOBiGl3rfLSwOHSpVxOW8GPLTV0mgclIM
bzZVEVF7nzz4nadyYuHkRFd7WIRsK0ys6KlAf2Uc1uljEvofns/IO2maN71DGBI+NgPvCjPEkkUf
jst4amJd2zW/Wr/lEbCUwUA7+vbzIz11voRLb9TwKJE1HnbtQh3lzPHVwwMSWFJlheCTLnLFgcBq
gC6ozo+GxTUKMczL++LGxibniClvHYFETDRPnaRHSGkKJJCf0R4109XDddwcZg/LgC+1W+2q+Ye2
PWWgwj3nQGiCY7kGGfQJikQqEIygaTHF9NAlUYh0r09z3UGRctAtePgUoQtquOKcTExUEg7EsvR3
nhhjFxREjTz52ivObSbesCK7udzHksVnsPMObQ3ACFbcaKAzqj1k9AMYjaPhvm7FXNJ2u+50Etjn
0dNXgLVMfC19Nc0GR/fGwID7H6YaShkDCwzsSWtR8Xaup55mtlY6NmGkqmcuEmpa0FljisvLDRZl
NuKnWCTE1j1IOq0vkmngbz8XqaVpa5NFcN/zsuQFDKXrZX/tCgMBuIDcTF0QE/KwQPXQHOcTSmqJ
wP6bSqVP/PF6roiUA/FZltNfRs+M6ZJN7Y5Bbn0PD4tE/ARZq5DubhAlztwM/C+EgmMzJS5wH3Zd
vbw5rkuqFkz2asweUuPfTLLGCZGOfv70Pl6PmTB8VwzmFBC8PHz4XL0xiEGRaCgVfHyYWbon3mO3
WZC11HzOROAh63+jm+Cg3KnH1/PYPnNOICaVJjMpvELg04YrYAvAexcLFzO3pPk0xbi9zkyMWP5q
rYtO9AMGiTqj3022hA/pBYskmQE7TlPu2PZxJDlcO2H51jTJLAwhT95k1TXLYRitmdvmynt34Dpb
shbzzSKPY/U2Uh281QknBpbVfNRS3/6cmyvIxY/+sw6qf81f5hLzYlt2NFSRCyRWX6nkyUybQhur
KRBQr3UozL9A/bFvM09EfZYCQ9rH1frKY49yB1kJnWu6YcF+HZeXMGmQWQCjDUSOFcrsvSBs9jnP
QKOwW7CbTCLDKXTXyJya9nRuozU5aqxuCmjY/6pB2hXaVaEKHeD0UNO5lPqIpI3Fw0n0y0IvFMRt
H/jz24+DRwB07jMz/czENG5tVkPsmXkrlZfKIMcwmSDQQsTL7GMYmpPZBtiNWm9o/+3BU1APsWwv
tSfHZkvDCZOHzP+8MIZfVusNh4tF0dyj+Mgs7DcubZwqqTzatK6DmztYriLz3fGCA1UGAsnkergG
MDfpgLlfzXuoRbaP7j37l/1fOTw1LmipaqN2Ts9kRje1wMXwFUSYLmb03DrC4xyrCBJu4bh+FppQ
dntQCLBCFHG2E61RxZNULpVIYKIAT1+jH3Nd3miySx2ZyV1wokNEDk8QXkg/uocevLxQxO4dwB07
Rij4+EMV/FDYhXngSk2NFXIqnXyiV60Ue02jFVjvbqPxZBjUhB9Hmz8b8vbZIXn49qNn70pF44mi
72H+wqz3LIkVhjAJMRKLYuByhYBmesBosRvVUVpXLAGyJoPaS7kbp/oPbv9gHAJzt6AZvGur4Qxo
DbjHdqlITVXNMu2z0hiBYEWEqHhZd3W6HJj7/r9wyIpEAuUZ8HbZ1dgHxn8oS2j9CJFBjEnf3PLo
65E+7K+3tXPDwrkOKJ8kDjSJfjIi31OaSCQlTHzLu9EZTsuAS4fnrO0xqhQ5H+FZdPacSN0ltLK5
MQn5aWYYc2+saRUSawoetyDLIlBuvf7QFE0liiE8BrRxNVuePRhJHypfdNoZ/rvknKD0Y5Upy7kz
mJQmRqfaFNjBk6gRRpXoE36Khnv2YVU/0uUNm1rWKP0kiY45DsyaWPZPDNDu21G2P7VrtkBB8p1D
x4phKsINuPKxQNWmYpg2Jhv/MaD1AkJjBLEsCdCbSrO/Ntto4f0WyyPPdEbfY0Ycq301+6K659JX
pBJ3SHoHikqny/3iNMF5vovPSJQeHVk3OaGqoX1/vQZqCBbWPmWlhXtxOCh28z6x4kXRkvTYq77J
69/OdFsMGp+Mn9eKOFGqTi7UIuzc02Gs/vU3iW/cqFU3isgpaPWcFkEZA6Lpg6i0FIgRrXSwutN+
891LQyLG0pWy7488C8X0GAuHRpsz8IkZ0SMIALGUBZyANMI0JmCeDZEVIfLnASCx8WmeXuTfRJXt
zIYwJfmPkCRrGat/MzjROKWrNuEK7JzurqS9xpvbzub/6pYGDs7Vo+Estg/RQtTxYDxf45oirjz3
dwEJbngwCvlxnqmYS2h3KbiTrQC36q+lqfUe9NP9RoJXGB5j8D32GkqVSm4JWImm397TlqvbuBXH
mZcAT7JItNr8HavkF6fo0rMWzEK38VF9CgclTImOTKkJpeHv7/tyhugAx+IhcWRNz4boSFmSG4II
vqFxc4xHt6MQradumZHtKRFoGeVatIFRu+B+0oc1os7XBjr6IJZ3GAqhGZ7flcbl3l1E6vtqp4oW
Ci01CH0CgGLIlrPiA8XgW7N5kZPeV35RGTT4DhsDjZqZptpHPYpI5eI7/95nqgbNTye1cx5iY+8J
aGrqwGy5Lrel4xU1JOWOPoH8b3hkJQNg6Kht5JxgphWN7oTSPxC45bbA8aa8xZjwyFuUgs/gm7Jn
gZ3UWjNZF8HJayeOeJzPSy96NgGtGAoZmIoQUKMoDyiB+p6CXt5fMt/6KSi4qmtvvyeVxtF7sIN6
IqM/qwYek6S7Jyj2Y7ywHVNsd+H2eDiZATCIM+Gl85BY6sguLanNdHoyOAlbc2W7XaGMp355D+n2
cXJ/+JB/rm+/NDmdBNKGn/WRmvXyiX/YrT2LLCLC9KioKx/o5ogZds9f/CZbp6DpN0UIJvbNQc9w
7Lr//Y7r3sg7YdVx2WgXUdIb7f5tmQ1Qvr5e3P7UgbqZHWN+bIWWgMcb/cnFB/UzNJCDvOU6gi9U
KtAen3hk3wc2Obqtc/ASQlTgfxhQnApY22+4MqNDcMvaSzadzEP2lu0sKdx5fuxQ6YD65hta3jCP
zIFpkLQVqMRerymi3Tin9QoQyfTGIIuWAZg83YShkQF3Ma0WQAYFTAoDsTP4Ss8+7LdXSihWGg5t
2RKFD1rHuDQq52o4EFR87t4epwN6mkQtQ1uxAxqWapPNTJx59xQP77NgtjCwOJaCApgEQVhYx+0H
j1V4YSOxlylk4idfo0+AcgcywKu+0SFaTZGkV9Q9wCMQfB2mS88Xf1gO7iw47iBK+xFv44eZETOQ
LkMZsWphfv1M9a7dyeQ2jYwF1qX/QWvN8CzW/DRx/10ddPoPAGsTbCxmyqjJGfybdbuVjm3I9bBg
PehgJ7x3q7STyLLjThA82+oADkBlckcJTXqtF15SBBAE3oXW454aYILjFKh5Dinb7PQsLPjL+UFt
1ljHwgospxeVHTBl8J4YLQLkk77iJQWvO3gkrJ8lFsnGNvZrkyVxlN+p5Vpt9nU7E9ZN2oGq2kj1
cddyOQhJuFsm/mlYS3/hW+GzDcPxCdGZCaj0ghYG86jvOWQ/VmXobYr06qT1ZaUtBFEQ8wHH7ULM
sw3rhKk1V4eG6AEE1e1fPTTyUwqv8La7b6Af7rpX01k2QaNpD/dSpnvf25RiLikUyLpiC2i7N/6Z
BkhlVOdzr9rML+PwSIX0kKs3yjcnLBx3Tr/TZdLEqRLAQEuAjJdtxlAxBznZHaV0oSShUif6jkbM
qH8R3VvhO9vDWnv96wRxLIzdHklClIIqvBY/UxoS0ti/o00aLM4KkWt/yw+az+Jg7gwzg6WbjasX
ahDy1YAnBjR3hhU+woCeqTWDCl6bh2LMV+xqMW0pYjlRyEujWSmYXv/aID7lqdxv/WWW2U6DtKL9
4ooTfrqMkBGqYZleJp9IvnOc6Cc6o3yljsci6I/MomxckHzybHNrBSVZHursQKLQ093Cn0AH0JrJ
GhfLx/Q7xnA2938Pn7OU8kDsQN778Vbt4vNk2lzN/02NiqcADyWiDsmpLFwN8N924i9yYvCyoCjH
oAlZzWMT51inaXcEhVwvrVIeRdBhDEjKaQukcsZTg/OvKI5I40KtQiTiIAP3lLN2Z1951TmuJ4rZ
Y9p5h4ZkAzhMhd3Okz9c4Z5Hucg4QSAnngVZCQyWyLaERBIpNfQQ52W2fcfaP2tc2TvKRwLj1wSG
cG70Qff/eENqWCLyNGGN/wTSjaKTpfK5eeNXG8FKEvffghObPQT+ZPr3OXkTBK+gPkH3SUMLIOW1
WL5HPiTR8lDrb1DgQoQdLUtbUdkF+zr1AedBkihs3jTE8cvX+dcdtiLjDgvKr4FH0J2lcFWPxrkV
Wu5RqVFzFN/Zr/gsThuppdy7Bq/7fgOe/lLM3iZZ5PHusGlcgxywwz2mNub4ZGk2zZgAy7gw31Es
6L7xcqaYKexGEYQxfrAqqlLjOyiW4XK1YfrTx+JG9ffIrhWMc7t6MgtAszGOAiP8zaZ+7SWz4nxG
eRM464I0Sai6F+tyexGvD4Tr3O16s8vX7wtc8YlhI647tLA39yPTIPMRVqj0OplwXI5cERAY8QsX
gUCkeuKQjEKG783RVwAz+Ml1trJQw1vMbyxsmPPr0VNgVe0SOw2IFZCOp69Eg6ohtFt1ZbmRRmvP
CmcliteV6C3DIievQH+3J3dwfcO5L5lmaTHzQtiC3060YOUi1CuwEsHECxH1cKBgJmjO8KvjmnSs
v1Aa1WpUwjXrjZw+V8K0I/J0+CexNVlylNNxE1qbcGZVmOEzGF46/nXQZNYMoWnaGMnC3AyrUmEa
yEAX//33/MnNrZPfQabb5CmbWeMfZTmXF7sMlQql5/9gnHnO9L1maD7aU64J0l846fzi/QPB1eDp
N0NRxOudoh93DvY+cCBU+zY3moPjahVKbkbOCemTKeLHCCrfdgAJNgr8N0m1DaubMeMvXEPAwwyV
YyhsI/TxdCe5e/PQjVR0x0899y/Cqot/bRIAtrWEshF9Ad/YPallEAeDvRMlL+0IIWhjHmg8Rb+X
zLsU9uKST0jqdujRUBAgpDW+JoDdOfwSePBLNOlFY5vGLEFJrBsE0pq1aEpq3Y7j+UCPEfN8F2FP
X9RQpsY0mD14ATl9qIASolbNJwmJkWKemGFTOAq3hYmyYAL+P3BdJ1qyIPnyTr0YiCCocgaBznuE
tnjt5sFFzzmju9Zvu7ARChdRoXv9B4Hjqu3dwB19UnfU5t+GezDfOLHiZBDXIxIRBery94yGb9Q1
7zthySVSttKBKMgkjbdAuCh7dhHo8fm4en8rQO0UNtWx+TxvwT0mM3keVe7tL+Uu778YOAz7V2x5
/X8Y+zazobI0o4dGWRlu0yZArswwuvUswTlXcFC9YmBGtocdutIfQvEcCj0z4N0jO1Uezd9CaSja
fwGH/FDbKoEEsBakRGsqGcZfEEzsWga+KlXV4J7rDGEQnMIiwNSOo+C0siP1a7O+jeugs3Ybt68n
+kU5734geTwXcHca3bVC7PxG6ZOJIFUtPqDkVvb/t9hJavsu5caEEYYqouCg/wQ9n+NH76yR8b4m
n6dLgqm46Lo7wHxpXhzjlQHXQPgZ+kl21gS9PNV9e+754k3vOObLhxJMW2jvvrqWT4D805okbJ/M
xRHryDyFDniqkYjQm3cAg1fMPlPPxrYD2NEqT7Uuc/MA9d0FQUn8vTykJD67brKyjcU0gBWyAdIu
D1f15EPhiOGFBi3hWlgy3CmihmPoggpDVyOJQLaKhl1YNjoC57D6xpki+1lhWPJPExPSPMqhvmXx
Qyx7TzsdTihbYvfGtgTswNB3ge6WX5SrMjkK+Z5x/CZwvXcBmpdFlneDSourBsCWXpxeA522jl54
pxjC+SIr2L7+9IU72JCyQej8ltPgmQNzVrqP1bFo4w/GPl/1Jv+PzSeAQSzfMX/SOj6jXCg7Baz9
3LSOaOzpmlvX4HuR4iAfcTs/lqhyf1HHt3fKnBguaZyyDThFhoNpLNupGO1YPj+70fifKcbSnezo
X+x5TEkul4Jk5LMy0Dmmt/nPVz20l4e+lfec9mvgF1EP77aFd2RbLqjNF4HpsbaV85W/iYFnDmHf
DVWOf7K1lJ3pVIKk5n+a9802A++1+Z4US8b06el6oOn1+21TXPPMuZbUgmZq2WeZ7+9pThOPtkQA
6guM8ScRd1N/IjuPaeMMY/91N6fwhN9UCl5Wcy3ozI5cuxrjfVDEsqq8NY3SDfi3+7QVxknp8Ugf
Wi7Aw90408ILbQHNOljRwn2NcWQy681UF77TKCwaArPet1tk4Rrr29oWoq8/JfsXJcCVO9WmvO7D
uLk4nA8u8kKDHpbVKdEzAhGX84ebo3uWhX6ZraIzPcc83bZMvl8mDJp+OGLm23ke2GZAcW3sSojD
SgaIgtgiQb1A/9AqJ4wKTnz5sfP+zfstpdpduvq0Z8aqNLeUT+ZrhpdEIbdg1XDcd95mKqUNigr6
qB6hW4bPs+2us4JddMV2GYtjnbxnhioQLMt2YJ1+zRjZEuxhqhVKPzulRQtaV8nZCBkwVgPQyGnn
9Ez3DIgGokX/JkL5BcJNHRZQy+iHKlwdZKVV8nzbBig0vYKOKj8ZkRvPN2LIx/p/KWkCO6f58Kq7
aMHAkOu3wWXkfoSHlvkAyvZMX/Qte39GPJRjGiQ94LoVMfKRXTLQkvxnFdZhNG6lpmZRE1bzcPdj
uNqfw0ks7ynnbsuOnYJIFvK5jl/s1W9WeYmtcwds/u3wj1Gm7VJ2hK7RgqZUgzuIZnIIWYgDoiCo
KsLuyJ5B85fxNM4AGAs/8WNPy0Hwmm/389mdgxMTtv+UZbJKYja+O99lO0OehGdP2zo/yWOQdxok
DwdZS+DbaZRKctZskXKsjDAiIb/1L/t3MAjJIH3/qAcKitIMiRnoGeZj6wKiLnT9nN3qTgjGe4CD
f/DfWkSGLYSO0u225xOH+lkjPfoySNZyQkOnMtCaPkS2C2y0xkDi6gT3+fPmSDbUr9CINceAskaQ
2kj6C2NLEBmnoCGvA8sr9ScKOgQXQE3PA4xoiuoZGJhZO0qC011mWLkRQT3IZz41MoS8BIy2hwJS
zpWZhvnpNMEYIig/KJcnuaYADUu3Psh0a2M0T4jJyBAzzC64irIE5t7RyxSptTui9fJUfm3XwuM+
MULbObgjVlkYVNBi3f5VFEkoCoDf2yfiF8n384gLPhGiBIj4zrOEWTDoC8wG3mgJS1VdDuBjfOyY
7RcJdZGL2XdWvxbPqJhTGdSR2OUWRveX+vzw1mGrLOvpUux3iI/1epsk8zhk88Wnc3bot9wXgjS3
0dsYNRGgKm4H5TJSnVN2zAdS8DhNLY710eQInCYUo0kOlh1JkKja6uZ286uJWHAvmwJVwxZUQzkn
nDl5WhAqweuFbD1XEQVSfJpk9m5nH49SVHu4vihzYnBgZq+auuTB+w5CxUEZfST3zcjv1fJq2+AX
opsRf1rxZSXmqctLnab1XQBoeAt/8PagsCS/i20yLcTNeSNFEja1f2Powgq81rYoQVCt1gTZGnvp
IGry9D9TtOq9d3/zBaOvCBnzw+Wr2QPUrR+T8TGzaxTzth80pkvZpzoS/9yy6YauaUBYe95fynk8
FpqerMPta7P4T8C2dxXgy0t0C/BdqxEbN5moRl3zAzwIOkQ+v+H3pP9UbVNIsFUj1suSw+ucW9eC
1RxEGBYFx/XTeo8eKc+hnQaK7Ab3pn2OcyoZ+3dgNBaZXKpGQtRPRT94b5UoKq2YvzfcCAMfJ7SG
CJYyo7ZxonksIxbt5d5o8WtdOcEZJdLRFDeuZxJ9bWkSs5Iq+c/QsCU3uBmoGSxlaZ7oK5m8P3Qk
zqjXsxOc4FjN4kwACiVbct/vjUxY2OiUUpfz1kwTPADqYEgV79Buux/BKfft0+Lz7YaR+U7wcuMx
+G12pcMJKgxSq7aZghDhQ1f+hVkEAappfEV4rHGvEDY/Z82ZnJSSsRE4TuALeh4vnTDVzHvNbbzi
CJuLc9djdXUBP9GKsqb3vWKFwJKyohBedAn1pGllOZHpuVGZhdJTib8nqKbTrjSH6mBoC8R4NTKL
06L1Rn0D3mKZJFgVqdwYAervz5szVquZttDuhqLXBtol+dSLyNW/mbiAYYhg5UYCPiLL3XZZBZUi
0i1cAHzLwPcB6UXy1ExOZJKfsPOwb1Dw832cKuDD3MSM4o8rYv45YN0Nz1zuP6eP+35sljhZgsNK
Jzh9FvDDevOtQ5dopD5ivwAY9TMlQbA4HXvD60M4kZTFzxLVrig+VAEA8XQPFG4CVHGlb0j0E1Wh
jELVUjWUJJqCz4+9a2ur2f1jgbAiKqMcCzsaatzdhpFEZGCFQYPxlUSZXW5xCCaWKzctnm5DakOn
6CpP+CGjub1x9iPI78+fMSaXb1ximJOCLiSuXhidtfYVq0AOPk6qUMCLQCUoI5GDEJgwWjWVzjKW
iNUutV1crq7tlt4yu/HMzLf9E1EZPv9NIOi/M5hSYkyvDXzWdXpNYboNxy9+Vy1Mc3BeEKCfnP7F
tNO7pxRVQvPWSrW5jAqTTI9KWzoSnbsvLmPuWrMZgisjwgvBXy7FYP+2udIMcj9pUZqRvWU8rNGn
Lu6aSQH+aOw+G98m1vMpVXiMFFGDMp22pVWDhMFJU6HJOHT3IbT2Y5Qan0ukYzGeTdV9sUWGkgbm
807AXsz7h+ACLrEngkMKSpkTIOKVpC0LVnLTEMIGheMga2SOYukHJCPQZiTY85cd2poMbLRyQ9hp
DSccs3MlIPzki6bW80ZFr4OU8xFgxCKqALICAyNPkWfT10cX173jAWrrWTSHRHDwrf5ufLU09iL1
GVc9LCl32iXmIbNafrQcYvra0AyzkyyJwPJizFqXohBJeamRu4eeitB7+cz5BU86yw7QyCHUq/dt
/jaCPIhs3o5pcEvauo30r3TZ0n6pQXuEu1CEKkpCEnQwSbYHcyVeOX7ydvApaKL9nVqGio43+Eqc
1qfo8OYNJnr2jxQMl3o+/O4LQtynU2XMAx8ecA8wyN1Nsi0kX1+xbGtaBAaecQPeHqehtlr5FdYh
uo6p/SHruvUNR0xsslC5DKi5PXyFgXG/elqX2ihJ0JmnO927sPwPsUEtggq2jJ1UCWyUguInGdg5
2AnA+CvBX3lf1N3ZT1tcL/4KDWrMXHQqzpO6dx/h/AtSnds6U8YtbG+LDKOTG07Nm+6u4lU0WhLT
nwVf/vL97WDTKIrtG06L5T9jYVgCFxFFQ5lRvgqsmjFgvBPc0AR1xUWS1XdJ2OcTK0tUtJYf2CmM
ZryrhWeNXAeh0TiKz8nhmH01NzDTwwKEbTPc0sDjACM1FK3lhh0OYsmyfO5Z3jGzzVDG23ySJzcD
MoZO5/sPGgAcmVCs7AJ8+5Q23flAq7Z3Q46N3CPMQ6QKgxcpUgC9AMdF/tT0bTCSVlz73BnuryCo
4VMudXnqgQnLWeDR/s9m8dVXlm4sWpbXJ7ek9uV+z5Pt5TRwgBJf+2p4JM5E61A+yBzlYhyzLsvw
NIKnLAnSB865hF4JD9cUqrzfRRxJu7mObXzl3l3vDxqbM3giWg1l77EDzOJklw9CqwSd7SPgDCxt
nDulHsZSShLgjNY78yKn7ye0/pmqt1JMOt+y6YGBahteJjDj8cOobppl7DwpyU4ZwbC4me0kIkRn
KnKZ1EEK88FPs8hVJhZfHBcKIM7IjXXyIFkIT/6BhQAGRw23lii0uyK/gHORNBif6C4Oa04WeVI3
70iIYafRHIJDO6gTDqtJSJNx1D2LCibykf96aCFhPYsdy/p//Y5pjTTN3iQDRdJJK8mRVWc4UteB
p280XaXwZegO+SIse9FTnmaBlz4tE0fJbO8osIvFxw3g37IY8GpOQ/k7zl/5mZoXRbuLUqSbalme
tM9vGAPyd8NntJ1GJLroQaxLgKJD6384iilwFRmkYoL7UO7jgX9l5QpckP/XIUDe5CzPQwMX8WHl
7Ezp/387Z7XxmxbhjhR8cKn9CGgHhuIMSkKpBxHZBG/6SeSfLgs8nTIfiAAbf9QiPmG+Js+ibQy/
0R2fqltAdo6MPp1xdLQ7KG+qZW8//Ii6rRqjGTsYlo50ijx8z6sam+6amiUpFWKJy1qCdNnq6Cmm
acnU8EKlxaifbAgPWUKLR4/RggxQhkx8OPiXEUW5NaoAdQf8wKpP0g4fe9uf38O/HGhJ4M2Rgi2Q
Ix+wMeILRHo5g5GfgEhNvgeDJIzbQZJtr8MfYqo3QatzN5Rt20goKwNk1+loEAvI9TYZOAnzb1aB
tBb7GaIxVWxXQeQb0zN05JNG0iAfNtwCKoeTfcHde85UCANTqJkI8uu7PId7YyNuuXDhQOwcuUy2
0jb1KVFGcNIbLkZL4eQ1nHqs23lTQSBYlNptyK7+dUEbR43ziMxPDB/HcwVDavu8tT5rSkHFVOAI
pxCJr+R7cU9c0o7k8C7sBakTkyHC0IuQlEzdWiWzOZa9PWmlut5DW6ADLmc/9n1ipF7aDAYBiC/h
VBhb31ZsdppDZtFpOXVI+Z5/8qN2/x0uTWWrdcy3fYEXRmddjfO+3pTiXG4ALDX31pDgyPSHRKRs
bDB5nIHOXvG4Rmxwx9jb903bl/Jcflxemnnto3Opo2KWePj1xeEI1nSPYdVAJH7Z03rGkvaXBFTW
mkZ33gMSnxBFJQ8xBEONMq1szqqGtxiYtIA602sqSajqXrLMpIw0BREbuxfBvreQfIU979r1+WXg
h3C873NgO6ICkXTNqeZUuThuZTNqhEIvDOKs1O/D7ZamSadUvgglR34+JxJij8NjRaJnRyoQfu/c
5HqWeZpgdCB/mDxi9VRHoiRwujhQo1xFYIcdA+AZRIq3WsszbU0/GvOes1iuCeAWS62uT7S8Ftl/
iVff1hKbuPKku+0a3OI4MgfjCsE9bXjjmZSA0hjnvnJ5t+eXrEe9EMDUqYSjIWGMuBiFzmblflPJ
/QIkUmeevOCHUfvwTlh8pJm4qr9TUw2g7/dAqBdxUscqQ4O9W46DRH8uPJb0UpYoFa/rFHoRard/
k8Tq8jgBmGQEIrpErVSN7CkNRZ2pzIhWyupMxL1hWoRagRUUdFvoZl1GUeRreIZ8WpZXgXGqQpOA
xNfRRKk8mxyP0nksKdUqcg1g4g3ukbZ42138iyM7InGvnuKQUkpHX3ZNrRVZC+1vAut4ejL/NAK9
LJqiaCW06PWCuYitnMUPDfl0L3OhxmxmX4NM2BeAEd6q3PCO8bJ8sbaJCa/3txTWUHlXY66y/GW/
Te6EXSnmoNZGC9GGT7INmvMczvZgqxFbxQU0N+i6u+0z3Qry1x9+AIWHeSTKHccrjvszr570UTqw
FKbqJ6IMNtZM6oF+Y5+dU8z+WTSasuGAAWUla5vqfROxHWZyzC/2puLTIQCVdr18JL7aB2NrI5Nh
drS6QnBJmQIddvyuyO47qVu4jz/f6WUxTRc61a+VkLZ6Fw1wQrMMcDMXIDDuk9Rhocdr/3rtu4jK
DprzysEMJfjgkm98eHPOhNl5uZK4USoI1yXgSAfKEv+2HMqdL86GS8f5AWB3vTRJTp9gYnq6dv2V
GASMTB0q6rhl00mIiRL5+TilpWca0rhMb0rV1PngWaBIkDPCcYRneKZLX0GIuhjRklbT1STDDIux
hdzvUsyvOEtueqLfrWkpiJnOBOt0B5pjANlE8LxIskS/42K7qoJGf7ZRQBo+zhzCdZESQmfFShko
2jkGetkigVh0cFzHRW2qSTSiJ3VwEgaSE3YSIvgpg40oVAOFkx6F5E7NSk53KsH3jZ9xdvNRqCZ9
81NzMbYUng==
`protect end_protected

