

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UYl0oXbWx07H12+XLY7LSDXLBZxYP6gTZvYTz2TKJK/HlMq0/MaxTmoFA++KzdPqQG+aE6ZPQ+qq
Uf5f81Uxgw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bEg0+1ra2kVZdqsGzhpfcP3LSyFAfoGp5V59eCFSwsKdv16KOkBLDiHpDDmfz4FuBKQxM9vHP9YI
VTTP3KvxWu9q5eBe18cRw11tkuJ61s4QQZID5Pdl7K/z/J91Y+C2pZgC4PyYfdbZV9nqC0rqz34N
t25TMZ4X/3isyExfaM4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uu9uMFaVElOirR8H2+pn9gEMn17E//IYYznJRRoXYZmK9rFyndxvWxzgXxJnpmdqmEWjml6gMm/H
pembPItxQCeo7XrM3lTsic9mzXXAieyH8uZnhARAVJRKdWx7M8NVCShTsM8b9SyZmEbyJbc4S6Ot
QgwnO11NxnwCoi4JadA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mjXvcb09NMDr5cbshxSED/yd+I/z4J19W3+kcWNP/OCSlWn1szLbF7IO8Fo/qEP3dvSJRly/ZKmS
P9xe6HqZi/Hq51kBCz4qioiB1vvTlc/LH1RyHY/WLqF0RFuHmjhEwQpdt4Iq9HALjkDyoFAQOLvh
1tU76/82ig93joc86dKaffZE7U3TM9Jph+IFapSuSYa7IhWH8QczB63lTMnaGHkoVrByWTXAptds
d2R3ikHwtMRxJY499uEXii1jFu5QI26PCikka7w1lgU+SjOvMCKSRdZ1iUl1Jat2MfiNiCqYAMoj
DlISuFAyw9808erW2gozPmJueN0p+foyMN/7mw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c/1c469blILitLPEgX86SdGoVdvoyvD+/mS37IQOELSF9DiZ7DNf22AjlyJ801EIuF2kDm/eFZ7P
QeSl6otd//Msh0knUY7GOjPiKvZrAqibedNiMYmuhgjyAivYhuuHW/qzCXcwxk4zvdSD8qmkBkow
AoGHtgbXvTQrLELWSOJ6kJZrrsBQXOF/LEnLzptFNvsA5mx30A/EhQUwiTWhLRCs0+ZmwoXPja1b
iewVOs+yzFKZxKCXtAslkXwj/v5TAyb7wwAWtv0TZRZmCPLXbG/3htYoj0jStM4a67AxbtJ7ssQM
lCdCllUOr0IzrU5AZgmBqrO+RYeoA12X4rjPaQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hUc2uWOKrgaR6N5dF70TyOCK9ofPYM1/2lX+qEswJVJBduhXVmcxmi0OfBsyfbBOXlaiN9aeep09
buHtyIvGbh36KoOH58SMb+I4sCh75XnlL4Nsd1B7XSIJqyPQs1i+foBbthDqV7JWczDAdgLzhQUT
29R7m/ow9arPbR9LkWhDfFTDRDdhWkgTK/i2hPuXpSuh01iwND2tZY4rwI0aVM/Cdm3eNeMGd3To
gQc1cJ5rut/srYm5QBf8y9aMmvnwM5epeTVH5j/o+D47veCwWGXWno70XbYsJbNWjoWMlR/ARJE6
E+ra4UJgO17qX6pHvFKbOdqIVzF2hfYgExvVuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504800)
`protect data_block
17K6P5WoC17HcQasQpJYbN1bLLMTrs652t5GoopyxuEGY18KHC+/bWfYvu12UAxqL9yglgCYROex
ww6uRyp5eF6cgA5bzlL3ZwGzvAcNFZSyM3LK8fHeBqrPq/GIGlH359Rxmb+xNF+8ei4IqgjtNXtw
Wdi12xV3HbN23hwEKI72fNZOdY3lquKkCB5loDplgwZe2gozpelzoG7BUafkWun+F5PgrK/X+M9z
kvuXFcGgyCAMyNka3L7gOOuVsFPtagEuFF6g47J4Mvez5erLcsw0bzPlXhdfSdacdMsodr4TXCXC
KvfJcE4HrlgopyF9VRiIcAPbQcQRZ5ZT/QowEWQbywYkoY4SiMOJCThzBIrWJidc0RfZgHb4g9mk
u0KmyqEWA+D7fNNjTsgcfCS98Jc7nVtOa+L1OznSBVjR5dFNaSgzev/6iH9VD4d57GxryhDxPnl9
chAqyYG1JMVBb9Ekl9PZgZ/8SrDMCaT0OBwY54wAM8aosxgwFwY7NAliKDKaqoFBNXhXbI9irLSE
47d21fjRurDE+eF3Zm6unJn5RNW1CFDSNd36C1Jcl+xY/t/XaGIOsYmvtRyn1xx1Zy7t4KBRTB6U
+1DIWzLO57vgXsyc3cz0VH+C9F81BQGaz7jX2cQhFdHm4cjkycDQJ36hFhTBU680F9LRN14sffZV
BEKVoXLVA99+eLe7P1JHzF19LTmIDiDBPLE95cg5EAeuDSXgRwmHVAPok4TH2mGGsg2L0mr9PXln
WOcsuLnzAeGCOgiZ6kwOo0GGXqlzT4Ik8qpKZ9RhFZtiDMRZ10XhfOixqAqDWIvn0Pa/71ojqTT7
Osqx/gfEGcmPpoyqiTW9819/HeknLuxWY/jxRhWP2EHUjLC8jMmEUsSfDoLyD9hOIBlxytoW2ksp
5KaOBlsiqVssLwxHcwlR3rnIWbrZP7IqLkWtXxZDjWS+Hkl+k+g2gmHb8oxedo2PovZS25/Ms4KD
dKKOOZXjd9/7kTrCg/dNFM8/EdXj/SQPWIcL53VVx5lWprHKRyqkRxE/WcH+goXOCwZFYhoqEUnC
gW6XbRO39LwXnKUIwZmv9Stp0fVBraRzgVozLnAeq3b/jeNhi7dmiK9md0ge7xo2ZM5bN4hFTFTG
8cUSkhhKYcV4i0X/SNNIfiEk+3NsUqdA5I0Mv39OpOmD3qR6wEhx2Zv8hwBhhacgEWPfMZkDtWmB
f8eRewme7oPTPXLUjSPiW+3GyUuGkyQw7Fj1olcom7tyPdYDzsGTTX39aDHF0DMlp1V9EJW6BMtq
INgP7M3i95+fIG1BVKFHwf0FLntNylnhUgruyOrdt34Loh7SLzL5FxJU7Qhq8EW7N67fs9hy8zTP
/w+Lf5yLE3ivBgu0DlPa6I57n7ZjdosSfdZjLxzwkQ+MStVI9+oTGkCNKdI0rtBIYJwxX221dfLd
eEkCxZ9yK2Ic9Zfz/YCT4AZkrcbtv8Is7ebnlwnLe2GeN9CkSf5x8ys6SwCDI9xO4iv12HTCJlyR
HpFMJFEykzxDRnrqoizU5w1oTHPyO4Kbhrki+f6SWvNolYdP+mCFEo7flJJZnd8+4CqvhCGFIhzU
ge8yvmbW7RNjhLm4EoJht4d2JjlFTCjE8wEob5dXaAOYghqn708JjiyVIOL+KxuZx4BXS5Kmp5yL
YaqqbdEo07wyhb4mlr9k5cwtYRJTVARM73+DiHlSF3TEBWuSCsIiimul/iHUNCKu0t/CNfNW9+O8
nAURsnaCKCtxfV6eQGmWWGHupRS5oIppLMOXYWN9MfJ7fZt4LRv2T0d9ZpaDVS3Ck6Wgu3gOMhB1
Ig02YUT3eGcTVwZnrSCInonfL5viDEhCmGY9EpNpqG86Xz+OPOs2Knt1EFqLiL62BfrTCRL6Pee6
v8HRJSpvJOWeJTIaf1H3EMsWVyNoNlsBBnHPyoZ7yA/azikats/R9eY8VlwgjpcjJMFAZEvzB3GX
JUIAs8HstO2Ul7z0pEFX2fsAXOcObU1rUFekqsbI32wQRortcXA72dNWo0E8sEKVv8kmy9mIdc81
mp/d6/88niisgySQIhz33UNV0zSMmwtN/S40cA1W6wKY1PDw46VRc83lUASWg00Aznv0SG4UAG+Q
n9tjcubxj3uwrLk9mv+PUAnXZw+iFGsfXvVNhM/RHHhukmCZ+yzO+fjKEm5mZSaiKiDTyzSBsapZ
6xuaNZ2RQk/ssrBZVumgXdHWoUAc/nJsS+C0q8iIHdpy+GEcaPxrSWOAvG0tBjm0oGF5s5O7K8uq
g5+qh+u64EcQCPj3OFrOzVqvneTr60QIEsaGDAWU7sINE4+g3Y9S1B4bEN70C9+NIxrPZGEZCODc
/f+s9dqdppIIgKxgMshMQ01fwx4Z6Md0E6qH2Ufx04DC+xr3IwyNfodK7L4CFcJHRLcq0JwnFZHZ
JbMs6tYI7ardnEnJmSQBAYLEEsunV0o7A+auSzwgjfshc2UXfXuml/Lv2KIx+pKS+ihsp7GaOxSW
dFcQFbPeuJpx6CIqXMVB7QkvYox6hr4FVRpB8MZ8ZmJod50HturfS3MVhnYYLUz9Og5bd8TlnGHl
ctNsv6+kZLh13EV5lhwsMBky3H2bdLlSns3avOhQhbamALeYn2nRhSScp9UjwYV2c47rgX3xEKa4
X5UVQSSaX7aRZfFl64J2pGjxkc6UBlrbOJAALsleCsWY0yzaVBj0NzHW6YFVUtoeDZRoWk3g3v4m
TvZwGDIOkVJfKqbDgz3w1xAjoBzqI5NAGKXhgnl904UNnGuaznuCSSBhj0ezaDIVJGbXcTX0ISOr
37mlVQy5J45t6X2Va9Kb5rzlnCmXZERJX7CoPCad917eP1y6qwVmMGJy+NZSswmsEe1DUAttV7Gm
FBvTjeYEBVva9eMKeLByHI8QYbkfaiyQ9WDjvOtxRUcAO0aTFXsOonLfL4WjvXR99VNJMl0YIe/n
GzWJ3dvXwmMHvY2Nj3bv0jPwazgLUjQOJK/fJc0sFvZ1JdYbKddH6rmeR1PZl7TF7p+2uN4PGLoh
zNRfzne2uCJmWH2FsQIbz9hgCXyPZ2jgt+Nsrgj2vW8B1o0DV3c4p8fk4yxyXpZ/sAM8lHXcGwPQ
apvbcauMe4B27hD1Wbdgy1DQA000MRv0DtrMFrsyjnMRbhSSG5SoFFdTXzJBXdKmI/pSFc/FI/YK
YZBC0amXmfzDA/CAx9SEK5OfwdKVZCx4659jQoK23p3C+ZBF8WxjzpYNuypjqhvCkvkLN12wcrTl
mjOMOcIKYYOX+GMkCYJWH7gcYPyuwS6R2OGfPkMVAlI7r+m4WvJeTjruDR2ufT9zY55gVcWRAdM0
9k2GxmaQZflth2/ig3gqs6VgzEeqHQI15GY1QL2Fyxgn/insv5RezFDSUIShDXDSi6hffp6IRtCt
Td+N3l7BDhMdTo+Dgqnqw7g0D/eCeVfoLUTFr5AkGDF7ZJpdQRwEAVAy5V3Pc3w22QXkwVUgdUvX
Hsq+TrVy5t32OIPpe9gYMfThnkgmX2e0bpnwHw8mqwIEOxaRG0XCJJlCT5nJrV8bhCcvbLKrawpX
IFp/cHgsbaVockCLWMgOFmUgQ3ZulqoptMlkeP8121bhwQgSHTCyovi5dyq09MvQwgjNbdtv6FDt
i7M16keQ3Ztb5o4M4I9IChY9NLfjW1MQklCQ2INjtgSy7GmFqMubr1OCwY1sB4UeJI3v9apOkmD8
dKhk8L/oGhGxWFIYf8K03JQy6R1SaKG0uWKg7OWpX9swTCc/1aJ77xlH90XwtjsyuXaAxQIw0lh3
Xfuj+aFKYyaEy927WH5re9AQBgmMcuSblXWigJLYIfK5Y6wV5d3n67zCDbRvul2UOdjDYdOiyA2l
W3hUhwdwyQreoaC90LxbvXyKbpR1tVXK9llRRUIC05Jckukq0rJmPXPkJFpEy3r3uMSC8YsSyI4w
73p5NfgzVvA6cMj1XgVZkZ3Tz/D0rEhWC720XqNVigHXeLe+JeBUg+hYS/79+nD3EF7c958wgPQr
dGAi/foW5ZxMnSaRYfse0Rw6lFNoobUry2ebjAPScbVRmQpLgjbLSxiW+bPK4xR1rmySbatge4Js
ea5OH38hdUyRRSYxNBIHqpxMx2iF3ZSCnHgc4EW5/gdP/c4dTSPGvjvvIaPcT3r+f1mjI7II2FJ7
M3Xu8qBdxeXWp6sK5hRWl7PLmRc2oOt4dBf9LskQV5A/GUIFgrINRDLeobUszpraWUHvg1qrZ1mI
ZCpA6xYOnO9sb4folYQNMKyYiPg9EdLGZGyuw1muOfksQjTTq4jn/dwzL+4mNR+68cfDntjoYhEQ
WlDyiEp+SIke7UES6KzHuS5lxbrfVXHwR+mWe5oXDc/fmEpTL1NoEcW7sZ+J6O050L+tRBsCUfz2
zRey753Xs40+IzIIDSN2nhpLHFNvvMZ54xy9SaCHXuQ9K27x7surN6HeuncDTxNBlypB+GdLaMzl
KRQjTvyxyilndgMgAPl2xny07TGjtoYsVWsphvZ8R3IJqVSV/B/y1aq/8kAiyDLULAHSoiKpq/em
OSlcieVik3HEyo7mH/NqIgf98olIdeGf3Cvs76czKlygwJ1Bd25eTqQ4qt3CZVXrqEtXgX5x8Eng
XfIIEFSV3QwWBVhYDQOsOYkxuQLRUht7E+wMWKwKKxhqGyFCJjnk6mPzMUE4CVrikIaoLj5Zjsto
/FmTXrnSfo6AmCQJ3yEFrI+iNat4kCQK9oGIU60WlVvLMjdugNSJ/l4iEHWFjdojGsv0wcKDLAmi
BKKF3M2WlcL+corNqY4fi/gq4Kngrp9izaDDV9lwM5bznC4Y7MFGJldz8VJTPgFKV9o7qefBLsHs
WmwiYPRVLJLo3kxshZ9ymw0LGcS0YmBPfCkDOzdxgaJEKHD//Nn9C2oCR2+6tpCSC76wqwUmD+WC
hQlYMftYWUJcNsYQlWxXMdXYr03I1+h7xFHP3Ipc3h9rmPU1U+ZzqW3/8PBPnpk+84dUfnssXDHE
mM/z1wjYWi1ltGF9GrKwNdWtc+jOIz1NTWetf62HFDvjKis2lu4WsFajwh9wUNvefzVUf/k5Ncel
KmIfgK0OX1dASfgMuA0ntSPIEXveka8G/utuy9QRWJA9y8NurSVzBFctEorKk7U3MsPz+ToThyJf
YXu6NAFrZmzWawTjgW1JUsbIrP44LcXc8/H2CKw1oJdojMbBTRnxTQQHgOJa/0ZjKmy/UxAZAqfp
Tijc9DX/EKTDpPjfN8NMvqK1aN+tsPTrxE8G9ouLehZ2J3CZVQB6MFCKl2iw2Gwncb5ls7stEpz3
5BdCly7oSaARJA5Yl6mSZbyxDEuxE53GTbMQmxXoBd3VqApCJI8tjSz85arIFDExdpoa17ZBGvnj
WZgxnyv0tZMoh2HdKskDvOVQ1SsLJm8nex8x4USmAWyuWgB6l1XLXYCvR/ys9zwchA3ZvuxSv6yX
FQePGHZDVjlLiZrsEhVS71pKyvo8dD5V8eKJL9/DnRMBIf3rd5P5QQZ4IVCkXWgx+jmfkJwM3kG0
D6lp0+URa7kF1ovI9Dr3rQI8TRwAFbD8Yj5nHPLC7klycgsBjOKZjVUNCoK7yKMKewSpmizKy3bd
r5/NfyB7OLA+irmsQuOggza/F4i4Q1fB23T5JsP6Nu8TeIQMQYkHsl6Xe/l6lCWq/uUpHjkGuSfm
k4YJ60kOPSQTSz7nZjOtPV6IvWD/vuxAtdSSEe8cez2awsJY9AmWPcWGP+CpvUTKiCJAZvVTRO4b
tHKdkeaAXpjuCHFLDxaRqlEAdCFLigzRHe2rJlyHmT9+Rrxi+AuI1ddCKeaBMDvWVxgpwW1ECkid
TQ7punaaKpLPz0bndBDWATGbsIBDWDUry4SGxTVQeQuOQ5YE7sXkIiwhk9eraH3XoH3/CilsI3yb
hCIHh1MvhYFJBqacOz483//Ep4/KA48Va+YJLsOrDlMydvk6XH8iyXdizG57MAgrAzIVWD9eC3eA
ceY4uYu0OuzkX1Cz6Wh0DH+qt7puzGjiL7+fhFDARIQRCse7sOusCn3ERGhTRYdN5Higv+cSgp8j
nC6FwhvwZRNoCZpo1c08JyNJ2ZzGinrvKGyJnCa8pGt29dIlJQ5dc+fji5UAVhn/PJHY9vHI6nf0
ghUF2oS1fVe2oeSDP9XvqROVlaRw4b4GsZ4CnAsi4tmyXjmmXQVkeraGROa6noQ+ufay6JuGBVFS
GE0z4AH2jvxv7/HTH1kUxTxL52iEpLDxxx2PbjkOsLC0MQzgWmO7DRgAA1TLlbAWzjY1d8JaBU1O
l3jeTitM1agR48s/y+FWrl9gk4shi7D5LPD26wCHEoe/u2lLrgvwvjJxzGxdxD/ov/tpzwZuhRBd
uXui/ssqZg8zCOR5YZuWDLPTGkcrL5urflKUPJ07jeT25PbW+/ACUtaffb/0VDBjXk0j73l+l9t+
eVgxploNgtl0WWOL2uAqiOQIhzDwEkMT6FZybJwoIf6GglcHNkMhTJOF8tVuteuDixKB2A8xnA+1
rT06Hy88RDmud64bnoUMVl3aX1ace07nMEcvEhCmCY2XUEQxAZfKUApIlC2HP+oNALteeGyaqhO5
+Q+dfJcmKviJ4MBA92xC748ncyoHLu5xSXXfTEcxfiqxnyrLnN9gMieoarq3U5W7h9MDyEIxX38a
rEgPpON/daD4sLmL9TdndmF+7cAZBS4tfzOf75PvCsXD/jU59PIF5KspMK5RoGhBZJs8HtCT3mur
GyKnZiqixGFQMdMYqpIXOhHgybg7r51p3/bxEoaogo+ISuLm3xgj8G9FVqettJKPiQ+m43LRPejb
a+8cdmtErvyoxtC8ewCeEQ4R8GBr0EVwI+UgeGtH6enczGo96ud/akvHXlCckZRVut3ifkmkPknl
TYJG4CAydu1ad7fwnGTaSnBrUcb2VBb6zgQOcO7YEOWbf8DKxy3Dr0eJ8DxzMRuT9KMMUnMddghM
Rh2qk5ItOC3luVagEoLG2Q1gftSj6hQPXDZSQsJ7erq8NbRikmzeVYvxUw+0oTFya5WKrTV1hB2V
bEdJwy4ImESDVCCkd/bFK8OZR98FHBuyHabIBK3f7o5a1vpUQi8tv9SHu5vqJ4cYA4Q7y155RPBo
VmKfe1OlFSlFZylvITnLJmA0bUZ2YfrYJPR77VWiXpJCCzMS3/J/JZtNqFUYqdarenokLjy41Xus
mnzZLiSk9qGCaAqQw/WchWTEykYyvWHIb1eHtrutLTcRWqzizFde9QN4GEEmN/ytYwHGN8nnzzIg
/ZFcuGgOnGmvrZ5vAvOUncchyg7qewvOhYRmBT+XnBISjGlzQdE6qN+81aHNPhI5vBj/tcayq4dV
pagRAFoYJxvT3misFV+7v/L+0sUGn3N5O54yBIl6l9Hdc+a6AELVZ7wl7e5NXcRc6KtEoRETjUz9
QFF3VYfmt9S562agSQlB3krTFOIdMcU3aM9sj4LGX+S2GDAbsfYOMtSjZP0/jUwUJ1Yy75e6AsE1
4jVhM3pheAwgOYG66A2GRl0HAxycVDegRnCWcexF5hiaOQP7e+3Yt6BC846k03o/CV5JubHnPCKf
2/sEL5JOz45SP6yWnhvtpXUKYK66QasZxU7rim7WzXEa5eeGMbQ8FXdbZJ+HYu3Iz1lLcRTkFV5M
lWzyc6fPp1TbeQoQF4Wz/yap58S6bSXSdwD+XDwzatOvL+08RZI+dWON+GKG0LAynh6SLsZ0T7vv
mcU2ot+DhQOQIEmwG3Dbc2KT33iRTXHJzMciF/QN0dg20B4nAgwxJNHl8hG+c41wJlvii7Vvr7IO
v5/i3sec7pLHAB28OaQOkC6UGsr2rXE5LUstwdudchHmjIL7aFOpTFsA7tONkUqnXyJsAOEABwnn
mD3QmwrtJFSHoQnhCEOzlr3EG2wX8uNXvSS28GC20h9xPenlWecLPyru2EuNMLcTcT21tb8yQQdO
9xyD8NYy+xYAQs6Jx8CBswxg5gI9XNPJjfsEI3WcWIOyosiaoOG24PkcIsyDWxS6oUz2WmuUgz9b
qESjSPByZDi+4dQW9aDsdoTBTeTySrVMp+YGWsy3uUCKbuGFUpVseBsOecU1EcCR3Sn6azM7/BbS
oE+z+bcPra7tfCL4AwfsZEh4uDNmALmDbb3t1gz+lidhQ+K7mXz3akKovpiCes+J2LvDVXZvEadd
zQHDlsbnDZA5710ogaIl51Bmcu557J54ABy77EocG7z6RyU+XwsyW9aOdxT+/RcsxDLLMhGpkYvA
xzWnb4cEe0HaEZeZhfCTDMvU86VYwVgg8heUWB2veATVAE+HC9Vzd1MuOo7vadgg0ozgYWkaipmp
cNY6mW2gZKXq0w5zkdYSiQVfxu6YYkEhKFjx3CwOFt+gp7IVEHimIpE/Y5L9CQFtNmVpjVhboN8r
yWgFjYXlDeQl9aSQQQGgwiRnTyJAmzNA0zxKeM3sbkOs+TPLjT24XFHKW1WXimefO/ItUGEYCPir
O07b2MEgeWZUpU4WU+ooP5R4WRS0rmwBf647HdJCtElezgcURe1TLIcWl/Q6Z8dSP3xgc2gfn8Iy
tC09qU7/u0qGt1qa77YWMn0IsZGXw5PGhRr+llYP0LbPmCHfGHuOL7LeKk0Z0vBav/cW9VdIWYxD
CjJf7sr559PYd5g5wfi3v4tYujap/PFdQ2uVNiyt464qy00GCJRK3S4kyi94W3WmrCh3YKZ/mhxq
n6HxiCwIsxWQSc/dQ9uJTR2mCaU+O2bCRm7nWUvMx4cH897S1Zl9EwGXYAezQU/cyOsXILZ/Ity6
Xp1JChl41WLXCZL0mHLPxcZTQ1Pfiqu3pVk+LmrUeQ7Nb0KRbJFONeEsSf/pbltSwVAnS2njLYVw
lUGvS6ZC8RoHjsfKQ52ztgUGa24IkTXSsDyKIRLxFUYsg+1jv1boIqImMImZCtdZfOUCEUfaCcV3
WKcJ2ZH9m4ZvhWgj2FgkKoroSmJTPXst7twh2kllwd3BWJQZexRJ9JhwMKhHCbgH8qW8nmnJjpra
t0RjsUlnfjdYvVTsWwnRi6aAbx9wcK//B2Dea7WdlzOQO7QpG1gVxqRiOuLG9rpcjIT/Ra2kgWl2
VHwNCONHppjHH6H4Gz/thaBSkwT1OaK0HFODygjGIw7nJmfiYzyclzZ1kjsmHBgROozh4oX+FcLt
TF0hJjsrainlU2v5bdg8OQtnyT5U3+vKee2QlN1rRM44clFMkqZ64G4CzOuYiNYr1aYouL5Eu9D6
WQOSdhmYlG/rEgi3oPLFfTG0xCUiWlmLJwz1m70oDAb4a8zeYJ9sYKBzuCCEE0UNAQYbvPrqZoxS
hThNjcrSVdk95qcmkMcPzc3krPPqItxrxVmvae9stduOZgDbvaSOPzgKu/MBYmwSxc4klerYH4PC
s1LFTo8KvDScjg98g97M+YsUXAhu88o1aRwIu4nt2nbb0JNfp9nsOi+dq0T38zIt5zDGrx8fSpMq
yyQPVN7zO0AStvtntgpbRoWDnh2vyJTIH7n9o2v0B6IyKAXiDvDpmISjUTa+MF1EJaT+kZqGPEys
1zf0sfp6OezxNbDSw82vxSPtyHS7nVWxoSPsEx8pDaoNm2CZwAXD3R0stYf95FvQS5XEapGsSLeq
IY/5/uPsOJDMcBF23Yw4xEsH7T4oBOuv0MPA/lhjXmlc8OR+bFMtTMqTDJhRmJpv+zZbpOzYM74w
UD4qJn9509CYw5j86fUNR069TFByJQ26vAAVyUVIR3rMjsSqYfvb3mBow4qRW3kDcXE1UmJQ7myo
4vOUCePTdv6PzGozeBMMjyLZkODH4vBmk5HFxv5pRvho94xKCTRhjiSfQuBdgd5cVpqL73ze6+WT
0UOd9OKa01xl8frMDprSS5cSbSXdrzOyDyPQmzbClMDl9fXsQvTvL5vBAdW/4k7jPNutZtXYdCwI
V1GrRtkDvsxwIzVitL6hsXQqoQIrwebZflriyLLDUwI+VyWXPFDGx+fW2QwwIZ0vAbHXhW90btzg
mOK4OAcJL9PRVVYOkhoB5HMaVwiTECV5HSM7EkWPSSo0XPdw4+KndNWGGjpa8QBb7ZNd1P2h4veT
8bpO2dEUf+Ph3xXls9E/5meBQLhxcUVX3WrLumzQ1e86gF0/Rd2kukzMjYBUxf6Yj3VsYFt2iLDC
tsn0hSRHyCqSXeb2N/BGkD3izISiJ0ObeiH8lB7YuuNuQP2ISzTNnX0K/HxbhIhQP/OBRNLI7Udw
bbbSlSIzhkeZV8Kt+9FPnLrLE0QlwXfD8EgQ+dY2KzE3J/5CKKh9bUgZBhIXDC1fguu/vjGoznPN
PG2rbwIYnpp2V7xmhCnukQo2yatWLRuAWaJGOQ9yYPzKuPwPepTE7gaX0aNDj5ezArZO7BXKHRXy
JU3EYbfyvcx+qo4+GEhfa6USdsHPd0UyiM/3W98QZtS9Up3SZdXVkKY3HYKuFbhrfIAD4dg5xwVd
2W/38UqF3FqXoqGQ97iz3OKJ7/bl3/WygJNMlfn6IPr0bRXm/8IV93ODYtd5c/q9HsyBvIgERmwn
e4wKkbvckhahD0k7o/LHBv7hA3e+pKwQbL36GXFZfj+/qVagyTJDWGljhM3NRsYXhH0jwjTvRyQ7
LV8k8bpOfV63WGOQbJBc0+QZrxP+eFvEy4F7DLSQM+EEmm4cS73pKNoLBoB5dmYpY71Jk0FS69ZM
H1bEh0HgxY36Kk0a4i7gN4YJqOuzDMnKhgjk4G20b3LPIJLlV1xC/9R+PRVadJuhu8RrEXTto7g6
LR53QkEdt6F1wlXBZEqL5UVl3S/J4FUzJL/rO0S9R6kNPE4tzCaMbVCSywuWpfkjGiHhY6kQSHKP
uEK8wIVZ//s+Pm7/zhV2vl62Hi7ECtJFTYQxrF4F/Lc/86d0CpdRL7/6mQqwXpTJpTLrJG+L8kxw
UNiH1qkHqWLWcZMwiAT0BRmdF15s5d940oRY/I/p/Sw/gqCs8+Hm1IB417sGyH9migNmt4nT36Sf
t/u/O8rs/lvEnlwT2w7WUObXvcinlSTQkMRTtZKTjGlJrnTyist2opdJAim/1BjgJ4bdor3268WA
dmSEN0y9iG9sFg16weO3b2BQCDCVOdgDPGZTbNeMCcG8nBAOeOThLIF/CLfQSo4aCaaY4JWm5G76
zW5vO4vHbXR6Ni/Q/cWkp+1cMS40HXWPHGq7hSQMz4kJL0XFeWknA3sYRJae819N+EozfAXyAFzp
+EINPLAy/wWGeWfYuNcVKZvn11pqTg6d+JMqH1KKiCFarBRvAapaMVxZn8ri4eWPEjuXKTBDAKwW
LVoWyfmIx+xuSesEEJRGyZLk+8vKi8j/wpeHS3JtiHClPrp08sbjiXGJIK4C+FsMvSrKHvpZFA3a
Erv1T+l/gj/cUKvJXD1jPE9wZwiMC1cze9HAchgTMXXbFlFWZfbJMhcJSUjpEJoN6oxikuc2ZuLH
Iz1mLN1H90vYMfHo93nVKw25FA1PKU33tuLJsOrBi0tfxORMIo6GkfNcOQNqzB0IGjKwA7zwnLai
f95rh6FiwG/d6Rr7HntTnxHC1SKAtS1qmzjpqdC7g1sb5hJGv6a3yngl3FoWdnjG9/onIo68aKhp
lxINPKqdpqtixthKHbjhwdETMvyucweCk2ZgKFc8dBgTsZY0oswky9gqQlnJhFTWPbF94ZR56AF9
pvkHrH2lHCUWfud208v9OGDJ3ddCH2juxCSeFig66xB7LBrGX9VIy66cMQMCdYWXCiX0vuYjwThc
9JMeQQNTkjufZPc4L+NA3aUMDp0HMXiMT0nM8XUxCVzrBHeCdrCAIdjz0fWOnyt5+P06rYvtKVZ8
oKYz2P3TFQNcttPQ+oi3Tqd5E/2UkxwrUA6vQl66K1KhErVR4Iz9ORccwH8OVaWWnuGJQtdI28LT
mxpgo1YeRQtxmOXSuXCqQXzGLr8gdgP1eqlQ6fxdGsdmibgZ9qE7mJF3bMhQLFZlx+aEwoevVZSl
WPMEHpM09nzeTEuFxrhYJ7pF/yBMQ7+itU9N4itNK1jhauW+Fk5X0jlzqzuaZvuvEYaYqh/NiWR/
Sk2BN8jrBmgxpVgcamoS6Tz9+N2X8UXSiLMYlgpS0a3bcunDaPE/90eQDR2BY23nKO5CWgZBTeh5
mGKHCGHb38A0BYQ7wqimdlaT/lrqTmNfOmNXBN1Ndo1V4oC2RW9W3ClFc8NWO25EE5xXETH3kiB/
QdDwmoYRCvZIALHi6Efsdr6QEc/5vQhR2LTSTzzYzCRzQ4Xkbp+1nfvfoIkdGjdFoyDTeWFxI8K8
Yc0n/dh8zNROI3OI7HnoK5tfHFUoniSqEhSpL+nPvKusgQOMSzmIZ3xfhgGyBi03X4JnL23kAucM
3rR703cCrNgZqqNF448QIBqFaMKdzCHG1GQV5mucV5zBNLO0tGbU3SYXuCcQTs9VvasEuEKJJHFh
rPnaq+m/GeHiaqcpmCOUqg4rdOlIh/tSh48BZcwBEMnRTy9C0kEy71dh+lJ5bdtRJvbq5Mh56ynU
a3uTSRwYoAqze60rsMduWD7EUK0zVQ1/rkPgqwl30DK3X7LWk1KQtPJyzSHZlhtUmHgMB8o7Ko9x
cAbYu9B4203pkDal8ujgHhlBKlbpy4aMSx3zF3r/X0gD8l8VcbyRFjN5KSxE+bakdE2urxM+9cjk
ozj4xO3pcUSjnCDgIpmc+G1+7h+VRRpwBtzDGudGxL5g70E6zbXjYZOQfrnMFd9KGm2FMcAwpwx/
gTb1Z66haqv31Xfk1k+yP/4rfpFVUZgH6JW5HkzURfJx6Ukht6/4TGAYQujSEKT62kvD1ZSSnKGe
zw3IB/su1skkgu5HWwF2BJ+KuTqK+1BtP/pSOC1sm2eM3JYQOiUtUJ/G0djkOfdmpGRqf8BNK0bL
cP4NbFkQbz+lUqGEhu2WCh9qQe1pi1XaBSY5Q64HMpadOEMG6mzyyoQvvmj1O8zC2akUDrXr7NqS
zXrYu/rL6HbOTCYrWsS0JK27EA38zAwYYe4je78mDqxcWHWAAaLS9/yXpWYs6Feul+tO/nQoplSl
5fYTX6rnZdwxA+Hk3FHyPl3zUAmCcqm7JsBnzEAqTnnytB0AdGpch2f2BNgP4iB53uZQ18dU8JjU
M46jCZ8UFapCs6hSsQuSt89XamhejAc76DwRcyexconiqWfX7bdEuGp5IzJTZMm8xWUMfjCR0Qcm
3PgDTxL9OXKnAfb88AcsDk4htshVhkQ/SXmrB3tYCBcm3CXhjc/dA7CdrRsV1VkNHedhkjtlhXZv
0vTYLIelBDmtBDmiGy3v+8pBxvcVuIknQ5/LcubhlzOUyd+0hXBjw2H1YJgJ3tyalzGZRbAze2eM
ziHFXCVp7xh+/l+Y5ou6EGGkaTAuCGj4oHaAYz5dnlMkSe7I+WuwL8cFUJEUeuftjGvvPmGVF2Bb
uRYAbsGJjPswE/RO6QGdffAcLE+lszEA31K90XdOV9zo3YK65Gufk361zqMKnfBq7kqP9ZqUr/q8
FckPbITbSRoLv9fCK/2qslj1hU73KzZJMwhNimZ/1iLb2/X5jlKdaK1gOEDIy818tUptn3Y1ZFwu
eeMsIAly2j0uSDbR3I26jAi8x8gkA4IVT15iLPD+7yrpdrTYokqjcQY/vmG5Zc8RakN+EIvgJweN
6hzevGsF3uGg+o8lCVNyoH6oE4AXbSlXooGWKvvGF5P4A7SFeTaurslHE00YRDw/QGA40H+JkNwo
7nnacTSA7Jmhg0oo2uWppx0SktQLxSiAQV5EgnqUT05hZsIQTPNs3YbFRcU/6Q019+0xBVYTVay5
nFSqnpY9ZpWukPmuu0oJe4y99me2PJiDJNzvG5u72nghDWq6UJtwx6RsdInOG5/qgtyVisnWrkV3
i3O7d6qhKsstnWzFNtARdN3gBIdwduuoSZqqZGoWmSgXVVYwDUN6SFNIMeflFoDWSVEjd6FXUJle
j+7FUx0Roq9EyydzjmnPkSfUaGmtoLr6n3LZ8jEb5bN9LV4WeP5T4rPoIbN5r+O9F9dHgCU911Zh
oZBubYnHBZn75BWMOOI2wfNv5CNbYrwdZu9cJku2ZQiCL0FEkV68O+zHonHfiAD1q2jjBmCJxyzS
AiZ3M/+8FtDakBBE8lWPJeiDugvj8MVax4kl/fHuEOvjqXoi4FlFTYb0mtVtSmEQxP9jYZOLc6sX
g9Beqff0rbqy2eXcPaj7BTB1spS0bbjK6zm7Ek0GsmyoyCDH93wutz06EGrmgBM+ZRWFxDhmR7Tp
1DFMeDfxyvqQHlXwM6NQZdwzXlAsvZrA9fXhboEByEN5JoMqtUYT2OGSrB3h+6hAh8jdjafRedA+
yu9uZ11Dj/LqZ4kyl1VcrUY8P/mz5PpmCseKfHhTqUZmlQAkM1IvnR9l64e5PS3EjrZO/srbZ5VE
a4/3SycbdQRyiIhJU/UZWYYV5RvTjkNEhxKkXYwZlkNTqAeqIWxirakliGDIbnLCmSi45EOWLDRO
KOCrizJ3Oq+hmnLKZ2a/kwkcmmUArYoU9qV8xQ3gP1hKjnzThhiJ+M8JOmAZtJwSbdF9Tdzq9ak2
K7S69Al+ztxk9Bx4+WHE3eSRWvasvwB1+k1FxpsHTx8BFJo3wLH4vVRenBRXfsRcB2taw1xoslBO
zzB6pSjBAravMSnUPHYHCPd0DJNySJv2pmzIqiFCEJgj/9X1gOyH6xYUhQJ8Plh0AIAyHbZtINa6
h6RG6xKyEjw2d3JYHx3TEV8IC7QJEZhNKif4ldbXkBxK/rHshZS7OVGJ+kedBYIXeH4bat/GKsvz
o/1jv3uaHEUYhJV2fWE3vw61K9EPcXGlURkqOVrhJ3c96+8j0e16wEe3BLMDf6pcCT9Ibx6QNFrm
Bz2LGOyzzgYjn9mAJk9BxVX5khlEYf4xsI+jPIiG8Ng8y3FB+rz1e6aVbl1F+zIkzumWz//7ThEY
PgTkKIr96JXE/oOTj/UBvQJRuiRWNCaVb70gJiVwnXikMAubo/Bq+yo12F+f5WBsSW1QXG1/zi/K
PlJm1R42DIKJSGM3O4zvsmNQIpDSalqLA6BLbh6Mh6elIn61nAVht+kvmrnYYzKzyHgvi70x//uN
AWzhROddHitwBgQa7ibwSodI9g06q29jAqyxnSCpf9+D5rW42Y9YC3HNxQTypIwCpYN+0GtlJvFR
IjkZsFz9SrdZc9EAxXGppWY5kB1TtvF3KN1QStMwYcFQJP7XG7ITjqxkLPoa0o514Y+yxWoPkdXR
kp8Y+sXxmtAbNF8vIlNRWRI8O+hUyQwNo4C4C9uRXg9QihE0ZgZycMU2/YcckugmjT2ZK7AnfkmX
d+X5JiuR2IOMIXkix15OV2dWoGlJ15PeDAkpto79c2nqivdpUnglFR7egSJ1eUZlWbDDr8uAAx0E
7og4YqRCjUObCt8rI0JTygRd7yis13mPE6jwa6F+Uy5CDWlX1G2MADkVFSPqNhPf15B9iZUkqTRO
ghC8AvsNRoYlulp2ACz5Wml92/eLYEal+92xdQSZhK7u5mASXeDeU5USSHDrrqddq34J/aMd5PUv
xLMlRABZ43ysYqsQC6XROE7rK+DkCG+HHJlsGHcEsMrdzMp3C3nmeCiYOYnVQEUNMfmRUnQjh95f
CJwMF2yPIO8L2+gZzJaeJX3oG77PiwrUEpxIeJuatPzgzYa5NYrz6IUtV5C8FeZ2EKQ1+PcD47o2
EM32vYXylv5UIjNwtMajbJZ9NAhHoBtkh32rSXKgmstDAGGuD3V6HnzRru5nquC1c+b/AX3zESoG
mYBuTvi1gNAwOSfdecBR6gdrCYTFQM23YD78Q+P/js7hXwsxNW3QHI0sMY+o0/IeJM9ulf+V8Grf
6/XBG/DcCLsK72vNXI64S4Fwwxcf+0pBMEo6EVsgyTBGryS4PRZ4ugmDMrvxYYutplSHoKxzfBX7
DhW6U6pjlFFI8VIItIu8Wrqv4C5gvdGW6IONSOsA1TJMRLkxRkhSk8xWreMZjYN3D6LN/cwQTPie
jB8cXXTjxn773At08HwLLUfHvdIvJdfKnftoRKpQfcDVOOlIcPxpQrc1UTFR5yZeTr6H83e2TASR
7ZDZ2fUgjjV2SA51XQOQx5zbg1/TKzHwDvS0Q1phJ938u6y0Qt5yDrz7oTgAIOKFei8dWISJmJy3
jk+R3kAAlFGjohEK6/rh9nYTbRJgP0PZWo+P0+ENQEyX8wzJYAza/gFk3R9wuzp0m7+IaNru+lIg
SsiupgM5zGmp6frRpEETKRlgT0VifvXV6URNfej/yy+4WnDJTC8cYjQX7U+UXpQrYeYgrN4DJazQ
M8QS7hOdegWTHm4jKlPoP18GNButB3X5wBcPas2zey712hpTofIB0ahm9rGLapgmPt+xclJ2k7Qu
bslSjAljVQ/MD3UkqkT4ehBkTfWFoW6WGBNbLlLpUuC+h67oRroodsvUcsaBKonyHKNJrJEGIJg+
CQuqO2P7SaFXejBIWvUmyyoUyYKcWk46x6I/d45vbeWscJi62TvxNzbfPky1eN6Qpc+W2F+5PyAF
z1Bv/6k9xzc4X2oRZ+mfRl/emqCopdU6LXWWL93NHthieXk+Od3bF0jqQy8T4PzwLFYG+zNoryjX
+0GQ7co+ktAsGeC64eIf32IuJ1rn/hKbVNGXiW1L4zS+WGkiZLSnapGVetdMH46tstQEfRKJZ+S8
Ynjp4ayOKLADFWJuUokQbkcFg673quet06PArLzHpSO+zL/cDsHMFxPla6kPj/Ud3WrTsu4RlH0a
KKzHZ28wqqAjTyD9ZKA/e4yXnW4H1ahJsKJbvrhobj6jNIHE2+R1tkbG2vNTnANL9SWrgz8Ks6Ao
2mwH5l0J7gJ0zCP+tCjt1qD5Xrio5YlHp5CSUL3LRv96zG+2b/1f6p6Vnznhy2s6E40jlNcQm9w5
YrmDKGyRst24yhS/fQZ8g35IBxDiZWhwsQ5QL7rPIhSDtU88ZhGBCUQhjl8/zg9O6K4V5zZQ1WXx
cDa2P1cTJ/v6k3R0d3yYFZFdv0wmGpK+iwt5mtFyzlZz7RDfWEc7MGoarB+oZl310HCGYORWB89W
NKDXfDDVvk5Vntf9fzqBkkDL9o6tqm7lITbsijesrXT/dXu2kvMdvJeizIZLu12GuUQ4DiFl+pZ+
mJKmLtAxDgVZIpMSkGPeYKdo8atRuAbVd4yqptXh3p6NxcJplaOm2gzmVg23cSBIOT0PGF3kN4F1
mVIpnZ88w8FMdpjenedL0baznde6oO7QozGCSinIU+jiJ+vaEJJiUlprMG1miSKKr6rHTHiSiKfG
CP0W0vR4eCVIuU/F022QRNjhROcsf9KMpUWu2kQCE1B/rxd3iac8Mied4Z9DxzkeSedBZ7nd4is1
a5elCkN9OTIo8X7hPSJL2d3dsJ6EhptLhdE6Dtao/z0tuQFZ9xMgSH8gEyX0eXaKDjWY0rfxNf4D
4NbKSA/qEUVDlFnszCGQG7kGy3g0j0aLWh++N3Tz7INHPLmqmj8GaCwgl+CBTFUtJFWDnTKd97CD
asU8pbMb1r84NA1MIXxw99E0ZG9rcjCEg/tBonJd2Vo1G1i6+J7NixR7zfOQK74lG2wkldfBe2NZ
Jb/e7VPcxvPCVJOm9fDmccIi1noBEdUAoiuB/IbL5WZpdmmlwYqkCgP0f7W7hPAoYpVMdUDHhT5L
HFoiYlz/dEhfCi9u2e1+Djv0thszrtHrgyoLatK7z/0UBegadAJ5azY1YVR721CpnUm8nCUY6Bp9
hM5YRxUf8fJqef5pdqkH0y2tW5J24QCQcVUoS+rssVMJkRGoPiygfbsnhquMZRBg7cntmMnpyKZx
ECkvTKJES7fMudD85WnyXvubW/WDIryXTrfxKW+C+f59OJZfg3V1Tkk7CL4uJejQYbGnCs99K53O
qhUEB+YLkfrlbGV0wQTlNrW7txJTWWYYs733JeTDTNnlfR0lXLWod4KTGOaD8K7vQy3aPWB4IusH
LtX9UI8QlKWfz8TTwl787R8SJmsc+/lbtttwgR78kb7vYAres/bDygPLuZkoSbIETrnzwgQXX8rc
YcrwEem4zluwMQ97KjfzxabpEhG3pH2ACkewh0/G0Sxjg1jxuX0gHQT12bBEH0NxH3MZ7v1p+r3P
utQ9ZH2pA7B2Zd2y/pXN74doYkfDnlaEp1yQx0bCiLCbe4Ge+fdgcU+7aFjc07K7UshOk5SMpDMs
j47IDxquaAayGu6xAaIPIwoi54x9lTzMAr63pSg9UxOwZC9p/cel3JWQQQUn3/4E7yLwWwHKIcZm
88sdhyuT897jPdncHmQ5aNRfVKMJLuWphaHb5dnNq2LKimFr48jGI/A+RmF1oynmXERijKCmrdmj
rJLhMH8pGNBX13i4mNax4KqrEDlXYXzn0A9bLWHwgI+bPadjxFjxA5OgnCUHhNSTDAF/3twTYGgk
1ekHkYs3Ow3oQUgSlr33IxokCVUTXH1oxGfTIW68dlifY5Vcrjzyl8dozPV4Dx5HZUnsJrU5ZY/O
h0UCw0Tdj1fvy+WqRMoXNZQRo5CxD0GcLLBfw5Cia+v5OSmacnSspaZNwbZYcbaDo0MPVUz5vBIW
W6Ky/EDq4Qt/Y5MVLPUeEbhhNGDaNIcilIO/RKGf00HNcL1xE2jofSbtXNq1O4mEVnrT9KC6BbWC
3UYZ/8yGxCQjtobtbKeumQ5yYV3KvqBsRi7xB5yEPFpK1Sv6bIX2taREgrdVUX6GjJbRheZ3Jqcv
N0Ffo2Kv/5DEyfk/Q3TxyhyIqc4JxZXOZsH/P+YIccaH8qlq+9uQD+AqRhsXY0V7OzmCenBvcJ+r
FIO7gM2cavYaP/cPX2v7cGB2+Nv5dOj4K/W+bsHcEtirgjobiAAUVPA8M/jEYrGnitEOIfLcdue0
reK93wHQJzXWQXvwk+Gvobe4shYapD/O+nShP98pFQCzyC4Rzntd17xXXkbc/pCmGdDJOKInkrYh
GNOYxGKBd1zki1EpjJ9K4A26AXLh6ssAOQztgCcFAyucMbcjjFituN9TZLQF4UGNtEkGyBl8dGYw
LoLrpO1GXEZ79Csf+gdi7Dw4LdROJOWTC4MfQNNsRBVPGOYA9eX36DBvbZxGwWjCpq06YyZK5ktj
IXoUiyyWPk0kMe6kvfS25UzQ5qfJhN0M7GgTHvJR7hpFZC4Qj0WnVD0umimUdCsjT0GstClaHguY
aSbr3sHJolcwr4+62m+18MbzNkzN3n871a60a61wCMu0dLxc/wNk7SzN++LmmWNoVvi6Bs6ioepw
HD3UCnDtNdDdeG3DDQCzInhOAHmvVvvfXP3NrimZgtnifgg4un4OJlT5nBa37rs1a/mz0eyZW6Ey
OU3zTj/F44umGdcOxdL236FlYUFi0QpE1O6Ahy+QKnWxNViU/jCLp6qnxUW2WLCIXKpMz+mMIs1F
NSCCQHL0+fRT6ndDxOnqZ3j0BgUPJrmB6uU5rWvncDH+M4sV0faqTtmKsUPR927KM2wz0uolrTb6
Og1GzlBjprxuncAjnY4fl46gP7XcKYfq30xdeWxWHr/FnSEVZy/GDg+QlNLbvhq2bOkDRxJCZU6F
Bv5MieqvHO1/5LRlRox+JifIslIx75EeXVAvnj812zHqRPQTpiXEB++YAbVnanE39QXwKjGLe+GO
x6DN6UPH7TaAN8uV1a0LEvb+g5BK5bS89jQjAaJs1WvAguAvvbHlZp6BkCC8gIrOLyzN5tKfPrPw
AXWiO/wflQDPr7IKvJqcYpyatMcG59ETJMk0FVUrUnLRV9djMvhR7vLzRQpfpV2tpBY+9jti1ZLF
jJe/B2k7gm3nGUAH823SPw2WE8hv9kRL7w/jkeSCi3QXFkc9T59jBX5ymz91rG97LdHRpMAa3pde
ttPty4S0RX8aBgdeFi5jMvRgi1a1Ex/P4wxUisNH9eaozAMNfM2QWWb0acwUe6yczPXn0Nn8CyTr
3/4kW4u/eF9SCXSCfCV9918TR/En61pi0ECTuTypBbpjzTe3i7F/4mBjY3s14B67D1vfExNIuMiK
w20+Lgwh+mNHSMj/fh9mM92uTyUC8F7kkgvPrdmwq98I7xDtGV4tt6o3Bxzk4hOiOSkVuOI2uebL
hxJMO3mJg2bpK5Esm+GOP0Ov/ijcBwXYqzawcmS3tgG0uoYFQOt1ruQxmiPa0toBE/igBQ8SCUFz
bpOTYWEZE1FoHe2EWLkbx/RQ+Ag0oEeK4N+c+4WBlFiDgHcsW3umDnoWzabdyZyUeM/qv8AI2lxA
e1VGgdhqn0eRHf03MGVsl59SxaV0soh9//W+ng/lTDwSyj6JsDcwJlgeEWOymEdr2Zdp6jqHX4Oq
bsjs36Hza90Ard9hDMltEk6wjfo4+4uhnmhMEux5ugIJJEUEJ1G7G97R1FYasKwgl1SAseqdM+sW
BObc1shGFGLUqo9BDa5EX4xD3OrI52f9H8baX0amdhnmFBGAuHgz9Ox20RK9rqaMWzW/qQYQqf1i
d4zcADqfc+qLYlqHMynBjfm/Y9bgb/13BiYVUcW05ZAjF1xxvuuQd6OmysenupGBddyipqJugpxY
UZQpPoNOZ7e+KqY7jcgavQ9grFltmEIMxUG8SEJ29jfq6TwBzMj0InDXyv7HID/ltsvYT+h1eO0f
loxOVjoc8XRNyCYpop1zn4pA+LdapjWRd3QFHvh4nQkDWKhj8KiTRBonRDQRbGkJTm0fRuakQaMi
RXjz5ikfoh58M9S87jgqdvOOOUUsW8GNA0G7V7EfpoWfpy/5Gwrw/Evj325CqTlM2DJlrF/bQotb
lGXd0CjJml5PvU/xJPmEF19BxnxlrM8hmwSkfWOMC1jYWvlR+z3s6l235PlTrSc1OBZWRzPD99qV
XUMmpKx/3YMHNKypju4e6C7z8aq9aw6TSYJb2EGNJenNzzJCzVcmx0a9F7GqLNfyjxAwj0EKgtOL
nvY++sCUyBlbgvkQ5JClVZGPojgL6KDEUAtezkxoPOcY8MN7aI2+oUn6eI2ZdIOBq0MY8H2VmbO1
Tr7ZP7DK0YC317Mfjj8Y3Z5yAXVbyfdWnJyYgi5+6Bepu7hN+sgnSF56EShJ98yczL5A7HedMj9H
MoMDZqTAgRxCDa65pCTiHtiMGHvyxlhrbGr63j9rIREzmHsxzTzU+aOwjWXXK2Y3uSmeY0b8+A+O
B4ND+3dl9FeDlY48Ei4LR2onrUW15LoUqTJASQHlzpCVic7uGB8vo+hVa7Lte4T+LUaaMqymVJN8
yIG3pG+i0Pq9uv39Ywro4oB2+7fLGopd6E78jJ808eEQKxKLvu9SVrscpVazSuZJz/TloDVornR6
qrIpxYcXmIcUZjU2eJVd9fHoY8te6Zr1gQrPvevoZQJ3XP+zzAs3AVw3cNHApyKe6DDn7Tm4WOfH
5zTtfO4sjUj8cxCw1ES1t62RIqcGFPxiWDFg7RCRiUjgm0NKXZYPq2Ktzq4L0HlGwNThVwaA//Iq
49pQ+YjV6qKF0mVa644wSN8EYFCz+HVnYYBH1OEUB6GbBazAerZ/libm9EOewOANfvbEUeUKQyKm
hF2C2kx63VMZPbwJMCsiNUmHfZ29Zc2xIVOg2Ki0OXl2j0WszfED9fSk4RZtT+PhZXZqlWL9Z/Ey
1hQyRpCtYK69QFkIvWNgrCWY9dl0KGipdhFeRuIHfXkvmYSUVPq3h3K1X1lrrno8aPtROoCA5tWd
l+VYVFl2d5ZdYTBoiyzxhYeMfv6itYqakWlG8DSJae21aYeK0imhRE0rmtEGs6Wz/Mc4+sVAsBJE
Z1c1wrWRkNfSIDEZNMzcYkguyKUxzWKnU1sJh6OZnbLCQoVH5rB5FpFE+5N1LFIGGahOeY9rFGUf
WJmtZaVOXLYhQhlOPHrqi7Igs+cYAiBTEDC2HM/kDuX1L9Av1EwJ+UFH1H9d8MPBaNnxUVEnWv2B
YQ/Su8CbCu9j3SryXId9yBux7vT0644Jg7tsmX+5/2ogeLA1wvlqJf22sKOy8E1tSi9raOXqQMp1
bMxpD+WR7eWSgvJINR8r8ALsfCMRQ3vZGdU5Z36tdnDJVonhNqykiGMxWeb7fxSAorIMhVVa8h7B
gS8DSDxB4vooT7Dd//MZOJ8gvY4kqg+zpQETbTbOSvt2hLRmxrP89gb+NvQ7ErbXsRqdWuiPPU9v
0BqdbSni2hAJN+KGgKu2vphuQt4WEJ2vpAFTCI1IMKKY+eP8gRw/2yQ4phIq1mcdTqo8nfJbm4CI
0MDTTt7MCn1Xe+B/W31xoBMG07AV8pYJ8ziqhCRwzadsDL3L3rw4jfPefCJ65VpyPlolRDhWUZoK
B1WONe/9daaeqy/MW5KDrBZpfDoRT/IyDeE31yCD1k0AMS4DivwXBSaW+YljlSXrJLeSEAVP+Nco
IGV/iz9HwQCvw3DcQPx2wlShPq3jPtBFKJXnl3lkjQvSdEtD7gvaIfMawpaEnfuijUR2dnYa4pK7
IGMP3vfrMylErXJQ/ol+iR9I0W93mHvaRi0CAN7UfTzwU79zPoCOEjj0opbLqiu3gcMyOFNMaJ5A
ooqTR/fs4GvN+SkV5IkUpW18ZXOobH9Xs2glJIxNJBY0a++989EoVDamUE27DI1sYo8PiTeOqsPf
U7NJu43m0yTbTK+nQ4ncEXskGtpKpKyO/tzDkQda8r6LnNivd4zh/ANlClF2dMi37X6argVro9+M
+SzFqqRRpoAs+GtKcF+BNvj4YQdNL1WquouuybJoNcDPDXdm0YtdWvcxkZFuuGAOEEHOSKqaYe65
uucOC1+OejPUS60b69OCiHSv2+ARvJrkyZ7Q9lsm5bEjTTin0MF9bykwCdiNS3GNLxjtadSOp6IJ
fEpTiBQaKHgy+M4AIQfLwCtA5si0DKL5Vc1M6krF4AEZHVhFO0UZVETgvdU+Fqv2YOrIlAfj2uf7
GbYwDjunUt4xvbg6dj1iHy2xjsETDEcWAqN8HJtUxu2BTZcxFsgeIRpNCM7cH5dmRC8dwZ6rGdIt
NcWaQGlfGVYr+FirpRKPEKWekFzJEsWArYrmowkVSMvbLOnCTi3zYUPIVIXj125uyzG3YSkom2Jz
qMge10d02+hGPP0AGhp6q80jWJhYCW94l5iDElzGQ9mrbpWxVQqINx7ut/iabg5C0lPL5x1P/PLI
zChohnMeeC2JYGtbxo90HDXHUVaT7iEUDAc8EfiDsh6XmmGambS93fWkKxHPRkBJUnypxC+wGIQy
4KSsRyvDd5Ms3eRrIpqktTEDqO3TV0ikkiahf7/tACMJ2Uir15WWCAfWBhPbqeMxcrtvDkKKzprq
Vph3/0/bf+o5/6ThDIx2/ddMV7VrRodFl+QZrFZ+IZ+55w+z2p/u7iJ4JMjh/P5etgGdmqB16Xzm
LxCCn7Rsuh2FL19wx7Ze0PG5Oh4gU5acEVtIhnylkTWYZdEDTgA5QZgFcw75xhG19XOwLtKBtJVA
LXKEA1+OJM0z10W05FuTd49sLUENi9ZE1oNUQn98t1Fc122Q+zfWgrtTXghvfrKCYglMWqzaik8X
SodN+XqmcSjl/HhFjrBT+pnJvZeUVHfrrR/OjjLjM75Ces1MiD5rbLv6WNwstat6uQQyMENS1aDJ
VDBY5xp+VydKY+CiCbygnKIBOqj4UL2HTI1aNglLYYpRr/9M8xqZM3Frh3v777fLEhHxMs5N4O4P
FlwreuegIMWi3wsVKEuWJegVu+3xA2t8kokw2wrK5Psk/0c4zI8bVKhTeQ+OueU3DOBgzzg/EOuy
IhW+tLb/0RNGC8WnmB9oCT8IHxQE8Y1qyX2wSlal6IonItpveFW4Psl9lceCEx4K97FY8EcIBxSg
mR1SVWOzLyrIF7BhjDqW/fZcovxLyQUrkgeQzh20q8HCeqdKg58CWdTOwCVl8SclgNJQ7dABrKJq
jESx7N2W56qIioK8HXze5ByPFlncoMM458z905hFETikCALwK5Wi/69/d4m6nlkY5HbEuom8KlLS
rG+cKGaEEhay9OXUOmUapQYgDmnFBkta//gYiDpOocC+7CGN8dSPGyQz1sL06hqI7rY5PFvOfDWz
JCjNig9pjW1cZbEHaMyXnSBbvinxdqO61LZ3nY1YqqGG+/O8SeyUbq/jh9o0SNfJ0pAJqbqBi/Q4
djAol7rAB/j0T+Plg+yVHhyhws/tPWDFchPl1PVoMn9oCiqdZeHrv64xnrytPUbVgCydH05mTPxq
P04/wxJkIG3Ma6ZJVada5BlePiBke2sN8bcyAFff0/BUm3Rid7U7a7o0wisKwBtpr+wR92U1wbEc
ocXY6BOWZJZaVRVDT3jwPhijDvmq8a1mOcSx2ZRso/OIhA8q5R+T6izEn0CtTk4BFzHkcV1Dcqb5
qHFH1NcsWOZKMgB7dRFdXx+W7A4OtB+IwIV/pBO1zZZakgcwRu48lWIgTnjmt4+zB8Sc+V1SBans
ySx+AAwhJjRofEBzhEP2vOf5cnrOjjHihzWc27ScRBd83181HT0HTRfnW87tNQYlCTswCBeDOBp2
ie9qwXp9sip1iZ+dBET79H+VK6r7c5DG7jVMkUWV6POLqu82PBkeKp9uYxSuyJIg+IAymFBhsIMX
1lkWL3ktdPt/C8ezlwv/zNU3dz92BYoBdL4UCdM1GkygOLYkvRAgsM1Mg/kSseDeuR6OUclvL7Re
2XYGvCIanW4Mf+jIGexJIEkekUPKt8BmI+TRZki5ghg9KECFEDFr8Sbd4V1m3DUdvPTSya7/o8SJ
GY2wp/Gjg4HU9Lq2NUzL5bHU5adrYN/N3kaYTv6TQQ4JgxF2JPEL3lnch+7JMb1zwO2Nhpbti3i4
f4TPU79K8dc3wrPgU67R0+CYW/89/7s0SsZ71AxK5wXUD+XcGn9SGX0or9Xs6vAwmMwnAvCbKafC
4eZmXdf5g9ILmxGIbl6t+ZnJjlQ0dbHanY6xVBhbBLzPcXZx2ftY0ZNEDjrYf4tIPdVXJpSGqQE5
G5k5/s5VZauUs/XQVXTO+X7yTZKoFx5VoTTVpfDN9fSz+E5ejVABsWSUGeeDsL0sFwLIWMJwWesE
5U76+7ue3JSsAVqfCm+ymxmNhubPZLGf4ngu7r8telMU63ovNblCqLZ6+epr6i3SfPMdEhQlOkMt
bo1oSRjgIYUtL06k1xVly3QnaoeBajllwFjnAWfmaJpqfbPPZIvzsDQDFHXIdwZCL74BV7GoX3iL
pqRlVM6qOHZNf9kj9idIKfB4mosbvsCTyt9Jcjgu56/PxhYW0x4859IJXyIfteTGkDWUJvFf6RAX
p8lMgppbv4Tqb+5VP8Xf0vlYQN2g6dCydL2J478H+gkt2HAuc6jA7Hk4wf2myJoIPk8o/IJEEupq
/vi28XeZI+eGi7PH1eIlZW6JR6OlFkgAdjfIxyMEBYAvWExosHv0ByghlQlnw9AE1QZJYdbzjs6j
SsqmavbsbJIL4V7lWtpg/aH2aeCPi2tzFD8o5TWWRy3b610/6UBvLcc97yQoK9o1Tz9xN00cXceO
pTYiNqjZ4qAkw/7+D3iyodtrDg6PmnTYcIXNZRVbPK1OBcWetqquHOtDIfjFypyLeURvTrRiSUBj
9nuHS1XjlHMdSdFaIyDMGywR3GD2oZuWSF1RTQSMDhwPnw1Kjkkg7YDgWU7C7PBjDyLQ+LkagXI/
IBb780YaTCMTbaMYtd000lJJgyQn/HVn6wUKDPeL+9zxs/TnYdJ+ShrPHfhylByhN59mqDiUoW3p
jlWbLBz8jw+i8naJO4msoQe7zZDNbLeqqyAgQrm6m34EfYTxypISYbsdR0roDrWZcF3fq3TLSoh0
dY68KWs0PGvL6JizctOA0VgrXKolVqlwG0pDRBamJLdfcdNXWpCb9rYp2SWA9rEnNZ2osogkRqt2
fcbmEFpb90cCrqtuKLmC2sP4sQh4u97yG5LluSiR561gLDhDh1xDYNr5f4wdjDrdDEK5AlNKLQfh
aOGIw77ObbgPVM1Z07oHV02/BJyZpi3Hca7/1a+IDCEv6xkqa68LeJT7pI58YsUtmkTofgUf339B
hF5UrwHZue8HqP7rmmgtXl8iNIxI2k2xU3MRjEEloLj2/yW9vDhAgfny8gIW7yEk41McIXScAQE+
6VYBUpUXJOT1OGVZgm9oA7/L6b1mUlc8iP2/ZYaNEq9retLXMnLy8jTAhGYV6STUOJKLL5iB5nzA
2nOzXxNa/XvCaV2vOFM55pQ9H70fenOWUL6E8gxt77QCQ3aujtOZHEDB5qS4wcf976Rq9P0GbCb1
SIKo08aqFj4XSy6Lz1wGLRBWDR8X0ZUIJEGOAS2xHhjQoD0C2/BWHHFAgP7jTaXXPEWhfeyFIdMU
b8SxRRaGwRVLu0vFn5AgBnWBY0AJRe+YzYQuNeZNp+vJ8J1CUPEiWvDqOK+37zcpBTII8TkGDcCX
8C1eBWvWQHLy31RpqkkAIBa2Y9szJU//VThAynk+IlNKZds3W5AynNq08q15hiyqVJayFh+3YyMi
QR1aBbc8rNTrv/GhsNR9c1VUsyWD8bt1O9+E8IF1tLfR+rN/mu/m73Uxcy2eFfPWjdWpz+wMB/H9
ieTJkAzgZ50CzRYWIiFo5EeGAs7oORoQbCSR5uqhjeu2ZrKQIT4L60HHC6eL2Al5yk94VsDxbp8V
T3LMg46Oc9K6Do5nZt1+w6ccEca99s9cEmf4+9DrztImzuERheLzSAN1TE8ySmjcWzQSrB/d4Szk
gOhDHj9OnED0c5clwEdgPO4M+L4YS59P8JSGeVGcn0K6QikkyegArviVyRRPI+ZiFRfkDPIsxfWl
/Mk40JKMRPtVPt38cmN65xa0dtxhmV277+eaeRN4rKjr+Fc9c84bcXKpcdp2tV44lVpHMOp1sB15
HrqjR93z4Fk4iYw+B2MxhaIcHGdLC1yEnhRWUGDiOjn3PWdCY0LCi8t6YK+v19GTWgLO9HJYMyVS
hgq2XKvvNLPjWJkq9IGJMRuoyOpUBfY0QH6rsc02xuJYLiCd26RGzAndqmylYqJVA21yE/XJyAJa
FdhFPC0aC8SIUqoJCoAt+K0UGbHuscE78ceXpOmXFQ0tjTv2KftK5BUEL0u46j704pqGe0YS/xfx
VQ5+zKYvZfnvEma5DfbOPJtgVYczDoQ8dQZbdXFNBfxE8qxMQnDm3tYO1O9OsRA5B0Jjxs0Xn0n4
38+kmF+t0DsYXQOE8KqVkgGzD4kpjtUKc8Ed70hpdfsNyMHKQpQ9IDgCe3MAL+0srEI6F/oHygJV
jvfi5fZLRdBCLGAAYFYK5OlrUUXamphEAZORxxhK7gP6Rl8n3jeZtYm6jKzxwnEw5xoMCkICzjC2
h9uKzm78y5Fslt8ErOLibCQXSLnf5vuy3Fyc/NldO1VX/HCnVsD8c1hcuNSFYXF+1PCIQ+KRSy6c
JzH4KZvTElMx0wDLJqnC6tTgOCgFHS5xeO+Y3FURaDE52aG+KGCvrBcyVNrNWKHDAIxwXXkgBgiR
0ASN+sX2RFHpNsA2ak3ygZg5EJH9E9/FQE/u1UqMGuMbjFb6sjY37WMPMUw+q1Ro65di4DWFrTAR
n1CtA03UEMP8VsWyBq/GZmezQyLFhSJjoUmVoeaq4ef9RA/phqgCV+yCE8q8wf4fDqSw8F1KTnLm
9x0x/ktYu8zXxfw7Dt4a6Auv+ZmUEVQ9wVPhgqA52t+m226AIEDTdmi1huX+ksEC3ImoEQKt/Go8
F8vuxqFME8jegqic90Zh/9+HvZXSplzdfOarAnyXfqupKkfu+NFUUIhYssBc3N/qgKLyAmf66zC4
ZCbZm7n2MXpwImuWoKMTefF9I/dwD/YiPQcKAEkGgXICwdxsC5qX68aa7KuTOEEfpYpXW0Rcb44h
TNYUACjnIEzcc+fE9ARkAGdZSSuSvxNNZXte7TukczYQrHZ2u9Q66xXz7a+JPc4dqjyFS8Dixcvs
SelmMfpDEod7PJgBwbn1HLxYiCgMOCCeTNKfkteMC84wrOuC+Q8cqIqx6RCLCv8NTcf4UfkSDkT1
IGrnGprIVohLc+2ac7tzS6WOXA7YmYFRsPNNvlQMj6l0BBVSqZd5mjw1YaqSzKF4N+sJF6v8W/ZQ
wiC7QNBPvNDanCqq7VTudQYLnP8mI7Kgn7Bd8K0R0dFbBaAbE3KCjJgzkndn3mIG6PENnWjxq/dw
/6ryzLZ8QFb8n94vZLq4d3CREJasIDVqD9QjFEoUZpFHwJiIIysCmhGLeR9V1cvVP+ft4DIblw4C
Oxmz78Y5kN8DVb3P1ekOQNwLPY54PgGD/NJFC8xsoKaR8CeTy95zO/BwxdJJTCkG2Dzt/2a1GvKD
+EzRh1JWn0qrefPCFQHpbiZ1kXaacUy0rKIGsECiBRzYLBKl6qp91+kAkykC8Y9zIfD/3L2HSKHl
aFhIBZU4UDXQki2OZM7WjIJ3ZKcuV7sT6javkByH5t8xX/cXrEiJhKSmvcrPjqq0fIvHbpyo4foI
BwMvd/cTdrV/PfkgHQOjP5yzZRQc+7+aSJr2hT4vL+MoZu742WkTgEuQ5e2ui2YM13ZQa2xHpZ1V
TdDv3WwSolEO66xBhj70OOPUv5i+LuFHcE1Vo6BbLPsqtd6VH17KYOm6aIm6pvPrG6EOAiEPknk/
RidY2xHA6pMXJNSzasLit/v+fNnvdO3UBRxXziaDPesEVnwcwsU/F0gqvUAIzil5zkbtPpgRn3lV
yvfbx3RKFJA4t11wQqbqt+sWVFJ6yC/Oc2RWlxIFIJVzY+0iM5jwjk92/YjBtUXG1a0JvRsHMf1j
3vH/6cqWjAcSvNktpMZxDV2r6rylfFqAkIdId+BMNuDWD8eG4cNX2DORX1QIWJ0tpKI34utniuH3
D5oe8O6fBXpfLULZARlYkjjMWZPFPcqhy1W27fq7FGvxhJmeK4G1JnCol31Sx+fwNkkJorGy4LAE
uGTFB61x46x1WaEgd2tFr6dyo/f2btK0cVHDWgvAANaMr+Pgg33jz53ts2ki8h7czpCjuRTSYJoQ
9bdXHp+zo1IWsDgBOF6GtryPVjZtZAQg8Otg4uuQFDp49yuLE4d5ORdd162295AyS6F/zLc7Y6vl
kJOOOVXudwgNjiSVzI4btN6PE6lVzh7f5+cqpMH9cshgOhmYI54Q9MIeZz5swB/AopAis+Caf/2v
QKCe4hQ5gBapnpu2OoEFxhEntUzX1fsvq+1uwPnRqIioYI247milPRQSA0EpgpCfSNLceu6qlxH4
EgVsQkX9kk20b1aFlyN5tugzbZpVog0ZotV1pbSo12zw59OLTU63GGSfcFznckfw/KhSRwxw+u4W
vpMcRTDf71PI1p38KrRF/AFaqSHOIvWvs+Kx293sZ6KICXEfeqwLpDtGhOmEyD6bVmFQAWqm3GYS
uyrcYZbuxXbBmGP30inP+zNJ7oEb2e84s/28hU4OiwQFdcq/bk0YMnBnyiMRnF9naSTeSY7sLC7w
YAXAap96MM8ZNV7PdGQobeIu6mzGjUbD1aoeO23fDdPastN/GGapNAE0IcJTt4UGhzADYvyAhyjG
vbMojWHPblLC0d2ONQFeyOh3Vs/iDjzZppDkTPFmF4Lrb3YvjCualK5Iwa88BrLY5Q4Vkfp6FjG9
uWyBFdszDmBE6ysk/p/rRbNfnCRmN4ff5y6ZtgQj6Fr94ifawWohdze8U0fDcn9eaarvXZorqK7S
sKCh5D91BPNm+vETjgirggLG4b64ZWstbntHVOFx/nJEDtj/WakJrdCKUwpqAFBAXhNvBSxYAwY0
u6t7W9ZpMZcthVGlpMVYShVHr8BeuDljoAZvM3JEkB74Hc1KSnymK+SbWLbmVIIXm16DkJY9z5fX
/Lbf3yEPrkOqOYbmAlHnOgR05v9hu73KE+wLs75BDpwGj+l1u6wyxicY5hI5Kg2a+6Hmti5e7Uh7
XQ17syyNMH8DY8NpKF5xWUdeAIQjhQVDISWcL+HFFfi9ylnsmEcHqi4tFbirT1v/804b1Tc0xP8K
snWv/O0HOX3Qh+RS9j1MxXG16/mU/v8GZ9C27+Xz279SiOOaRg2LOHg1Uyxhb+BvVx/6nC59o59t
5337jOia0XmMajwFzKT39hmzFn5R6yiMoe0MmZiFsRlnjLb80W9IqfVLEfFqwmJ+TtCxZsAB8RDJ
qCOdT2oJbRkW4jGAObuEObcRKgQZnwj7shMX4dSls2AioZKYy0PkVKJOe8F9JNeabnPzjqwvlQwH
h4tDZfkCTe4WoIhkf+goxydeMCjGDelnG/St41xy/4wz6IPbTjYN8jWaaRXwZm+1LiuStCh6qeEA
Q03jRqMDZerfQSXkWALQGPAg5NeTENDmoZOpWt0L9yOFOz39ebwZIL+omJRDXJ0EcR41tLFmGK44
h1ZOgnKjWFNQ93f62UWFAYMXuckfq0wHxfknPX8fq8PS7rnkZus4j95j4vXWlhgxMroYzVfBMy1H
GSVIbbbpYvbxf+q12D6NTQUuBFMl5tY1TPneW9Zdi5g9xqY3sJMuGKsENA+hdS5KkrUTV3tSLxIy
o8nVWsevnX9esheDmkg6vcl1FBxg84eUXyoz6uR0zmamXjUwvkkYLsMGH2V9I8rfUiGdYj6guJT5
T91QUnyG6/a7YgG7KJYBQgIw6aTQrKHG3yj6B19qGNeUPYCezMLKkD2I3R0zKkIt10f0Q1JcqUs9
sYid02HJC8/Hjksma1KyfJfgk1J2Tlj/v++MjPVAvqpyf+fyeYpxNxz1flHBq3naq30ZiaA9Bbof
K9wTBfyzfcGXR4Pkhqq+OO1q1wW3ct6gM8LYb7S3ZiFnv88vprLmDtmggZ9ZQUfUBN5kuor4/iMw
8rCAdfLmMccjt2dyMiwFsXB+CY6tTB4L9lz3HvK906Z3hUAnTcsyRVPHD7dPE8Um79Btp6bvrKmV
zO3j3Gw7TRXRVW3bq0XmNOHWefpxs06OpNvTowGr8j1lWdlA7B0FBWeD++pIjPlLEeYnQVt3I/8g
xOqU3mHDXwLSuu0sQdAtqlnRvq6c5sCmL40tPH39M3MATQ9C8xtzUgb4EOkEKc1iGndfPRX5Ck2/
lWuk8PwxkJkgEuxB5c2zN30VrO6LLROqU3/TPYZLOBVdcRLMj0zupGvCGNhgkap2LEKx/uSVlLB3
TypJv0xZ+fTJlmprVpcHUrw6+dWN3qBfSMWuk4pe42WO3TcxhKJdoAaslnYGuZDk1iXkKVnb65xR
Pavxq6cUwsTr6YlqS98DRlpFH0XXCzbSxK0ou2wsTA3Raq0+pky3gOSiwLwCARVOjMIWVPqat94x
FWQWvCKVi5+DzEkVChq79JVAtvQ3b/J9aj1z/Lkcaz/UFaQpz1yytIpW4dPoiua8QAnkHAJBVdHd
utmFN4ijxW1gxCdB2ewKjzCiikhDN4k2TA6P76oAsz8MOR5FtXg7A3PIp2FKC4V/URibbTfBvXo4
fnKzLzdEWeKVNMEO6NSPlEp+N8mgfTE5H0NNhxMRhHivN4FKRlWsYwVxOxFEE5DBpP+wq8j68WMy
ufy7wgakkTg0o8mduOIezc7YLE9jzAoZJrd+4hZcwRXKI1Ts0M9Vu7TFYvGkGq9/fOiNGJ25mKx3
gEjh+31k8qTioT3EtbNKmQssS0ew9qJojSRdNw5aRN7TAzxA1tn2Xr3A382WNc+83GOXRlB7tk8c
IRrvRjO8f2EOGpBzrFY+QSXyp/Jgmsc18Y2qsmun5+jUr6i7e9UhI1AJTX1PMshJFFsgZ7pHEEZe
SooHDsmVunHJoEGc9S8DMGupzFe77NGMTt6Df/tFsMRPn4xzLWrXF9ssROlngPRqGNZljmrRhR5R
n4a/k9vxPGPr8H+m2w8n/H9WGLAbqiCFdlfuhXCk6RFHDFsZH+ngw24W1m5XHJm4WkoCn3YW6PJj
YZcbDJtrc5RzVnq/7JDlUW6mKIppDh2lEoNSae/yG4b/Er7FJg3955BeAmuOA8mOyt5z6ZT/RnyZ
pGOzpdZ3wwbaVI0toDCc9JxA423LuTusq+w5VMDEQ4qlLqRmVwUKT3RYAUOIm5mwtvN2EwCexQpl
ZZUbN1311tZIGkW7XVKJiVSowp/+uLUlMlFuA0hiwj6ehmibI6ZGYmsH9SL87O4hPbLFfZMBaCYC
zK2WZHKGFt6Xucv//YaN4C9TQADVQq4KdKmsLV6aHjfyxA4inVXlLWSJ40BFuAYKr8SyMfYoeVx4
ndEgZNpuKiEpddZknN8deaUP+pSBCbRBmG/5i0dVtFMpZC4pWx4uVHuOF7imAq1zkVhPdmcTxEwx
ZWgJEx/eUfUv3HuxZABqD8+cAqOFsbZRydjorQqhe4KdxMiBZoPbBHYF2C1RpqTJ07Fx+h7xWVcQ
uBTp7mrhwnQBVeWinrNJo+5AHDTdfUqcRo7JSRtHLTiWHLfgXprD/dfao6gOJB1cZJTpp/Fridg2
oregsfMxhHW2Chnx+OBk/5fP3ZNzhHDHtgyFJ1sxDI/BKqnblb8/18AhimbGuIhZXnDqW/cfafyz
JMKrEZdAS8lbrP+km1Fob6dHVVDmeSIym2jLpQ+wcanrgltGPhiJsM/hyZMatHEK7PV/ZV8vDLX/
rCD0ziYNitoju+7UYapKy9dM0jSZP5eL2z5RexL6mbkSNc9TvL6LSWI8N+xd66XwHjRgvtjCM2kz
rOmB2F6gSAM/HDWhI/RMSXLKQev5ro9dcRGoGtmXag7kzXBVwCz7TccOE+TrZDg7kakyq0foxYot
tyqPcIP3KlbYUg2hCWkkDQz0sdT7oFCHN+SO3JwteR6TyTSnFuRbRsIbdDem2j+iEl7GUQJ/kEzV
eOqRTPA0ddk2L0GwOmbzhQbi1N46HFbcbOHW59dUa1m4XBlj6hZZNlQ6LcJCjoXyzk1JEq7bkURR
tAspaG3r26CYgXA6bTRT9xJz9ID0ILS++i1Er8C4Cy9gSGVmlKfokIkgDkdTuwz0B/LtuSP0tiCu
ZcWcX1czSVaIETWvfZUzSN8S0GcDjbIw7SdGeBrVhk6F7w2whEo+zLbHiAh6jFsTqV297n4KxxHL
tbzjyQ29Ar4PAcNs0o/jZ++Fz0l4LGl/uFE/TGCX8nt2ghgy0pijgeBdXl9CIUzGPbK1HMaCrq5T
jhpUTFjW++YmDm4FcvPAIUdQVnPksNg6HFcGSFRYcTNmrpjkeE+BzvrpEt8v+cYYpITZLDaJLdBW
CmzJj9rzHU7sIvZs6KTM1xe35Twtnz2/8L4OCxV40RvWwuTsUY+Zlmwb8OMhUmKPyfZBL5g7mVLS
Ww4yCKH0XFKDNT60kYPSNV/cLMas6TQdEKHK7Ec1oi8gfur1kAhIgHqib2afZaO8XWXs+JfOSrO7
5sk1bW/Xc05+/moWgvjgmERL8xsH6owNLtCDjdTDcb0QD0iFNCrMc9740Y7iqkzz2FCNaARSAlGd
jWRgejN2WBvC1uv5xRvvQHWeddeRm5NTdmCiu35k1RYnKxASePuxcnmAi6nyNl1wIMt2VRtZtjE4
rAV5o0aShv3Cuo/eLsyR1GATu6kSrjXPWsS7e+HS7LBXkuP9V9skHxH0mGGSFkYj9LSvE+Rygon7
pjWpUFtPp4hoSU0UkrumMRLBfEOMlj4gkR1CrYUa0mM598oKC2+WpaVy7uG+5iVY0rigg0JtRtL2
GaVyKrvplmn454ijyC11iN2Xbzz5BYfAzgWlrELJeG374z6xgZOglLmumdQCmR9IHkF9gytXftcE
t9llF7oZ50dcrkMEh64dtECBQKuo4TDdZin1YZutLRwKyoawLploMiz7kT0g9gsfC1tr2VMrk/TJ
E+AKTTN9f8erq4/WZpZag3tiIwbsYhBhCCRxu/zWkhF6JUJR73JX/u0cTQPV6MNMChfG6vzJogl4
bXSHMThfooRc444V64EGyfDI67XTC9VXNcVd69wjtyy7xfZbNKpjFIvTVlg98cZd/cs2Wro9flDA
9gx61FxCVM4m0ptZGQPuCB9Cn8+o+R+EVUJa2Lad2xSzWTV+SMC4JtTXiAbrYImFw7oGCV7xQ0OO
KPYJT8HFyeIF3KUfwkQ1Rpo4+UJspvvVp0kmyzZXckmYuc+rcUjUizhJ/vGWbtV2cTsnELGOqMos
KputUjIRdaBcS2hPHFz7EteCFqe9NwzYM73eU66hhU6ju7oC7ydB2iiCMV/HuDwbba/8AMueqbTU
UKm5i9QWcK4fpOPfELvivsd9t0kI0lbHBbMFTqgtum9DYZgypPI1MOHfGbTN5M/fj5ELIiHJvQkP
eefYBQzgF1OXEar/ePH8kTSPSwwLYjjZBd1BJTYBrzdD3zrH3ZI1Ju9Rj/zZ3PVp4PPsK95KSBMf
BXd/Jn234tbgN/BbGEvFboT1l3jbFTDPuso/3cx8dzckaE6qAVB5pMMU73sY/4fAY4YHDvKePOsA
hqQ2I8eVfCHZzZqFhCv398P47bVPiWOEosqobbPaJ6fwTWObi/c1QqLflNHkHZVmyEe9DNYI//OR
t5LN6yzYTOzvtvsay+R//zsxZievmbLMOpyOuyKUSF4/jxypYRQ464+eddw51wA6jcHKexFw1zvm
+T4evfu7K1ZxXfOcXgclvsiEmTJS7vds4VZVEejnGsxohv+I/xrVkeX1p39CYHKXiHP1i4hc4akU
k/+5G9AbyGXqWhUwHQp4HncU0kniERZwS59KrltwAF+osJxRdWCc8Y4tVCoSz2Wm+AjToe8fvHvj
kB8zRkoHIHoF2IPwKFRd6CGmbgPW/hYIvXhdvbMVVYHLHo5QMVS4asZNxOM661cEARcg0yEs0Ya4
dC10d+pWw718qIpWPN4yNPhLSeUzFdmv+WKtHLV1i1kBJrwbusdtfbTNil5QlzpdgEoUm4j2Geb0
L1jG0kn41VaUWaA80dDTjksX6ZiGrP6vsTX+vpZRB7UU3kwFAO7ghmvYucmbnK8SC3DnRDx5haAe
lJ3cIiLiRbgOSuWRJ82QSffcAfXlmFvczYCt/9DwQZCaAKp2o2MUiqbI52zXCnKRuY52hxObr4l3
6HWEPRrf6T4By8uNaWljdY131kedWtOdvE1Pq0SN+33VdFIvOXWyxdAeRu9MbTxebj+k6DWGYFjF
L2B9djAU+9ypZSbHCjhkORpykJOEOImHF/hd3Kd+4Cagi62Zh41n3ZEqyyI2sYKuqXjJ9o9isKZs
1DbJBuqhojoZO8AEWZq21tjOAC981xS+hAME62bxfXxcR916N63mxvlCpWq1xJNUiy/aVB2GeyoY
tybwzHTdmqMwDDwU2/nex+MKmA71J/+WKzhbkyMswMSc4XN2BwXA6jGQccE/a3K3h8o/xq8LoZYD
8tKiiEEbzIciInXiGpBfREphaSjyZYk/Dp034HTyxJJfjvE0U82M9SuRT6bKQ38iCvdLfMFS2NlF
EqAH3YC/zW2l+mmgvKtf+WI9WvI8odFPTtAH/sbqBppDoYAVkoa+EQyJqndT2+dvsum/aIU03PdK
4g0CS9Of7Ya4+4Gzbw4MMcoqlY7GtqbT62sxgchHAvh5M7l/wjbbVOm1YKx9wzFFZP0y3xMfDqIN
hmDk2VajcpK2fLFsLD6MV+Knh0NtbV/PJxSwpl7BtzHGhX76qqz/vzBwbUf5ODTcaMGV27htyqIx
x0Bytu3SanZ/eonl4471v5gZwDmyBsWxjF3xjRgJNDC/8RLjfQfsb3oE/M00keha0uBs0YSTKq/e
lsPnnGEVI9+Qt3gWV3OaYXza81fLObmj/fLehaxvmhTK+VRZfskAvNsrdU2MsufNq8FnWWCFB+fn
94jm6lZbQICHsSYPJCXckAnE3LH7Lqv6saNYUBz6hg0ALgez7MJQh2nm7pOpe6lsZtPtoIoNKUQF
C9wBIHFQtAfa+mJQJtlxQxu8bqnen7oYrSnsriGvL4zsMnSnuv3m8QKF932TMT5gbAu7TGAM82yU
wwyXXg4amHCJ4Y8jn8ila0A0dWdTlySswhIb4wNVOYdFjMrZNTCS2d7qlOlrrM7Hy8aJxNCns7v9
+OkcGcmajv45K/EypuE57pzaoBTMHr+MrHab3QLlPBT086iBJZ2mlQHBSl/KGm6BcuggcczT9yPa
md3MifNoKU9/iTmaxx/L2pbnvMCBaZGNcjKHbmqnyra8w1eI0tr1ivfFA0ckzlAY+AlDaKOKB27Z
AyiyW8uFYaZkInAEHkRyzCsfaXg/TGhABknwDqYDSqaT7lVaGqwfngH5M4vt7nYEaGUDtm2NAICe
F8vTtqra1qUMXeyzH11fYYQa1E+GdXO1TcDy+03D2jZsKxiCNGLBJuiNYP8hpec51T2HgGjrkF7a
RAmXEBxvIp7KPN3z4TKQD91rOeN4Ju3OzuJS1lJS1DSafrfyUagxIiRwHdhQi2Xl4iFyN6vTMoUC
h2T+mXLLYlL4KEnWPBjg9gVVdi7NfN3j98aKvv1iQ9q2NGvjOJqTACmmgmjXrorJGirdbsinKF7y
4i1KObA5DBZGTgb114/ij3kvQTLn4MO6GLFzKIu+3NI3DAO66jfV+s1+t2KAe/P6SpHv8nqXVAtr
k53OOnY7XZDrFZPu+De/49PWPGpM1q1yCfA5878cBJpLicaa0kh9WwasFirXcDH9QOVdrGxMZxiD
eLzhjn9kwvNDwkOxOzD4PrUHJdlb4hng5yzNtlRMLHWfZn8ppr5ETrSGCixVQGiVp2WaG7Rycuur
0+Jl7pHz/KmQZmDJ5k7r0BtMTc63i54YYMap2k31X8005hf+OXKXBsBbnQizyqWhMVRLs2YVtPep
W/BCxlrvMXdxE3GBOrNOFnked5mlzIBu8NzivvEiolFMNzrlfrV09EBRoNGiQTFjgaPLS2QjAUGy
YJRtKgw3AaOND98tp//wA6ZmEcf3mSpFgD5VuDLTLfpFJUuIPds7GZBNc147AuXxIDblicVpOpBv
rgbnZwMbv+sN7zkvw3r8DykhBiC8lGqq/Im2hGRarzJYPepIve7m8bYuc0ihgAdVTG76f088ekMy
RB0jBRnRZWpOIY4i0s3q83RWPNGkjT8YFKBpAocZchMoifpZV051dYz4aKhrwNRVCcbv7HXkmOxT
ggx22CJ2vgmV609mpkusjs4XB+XeT/vED5l3bjHGIeWRIKLfEbAylYz2JDOFlbFB7g6nlbsZvBCw
woS89XtOFe1Y4rBeWG9MUVh7A1hl9g5xTclB2smZoFxQydi05lnf5sTqkG7p4J/Ka14wModfRxad
CRVhK0uIM4z01loBd7wY7h5d8wnjUlXZ1adVgJPIvmvk9BUFSsvX2p2462PwhhXeloFzyvt+/xxa
LJtcJJeOFk6UeMwANAeGc3dJn76qB42RUFeg+NaIrYp7BE1d+yNocSXCz57+vp003wm9FYtpQmbF
1BXooCwVVSrjW2Ns9lpSv53otNH6eRXobMlt2cjtSd9PijjtPc8nUB0KE8qUfKou965e3v82p6VE
6SKJHSYj1wQw5KAHIkKTC4q+E7YW43HpBiYEju9VzDo7hyqBC95wJRjJlWHAzoQtC3S4Ccn0pbF5
mCNQMkrw+60UN0RKiQd/jRcXMm7hEIpJcXkYRsj3ocQHnSVtgLFJm7UFLpfEfGSY7cFxoppmt38t
go4obh4CtCiSY4coG0erPavYqRTBkxmIllOGOiqZoMeRPXJoEPtTfoMSOZFe+9OVCKV2McuhkhFK
kDeINeGmhDh/PXaBrF8iIVmdnh4jxErnJWJptq4vGsURDElA7YvMp/FkmC+ci44bpb6W32UQc8hS
EAma3w4auLmLBB5XIWc7UGQwAubNWr3LpnUk1PJ3qEzha8H6n0N9iqC2rKwG3hIkBpvBqw+7gvrG
DkDZ82BFgnvw/nUxbYJAyEQbZLmz0NVHOZgR/rUMkRNo0Ox4tJ9UFaeoWUZ+1aew250ub/NEgHZA
ChftptyedZLK4Ec3+pzg923PTdqEGPI8/B3AnRd2PDYjn0Z0PzLPEGEwtlqvdGodm1D3/9rJaeD6
8WzMcXq+uSrjOmyNCjq9I2UE1qL48n6CZARPZhToyVcY/wt3U6sMWFNrUYO+VazvCHd2o8aHqphN
Ro6F5BfWy+6Ab55PT1NgeO5TegxaKODgd1yWoi4XSfuc3cTc7obavGap1IvHOKDRdX90+d1a7bgP
fPrgzNvPKV8KFogfOOJSM1etK9U+afWqxKNT05xDlrx5KK8J9B19fVswO3AIl3yr74TcvxJ7VUyh
kBUUnY0TSP9OGb8Es1SWjuseUjUwG2gB9cPbPBLHGy9o553IZJ8C6z940xX0a/MpXT9q3E9Bq8zR
56VhPE0rCONHwSKJryxjWv5wPcf4olcxzq6tFF/0yEgo5S43JfJv2uzj86f+e2UHBSBrbkhUPKOO
h7D0WJfsD8YNWZ0mvMn3utkz+qvzsIE7CzKQed/w3khUcwoLuQhChq4XyRREBhdxpqnEPQiIeVsz
Qen/l9Qm8zh5DZqBMzeaWq7A/8KF5lkMi44x1GcsM88qZZgCoEdRVyOx8hcHg4lnylZYwcyTP814
GfzwZgXIEff4j9nPhqli3CxvTvAk5BZeI1gAnRyNWTFgHp8ppu/YiGtMKOG6wBOixRXrlkZxKZpI
SndOTWQ6sYrWBFr1A+OfGRIo4Egdt2DTafnT2I/T3VlZVhg5Ld/r9OY46erfdDRLu0ct+31w/5Xq
64JShFd7LHFXJxsqQVtZ87MvePg90lWLBGxrko8SACg1/H19fmuKRFbD3tmOOY47VPLoxn5ofkmy
mjejuTnXHkYO808KdsL9/4tK2LN8WUSGFd1Zv1JzUoL5hMguDmw85B+xtdd8Dh7b3EQFUh0w6No9
IdnOZ/4WuZBYSfrxldYYxKsKAN8LJWZLcv8hCspFy7kn642nrV2jwVHgybeK0W+7YMXMf6wkZ4Rl
u44qyjrfRBTAFKF//XPKfqvIPhj+bHsqhKTVuOrLQqW9oaL4XQoYq7RET+cxIvFX0g6ls9oXQnR0
seUTO097oh0ASycdvWKaBVdcnfI4cN/nwdyoGbxA8+nF9AJp34mtN//30kh3IZZuKZtGIJlFj6KB
b6udJbwZg16POB/Qxc8n/Ms4vjxkwRQkKkJ5Vj9hcuNE+mvSCnVq6vzuBNPfdUVUAvl7L0omQr1O
xDtMmJAdBiDhoz6X6wFdQXJ4HlQcvBWTq5pv6pfkkcPyir6HRaG/6TWQoooUFRy7XsP/jJ2IqqQt
W14nlu247fIBeQf7Bx/ZQKv8sVfoHcdGTHeKZk5fuK8LsLDEnDBcN25AFpcPMuHzSxKis30gYpjY
6ob5sREaIrAKNqukI76EkdXfUL7HBjuFvtBZu2ePu4BX9T9uisfNqsf3ISWsg2CWqzDXJG3sSXon
QhA2x1AqbaPXZouXJUU96AiO6ILUI2aaAhHjPhK/sDhbqpqOtj0kTtHJi+PX9U1X8bVnmPRjYv99
r6IKm9Obvj3c6VE2NdPLCNUEfpppPS/5huryPHN9gjfNrZUPfH/caTsqNUVC8t5vMa2PQY8UZksv
eh6YK1Il4FhbtjANdmFC2X3lNg5ZdLcs5Bu9HGbMJu+j9/Zp4MLOXi8aD+vnSIOa6DFw69OU4dYn
ZvRSF9zA6ruUayCx5Suj2yQHKOyw9lLDvKkAzKIqkMbik58Uj43NY+5ViJJg4U0YL+wEAnuX+ROH
zg4n7xbemUPk7yDdCRW7GXW6g3fm+Jh8LNUTJiEflDdgYvIHa4MyTffhS1UuVy3WxJuHG6liaWcz
JX/EPZPkt3748bd7vZdHTy8fivEp2vmd/kCyXKe2IlXiY+3eji07cpYxhB/GLAr+yRt7yvQpQX3J
tx0A4AS7tIP0W+9+dJswUnpqloVsq1VeH93Qwko6bF7Wa15rwudokfcpnor62ct4biiCuoKJ1aiP
LpiU5UZAE2mvdBVDfj8+DhH1+IXIqX0R08ITzvDEPs64YLkYGXORBUlyhqcYLA1oCm0YEseElC++
12or5tsbdID888BGAsPw8Xw6NVGxP4MVqiL3Umw+b8QJU0k8p36bv+Ko3/63v13qaR+D75bLOMpr
N9j2zEwkhf9iXfPxVOoD4YjpVxBqNe4lQbJpU/xAFcJ81gTIz+FycAjFNV5kpPvFPOM8CNFi7sBK
3E+buwyp7bdzuCawedq+PkGjSSd1aAUuKG/w6LEVJvfLv0/gE711Fbtos1tXVZBL/jWkfztU5/6A
WXIsPD6cZx4rlUooOfyM5Xf5jV63D3/DBpecBzBKzy4Hq7wr6dK3yemaCCat5y94NI8cn+42VRGn
dN9awg3vqpDdh9S6+e9LlkjhtPRCbKn7NAKzhOWWqWidubLluw44M62+gOxpR/1SCrJ0qbDfD97X
+zMkafikkrhxHGoijTZgeyo9NQNUwWwfw/qCjaGrD9sLzNgFjhTzDCQoe7li5nK9T8lKvlA89jvh
rfbmTsiHWnBTcPOFN8HYfb/LLLb9nmsVFZ7C95u9hKK6ssvTEo4hbjCJxPTy6jq5uQqJXFVp46Uj
FxtJ6LiD/4zmTrK+mUo5KAgyyqeXsE1jC2dbMVwpnMHs/AcIRJifawgOBcPIxyiPxsIovOHWFFXw
2+NTpeXBLPf/L6b8WNEIoMXgqH6AqHHxfbwrBYhyXNPZOpm3Eq96RlUTapc1SCqMCXiBRxywVu1V
SjNaCR0cz6jWte24s/OrHdQO6YkT5LedfeFstZupt3laTPdyc84in2bvrbwBUEoEbs5CDV8w5JAa
Yce/9y0JdMOVBcEShGdMdpyUcMtlX+wkvCglLl46uv5/8pL8JPQk3XdVH1R+coBnQycfspRzpBvn
X84G9NctIZ1qURG4SSBH86F9HOdWtY/iXkZADvALvRujLHOHdBCEQGuR8eSIDOOp8FeguGLq2Nui
ZDvhb4TaSWq5k0kNAMUo1jUvZt6y0ZfanN7mjV1uNn0vpl8VEv2KrIP71Xj3XdAMPGqJxA951WV6
brEdkCqykXIWzl+tZudZ57nHhhroXUy+9govAv+VncFgFs975Tia+K3WTd25kJsZzA/fUxn5Xko3
h4HCPh6jGggGjp/umeIgH7aNQd7Lic+J2BveXTXieqmChqrNerfMYKVzMnTWgyFYm0Bqh2rmVXkg
mMVpXRj5pTKE3YmQFziJ/mGBxjmesRZcZGBmJcrtUlygexIXbQBS8slC+PudQp99jmG6eFt21LU8
SiwmWjairvtAuXJRu1AkIrsxGoT2cWDofKt3qLT75nehLupxZgOogTsrM6ZHSof6j2N1xsznItj6
wvYBkHrfFgA2AlkNtoo5T+LdW9eQivy/A7VTUEuQ9tByIqnzWqu+wpHZpjE/Cpve8ocj6kXCE/HD
bylUMH0ktUenV+5rlOHRRsvwIEovHxcB73styd7U74oFyXlZIxWYPKqNCzKprBAkzQqT82HCzOeR
ZEs+Wn+LinHFdj79MhZ6dWwrid3Sv3olzOt3PlH5cPvGioxG/lhW4/zRVE5yQD6k7vQhtTYukQMA
jqejOq3uupowURBxVMYWOdRoA2YXFJwHTIbXW5gYZ/vqjmWSoGhVWp1gO/3b35eUClc0DReRDkG9
nttCFRcOpArhvxItO0HCezEls+RBztlq+Esa8pb3koaF5rm9Rm+Y547qB4zw6MwgJTCczKUdSh+L
GQTpXgLmRArDdCTuR3LjMu5bGKd2Bh43bJv8wj53i2b2l9nqSgdWAxA5GbOILtDd+Q2Rzo30rsRR
FKqC/ugf8plSstuwGHD+2Heh/9vv4vvPKGHj5ZM/AdRGaA+IDepmxXRtYWiyzWr8buIXLe0SA04L
hxtGbvHNeQvAZQztmQj1JWL3IlKskMJ0/giGM0os53rubnlJKbOv9tb4LRiQjVMTrJ16oh66CZXT
nYai+0cE6Tom83QacNqTFh6y/NezTdT98mxYFAI+ixzKIdWc6m5QOALE7J3y+PEEB1RaLDHSxgeu
xVZEeqY5jtO6bU0suHMsuy705kH4gVad+WYdbFYpZi2Yc3/LRJvh05c96N09E0JXmpo4XxyEDpA6
uQVBtobZqw60D6nLX7cjd8KwFPJFXayeqpSmphfms/M80wYI16DbtfTuQwWXN+y5hbLnW4OHqhiT
woNbJOzfvmWfu9Hj6oCpQlE7OTKeQsIjOgwupmDbDPYsicVuRCGOtdPOfxkPsZxRuYM9SKWavOVc
W0MOYssBpyHuW96J0lYXu1bci8rp+uamiEzJvLb/YXQfc9P6/FOnGlgA9ZSB6TWuPndhH26wtQ+s
TfO0C6YXiGkGHhjCvFm1CMZW8hPMbO4Pc8KSZvv1Y+9uXOXG8Wz9tE2UXBco4pFIyAbz2GWIRSLg
f+3ewyqpJ+5Mm3S1Q9r0ucbz9dLhCY5yPmjdE8N/EKLaVjkWp9rdHFhpf7gE70eRtIfYBuaxE/nf
N2hmGDfayhQ4jzN9Mj7LSAR1COYf2v67hgZ/YDnv9pGO11ls0oHNjkAbFcEHpIuGJWSzwzGY0MXj
Dp+y1wavxgXDBZ4KOhTqKsM9uhs2qtyUbO04k9LG0Lqzbo2BXOVVBYIkJEj9tIGQUSO8VrWRETWl
eBQjyL5xiQp20pfWLdvSRHBW1RU9RvXvL7IyV4LlT/CBJJ3K3FOV23aG9ugolHUPWPuwfLLinASK
2x5xqTdhZNAFmlt6bf6hTI3FX6K0eSGw1w5wgDyGBQuj1oVvDdr23JQBcIOXvQnoeOvkz42tVbun
q+zZB7ARth7DuOY1sN115nmy7qn5dmx635bTCJpC5azrbLyfle+uzGLO78VCaqRYFaFAR3hnb/Aa
r6XjGcAr8XjDIE/tyWsLSGHRklAO9Ab4Kdh+bElPt7kgY+HExiNegISJ3Vj6XRNyw9D3/sZq7YMk
YQiMm9NBxCltHwfiEmv9EvxxEpQwZRz9HDXG8UfDBKuGm3lHaHjpm/e117mCdmjuqGKdZLZ2pv/Q
Lj/J2xWnrKa9WmJQFP8Zmr1tsDJEdgqmDzjFSidqGViITj7MC9TkBD4lUm8o+uSmN0/hxorwMZRf
ED61uUgBs1vENWPPbak9NAtDYcDLBt1+ZNvIA/KLVl+p8waTh9DHFL78mh0dCc/6jZf7t6qF1dEx
+XrHjHTyUht+0jQs1O+tkQpRdOL8CeWifKgu3zKiAMtnJmIMDQe55/bPWnE0EA7EwvF9YU0J5JCc
gNBCf1GB4BVu7ytH1kmDyn9Yu3ByO7n10ufJg1m1JQhOlP092Wz8KdpjxG0qtl+vJ7tSD49dwV2p
rEUwWLrQECeKEizZczhbN/zviJx8poRFFHhCrxD+AaPsR/LMv4ykxz6pXP9Usn8QfeZDOgdH0PcK
pI0HqH9tHjRWvh5sXaGS6CuLT7ZkOvbPHTcb6Xfjdk+bgOYE9mvNXCtZnTdY4QM61uIXEPPL1sXp
ksVW5zTlzqHpn9TWss50t8fbOMW/3qmgHZYjMwgXS3Vmh30LFT0+OekyDB8BZT30hFnTsIC7lgcC
ApXizTMZNJW1K48DTEG9ThFNYOBI2vQUGCDYlX0Lumxbl9dfBoA46VlWmUk+Q48spZVIUnYA9wxx
DE40Wzv/bhyqkFk0g/me9FhNc7dQwWNc3GPt/niuVvRf7yxyGVjjU9hVYriLP+3l6QJ1j8ZQ5G40
6f86wOuq4EuLDXq2LxUf6wiapfnRDB0zhIbix4ACnY+zkYA28/v4p+SGlv7jyFZtg+EX+eaFSckj
LFY0Xyl9er9SxfLtCtn0qIxmJopEgQ1nLek9vTsYy84KM+iY84CgbWgE9t1sodpKlWBamz0wm+3x
xrVSiY0IOLMAOXqfKhWpYjK4joqrB8OZLNYmHxhkf7mhQMPNUzdLgT12A2OtMEpLebClzAIFagog
1C5VbI3MLc5ap1JerK+lhG2W676XsUsxJsxdBWHjjeo6TPkV50f/aUR6lmXEdN3QipXtC25GLIqB
I06HtkpYQbV2Vh4Rj2llteF0CgbSVljClrrSFq4p+UV65CpVfUw7QKOzMj83e5rZrHObYM0EYejl
svNVChmWhxdAOHvIS6x9tQWt2ECjSGWu2iUK5Nb+M+D0Tfe7vus4N9nMIuIXGUV6mZj1uhbkwPsK
LdOJ81ESW+opGKGjj1BiB4lyOAwt62EZvk5C4YxcfU4UsHQDPUPt22AqPC+XYKkC5fqwsgw0FloD
aUYYD3kjbNzCdAi1DfyQseJ0j1TFJsej2kpbV7mLcbGVZbJA0zWDTa1unVzZfs6BKw0wCM/8qyFE
z9lKlN3I6f0Lr1NL00eojFvqeTEpAZ86tsUQNlSLwVQW4Erw6WHpidGP5clkH5Av+Tw0HRF1TI9t
QPtPgeW1ssKS+vnRjMriXYp5XZ/gal+YeoEmVGUZEU275cZySX4/llMniN9qVweD2ggzPYECY+2c
1rk8NjaXy6wjD8Khq0TuPA1Hhs6Cp5zl8WYooCek7MGXrlMUSTaNJOzPPjkM2FspbCKfY54ZEXa7
kD8WTAEo6b+SuF/nP2RstlRX3ljEphpa6QzRj2RLfxsaps4SQFZ7mv1hdzfHWNwmr3UScgWOTHrg
RFWCZH9UWgLgVD0T1yRXI7k0DbQ1WLyrmzrN7FvHY19e8J4Sm4xcMmpToCsbCiZy5j8rquvSR7nK
zGjV9jL0esrcigctgs6kD3Pf7WoacOfLtkp0pThxwFdj+bW3S92ndPopvlWqFj3+wYXT/qlVLOe2
fngAwO2VF2K9UGRTuWW5ovSj/N7sGAfr1yU/AcV4D1ECJBPIST+J0HGnmFupq9UOYhurhEMFE8JG
b0GiBFHDxO/hy9ZCshdwh7Y8q3FApYCDIaP3GtiqMkXkxg0Vg0WzeE0GyOILvnJQhJObpJ1+q8F3
MngPegwwsxdwHM0b1lOLHYSpVV9huNmFhMP7XCKCrnUA+xvXKls6ZNXJPBkDf/xuPccchwJi6Nx2
SXRPx/IBrgJ/WOU6hvvvGpkpCKoBC0AfqFPGZjaEAIIVbviZRU4BNngVD1ylOx6T3XJvfH0TIgu3
a1fru4OBTJ0HtazIqmuldyY7tMnQm6lw9e/4gRAhMPcdZtQrmIBp91usD7dSCgtxqDPlxu6qBdK/
QzJA4yv+s3gWNHDrkAKK7H+YCms80A6GCLOxsTjM0MV432E054iaiebiiFCaLZfYjEM38O5xYlyN
LrjppfrTN8kQlQjis9H8Cw9yxhtloUNwbYJlZ5zXsr+WdhmkGE3sBYDFZmkOOJ8/YS5CbG43acpR
M0XHqsn2a1FZR0wY3JUJE2pRnOwyK6JledNVyOoVNvQ1aRYbECMabp5wkYtx4odwR8h61+gdfhaJ
3kM0StL48pmxxA4Dezem/G9V21r0vGyiNObXiDgH+g+/uQlRIvl1wSSC82JMoQ8lK71cTMrJxmwX
VBdrmUHjzFJCs0ZzM9NvEZiKvNbnMB6T09GtEq2K5RIGVhEUmBATyG8fYAqwiuyuCkjom7NPOSNA
qMaSFKTEQmH9ESOCkhf3ADr7dCT0QdF7pXdZvCuq5Gu+gaDowAIhRlgfc1gNFvLvq/1SVLPFCovP
3mdr/incgoWFJ85A5eKJwHqE37YyVWIy39ZQPssql0/tbGxgEuNUVxTTxKiF1FKHD7JbtqqKlf7g
gxBy3R+axmJDu51uxWV1w9QSajZOyXgQMz31biDpDa2Pvg1JZmoKoLCM1RjW2R/SjzfQUW79y7Nn
ShyXRXFCn1PETw38jZnS/U6f9e919TPAu0ToptxnuC3J3a5z4rydov+pndKZNEmu6pKkuAtLXIi7
oZk7Y5XGuj5GLOTUBuG1S5tMhC01FI/tCxX/6OQqd5CFIx+9arFst/pgMDoPMpNs8Pl5zaeRCE1y
izIe5MHODWLqUzHq2Vlor22D41gu08eTEM5EBdivd9kle8uc/n0kyEfiDZoFh5OSVo6a6cXCQ6+2
DmXByHxgiu3DPkxvIsVgknDUJS0uaAsE9p0UU+XvE9I/1yrxiOlUZ/ujwV7ZPKOBmCVRXeK6wR1x
ZG5SIXCC/e9IaqlpzT/iH6By7XLqOcRAKx2/RCwTZR9Ej1fiZ9hbbxyLxJlHNjT6TdN3kufaZcl9
5KpQ1KaKKHA7hEBan85ey4jzyZuawfgaepGOc8Kxmj8Q0mXlksjJb6aTd02RMTAfrIFmNxYr5xTw
Zml9bdiA6Fn662QrE3IrKRlonTHJl9RcNKLZr1phrwe645NR5DHS9ZLJjfV7V3/6aV6mcU3ec9q4
UEIFplS22N0MXjtvkJnuTJXHupL4HXQi6x5FYLsNosLx3iYfdk3GFOHrF16bhfq9nP0aenZ84Umu
2XpqQ7y9O2Re4pzTE4mWTQUwKg3/0YLRuDEVuSX8880O8Vt464mOKJOlHzsT0iMcGHlP4uG7aON3
EXFpzfclt2x8I0w52CXq85kdrdkanAXQkMt920o4AB6/vSTUWgOmmDqx692GJdDjHumccOs//iwU
qJddl/WVB3OcDvYeG5UBjTRuONKU/YGr/3zLn0etHefCAwD3ZkTXGNfQVsK6qCthjxQgJsyQzOu9
yJRTJ60k0NJ2Ru5N7TegjyK6qk//dE+SqDVJq8a/9TwlUPd3fisF7oGGeckieZUBU6lYaq1aaD9F
IxKPWYUJ9eGGVe/Dphap4K2rLEgVFZEGxJa0Kut+88vJ8DO6PAo9GxP01I9FwofFoE45HkpIFeUR
8UEonb9Jni9zke6UExW9/VCMPkOWo1LgNRLxG89fFR7a7Y+DHBRJW1y8Le1gtRqQ3h50KsQChkzC
XCPSspxkj+1byPjhlVTQiB470a+Gauy50gHFF2pQcz0qsT3Ao4z/NhBEhQzRLXlxGX3fm2KGb9UI
/fuSKGPDhyGa8bbMVp62f1FmrP3k/rVl5QlXXofW0BuEN+lVxNP5Lwn4okLmqG7SBT3nr+mOgftV
x72IDJFSFMLOzdyTAakk3rt7WHlCmgXW0GLRzBI9V3PrXSuY/AHLvOylW+CJudryJfHk5TWVpNRN
anZYPsmvXlKq9ptOdNpOL9i7CIiB7z9nRqyiKll1Tbqbn/TJioaA229xZmodSeaU4BMnwpXCNr61
0nKjkwBEvjRr7Ozntjam86qf5n5q+Z4AW2yl8t5xD34+NBsI6qTttGg7vh8Ov2kkgjga6fTX9kZZ
XDZcIduKniPbHrymwrAGDCZzYZz6NseO+L0TN/Ndz1BoXyyn8rOxDuYKxD7ZKO1wXvpSGJXTQzzB
rLhwXk+C6Ezme+6GA6saff0R2Qauzp9xJr6QFNyf7eBDN38ftArMJ87+PwCwXw4/sBaO9DdojidC
Xzu6WRWD7i/9F4275vHXAww95PfZBnhCfxsvxGdKFP0WXJ7OeD27VtXlSVBMtkEzS8X+fN6EqZb0
ElS2Fs8/farngwQlQ+iGAYaxN2xNczZWFdY4updHCP1MrKGYPnOtuLMmXptUhs0wmM0fDwgg25N5
9+xdmlRnX9uXLcq2zxU5KgFLn4YhCCHHBjhuQ0DAsZkNJsgrdZWvjDriE7MvejwBzHh+EWjOXUpv
RB+CfzpvCAEMKaXSgErDUs5F/m1cENzWmS2wj+Elrvx8RSl3IJV0Dmc7TVxoQMniPvyfEiE0zuul
wnyDsQVBJ+5aIE8wAHSBBZi1k6LOi9Kcfz46vN75VV8v7M+xfTv7RIy3CG5Mdhm02Kxtuuw9OOgb
yKyOUn04U0mEsRx5fz6zVUjXbQ+DG91Ahg57iHznT+zuhfqjbo3E0S6mykRt2f4THxL+FWhoOgR4
xeqb+Fc+Zs7bzx/nLpENoCdH/tge5cOwRxo990qgURB7LKIFW13uqjvEBp9n8wXo+GzeoeEF/iHk
ntKVl+QXCpNsYZ6ejHfiexek6MNMKtig1LtmVuOy5+GjqI0Q5LYNid6bOUMeDDcG1VUxOWXDM0co
zrnKGZSje2CqyldOUjFEXz4vJHHTU4h+KM2p26OaneFC874XCQuGc3/5Wa/g3IL/r/rT70O3qbQT
q/rv8bDw1FhNxT89a+beX7wRaA/oFGjqfftAh1rwqIKV1onCjt7TF5pljBba5zPPBzy2kqgZ2W9l
bTySh9FlkkS78XpxDEDbrFy5GP+xdEF9vBI7XUN1teGI/A1Bf/KEPdIMGqjl1ycF7W2OJJ0vPCN+
l/9eN9aqzVyozDrNsj/OrAK8D5OK42ZMSifi1TUJhRqSLa75t4bJAZ9mKIQgubUDyZhdk6uJjfEk
0VrnJoFJ9gr4zN5srFwXg8SCMDwJDgUsZ0p7ZmNrv7meM2vdGkas2gKDq5NwpZ91Ftelms0mrkmr
BHZ0SY1DFqQPAu5HqCG+DKwpgpCokptULHx7doQYjZd/LLZ8fxvS/6RG1YKClOTWCfrtcRqNZgNW
XAZplHvc7ezEQ/s5WfXKi0ZXgS3qQamzyYPQmHahEEK6FBUGnCLRyik/hkDXpTUeRPUN48cazBjz
BNPzWSXAGJROSM3whahGwMbboMa8xPF8daX7FTvLyj5Cbd99q1hCQ5JziS+aYCYsxZoEVbkjHOpE
p2+soKHY6fzUVcjv6f5ASPjte+MiXYwlERZJckRSUyhkOMZJj4FBSLEMAggs1bM0RPzyAxfcg4U0
IzTnPP7iFvGT25mSlpLYNAFrGarDdJmVIY47ZXg+VnkOGDMnNUS30Ng2k9RGeMEZ+4Fn63Y2Qgfj
3uIqHvFehkuAcUih1eLzbPDzUqqZKQ6flQ022m8WQOuHVuOWqUEctt9A+L63XEL/n8vMPhUk7WbY
2gu2t09Cr1WAXwD2lBl5aOYIKRQuLH9t82yClgLa/rErUUibgaXf+yB1CF5hA4EHGMd1g0Ty/ZoR
mSPCX/DSVeVoJ/m6YPcDnsc8aqN6/9vBTQessh/v/WqppcJEtT2IROVatw+A5nY15JsgJ8bxKpvT
e7phPUodWu65vsE00frU1Oq9IbX6nJ7cV6tXrMYIWxH39NGIDtIoGa0rOoRycmW10oBdiQECYqhE
Dqj4c4D0Ce7ZyoSCxgOYrg1zHu1jtRRdfaG8vvHAymLA2RReFe0RqTS3aJI6WZhc0lgd+PN4s+3U
8yqyhh25s4nX9oFuZiWHxmj9o69/2jqPWBz5tHLpF3k0tLZjlEEol19VVx7nGze8uuBJpwt/HdwE
a3D1AziDj9vjpyfJZgDjLGdfRzuKIsX+3OpAQBa4q3aD4Q/P62E6uKvEX3gNhC8pjNMyMznl1vI9
whGbO3JN88B4K6BeaziSDDgvtrTlQQJT4P6kyXeOguTP3su2VbEsznadc3P/EsdwZYdQNf89T5V6
22VEAyf1vaUrlMXMHD7P+oXRwKfX8j5+f5z16WZS+EXfVpW7sS3rq/1aQ9U+UAkzyfEPY3fByEi3
z24eZoAtzGBd/PTDkYjoEcI93MsKHZn0jQZX6MKTojNnDPp3sGA1hY+RBZ6G2aO2ZBCflCowiaeO
83ljiN9xHNOoCy0Dy4f5jzNuAxJ3aYO7tfsZUApa/TZ5B01JZ3MGhfOCqDq5wxdz6Ysg5baTzhjE
OI7YmH/H6SOIAaq0cQyr+DxgOx5XMyoLDfkWXNVmfaOAOJAWg+Tf49m1uD9AkONNT2PaHXe9gPzC
9rVqK66jGYd8kBUZrXhA1yYWYgQ2JTsW9kdQiyDsduA+gU/j79ZaR3kkcoxKLDrYgSGuRaweQpst
aokkQiWBXvyq8yhHzYSwro4Us52CYWemz+QeiF0qkvnqIY6naQ3QMBQJdl7qThhmTcM/f/QKXIVc
rCIyGJNkhv6VizwcKPEmha9COvvgXnw2p19zTBsHaBx98YRx9cQN5sd8T9eH+mUrRrE4jHnYsamZ
albTdmFerqk3JuTCHWg8kBeDxJ++OkRVbMiXeHn33Cuc47CarH+vpf39Z7M99ZJc+EXl5jPGkCks
09MKvsHo02o0bw85TTJchINUKFfzJyeOz5X/UMEFnoSRNzxdReAFEmGgc+QNXEPrNJ6rX8RjaMeo
auoVg6bYPM7fxVGtcWCo8WvLcAYe/BuCj7my3I5bKD727eO7FZyfHCiwQlc/lwDNI2gBmR2V3qSO
TsEVUqYqyCQxVDqfEzcs3QsRXcH03elhMJZrtH+eU956QDJqxYpcY4n+NIZwblUiO7ccDDSu8Y6n
PXyHBcZeSBrjZGLCdy6KZL0lRLLxMre6oW6e/BQ4oideNi398mKmn62E3TzoFqN72c7bQuf2nCWA
yeqbSET41vNry8vAq9MhYvjrRZPnkdo2ozYo3xIHFQKKPPzC8RJzpb8aBUj6pu0aPSVCXWanUVdS
czgETn0B0iGlxjbOGukomuphHILmF5RPjMJZo0JEawp4DhhdkvTni4F4CnT224ObbaxLTVJcozMY
USYTuqD95yYOFWXNuVZJM2G78vmruDikqOZ4gnYGuVtEgYPYv5ScQ7KzVsnE5AUKii6s2gbxPuHn
tz9DEzjFRP4Utn5hjBkwtTnbBjkIp8LHFS5f2ctk4FjdVIdC2hogIrZFTu4ShDwApCr8hg4PWlD7
OXBh7+BceFaFM1a7JtovR2O5eGcXIQHYSJWRa+NnOd+3GYGQfPaF31M32B3aTsNjrMpjvOxSqcDa
a9GexqBAvtPWuk4Ph7Rvzxi9gogS91mymyKjC5nVdyRsGkSJrSXsQcQWJtLVe6rKo2TpiwvK4yh6
6AG+Rv9oXUryVddHr/8p1O2DM0NUNAfmjihA6HL6e19HLfpwfqweqe/ZR0GEUojUIes9YIFteEeC
h9XExcBECf9vA4a4Zut3oentq6XrNlBHwkjuq5dR/WLWNhwPpLg8b9vV1vwprTKWGoIXICuqt72f
swbtbrh5iFW70IXXVnzu/XqZ2+jPDVxgggWv5kQZxpgLrqzUHKALOOlwBVGvd7fMWTjhc4YQe1wd
nmc8G25igpGRaRPVktTTdc3JDM8uz0+bPpbMb5mZ16qeMSLmz3ig+TrAOCoYN5HYMzBaKp4pZQ1G
q01/flaWC+m0FqgdoPyOZ2KuxRSkIqvT3qyW98o6mLAZr811XP2r6E7Ad4NUVFILdr6zJbATwdgX
p9n1GRtwFfbyfBdeweAg4A9YfxHY/WnhJ5hhuf3WvsNcjOqArRypwbj4qVxltd9kUF706+9jMTnV
Am89P8OXB9WuI180jiJwq/jAXbcmQaXQDo9Boe1+I7wvfp+rN5MlvzQwjVk7EMU4pDy3QKL9E/31
Xu4G0hjyBfO6HRNAQGzkB+ey7nEhGImfd+nSmLyViz85KkymHcdrniZ/UZaIQOalZEkI7fC8pjP0
bQbBMJEovzoLcLPyM/4oLUfgrjzeL3G5m0rjrVRhJkbO8sD4lgAsQICAqU/9OF+7od6nqBYo/LR5
M+BYm6+g4M0tzSgMl1B0k8zLn1rDU3e/vlcOnJVU4h7nDNCdpAdy/1JGR7/+q3zJGHUIRatY7ZiF
RDlpUvcp+eXcnNlG5XDR2kYPPC0IVmpgcq4DCkxpjVI9nOLppq4qtTEHxNBIwbiSgoubL4WZfAt8
2+qDhhPeVQ+zCqT78gvQnPP5uaRXIzHc481pExZR0BqLJWNdwo19J1VIAexwirqQ6GBHC524oLOU
zRTK6vw7HChu12j3kTK27hSU2bCcveMrNlZtLGzhGUPUBlLSLXoJm33rcUcRwFEhOWs/PFSeJDwg
4ytGjZb1hxOctLxAPj2Nt72AR42g+b7VA2iCPR+Mx8VIgv9TFae0vH6IBY+jYAN9SZ0/YtuQKCjq
BRT9AIpbAV3qAM+w+Y9z7gBQVMJv3iif7l3EoaD036x6sm7WQc7nIgaThGJfGHtPsjuzTTRWvErU
kvIcyuqOjg/KXSDdXd4K3G8ipJnyA9jCD5ZIZsLXKNiC8TWw+1MD7aNkaVZzf5ouyEaIQextBaJz
fNfsKwXEPmnJSpAJqF5IsfyXWc0BUezzQXNkViUYCUygX2T+TZaOOG54YcRdn2rusOuGgaptQ6yJ
K5wdGN657AirFHO3aZ4HHkK0aoxEeCzWjLj5Gj207uSZfLbFGikQtdFLJvizR2ipT8Q2rC711Cp4
9+gsTpOu/eyEZlQZZzGdciJ6UYRNJCqtD5Euanwcx1A8gZryIqzskQLP/rWqxAy/VOH4tl5XWMO+
aoB83RhVS0iw8dRxr14+hmoZyKbVZaoQ8tIL+elfVVzXpbPZJKl9dxDIiV4vfZ7oyKBHtB2TBCyI
LbDerCBGH6qcyV6y6BK8Z10x2uJmWb66cKQHlXQw5ke+tuRRhwDp7iSNox2yjDLZPL0quKDKsrBH
uBBIB48eWNymjLGiYAC0CcDEdxrqkJF5/J1m7fF1koKO20N/NMMEsaQvyGN6yyq8JG8EjakyH8mV
lqyZ7B3lMvGORXoXiYo9VgC3tZLBKV7VxCSiNh/ixyV6cF8+0fbfqPYAe/SPgw/PUE/wjH1w7L0d
q5Xgdjw/396lkPAaA1yxW5ofac5T+AfhuWbbwyHu/zUh/he2KTy5qxEAbiy/gCHD86I81bUfS1vs
pKQREfQiE7AIHcshTxrNrEQickJ7fBTODcO1OqL0uL7b3B6AaNlCeHE+K0eiP61KNJHMaXSCdX+T
1AeeDRV5zjMrgR1gp+6vtDhG03GHpTZZ+iYFrrXweadGvZ+dMafcWcZ5hYa26x1xi+lrqE9ULTmP
Fr+SZaf6UJlq7uEXJMXPXPERTuwWz0cDJ8tFla4Jy2hCeZEyEp6S+pVN8WWApFeG9QTfACgffMht
kIyEQJ3wCVBSxONN/jmzBz24jzFsQRSzYYJRSy/2vSns/Fvrlg4sdrtHjqpcHW4l96m/wLpNMUPR
20A3pTpRpcZUo0mWGsB/MsmVVQ0E00Y6d91LJ2fgah8HtdEtioSqyS+7KZRQYq8hKigcLjC7JdCb
oGiTdJqy0KNtVybFoShkUMvMDX159opCgI1ugNWthwvzbYngcq1ygrlw2VdtiZLtYBNDMxhoUfUg
ZhQ8re8wX1pFnMB9gV/+EF8UizHkJX+pQJFnC8l5zCplPqLUg5hQwkWZmZU3mqtgPjNqFQhOtUt5
8wR/SDMGSt89/qqz3uCj16meAsE4JKUEwDd2a7K3C0f2C9oSAe401l1CkRvkjnE16jQTFfHvoyhY
p4BJndZtEK+km14glDprufHSMF+3Emj/XBpDJbxva7QUegaBT5S0GcMm5ksEXLGY4rNwEkdR7tzX
HWCUdUvXAU5Z5gSPHURboL1CElmWkMiRlLaC0cm6lSiKLp8FyFx3rD32D5MSCSE9tJm7jnwB73Fn
1Fj7YyURexotOoEWJAhK5oCA9WxLBAZEdQ5h6JhS+7pCsSewLGi6GDRPxirisMua/1WE7d8OPx6a
qLPCVw2wXbHurMF/h9fImADzh+KehOJ2C7KQp2mTiVrdsq5O8HWxXbFiE4jdeLVQQHREVF2aWLJv
pXiWO9kfcRFLzaJx/x5aj1wr3/T08ExIcT7g6L+uwuJa1I+F+s+1y6MBxfwLs1Ylk/9puHhu1u6v
FT/xwsantPqUwmgwdVT83TrRwq8C/7Zr5U/4pauQFFfpim/NCJOgYMN8Sn5K5B4jd8fJ4iCCVUnj
DAxTO1ApfzS5aKCUeyQWkUA2/uKPFLJrLLfOl9i8SJ+rtV3bU/t/8cdlCXDmpckC3m12Dit4nC16
RBmCleYS0fu3ftHnoV8bowysVUDnf/Z2zNnvQ4zTQjHAQ/xilhtphlMiZRxNTwHGYy7yF3SmZsKL
DUokwXUmuM+UyPdJFRD/7y1AjDBluV6MrcQd0v9CWiLe7/w73h0HHxiNKxbWedGmAxyo/Q6UMUq1
+jd6WgCeEB1G67/tFStZ8yFzhUmOSASgU4zR1EAG5cTt/8T/7WIVlnANTEnUo979tsBiZbDFe3JA
51F5hfKB7LC/DyxtqxD8TpCcaQlDbDcFVXH4Gf8Dm//xgnCL8oeKhOuJ4+k8v90DZmMZk/tAxNaV
oSujhGO/NIsWBmSaqnV7Qo/KnviEEzrzg1CEEwMEuCYI2aeo7226M4d/Q00ZUkWc1WYnzN2n2wZk
bNDtMfP6NO+IXKaX/NSaJzUnf9jXibthhXEsqqCA2kLsJAjhO6Od4kem5JRy8+MYYLyvkvGbSH3p
o993u2kXGEzpEi0jV5ndYExClLqN6h3Xp2RkxvBVXW9HKBzPl49y7CEDeyvce06HWMpC52ncFGG6
AzcWloCfs116+NZTRroeBlzTjQ/yw+29RoZkida5lVhFN5TxBsnmms8tMtJQCzo+CudYIssA8CTM
IWS317/Ox8LOJANPNDe78aB0ZH1V26kPTMBdNraIimT1qLERKrPopUqJHtGjH2OUb2btqK5zpEqA
y+RkyeB2p4tBkpD4vgP7pvNnHbPhkr66r3o9tGWexKlOVg104RivoT5sV3ND/TUFmFUYCRNyuUvn
lNvHeJMdIK1hA2BnoGQNI5QoBnQKDj9ORB7Z/a8K+1VKpp2SIzIhHn1y2HRUzB69UpRHGIKTGxfE
lCvh3Pjo9X6tsMp4Ohn8kDasElVxU+nmxQvD5xOpgJXhFeCLi/IRWyqBE0NvLO9Jp6OrynlkB2J5
6ACjmt/ZDjMZaPEOrU/Q4yonM8b/2l7bm42tJI4wlo/pNUoMQApI/1+TcA4LLBj1pi3orUERBmFO
EJnHq+qb/WbFR9yQf/chlRqnjsbglkFw5JUfSzlhOsCoSfVCcyqjDxzaxtEJBmuQxMlvPjVr0tvt
dagDB+DU4s1Fl/tv1nuPuWEJ0/Ahauv1jY1vWolCMrw1D75JShfFrOdbs5M8gUDwdsaeXi18Ffw+
eQUsJMTzFYylvTFGDHk/Cmf3NWC0ZNAg/VUw+h6ZOPaFSO53Ad1ua5Q4v8nsFAf/ly5I6y1PJSyk
a0bSnEfV0G/0gxAjaCaKmz+tsTK2h8tesH14Elf6Y3UbBtPX06e2NEgnzmZ42L8uzuBxzdaMxLXC
1KHSgZluA6KnaDMOucyYuXGubkLsgQs0toZUZ0KUrcNYdR1jNzV9Ic+D/5DeNEVMvBOrVwxe7uvg
ZMAGMu4uMq+o2HpugqEqm3Wt6g3TI+J6nInm2C8wfKyFF7Vc7AhYzWvMRv1qiOSkJLmk6wU16ZMj
OCtjDtNQn2Ig7iPHmYgUZwyEWLFby/1Uj2Ukfp8rQNGFrEBy1KKHMrl+9IpG3jhCoH7GCx/A6AF8
cd9r0wMdiewkUqQhEBD26Tjvo2wVAS4n7gRwAqyRmUO9j/WFv/zDdNAQPMe9p22FpWkVPXOctKhE
kFqe03jv6JLM3y2XPB786IL5nND43NFeFaKp5JgY2JVCSrEgdu3VoeOJxzYmRBwXgcXJ4Xc6IVUb
B+78L87vfNub9B/izCQ4oRHROIZ37iClrbtT16AbVkC0OdaSNSXN/pvK2gPemYp2cYbBsgu1kA5E
g54sona4jodf+PVP7qXmAlHJuajTdVuOKopRyG05DydcayRnqWBV//ZPN9424BmEdNgWiKJ2k7vK
gBcMHnnfZPuWY6SD67Sllty7xUFkO4PRx8RBJ6WltRmmpLQZVh/X/w1OoEnXWI9tui56IXt7sMof
vfu4RCq8QCp6qaLHlOGzpyiUWQStAoyYBfKttbXo7Ml2akE1SJfSDhwHwbJSGUOsxPGiTAyLLT17
5xvs1v8bDyA7cGpdVvLpEq2n8BZvI5AqRxgVlolHATSaRal9aafN7rqXQ7Q4+Szu41aeO3pl1awz
VRoX1nc1k7A17bpJJwYdvkD15Rxd2DlExnJjShu1klC5k/t0mrdhYhY0k2PLnflnQ+cU/wTWwLLW
XmfRB5EY44LjBPjL8Bdw5nNQAqTik2SN0WEAOk+WHZtu/W+bpfwFG5oaHBeCdw2uS6KqZpnWRbN/
yrw3kRG8UAOWRpak6ZGxkZJl1yuoFbaXjPEsKwVT/vIGrqIJ6D9GB5ayC034pn059IBxqietAfE6
t6LCVNl/CHBjBjZsPxTWAwtcQk9IuZTKKSc87CxSO8vlh2jgFqymqYQxtdX7cha1pqVGQ9yY5BMH
KRM3iF7CCOQeRu0wpYKlQ1W2RCwmq3Zg4nwpBIowLte147XJb7TYCvLFJbgKYwnASN78aQBAAL+s
cBEcO71xcDxEKJyT7yjZF69ECYqb0F5PRa3VSeL4i0nEYnVMVUoMPXo2MsVFZ2Sg3cuNNphrzEDf
nYfmznEFz6tDgj7ZYJOhkWNx1DqCrCnDMG9hUuTbChqCW5+o1cz631hNTZD5nq8UjuPHMdkxVPvh
o5u/OYyWnuoqeBLxY4pCzs/Qe6gtx3tBkic4DBMXykMZsF/qEln/ZM2BhiwfDOBnhDPU8JCsqd1O
A+WnQd9fIPL7Cmx67AvuBB8uLy/x+XypwGDCRWtHH0J5CAbCTYJBQPjU649Iz/Oo8byA6WzxZaa9
VXrNv5pfiyO59TQL2hoxU+FCpT++y5jzUGjXfjdrVsfhDGGntceAPgdhFfexK6Tcv84z+Em4GPv+
3U3MiiyiTAjUY8B6WBKbz8FNK6RjXaQmXkt/QPQU0z4UdVF2xVNI6YKQiGAEIH1PFz6rcnVoKOOb
pElqTUZd0YI/i1EZ+BRn2dz2QrseE2ZnIHl3draNdANtwKTYWtTvGNBsDWjEGFcr82E7O0mEfVXl
ZUrVmw8POPYaCCcD5fmzMVvXZr/8aT8FABcYQA3ByteUKCVF24LI/OI9460WetCi+/NtomA/UXHh
G/V3C9HHwhzgcsd3DnIamRD2SM0/jUaCN1YxCjZBOK91DzucGMYo165DMzYylrVRvicDs8/dbwj3
pLCtmiqyA/Lf2d6PI+uDGVFO7LyXI0JnYs1Sqyh8LNyVi3X7ERii4u2kU40li1VMRAVrPDMT/5zy
NXLbSbXR0Qp9ZCSv4NPHYospj+/I4gByk+l7Utyn6+MYmY4Q5CDu0xUMN8P00ZUk5dEz/buZ71xZ
synxV8QuT8YH2fBT+0CmoIydcvAR8NY0HBpqoxL3amP6FCEFGZcPuzw+5MmU7kWv35b2fFyhAPsD
xsFTY/nHpGDj0dsJc3wskyiG2c8w8qQe6Sb+1EzAhmhqUssYIgsAeMxkc/2PU1N2jR5gtA8+vrWY
fetFXca3Gk8AXZv9Vh4AiuvgeUOURvrN9rVMuY6vWtvFqZyAoIT4unDE8XISAGIoTLTdRSMKNWTa
vGz8uhBoydHJgrnWj3SvIOTL5Blnrn25nA7BToGE5oy8Y6cVukW24ORGMSWhueP/ETNgDZQ9kSo3
16451/WYtM0/g44CF+Cqq0yWjB21QVGOL9TyP+/DI01aeas+4BsyaWFt7Q8t5J8YC9WC4lrvp/rB
ErbTGoaRWyd8p4ROKt8tF4G5E66abfxLD/tt75q9yuPooZcRiYKSsTzdIW88sM2Q+Wklo872gLxU
KR6lTH1hnvLJnUtS+v1R/+IhbxvPMoqonPTqhcSXWtnr+eQq+457cPslL4r971q3RSVlDeTlZ2fa
+fBn/jDX23TbQTMEXplvS9trXv1F7+wElpXwSppe2XxDN0hAdZZ918TvnyWONUbF4BVNKjqKhfNg
bG96D8ja0NFJVCvIMvZ9F9bRQRQXH0o4CMiSRxChHARrLfFT/B1+vW1NfqsBS+1aP2ueMXR6yVdp
L/sy4HgqlWAuJaMes/uvcc03PbZ6OtgT37tqoR0j+1YkhL3JKzBGxGHXkRxH3Nz0yQH9aHaGvoiK
4zyOQX5DKF4Mk5Mm7tfSusJbdqoNCD/azaET8UVVcV/U6vEI/oV5rFAoR74EiyXTKsDR2oBmZcJQ
UlYZtTCbGQHWAICQuJLLJ/DYUV/bLzNeizEWVMag+2xkf0Cx6ALvltbYHbl6Uyed1L6lt8uS0jUx
WQJDt7bh8v6gciQIL7TMhLt5Kh+sqhvFUkBgcUSTLx9tsvwnl9krP2/qZSb+onlhByI5hGMKeR4g
/BVSUl1Nul/F61UTYHVmfG/cLrh3enxr2n6r+XJM8j++uOqup0rqR+UDHkeTdWyyeuGwm9c7+KI6
+tu2UY37Jx+zWPxaGwLzEvX9WmliHMqryQ9KL85CTvjixZwbMKz725zQHpqJoI2i8gi+R76b8RmF
BnfGtySKIK43JFTxgcfkfEmB8cHFtjpDrq7l7uKaeewrfIUu5gZTp9Z5MdIVUUjLClQMH0M64xP4
gdR2MR4RvIeh8nCH/wb1JFYu4eZnZpx8WzPqvsdV2SBydJJf4md0BVmUE77SCRgykXLyfoKvwWCJ
VM6JXj8UmPxf+W27pt7kXXSGNBu5PpJFd3AfuNAvq52r+JnYC6aLUj6Incp0pfGNU6cCkxb1KZbO
g0bMsSYVw8kgUeIf4vzO19SQW4cD/XQGtz+IA4NyOgoxUxDyyU/1YrHRtX5YT8X06m5tZ7+Al0Kv
YY0t+vN32c00uevC0ulgH5OkJqtSymKB7DbSsvkIKKBaXkA1WF6X1Kd/7obmlClv3KOtZzilqfWn
FT4lpioTm/2nR1YgKB8NrGuqtnXlVmVR+yzbFMVjmvHfbo9doGi9Lir9oaW3oEqONq2XqxxmS4lj
mZA6z5D0FE9kdjmsJlffLb/xB42n8yulCFyD8cmxTvNvwiKpL0qEw1f0pjjKdxeoCyGSMiNux4r7
4ovXlYhimxGIoCpfhH/ELwkZ66QiIgAC7J9BG7fvFY92n4Unm+yXzYzdrKW/w85PiWtfMsPzi7N3
yudDVPvZ7bV+cENKgwG71Xrm0m+vdbwAOYN0RszMgHDhyhc60n7Jix+k8zC87DHUdu3Kyls/LjQP
b6XThFSAsuROoF/pKQ5OyLQX4q81ucPyjOdVdB2dqUsrQf82SVmggrMrldmmoVPxBMFJmWNmMd5W
hWF6f9sQ3P+Rw9wIf/WKk95Bq3NAeh/MfZNQ4HxmdPiULFcrSgZT9pjXSgQssLz3KGyewQyGYOsI
DqJtb+ekYP6HPb3h7BoAc7RXZdZ7rzwOTq8UqQMgUXVjqCDlq/OXRAOexA5Og5Ac9FTi6W6ayucB
lrUP2ztXvCBPjbwvdsXdaj4T5+xiFxW4YBzmm+31tuoqiv9LyzHCESoG6wue6mbyBUxsEFTH2MKQ
hhCXlmEb6iYcvgVjo0EGDK0fF/oM53MWl8oBrVIWCUNK38fZ7DetkJERKh674Jlsz35Zadx1WU2d
27xSi5S60nwHo6nUslrxDwZtPcbW9Q/qDLIaDT1l1a81shf8t9AW7ySNpGQ/aluW71dnMyioAAI0
esdsM8atCdR+cnRJq1gltRkSh4jpv2UtVWkJb+hjeN4g+TlVi941dDVpkQOedcfYPn2oR2D7unBk
1XybL0peV8Asz+eYJJgTcHGpIZODrHjnfa93x6FsrPWx1V/oBwu+8To8QjIQ9/ZZBq95aD5rs+Lq
qrOjau/lKrsdAGJH+R0M2w1SbbclvYGq9RstkvAshc6L5fyZw0ha0VYwC6Rql9IG1HyDz38i0m+m
7KlIKEhCYiS2jtqZnhu/Hunz3BAOAIYDfAMZGWWl8V1LXXBSe01OU5fDWc6pkW1KHlQmjIYpyAXy
5r7WnghVXdgfbFfe9KuvCBEBB7fXwZIDeZvjQU8TApCbZCQYXYe+mMmGlc7ySXVcM6fphdlZLXLr
sDgxssWyharYii5SXt/UijUb00ejp8rgyWUNOmf4f2RUECJqlfm3qaaOE2uylvsH56vqkdrnnRE7
AXD6BFRQ6upH2bv9jBpRqBgsir86AgTatjuapt3IPWM5Ds4uIvWLUQhM9U8RB0G6dTwcEB+t/IO6
m+Sp4YgCX1rAMTvVjvTdK5Q/O+AThIr77LwoBzoPhaRusU/y3PWlSzt88CKW2O2sgOUAV5JiiiB6
nz4oC5nHwl2KXFBumpxAjeFT+15zfHFikplRHIQhJlTQCVnRYICcvMrfMMDHxVWc0FcLcSudkAPS
9zAowrHFfrMHqXau1zhWdYxXSeR55UmkJw7Bgks7Y8i8MggUcBnCTssjDGuXzh98nsTqEjkViwHy
KW2ftTi0UVyvOkc4T+e0bZc5yCVICDTs0wt/YCLE7/fhLezKgJ45/8MxBG7A2mdNbpVTS8y6ozH1
kXs9t3OY+aCLy7CRi4EghF8SYuW/UpH9SDkuBI7SmTBMLXA8Jy7svRZT5GgsbvX+rWkjAg8LLjHU
JxiT2XwFffbQC5CPTNecMGrdU/1BxiGtt6ElEeZMfsogWjYErpBXdHF2guUsgj/4rgeBonCcpo5C
y9An6yloJ0SXxjT155ZwbtlmlBC/FPLgke/k4/HYa7QwD93Q5pAgQgIbD+cgiubrSSzLFzBUJTt+
WeXtyS7BaKV4zNTcZ8d3iGHu6Zpb5i/zDshXekvCveO83EMt+uXqUiOhqvOEpnaOe7wfLpOsZoLj
idfUonATVDOdmbzGGVicBfHgYDGGLg9iBEo6woSCslig5sR5BI7Ljfw1EzlN+KCoaMcRhLKWr1lT
B5hRNPj3tyHz1zI+iXVcJbXXxMTz4JuIgh86hEd01//iqZlomtbY3U7XhukgaXlltRPmmXjK/Vvx
x01Zwaj1yrfEw62XzKgmb10JHPBS4sRtyUexNmn1FI67Ci0sBaV5Mbcg3jawUBFWOIJXRerouwCB
Sa+lPU2GREOk03vOk1h3pCKUHPXv1kRGKhHrHdPfypz9vMTuTJQ8U2apIEyOtG62FUuPwthTqyqm
Xr/DAeFLuGcJZFI5CC9df6jvZskvptGb+hPvghz1quBo/LqyFmNT2305GZXMDOIgtS0D6abFY8B5
IxkciDNg4oq+UV+knbLlCGA3viLF7qVrm4SHnt9FMxX5Cgru4ms3ydWmIL69PMRaN3naguE2TiTl
E5VZ4l0O+wO69/NBl8taX7ytycSzkhGewADpqrs8JMcsv+seQj6Ss2ubbpTkHo2rH7ESjlIdDE69
Ie46w3php4WuVIPidxwwmcn1/3w3VRrE3b4ZPz+Z/k9cEVVkt/DushlpH/T+4AAxWqYpMmQS72Ck
Ofd+HMQY0Sr5a5s6mgZeXt0SFMxmtiIig8zvrtoDRGh7lf2729RHLHb4ayRQ1iBX39ireLKxNLlf
u62JdzZmLPBWgqnc4KsDhAcmVg0Jy3Ox7ZFGQaadB5yd0TpKAhwooZchhHrhNvBpaXka8BdIuE5V
BNYkHflY55f9xdwoh0A9OrrRHc6H0u9oVcxDtE9qk+nFc8yOxJsjS3tfFIJAKq3v1Pz7dqR7/zk0
WYLjHR67Lh1q4w8TiS6vt/pYYAA6zdSnTrYBL6egBX971xETvwiOvnD3UOg1Nj5qUhpuZtPECO94
+BKl01a9ZIZYCVfV3BRRCsx/n7lJF8gJJhtKqyBDNLct3oinuw2u0y09IOYHhvAcn1xVl8oc1srb
dgaIHZNSKCoOrTsawWfF2hiDQuI2QE5t26JrLwtbx0IxGrGwX7yTgkc58ozaYb5FUvMJ4NxAsYIl
4PJ60A7zMs8/jRD84cDezy3AXlT7jHf2UeX8xY5tXSYwPO80KEUN2QYrpDj6DOC4Ua0orOl62Ekp
gIq+VMInqbdgtU6C2jXrRm5nN0uBjTTGWVmf1Hu5zHaXgdD/N0et6LBij1euJoA/P142K7t1QUaJ
O47+AlkEhGSqnML5wayuysEmfYIgqFzOY0HnLBESqj8wNJUyoHhdnzazrDsmmbmifSKO9ssra/h2
J0gCHl41RmFlxpiaP8S/TU/iZa55WlseJbdfqYqMbW5exrjNLAwzkGbIPzW4HUqybmpINTS2eYH0
Bb+LoTVJ511HzA3Ix85CcINxBnOyNXCpRAfaYlC8cCvEL0W5tPGMEXj+73mRuxwKrhGZ62LRkvYz
8d/UjebOYj7UAibMqJcrsDA9k7Y3gXTuQsU5U0F61DZIwcZMSMEWMpdG0TKk6fJYOFV8roZE1SSw
TGtKd2MGbjFJ+jCK29MixCTV/py2achc7NHTHTtDCTQiWcE9Yv6iF0RSBWpXmrQPEsjpO9B7imXZ
VJzJHj1TBpdM70EQ6N4eQb352we0Ub8/7MxEBov+0YIYMeWJA0dhzcgPo31g3kkeXE08P7nwcbVX
EeokU++d8cEcGY/BClvJMFJt9w0FdH2h41gLfFwxN7IZtRefSGLhabSnm4pHrfTfnw75Z+XCw9cI
K3FEFKRpbmDJZBVyhsFRaAYll77gBOjyejZ8FmlL6ZCFcC419JwgMYy2rjbnpqKHPwvsGtPY8wFp
lMRtO1I7Noh7xHlRhmfQ+JrJVxWVWRJjRTis58BoAWzSa+4HpQbqTWLDujvLN/8QPMmvF/EKghPn
a286WyMJr2KmnOmkCvOJWwEAU7t1w3CEGbYo1EuqDwJ7vp0CNfMefyeWZLDLpzqXOj+brHy6sKfV
XLQG8iXpIsSMsag4X9OhzgsQpSD7bDsFU/DwuE579L1+xm9OD4d+pgqaLcgcLO+6LG+ElH5Mikqh
I8H6KhVgWgp65VPw8kEiiHRfTbF0gfwHRZUy7SIKuex8VHLMvYwcEuRcfFRIKvXBCro1elpYJgq3
O4mt12ZKUC/efMPgLZgqaGZTkxHOCWj2IT6ZPV9WAgDV7bv/NuPzVR6Mz8H+p495qWfCzlludnly
094PqGlTaEZU61s7/cSlo8ZaAgaK5O0gTJtGFrvf1XNIgYdNpTdl4eA73PEzWBpBZIRajy2Zfpsf
kgmQLe1/SYEyXXQ2vj5RL2s7OD9v4zSrYaT0Zn65Bw831p8H5DF78JQsu5l7dSSB+Io+zQzVTo2U
SkuBRs0b/5XWmY6prBwM8KqDBzzouDOd3zzIVICfIEpOjCY9gF5teRby2ieRLSnH1celEoN5k+F/
EcuzD6Od2MKN7YqpSgDi3U+W1rjLdC/VFirbtdP33U6Fl8Jj2ido0l8kf1R7ajMaZfeQCURDY4i3
Nu55aWYLlSXDU+sIa3nyacLpuUGStz1RC72ah2+mtAQ1ctp3A4jzSnac9arC73BhRGq1cl2Abokd
xC56P7FVPoM+BMhSsET8D3D3PGypvXBUiIS9oUj4jcaUcCo0ETXytm86Rkvbj7xlMaZQvYK9y5N5
Xaq6+2MbDtT7JDKVPJp9FQVX1QWgglBu5Tc3uENApFyx6YRDiitPKheIXz1XYpsWO/V2LpDPsw6E
BLkvAMoNimCotbACoDELVOyS2q8BzRN81y2yiVKSHC2t4kA/z3dxOobBm93Z9s0IjfjXtg8FEqG4
/iBwWKRBpi+1sDx61yLuSwACJHej346Da6X5P48FkBRhBRZ5bQXl9erQgZ6yh5sGq2uVj7vhc+3M
D72V5mNlKMTqYPCWs4i3rNpnmLjQgA7AUKz6roTsUQ1Q3Hh+h5fw1ya1xF/C7r77Oq/1GqGV7PL8
qAqLw64I9w4UoxYNlRrPXSW91pN+QKqtvrSLT9+OgzHPnqazNuASGjFrZ02orsbEouJblIUzR2cN
KJ9xzSezp893RQ/9ksoTofJu6poWP0gpQXKJ8kRpukpuky/NR6chiZ05FHetMKZBdGNi5fcF2wj8
fZ7IODf5T42iUYaSBtj6mywxEaCv8Dwfr8VBMmDvdCTlzaqnZvQT/sTo3PsGI5+TARfbdfLAdC9c
eomFHwD0dhGpVVrylrNGVENtWx14uG6Q3Fb0RYU+/DV2QMp4Q8I+GxgyCoJGH28vOEFdkbDUc9Eu
sijzUmvvmSbJj6f4kE2+0/0QiiG9k6quJQY0fUwXPNfW/Obr9jupaMr/2AMTFUgFGskzw3oglLuM
1hxaHaPwDHD1e07Bysk17QFjlqTmRZPNB/IBSRQGMtdfYtGqSeh7XC74aaMpz13gB3X5tLhj7tp8
eGl1VnLPV1WYz61fGPWupqYQDhnSqh4e9nPgPkiWM6X61/5bEor0wjG8iutnpWEAoD8rsWLqe2Y5
iyO3nqcyEvo75bLngo5hmsuUSx/5yFbjYy3OHKNloYJP5cYKzdDQo4QoewEbPzwJgCVoFT4aUXAN
2RXQ8IAbpimtGW48KqZkGCD2KGmAEGh76SirkCSumWWKbK7kJNdqjMkzXnqiUWrprie23C1TRE3d
UDe54X76+ziPCueVOMzB7a0xUxwLF/NGYwndV/FxR56At/yDi1yhGkoEUppYY1ATXhD78IDeItkJ
wyIHHVVYAsHv59aO0zPC89Bo9YOdCu3nn9nVmSTXNTccXG6luuICi1GzFJ27L9kGyi5MZxqRRCDp
xru24X6n6tb76OYpUzhvZRX/Dl7qo7VZCP4gKQuj/LH1JxeeZsQMrwHV9yf1YpiqSAUo0L/XxOHD
DN0EzIbUJgCfs/MsznpdtiTRFoLDR2wH4xfOAqxLEO7rwrkjAJHCNLKrn+XOZz76wKm1hFf3IqFq
DUBW1Mtvpn+CrQOlQRjZZrZaXO1k7qzB1NSLPGqBKAYz1mH3x4GQunjCbBjOBJflTkkp0pF1R2vN
LHxciNw1S9P37j8Z1So7nMFcB2XigXNdSFISQKJD6zm6XmTTTFQ77f8dUhSyS7xYA6Xz5p6dd9Lv
ocE+FxfuquUnxucCTLI6KSJehQURagWSVgpn11KGfanU9Nheu/LPenncSjzo+vdZEKxre/ygYLOb
G0T2eTrKtKQvUGLlo2OnKmqZkF6JYASM1tuvGXTidaFNaLQgrxyWWeAL2v0fFEEvmbcmcSpttH8J
BAB2ECsh6wFnhJIF69bSHke6vqcoXHQdgErCHrB8VqiydFIXwtJcyOKutqILyh4KUeXHC2aXVInf
66vOVABXysfpumgiWFz6Do307QqvOJp01sGRW0XhZIpGmhsceDO52dK+a9nf2tPg66PNn7ltcCUe
JPVl04h4GeWAix5P0OiAGIHVwlG14MXA4bMUdca+AosQh16B0zk41rWYKTG2R2D2FtDQpXgBQTsJ
uS1WP9hdy6f5nS3mptxGPNbJQq4X3opkqgid8qP0Txlb42+7pcxK823lKdhKFHieIhZpD8onwdte
Gx2rRwmR1dt/T/lZAVVUEgGa2yM8zGCTUs0IZt7ylsqwUYAv0+4L1jcrw54AW8opP0NvxykHXiRY
PyAXq+b9xTCzEk2x59Y2MERrZsaVYup6Mq6A5ab1AZN7HHiw3utZC1LXRel3aNonXHTzd/S82D7v
rYEItfdrRqyDIDiI/AvLvlt0KvnA8FcxGFR71kAtv2LvPh3BL1EEdtumGEkYbuCEKeFjJRMH7EvL
8SbMGveeDvbu0rSChDeY2F0rG0y/Ag0JzP4Fl/DbSq1dHXGbZMZcmbqAemu7iqPIqdjjSA29ntdL
pXkISm7zsRI8wn2oWlm9P1AlpgVc3/5Bbin0AnypZENkhvrdmzpS3ZBnNNlFYNyPVML+pcB7L6VI
BUVMyOw1wZiwj71DxaPKup93M0AFxasVq9yuo0OZKwNUW5mdWfbfDX8XeBo/Evi/DyNlQ3T1FgFn
hplq3LC99IG1KC6pImCUCDeSAFTG9OU0h2repcrKtGPQ6hynvxNgaQGPRLRVArHgAbzCBbq9KzcD
KDofXF44BK5zX/NgNDECUnMRc4QP8oM4i1sIOFoIMOk36BDWDywBi9HGU85+LpqBELQk49ZZMsZU
DtvXW6kQaD1a1lOcVlD3wMo5qy2Koo4t6BBhU6wedVpDJ4/wjZcv0Zt3ECsri0Q7G8QOlqns4RbS
5lLbuffL+q2ocJ3ODA5WsRjjlPS8tXYN+CqqW745SQd4VmdYGaN25AMNH7O2B2lF484gDoZdB4DR
7+whglYiJJh1KQQuncjXu8lGK94GzdZcCFQeeZMtXag41lqDY9VF1tgbwaos++vDVBFiyNooLTyQ
OaORMqvtSvcclPaPssy6qm0H2qgY3TrCFN3c9MSEIZzUZxZ6mZHdWhab7AfHrcEHqKkF7nUcyLZ2
zp1uvBHbWEXHMxt0uiWrveDbMm6SLEUXmTqIwwzUHfW7syK6E4Wxa8CAqt5r2+LwErwuXNypYFif
apB6yUNVg1DpOWpNu4GM3FCDsdDaG9AvAwMXIncDNsH9OgkWSbo89Uimj7sCdc1yLqzuG33t+Hu6
PqHysm/yOPSmC8dm4A7PtsUn7TCU4srL3n81jCNQeQMaesZ8reWGOVYQd85B4C1SOZ0j9myVXkGJ
SnnCEVsC4yQ/1bQl5Yhknq55IWeVAFys0Jpshpq7jKtcs/r1yNM1yavpnNxMFiPZmYvFW1Svsrlt
Nt3Yii6pp5puivMF6qMlk5Ox/v24mxxE6G5azjV92cw2KKlEA3EdwINF5Ho4X1EHCsJWCLAVm13C
ooyMqv10RhPnuwTfIo1JxqdtvF6KSKq19Toh3+mPxz4pxA08rp2MZo3FNIpYxDtzc+gM2BRUiWN3
nS7xi3q/flzNqyG3h54YTeBIEQAW1ZuWz5O8yOA/1tsyM/td2LMvhEt8T6qbd9L/muW7IH1obB4b
hP/X2zUo+zhW5Ey9gMC+STctVpXx4cesVc/S343nXrkp1+tqhLcLaUBPdDQ1skM59zJW6ZeynuiS
Kd69fCtX5yzVsKU7lw7pb45nTuBLjxx7YvPmkdJNNUCFNhfMhNZYpN5iDT6BrRpo0i219RlcfwTJ
uNRkuRj+Aj+ItDp/kKwTWXYkBZTHZ1UQmfOj1XC1nzv1PhG0zVyr1CzzkVJorvSUQk76dslvrnkt
llRTmAaPwal5BsDs4m94W7e/RqQ7Yxsy/ElxbFeKu/Dc9r1wua/izXmrfi98K+63E5EUpFwprMG4
sAVlLPyd4piTa+Zf5jkYQ6aO0xMnkOiIqfpAN+8UUAZCcaEJqsZJGtdd03mPiZozoc5pgqUBkNwg
UVJzJqVG9EgeasW8OS9LsH/Ua5aT9XYqjH2PEjoqUz1gQRe/mv2XI2vYH1B1Elu8/CcRqZ1kNguZ
dudVyS2kzIdXRx0JAOdJz7d3bHymZ0X6mrIWKnp/V2aiPVL+1oL9TDIGee9PaJrzSe6CDf/ZaL/U
l10s4oAJKmAucH6L+Ax4sPnRmOr1h6CLVGeO51HcxiCMRVVLdN4z3Nc0UbkHmBN4DKLvwhfQf4Pu
4Iy+/K2GDtbXJZ3KuK7ota+3ELRM72HSlHYEmkH+3qWW8K39QHGh68oLGDiruwuCTye5yPH1daGN
Eq4Au28NvjkB5yqnbR5oiW+bDNqZC39w97A1YefVJYZoWo4+y5POLZpu+L/Sn5Z8CadmxUA4+i6Y
Swzf76HlijhtqveNGwgCIXWMYsG7cdggs5zkDtFZcVv2luv40LJLqjqSadnNFesZW6kLbBbMiJgw
qe97JedAEkRFak5R1SCVUmkSQM+tGrcdf9lbRuxG79szBakwy5YohNs2YbDvz3P776Rrna0cBsGW
YD70BvLzxgmLQl+PJEejaohxnjNHpcddTGrgJuvl75Lsr7Ny7jkkfXRABTre0NmHeD7d++jZPmBk
iGiVQ3p6ksxibh17emhtHDqAVzg7rwBysd03r1jb80aUnAqWpW64vZI9zlF/9NcnYhy0yvIMq7dX
XYKD+ZzmXIUvAFDF8w8rp6PEt4yj+dUg11473y/xx7OoJo389FojlOO6dFCuV+WbPi8ZRBn45h1q
ps+7GpaAiXxZwxqaHrog+SDu3KsZhHXS6BamP1F25kYVkpYSQvaZKbZtmfSefwkTtf2FSWx73haB
90N0fjtZVAn3Gu1Eq7pUQBcqc2zFQQ6hZM58Qns/nqAOKids0Cm+XvAK6WKROJ0hwpaKULDClZIW
xVkPC/vRxdyrr0UxXwCTIKW/VvupructTrhPjHTjQQY8cQd1hl9SDByJ/kQgVRPbqurnaY1Oq28h
xVtOTTKgj8wwhXUObsXpwFa7qSLDt1OOHPkk6XnZujq7xJfuNnYXFWMlCE4fzxzRYyPxYaIkKKRI
5t6z8tVYRPWSCB11RWNTZGICwbvtIvRDpZZrvZlfpvA1mE8bQfcf9JfH8Xj7dU7gbOml1T6YoQ+A
Syg+AiLcCW5TEzMKWOf8oA6UC6oU2bgyGGrIlnMVpYZnS52AusD3PluVPpzYA4NmxFT2MgHwgbIC
5jW1JM0S9F/WgWlhQehxO93qeHAcz30pipnaG2llYviERAixKaIlvBfI+uOCZbiOXit9Jk6Yg9h+
QW0OgNOhCTbgJvRU3dcGsZq9EETUnPZ8WnIRHRZUNLMWXcuW94EYj/+qYviDYQSSCySrtxvqGWp9
UHZqUsLGsnKOS7vnnDVZAto7SxJdVh24NwiJdzmfWHgeY4VHPPgq9xuuydlySrVqpqqsB4G1ReK5
ImPSxCgOYvEA08ZwCQvpic4bhkYivfKo6wXK1LcJ+S799TnVfqekbjnmPhQh24E6/v69VQu/889V
M4UYrYvkyF/149g1C6NSrgm2fLQ7TgYad7XADDrabfMLzo0PJ+Fp9lfb7ixFmRPcQi5WR9mvyhId
0oIy5sUjptJBRUfDfq6O6aCxcRYpLqLAe64ISn/wDPad2E9E+kRqig5QNRMr2BuvvVeroFwKCmQo
3kvOVfoliWr4UTEwEk9K7qwM+J5QHt5TfGxLdnmxPhF7sDRAxatAM11US73rVIxfSyjU2J9YTcWx
maeQJKAj1HixxwxRkeyyTKbwnGRRfuo1C/Z79rzjBxehmTtvJkBDZGVsrBRpnfXuq3O+FonXpCH+
Nx4PN3aHgBtCl7AD+Pk1VAxqheJ21o9oQgaPmo2lywpw6Lu/0zAEGOoiEaew3w/vWJypcBkTgFD9
a+fxVDoHP8w2QIhIDoqQu/R8iLUQEi20lJu2ww5vdwzPHFaxTzmKE8hfzS0sIOu2zux5KtdAargi
dQZwSlBGzNXgeYH8FUe+i7TVfB+2c2G+MdaI6WyA2+g1TFdoUhjE1zQjw8y/DC9U43Scml1lDTAE
qgJaXVLszSsDw/6jLoUXue4Q81Infm5bfvjd7V+Y4nnuLXS5OEpUqmx82lmRZ4RWieC9fgQZBE9R
umqWkUbU9p7gqpd1rL+Mrx+Duc7d+EUsP10Biz42+KgYKk0k40KlrFFr32AqHrnu0NHmOIDvg+IL
04rn1a//blsuRxwKvhHm7XvaTyWWJIuj96V/CseB4kDQc2sJmcv0y3ms6Xc35NT/1kvCaT1ITMcU
ST986uhltjCRArN/6orGF9MMOQe8TxOBNsXx89OMBSzlUfAZud9B6zDFxyXtZhfgH6Kro8CikZnT
TAnss4kjqXHIjKDNgSRWrVTz8aIetEgvK/aWxgfznmisnqYqOUkcNVDtkeobDwWE5/PUB24vOsBm
HKIn5Vxwrkcsaf2wGhrhLGRz/JTFheRj1Pk1O/qBNFbI56OxBS2pUl3ii/WsTkr9nkKslgfqQI98
DV4IvbhVrA7vLxZ/VB7Yic6cQb8Ye1wsWRj1OtNPXWuHFuOznp5lON3ePxKjIFKf77Zg/whfHZy4
6KAN2hre5cxWG+gNoBPK1a9Jk09ZgP4sGniqBVyeW1fti2vQAxxCRptiTscbWZmsBxquSFbYfI/K
L61p0D0l/XoXuqXv2DW/HzyiMArSRE5/w/m7YTjhs/aNCETj/Vg8z4pMxaN6s61DVMhHkrHSGxk1
Cd1KqSz1IJINilAZXuzmT/LH/5lhGV1QtAlXkhJYEkwiB4fgxz+4zHQgwEvEhuS4DYgL0aN8HaAj
2VkJWn5PqkEfclpjGB16THzP7UqWsOdmW/DXzId7UW9/Lu4YotiEEDXiEWy8Vn9jZ4jn3M0lBiyt
ZS3g6yG3V6qnSqbgghSIoFfA5u423jSmnp4ZQHzoK7mlL+e9bS71zkOX+9itFWKIb8imtVNqkQDB
xxwIox0XANRE4NmZTI9kVHumsZl4PIuAsw+8oWWUvp0vYAl0cS4MIVBZcaTDU1jojU1AWUQZnmdB
DH3OoXz5oIB0fGdGBShfAwAuCcfERvDAwBRoVlMREgCOX4cP+kbfe0pfheXaT7oSTx8a1cAKk3gD
vO7nuA7Rd65HQzuoBav1CNlAjg8aze16g1LUUMC+m6BsSGgwr/gBPWXIAj1B4hXn8IlQm/gPpiLk
n8myZqLYdkhdBukZZMZQqleWUqDbEZCBG7IQTARIeLWRcFeiztNqrmypqCAgeH1L5jHb0USpcTj+
cwdJiZ+Cil+3wWtpVN6gya9O0GU0HH1OKoLzBQdsTFpN4Rx1lf5p2f2Pfoj77uil9k4YA3l1DmnJ
unoi5gxqhj04K6T2r5zoozzhe7fFB3ZZ7WiNY+J9Q/L4nBuf0J3wE4cFSExP/eyIAb5XMhfVe75T
Fk/GLvu6m/j1cNcM6PRArGIyOikEP+yAITNzkI5EqiWHyOQ0dXAsqxHBroUUhao4SAt8RVutCL/B
1tkLKfXi6///DuzEm49cq+TebhVOQW2z8rGf5l7+wpjJEWu1YDhHtE79SCg1gEQ5gzi9YX964UHI
/zJxfSIUsShCGjOBle8xt8zqq40ydS9w4qbQqQMLD2iMPkERTS35DHG8Pq6qUyiHRsWVfnLQ2qs7
GVchHJSFawZ7cwykY2rtdjnQnV2hbKWKc6MBhN+0VIQIRAdYmzgaiPvkDqdDwizj8Ii83+t1xhkS
6oxuWtoB8YGOA8dLfizSmkT3wm2bfYBNTLhD9gD+gZvMZAQ7qQ5z9GlkSo63ghBPolcbem4qruQ7
s752W+1uvHl8LcO3Eoglnwh/8mzaVytg/Flu/q2XaBl5fHSkgumrGmjHeQL7OQOCX76A8mwsISlE
MOEcIjuKsDPbjiO1ajrr6tCIXSD6D4i5ATBUsA57TCcb+fUFC/4AcjT1Zb0r0nCSEPEmAQn6Rgbi
QT87P//EU0J/JAQoqj5tjtaVMHO3qDKTPpt4wFJYNoeiTP6XDnN+xnfqfIFOu2lBdjGYXqseXzQc
hU5qsHTs5ZJvqXkCkCpNOo3EuiayLwILoMLQZSlnqRqMWwDHWu4SmIbukstd+ObQnpIQwl5hh3LK
1Rqx0Reyntcktp9V7Z6YX0eDOXGS3D6QTSHmQnar00fu+ALMY4RgN8GXzRvwgJmgYUfx19SSLyWf
VsmJdNW7p/J+gCwwodwggybv8ulsOzzTbTq18lZJYvG2RpuUR+FWNH/i9xE1XR45PBN2zttC/F04
7Qotm0kBZmdzQHNbdqq9HdqB3dWnEXJycayeR6LI6sD31VPCvo6013YTUkMkdCT0XJTo25m1sNhN
Ynbv1T43Noj6E/3PKbyJQsKp/6Edz7IuJVW7HDiSJQWv3nNvNf6WU5D5bs3UF0H05EYMV9MVFTTu
DPJiW763Y93SnYqUuAuhzP6pqpyVeShdUXAoa8LaMMtGx4A6arx5YgZqNtlc3DUoa56oVcRjzBhw
0DQW6bZE3Wgs6czv/E9SIc3/0abFoewwo4iwMijzxGHOFMzgiCzT7rJoosyuIl4WC1w6An/WcTs3
9RpQavQ1xkRCAkxds1gbhnLY6gzlkbUPd5xyNGuxvJRrKMmERTu9Cq+yL1YxEse+eJR9Um/OwlrO
IgFLBxQ12I74lkLFgrTB7OuafPcwkS0FZaBX7iI81XEuLIryC/gt81gtFyhmbh+Bc6cWlicR9S2W
o3wEzNr9KO7RAxOzf8a6aP8wnkUloljCVmJ++L2Pj1u+hL7mY0q0i44aSIEKf7p/xhiv/lLMjFxe
4tItYsraLGot+6SGgWaZNdnNJG8qW4ofugKHcgLsBNzBtIVqfNywapq6sAnwt8XAc1+cDY3Xb8WN
ZzDXxv0Of+5NYBO0Uz0oHseq3wHajsPu+VPbI9nb8Q+gnZzrJgPOlHMCsQ1y1DmiWSZFY4esRGvX
DZu55Lma0jN/add0EbmajpCJ8VDUzTMsaryoveTimGozTgaxCj5rNWEURH8zL9buD9Y4SU2jSa7Z
mCe/s0J/ILJiz4yN/9ftI/37z1Ye6f4rsLmWRzMClPnliIP0dLzdawevlo22a9JBrYBE+U8dSXdQ
OgG89abXcvJrA2t26DV1YF9UL+9ly/DuZO41fkG400UPKtPxDnY8NoKONRXClHPftEU/ff876B66
WdMxeNF0KjikFNN8pW/zJH3U+uFDf4UQnIhIzy4I+YhXx7b7TtONULIW+xL3hXj7YjU5oP0nkzq+
cEKvsHdw3lTRvYrGXaio5SxTY+zDYSDfs9Y1VuoYlQBhKXhFNYe/VmtpeDUq8iPXeCcVeEOWyqL+
ZZBYxPav7aMTKWj19/oDspxKq66da+j/e7QSqYSXzIM0oHJKAq1UZXcPp30EUtmhCJpqEC9P050d
8PDo+9CsIBq8UZTf1qKC8yVbIvfM8MTtNp63zZKBlbdF/wVUW2uoFadkDSgR5oxhMSfjUVqXUMd8
mp8yvOqE02GI8IBU6/i4UEZVrUTF2lkoGcyucSRNh66kmCfG9QM42NGUndelIeF/5Ys5Yfd2Gk1n
GGEALZqaSG/8vurrTJAqoUFWXPGsCAaDzZEGp2EhQPVVaAt1bQbrsNzqNyoIZi07VPOPfwtCP5vd
5tQ53JDKeilIkMGrr2Koq/Sm4Rgrr+O4Il2hSey9kVZMDy5ILNTCY9hH0/+oSgQ3HP050+v4xRBd
5K3VmSoWkv+Rx8WiKGxzaVQwBowRKm4Q7ndgbTWxUIlsuMt/yCX0zi9N0k7Vfryg3BIFiTee3ake
X9hNz5h/TCrKXUuYQjBg50Q4FLtcuIdNo/Gsb2B85BsyThZl3UlkitVgvO8j28+0cj8dgS6FW8jF
mVpTwRW37jhADKfsURtkUtkcRJEkYyTeUJZLh3ymRWMTUBbd0xD3hbAmrsLJJo5P8/5sVv0AFuls
d6cfgRFApO2IGFCVh8UV54oi89XEpmE1x2TSE4aCjjktSXWtq6zXbJdH90i7ixunwtLFIwOVeecp
UZdv43eiVza2FxIxwdzZS/VCh3VPmVTIbh8dL7pXs2qI25KUq9vCIemTUwHRh+FLgC3iPwUekD2x
jOjYQznhNJZ751kx7XHVzIABJ4pkdw/UtEF96UcDLhPk53tzgTZBc7APf8bn807bcmRowGWbxXOe
vWRbr+DRABydSffZuXuqA9n4UwNW6L10slh0JtOdwnhLYCotUVZQXnrV79TOJ0UkYP4w2fAZ26jR
23O+wWPclrg1CSaBbfFqnV5HQZqi9Lxj/ljSYL7P5uaNhQP/QQNvmEwY+m43TvV7gHA1dp1oudcC
idFouz8qNSjGL2IUUEr4+6qckKmG+sfdlxs81yenRWIuDwVMYhcuiBEOjZ82YUdBUB/HFHDEGCgQ
fY44dKrbbZHcNYtTyvtdtm7vs90cQQ5TCb8qjF5TvukE2srKJlstRjPyrGbP/Y6PHCH4Rf+hIU6C
xhrR4Q6XVzBujsm9wt8jnLwcOgvolqZEjk8iZXxYkjKVlds736ZG7yssCIX5n5W33H3U2jN1+lkE
S23zlHUBZeopd+o6vu6NieFy264+9uqmrUTT8hjOnY75zyz0KUQqgUpkujOZwCaVTj4AopRuS2jr
YpcS15JGnIUZi7WiEQGeufk82BQlgt/SR+WUM6LLcWzBlgvZ3nI1vS7u6gOcktXGst5LEs8WPFKm
/7jrr/0smV4xyOW+2r9RBlqPCDaz+qsGL20ZhlDlUDhnkGmjANzrOLLJlI7ChukRVeWySwDnsUnS
fZjcVZHPeizKd6rc76zoybm/tIG3vL+jr6r362FoY+bHY8BrzXzxL5dp0DgSZpgeqnB2HrOpDihN
7N26V9g5Cl+Stw5rJSOtPLWs/2dsmOVzg5cOTJnhiZvlJKM9VOVQDdtuvlPpFD2s9GKSvo6CVjii
DQ0hISvlOoVy/NfCygcNBscM5ywU/tUNQQWOJ9ufSulRjR+83D+0aFiMusObqUWAQt1cmBJB+Hfv
ubY9xiY41OfR5RAJ+9Dezn2J5Fput+RLWWo0oAWTwwKDVZtlviasslwZ2m11bJGRvSzu86V3p18E
A9wbm6w13U0Iv8sw3no+lg9Nigh5tX4gJ+TRprv5XE+l71/RshosuDYXrSmsYUiGDilnjSFRGzQU
INXY3ig3vFtAw7FGXFaL8Hp8hDLoRDZ5iRo1iEcTW9nUD9Sgb1Q42lhKB/JZwL3TYB4jiiUOtnk0
OrONGXka8eOr67/pP3ml52B0GVzdRmHI5aIPEHn4LpJNXSAOYdfTwI51i7uGf+UAJoaJM6blMJBW
uJoyFgiFUT7F3mhVGlZTKHOEZBj1lVI2RMJrd5pSqz1RUbCSO1w/p7BkMO0UJauV5zjf6OKSiSwE
YEI6V/V3mMgx9g68zxCmK7d56Pg/FtDXNPtadKjUevNrB3j2mWZs0fpm+fp/Bl8dyjY7tIxEFM/6
A3KCjRVFm8fb+V62FXVP1Wcdg7G0wVurGJ902WKNMRHFTQP4mciQPKZ9vb3yXHyq1F21s34PaftD
egSWEtSIulbav3AUuAv5CLO4mxhj3LN7InqAqZF9xU+c7HDyxnM4NLlWOhlsrUIA4YIqPRVpnzFG
gxwQYDishObPl5X/4yA6dBffWa4fA0y9zPFfU/DH8/YI26Lqz2751vG1J7GOx1WDd8lHn0EMezKK
I6Nn4L2wVr+AJMw9kqPvKMNGPxpZVoQd3eXq8mp3LclXMbiHS+xBOfczDo5vJQQqsD4eDZ4ujlR5
7UXa0KplH4GDu8NqgSAfO34Svi2+Xd2teVb/9jwxPlzp0m42Ue4pDMcl1kdnl9vB7XxYbfeUogbF
zl8v2JggPr4bV+Tp09fy5l7kl+GeHoLVW7r1S+t0nohY8DGCH1CC0Ny9n1/LYtM96rrXtWxwQV1t
iq+wascS6DOzyqsYq/S5KaCMgEtv6pNRjXOUAur5P1yUCYpEKRgQu9ArT35Seg5BRQIqNych9JEH
8ZbTTWIZDKO1DZmeQdWqbjOLVFB0R5c7Jrmeng+60GpwohRH0FMrakB40bbFt4o1O7ctpqUgqaI1
HKk4i0XbOrGHuU9b2PMe2tfWN5WRMHPdgSml9hDWTeLRLTDzSCH81SgpKpYT0nF+i9MiDqlbpsLf
DOSmwIKZprPZa+YS92Wwq/wIU3u0IR+JcSShytDhJF1BBHuX1UrGYVrMDwgaOdwf/+tnqJUTu+RG
ME5d0wKPO5Q+6/biEmkO4jJ7YTHz3lZEZbwfo2VySALV1NRLd8zsLzeBR3mHITlTI2938cnjiKK9
7Am3PjgyHE1Q5AXsYfWMx16pDUnzCFveGnpTaNdnNvQnP9CVlYXelgG9grh8SWYqB6Namnk73r4f
o8DBlrtm13hhga1YbK/e4FAnouCSPqmvNTh/gYh5E+VZK131oTDNv6gHIbEVv+DDcqnyqRGpWZeW
FBmIKszr6JccShY6G29EtWXSpgIBjxCgQ5xPhUdfuBX59XZMlE9xc4mwEWtOwTlO6EZa0L+OkuDq
VOB4fyZsBQB09eRHpVfmJfswOP8wFhp/szYqIUXW7VRlK7kktmOb0PsrBmMw7ZhxYuAhTB+cPsSp
3S0dhi2K8g2ARjHHczZ1664KIeBOgfHeCEgV8wD7c4Wd0e9dbf0HzJQx46tJkrQl7GC9uAWFpx7j
HNpA4AlAj9RlyjzMBtX4sZ5Pwv7KqdxCITN2qEUs/Vb6YWvXuEB11jC7wMvj2VlKJ9nPfqoUGqBh
l6LqYViNjosAOk0XO60fhKFPdlxhXOsdZyw2ib+5sjs3fwa08SzTDyLnfuof1uHFNMnn0n3Yoz/X
RJIXp5wf3536jwiGocmJb3sm3D5ufN8WGAldX57g9F7xC+ohGSVPfXk9czlJt2wkFWN/9VAqKAdp
67utZ83IoT0ls+TU1FaBhx0xMfun0cIx79gygc1HVwvLUxAYcsnIKA1Gytlbo9sQfx2LTuCN+Bvz
p/LAcT4A4cdjA2jBSSPw/1ZbP5OJweKyDtuj0hy1kN5hNJhZhcF3Hgc6u9C4GGnkrYFeT7e0NXHr
8GNG07SGq3LBHQtrJ9/V2xbe+4FC9ZxQ5oJGW6JkKcdWRzT4JHTCNM84ZLXRPZ0motkVyC5D7Gbv
vAFnlMe4Jm9HXVMF7CdSBKY9Vp/+08e+8gj0PrJxHW5HlwzeXvSSW3Nu09OTm3Cj7nz0fOThNd/i
QFrXBKRDWshRNYPlXBiRHz4h1RtYM9IIQBuEh0qFvRSywAOIxbrRZ1Ui0wAvOC+Fy/qe2JQa/EH8
gaG/YW9PNB8st/OgiMscHICICL/Ay/xWfsajZudHFwhcXVlf2ksEtjv0rF786DNQXgCnycIEvKMy
06A1vEzR3CXZHAl/6x7erCm2r+lTMe+pYtPzfixWIzUqARnSF0SDQnLW9aC9XtU4mVymJ9PjokW6
Rbhf7rvfiDW7amjI3aBticCvskw5L5PCOmDE+As7wXqwd76h3qtZVtdGyBygiMJJpQwVdX9rvZI9
9fUyoSx5t97dm2dHp38wheRKZ0128P2i44IMcTyIKeoVy7E427ymZ2ix50/nmCvf2AFaU7vVFRyk
4iC6UORw8rK6oyVk3hf27rrcTRq4k5lO49y+eG43S35OstZeVA7Ityuia0/STUVpui5uuWGoFkU7
G1r8SSGrj5s69309zaqTfXu2scQwl6PEoxKEllBtq6nlauXdWXah6pLu+SbHPwf/WQYOygUnuooC
UAGzc52MZINPf7BAfbx/fHqdyh5QZp+sNJHapGjIS/PnzF6rmx/fHYZA+V/fwBT2MCEXZC4dpgy8
4hpl6YA1uscTjKVkWz+2emsr93N5SGkIchXf/6KuL+b8wCdCpErG/q38NgIRZ9Y54EaOFfBfYSVn
FlMyL0SLFJdO9sGDHvAHhiNra4KRUlOq3ROcXk6XOMpTEVBB89W1kSkX3XwbDubdL0wvFHhy/oDx
M4StZz353KQ0+M+gm4GtGD3OprNCRZWhLw/XkzIl9Dv+R+XHUjBdJvB0QKLsE0DAtqYwuWJ4BrxH
pNhU8/o+BauiUrygpPkC9nhLn2Byq7grwUDKPv79sMb3mL4zCcQEHeNc27IrgLhuJEGfArWtwYxy
YpYWeBZfremObufIp3v0b8ya0BWoGjMJDGCDiU+zZjzkH0yc5XBqRLbuQMfEAAayx+StZzjLR06y
HCyaPRN3Q1pjZu6YZphywwShrh9WaBuQ2dWC3wM7UFXvFpencPPo8qCuJvYPMlLo5hi8ILqcl3XV
7wrKVOVGItk41dMvzgHstFiQEUyMxLv8K2tCl7LXb1BHjemb4cKkpREMONbKwy3J5M0vbYlUU3NM
gmcywP8KugTcMlgbX+t9+2QnqbICJPSbaqo5LikIh9Cll6w0/GuVGHBGxLLXOAmOR9PtsjaQNRls
vUQVEL1uDYloVIzp+K1i8ytpbJV8758TcHAofFv2RAj+jErECBnl5KDgudpJ5Pv31r/bi+JLif2t
BWrDBoFaiab0lXctski1A6DSgJplnuXoZWftitQKCnRruT7uXZRlL1+lVZ5pOkYLTpcmsBw9b8LH
OKXsewfcVglY6/3NUj7c7ovwbEjeJ93TkjYs3c77UMAEIFbheiZ6BHNSGHyaVrDleBsBpcbZards
A+RMT/LCkbmX5w+FKlm0ndCkFcI56TyJZcRjdNj7t7oagRm3oLUAhJ8iUDKpI7mxGzywZ9ca6oMr
gCHzJTsoFF3PoIiDTUWPv591smYZ2S7Em86ipW8X3D1n1K0BgWIthomEKN1DdDepC70WdITAlZGW
YtZtRPIosLfq3f7aD+/jy2oTQFbp3tzy84zygUu6UR421ys2H/yYFVUPmRU+My24DIlNdEzCGEXH
zcuG+ge5DKAiq+GdN2+tLlKtmu+bqPWtF8bRNemuF12/Kd+1r2gx4014TRbnN/QzQnfNr5ocIILD
ZJ9vzdTZdDWSOu+SKD1fKAMKjimBsLi4ro+TVn0iBWZVpC5ApptE/ksDTVJMVxtFwoE+o3IshGcr
g5G/bJfTS2mm4f+9eubZlVg2SragyPFcbXuynw3+nB/Bz9ik+nO3DMqpqVq3m4+hgBiYyvc7sL49
hbtHU1X6Xh+U9+Kg63UThaEqjjYxyxf0hpIUo2VmxdFVlNnrYNDTQA4Dc6duBnH62QdZeku0R26C
p2+BUP9t6Oa9jSwsDZNx4WZY3QrRUA5+y0SZpiztVm+78BHLAZhqIrWTu2nCCH47c+X78gv6rAra
m+N2SACMniALRNfqTexgNipyZTA2Noy7I8lEJvX0P/biDN2F8RK8jFlJZNWld7fMd0+GsoOKgy1c
Hqm307FOUbimQvCa0XnTA6dhCsZ+Ae4ip3XZRNjFut0DnNcZloiF8L3FPNVLkAjewR5ZSQSeA3vc
SODFPkrfbfOn+Ppnf27lCwkuZMkFUdQQkwP91Np6hCap6quYrQ4AMjJJxEe9Y+A9xtM9H9DVbr26
CpReSsF1JrezgFVwVINs/5S0d4pIWqfEtZpmXHEF7NcPOSwLzL0tkzkNZ+QYr1e5LhatzwrdWUwn
HbGek+rOvAO3K0xCWSQCQ1jSGGt9CFLydjwQnMKqJCXD0NtReusqGI7VrgXvERqR4Rdv9Sys/1EI
VQpAgCl2koEcCZZXlUYSdggtEpU+hiVkvSLce5ICXSTQndvnWfIoJlYHb8g6IV9GaHTXj4vJPcZG
zDgYcN+zOdYehFZ6tmZco2lfj2uVbiyyzCc/s4oaSRr3AyiKKxPNMuKHHwsHZ64uRl8rJmdTggc5
SeG6g9UajlV4DqkHwoqtV/PEHgyHjf9mH5QF5SW6WC4o9o3aIKKnxugUFeyJDfJ0kJdr+KhHwmte
qBZ0S3i+YsPbjB8vYO+dwTO4zbbk9EMPEU0T0qwtEF4gVN9JUMoHFBU1ejN6oaBNP7bMeBHwQ4rN
NPuhXbbT+ty72o8hcBMFSVi6cOKYDYRBOZ7xjli4NIl0CWTHMmUjsSqGbcnVfizTS7sEYE7m5oGs
74QFzWq4kAg/Rx4I74MyhV+mqWMPCwRt7hCZlI2UbhxIwxNWDQKWpBtB3S86ngqqt36MX2QwNC13
mLNvEcLaDgT1GLfGhFaOaWoEwncodJBnQ1EnSg1+MvlE3bk1KW+SkUvPLVFTNgUnwmjvcRppcfVi
u12ibieRT8HOG7fy8Tas0IdtaxxCFWqLWMk3xROTBtUCuEG83rCK9kWFiCRSeU+lVkMI3pUDH3hL
JwSvUAt2IrF0vNhG8ZOPHM7a+nwmjuA8O4nUEL80loC26V50y09vs9mrW8J1CZnxvEZjesw8mQx2
vHklP74BkjOYbCzCWM43qmatU+4Z8gpZm1qvkbri0JioDXuNP5ZCYKHYE6YRs8GajoodMb2zj9ha
md/kCOat2OiXj3h/bOC3kXYliuC+m3XOW4iveO/nF4TwdP8GI73jrkJc04q422DW61Lqf12Q2HqU
VIDGCm2J43HmF/rP49iUEYgft8Y3+r9d4nXoSqa+F7bf0wA1yxohT6MAurudLeb57pV3ePcEt8Ue
gTsAIhB4jq02NTiXpMaijcgjJ4eoTGrKyGkMrpgnO1+2uHkezXRYycGeUclevMuytDydP0q9Ug+p
H681PGzKFKjYIRNdAGMxvQEIRh4uyOVi/QtX+Gg8kj0nHatBcMzK5mswsxL4uLgs6N4cvC6pPq1u
+LkkUzxyzADXQjKhe7aBbQLoOFsiVIKyNl9ZshEDBWlU0lxlznt7QOy5jnMQnH1TJMfC/svfaVWq
snd9QIZoCgP7SBVqIDuE2wahHklRQ8VYKypiFZtp0TmbGVFqbYZzkaeWduR4huMC8MpTjy+8Iqzt
Q8fQb5nVV6FoN0wxbx6yOAJW4mfcKcg3Kgyw9k+GpMsPWMLa11HVkfIgf3oQSOAvsdMBFlFYgAAw
XEuhIn/vm3IwGLfWufb3gcHxjIZKv1fp35GoMdEjJ0PZG0L/0iYNk9Jfesz77adswCsfMEy5PBzX
EAnMqIDlBOSdG29ZiGkuU2Ix8n/e+pgEN71KLVmaEpQlxM0W3Bt8RgXm1gUOjf/B2dCT4gRM2PPB
eV4fSBCYrXk0cfki6L+/bAM7hWmXkVED6sUIoTEm93BD15KT/VvZ2yrNYbuScBGWyvR6ne4pGpuZ
qW43G4gBe3T4B+n2FC8X22omMd/j59Oo8mI3a/vfb2fRlK5g1SJ9xbd+J3/bTQipjbsdv9gRxnSL
BplupACWDGVnm4r2wD35mvYOQxz6Nb5zqAv/fw7mICt5qPRYdatXbq6mvCVsvARuWZFvN8wsSM3Q
GVB9Kyre2e0ZYHBGUhpIzfWrIlD8KTY3oZI6e3URZoAkBipyUQzNebFOm/OkwSRk3ohzoz3yUmdO
CacK2tGo6kLG7f5duUTxpSLxpi9V6EbGXpOGwD6CyG0m6HruCMUbSI6bc0fZ0uabcsCMVaGF2Ay3
yDXOs4oEfNLHUQhN00LrojiAT3/JaO+suMFfLyJS+/dWoCC2cjsOigo77IxShIFrrLMj2Wu7xvwr
pgucx3loxyefg+uU+zuLfJUnZjjis7I4tGJNgeNaALEguJWzftUS2qqCc7QhpmsV/OocB3T5+6tt
fjJ6HJHjnbGkFGSVAkq+TiXoOyeUzcdnIflfWzmIQf6d29HVtHgJMSV1lMwQBwfSr9c8koZ/iL2T
YXe0bZA2eNqs9+Qx+TwvxcT6fHxwDACs0+/PFWR/zS10BmHHk8kVpuWxXLdrAV9AjkzPnXqeUyz+
uafPKp83+J+cQmUGA18QFIDDJ8IPO7EDDtf8UpoxMyF+uRTiU669/tdbaz5sWBqG8BtjlXl+18kQ
Z7qlK7AfKNyQeBDk8TGmSCwz8atM2fC+UjJ+f9KHSK8gPYJXt1o7CiuMmcO+AhWGt99+VfJytjrf
0aAod07mp+wOy+bPv7XteIXtnU0zp2lS3w+xZf4xhhQlV5oXWtaFxGiQbF7lgDSpdVijYn4GBiJm
MDWN2pcH8FKIRAAlrMsGMwr0Vgwg4/gi2QnLnYJNVGMPH52hZQVjwM7Gv8pqYia7Db0PKkh/v1gJ
CPP6UX6b7uud6aIRtuo/1g6EKFlYD/6oj6HFI2rVgq/IQVoDN6iCHqamWTnthOmIwRAnKxLkjd22
D/4pqvSRu6dI2DvC/i3Lo8hW/SGHRCXlxhu3MBVfG7Pc+xwvpxRKba68jf7VzLKswVmm7FUK9/d8
WydUxWWEqW9V1wA1wJvfASBQMoc0igRV+20T/Z04VwHZDmr84JN76cQbLp1dviG/cvZHIEF2/J1Q
jndWgTtc2T5Y4P2pNgZj7hK+sbfhzcNZzmnJvJhtN17Sm9uc/w8iNYRb+CWqStaTFbdtWxwIODb+
cbkgg9yX8q6YPkr9s0TfFPkeqO3pJUQh9XB7zQ7a/NssxJ8HEpeZW4AjGFhE/KiWkKA2F67cx+kS
hSAf7NCE2VsipKZPZ3evu7AM8FFgKYFno57QXslJZtYnMoU/tIRWNZQQISwnC9KJccHOOM2lqXDk
DhRaDPmyyKfljPFlvG3Dz6OUmkoqDhMuI3mERLzWco9KE9JBoKu2edSeQTN2cwUuE/aTnO1ADqAe
hwmomv8aexX6vBUw5pTYjF2dF86qU091o3n+54m1+imONyCibOrupD77okJNY/oYOcs3C11p98AK
6Syp5Uaa5yRlDQI5B6kvTIYQ/+oj91kdhfuzgVgjv1nizkmfrRW4SIoVhHaTvgkoxSWgqXf9TZoM
5+MeAJqzmC8v8KWZP1Cxy5cC9BsCouN9f3SjoUdubFDEfnONGm7wxfVNPufXZc2PVe6kp7cu26fa
42Rl1NTitX8+VmFxSpnk17Gp1PdvRBDFIRaB+sIucoRgTBhthh5JkdF+8zZHsQOSwFpSQrCtvUFl
i1vvJ37bqtHqxUvdQw5nGgYe9mar1BPN4yHUNcouVNpqWZbpF9uYL/vrk6nfPXRtNCAXToY8LvbC
u47zPTGtxl+CzdWvFsNs7Q2CiMVZFT9eSAWaInkNX7LMtOOTOZ8yEtg2uXqA8B96OQqGdnTW3Ui0
LLnYbREhnlDnwSLEdhwDN/k8/ztwE5H2eN/NN36EHAZ6ZsWnj2OyCsSAoJoUGpPYadZqlU1Bmi7X
ogGQIzjoupnu6PS1EKqZr3aQOCbnxdDe6E+48vEiiW+kCi/GECYIa7X6p282Vox1ytjJ8SsiC9Mp
lOYLeQjezGkvf01DBlBmB2xzIaJY9fbLJSa2wCs+PdOnQuh6/i5llh35byi9ApMjVqnO+qr0X0ca
xpmKXh0G0h1l9pl/93IsJYghQ/naNVAMzSvk9f54WP3ANwTSQihyAiaw4HsI8NVZD59f4eTGtuzM
3fiTNxnr4F2onkb7BWzBiCS8zZmjbFkOKhVRv4JS5YZs8rg/DCaWHeW1tZkGmZjK9Pw5rY+iuXOb
jlCLnpPRLCGvFOaeMSuwCUtclh36cSB3zPGJ0PFgziWOilyClsWl/1LDW9GntMAK8qU2qcF9NKYu
dIVLZ087XCp63u7H/FHxe6oxrda05Cf9F2OeR+OKYRPD031R5DtjnjzeN2W0J33HGTO6hXTUz7FV
b5vX+7MbwmNg7py7dSXyexY1//mHb5djM5kOdzcY95TwvOx4vfSiT/u/wG0FUclGBAgos6AafQLM
6dS7lzGPAPzZ25o2bGyhGD6npCPeS+HWiKw6e5eZ5vIiDyBogtMUKBDQFN9cJxB+dLWa7CA1T7wQ
cWFH3mPLq5sExUOirwH8IIDum9FsFZiuYto+zO3UyKeBU39i2Rge5BkoGTfujGVtaeZg/QM/7Ws1
tCxRPCORJZAPKODtnEmWv+nFiEOh1+HhqVjsUA4EtF9S9ue2JlId3qTb2MENUId7qe0AZpa3SPly
b6iD84irc7YzMVqs9C4XtKtBc/ei01Mimg69QZh/Px4JBIUPkVt/UAcEz87f7nsdSo1/BliCclO8
D9Qi1RCXabsFir3HnIk+ctAuxQI1H+4NhuzeEjQakkyQHFdZY36ACnu0Z9s2ePk6abQePsD7lPrN
QUXA2FzFFgovrS6pyXr5QCLCNDfwgca/77VyhXS/jqGz5ZvK1Q+2RII1KxXhIukGQUiKTxk0l0kh
ciwc8+WbJ6mFfBGpJkqSjUmAqO3IJrojC1qqyqT+N3rFN/8qzESRQfewKSk/niLDFI6TB54tRzgx
7ssP/MYGNF42PBoCy0reXWK7JhtoLzV7t/G7ZqO4YDTkFR3Rx+aU6vAW1KOB8tBz9Je3QRXT49GL
ydYgxZiyctzjpgfW7NfYZrzOwydR5ezDyYXHzlX4H+Xhy/h8PyCk9LW4116wgZ4TEYVGLv89EoKW
3fHmaB50Osu01Zx96qapGPtUcgQCc6j2QiYi8t4DShHpnZXLcD70DPxvzbL0eGH0XZlC8BP6u7rm
YiaeYwja2cVuc825mVaBUKVpa2gNvFvsivR49Jt33zQWc69ri67xUhYa8Hox1ygEYmET66Vxtrwg
HSgQZ/a3cBW9qb659fFcHDAGgT2qUMSPHWZFmRKky+60rNQV4taeus+pyVVWE47o/xVmTmIFoJmT
VVpOtAlN2UdmtyL/ingcWmsdlmWtO/ACeyC0mOfUSac+Q6RBotyK05xr7NNuwdcv7gL1wVedAuyx
bXFLxzaXCKTSL1rRrapSY/4BMc9v5QrxWpp7NfvKx/zT83CuUFCctEzM9/eUqZyTb1dCeA65hHOy
oh9OEEpNDYvN4QV16UCDZ3K2bq8iVG9jtjt/4eRWvNyzA3PjcNguHdv+0VO3NFGfJNgKVy4rkIYM
2H/GRggTL3+/PHp8TIw663My6L/NO6C+YqLXFgDOflIvUt53wlzEBGjOjwzAQVZssUiidrzWG2Qv
du6Z2u1Yd2qOf/a+NBjezNvFFOaPDjuVS27AzE2eWiOhrVugWgW6nTQyaVB9Nqd7nxzxStHnYMNW
QqeftvAwMypaqWCmHea7m/971ODyUJnNxxx57pgoCmcF3bGgVNyfKKmwyqwYxVEFVvKxXoMvIdBi
BRKCeR38LhlQ5mB+Zc206I1g6GGC4xjjyZnc14rKi5l+R91Te+xN5I6VQX04PMM8LfC3dr3s2RnF
esPJF/WBC6IGRNZ9Pr6oo6dg3iexV0TijAZqBi7OVA+lDeDkhaBz502e1XeFnvWlay0stqHhEULe
26QZUdXNF+r52/9UpVyj0IKxly+kkaoYykuhaclN37qEJHIHEIIG0Z6h+x1PMtEMKCGFc9GjHh3o
FteourLm2lWcvLmR2Bd0mGGgPMgujdbiwoUdvjkviTJ0VKoMVJ5ZNTW8MVipkwUok49whBISwIll
EFHFT0x6J9KOUjYLlqIQ9MHHORPhhUS9TLelasEHQtD4LA5VLhSjRWrTrg0RWIZbG/p3Kt7O4MCl
h2eL/mqcmX2D7pdaxabF4ckw97DL5EOK1maNUv1aFwauAFdkHnrdRg4ayV6uSf0C1/2ucXV8YxEX
JbEFCmmbvzwN/upS/m+yJIDMOKQQiJmqghyfKJRMoLQe5N8yvo4yJvRe5pqQJhaZwBCtmtigN2bN
LsopnecJzVcqHiQL0axM7RjS19F7dhXgVReF9b4mYJiOuzWw+6OiGcg/67Yx9elfQNZbwu2ky0sg
/Nf393tV+J359Kb4zSo0HvHy9gRbhKX4FRHNw/bMDZXfAEEbC+6pduDLX27YmeRRbPEs0p12EfIM
1bAC8fKymEMuQk/IZS2eOJmMGH/R/8EiogeT89eZRm1Leb8aEiDxmbixcLU+BkotIvyl46nXifT0
zNEH5Dh+NqC53p9IPvvXrqBu60N7k5k+uK+B0iFK+pi0fLtO3ppnqpDWIZZ4WDfpswhmbmA2n3xC
iuX+JsNoHVrLjkVxIdK7F5pzbRwRVMepePNV2E6Qtugp0x3Z3enQsLMBR2AqhZEZpPitoTl6cC7x
3zywC7Frm+UsW9384GrL0Vb9hbUu3V1JjTrwvEyVBPvtMsvS9AR8D0hd76hs5C70GwxTwsiFsNum
ESReWyl0h3A3GoQjyMPRxv5yQprWYJUz+9JcHnpNmJO2I7PvNH5Q1YZiASvzlW/Hc4sPTkXAZCOA
BUPRoxwbrTsUANVOIPy9vzkjgACEvaSaDh53x8iN059265KYd3pVL+ibaE5Y4j0EAbAng7bh0nZY
XVWzObCp/cFJwXIXkNUnNdbiAaKTG9ke92mKxCREtVcFhBFvLUkTUaSSCWg1GeYl3tF/CwAeea5U
m3ytSweX/vLsPV7Fy1UAlEtI+HKXMueGD4u0X5y55MVljwpPBho3dYdeuZMtJmWq9SugM9kiZRDf
wWhZKS5Sdf1j55SfP0VoWT/LjkWpoNyl9PmjXirahB6c8IoDOYRvOT/lvl8tzROXIzJfTJyyf4V7
dvrAXe3wFePxz0cGai8moaZ1HWHbf6FZ4mZGVwu+g+QLo07YxBvWeWnUdbAjFA7IVDeGmb8k2eJv
50avgiy6q4Eo313O7CEmDVXs4O+MFffWi7s44IMcSw10gZUfE7ma8hdKsFmPabTo9GzAKRTnaC0V
szvbm486i5ygvLRfyMLB6ZH/Pcs/F442q5zjacBH056W1qd17BMaaSsY3Zl0VI3KiCdVJYJcqPdt
U8rfqA6ON6nxNU93cPDlojYnLr/PTXIEzDQ0q0lgJx84CGPPyYTiGZLpLGJ3OaXpXOrM1ys8Oj2z
Xqab5rFugLmvZ+ERC5wYrJkw7eLhDPIXkseW6l/TYG8wE99K0F7tIWGssErk01nZ5fplZwMk8FxT
HmW9yt6/KVLc/WA9dNK6kPT56e6HI9pcoEcko8ZHF6sa/CWz+zFrNiNeEiwjgVSt+Yew5KO6w6dT
D2PfWp/yyU6Lre4BrDqKYnf0xTikm3lwFBy3GGnlu7fGajyT/y274KoD01KbySmK1rBWObUde7Sy
bLI7ucAwKLvTRxlE5Zhu0Fzdc13llc+tPxMc73RVcoD/3pByfgMdJ7+xz6CdISlxy6/A+yoSB3wZ
DwnAmDWjoHJwfA4P8Zi4ltbvKQEoK6SUL52KT5p36xTqS0yaakaw1iq2YwqUgloaRQz6IriNMtlX
l8pE0/ntVEq1wkRRllN+06DtI0U+soJdhX7CWP/rVsdYzx0nUYsJkoqh/WRVXTOp72b5D3HWd4Tp
kS/Zpou/LZ5nHIzowvvBQfuoRXewQo8Wpda3JhZ0H8/OQKLDXkx9vva6+PG+cWL2UL4Py/+s8F3w
uCS0FjIc0K1JbhYFwmWiZjHbUKGyznoFhkcq4skgabX9tURJwN9rd7iSKLo8x/84OeIUTG/9J0fW
633g1PMFDBjkySZnCYUbon2mqHw9VRlaYe0QXVN6qb7GoUFuAXeVvpqaBkYyyJA7ppFeQ2IJG9AD
KXqbmaZwQR9guXKgwPlkH1yZi34EWx/kXkxp+n+xcbU/jLKpfhoGgu8WNLRXEBBY3ThGqc97Cs6N
iTU0aIlon70HliYdArhOeHmYFznJ+Pr98gDJWy72qh3I80fYxZliFFT4bAhB6GHKJ14kKAsms7g+
avZSvbUA/fqVPm7a3qKNH4hTFU3D63POBSF5K7LPW+rle7acoTZZZKKvJmVeLChtOghyTNN9aMKV
SNBfSUR7fH896TgmXUP6OWmUg3QhcLdiy3Exxl28gnRyj4omKqeaGQXHcOh6yPqRY9PSBuXFBOjf
N+vZbY5V+tb+ROokS/i80kaOUi4J+dTrKNR3/MiMW3rH9OS8WQ6iK1vtErZsRW1E5EWYtEcgYFd0
mEMObPr9ahTkrA544jZfHYuxhN38OXYuiGHIfFGS8zVAcy0/8WDjtTtiOyQdk7plTX2fQ2VXDLNl
V54cVVGjp/T0IR9P220rVv05DJtBm+uwsfNW9l1+EW1OYW+5xJ9Oj5uJcntRF3MnGq0EEVOZKm8Q
+RCZ2cWHCZP/TRoalRAoLPHqOoL9/DLtxbdkj56+cmLTe3eLgaCHWaSywz8x12j1JheKElj2QTbi
qCU3hDC4UwC85DnScP2ESUvkEir6wvP+MlIfgjfPrgflW+dHw2DZa0OY9+vmEdvJ9pNff4+arpc/
Lb3GMko+NTfJeEufXsi/+T7FKugxXJVoaQCCirB5Tyc7Z8YETSwd2Yu6IfsppyCp/UuMXpD99tIl
PN6vhvryfh2P5dDHvKkJkn6lxyCmpWddRpQVoAdGIWnC7GZWCfMpvDO+lZrWdZY26jozK+sBRCS6
fyYxLyFtD3fxjRucIDwCZhz3mu7KdyN4Luhf6EnI+o2DgQw6eIEyJ5weXWKaykmebMfxNurt4enW
h6frUCGx/XJBgIHREL4+dyusQT8QFTaiQDEL7l8YpUG7k8R46nNd2MMGYavyGSb4CZrQlsghHLql
Hicqx2eGDUBlXA5Tjrs4IxmSv5EN3b67WfoRbA9Lcjpa8Xe4K8KMHZUw2yf+6Liz3JXg5riEVyJK
/jI/e7K3ULrnFmjXkj1PzRZBErJ53XVsLquETAShaD7htGMBCm+5wWcCE/rPwxyid2yoYZz91tZL
cKxU6fI7GqbQrKc/aJrgw4ITc8SilPsKzJM4Yyj//896vzYWPB1hN9QAj3U4kKsbwdX1tywxz3+u
Vj/S2bnbsSb2RUHiDzoIiS8LrAJ2iJ8IGNar1s1kkIQzbZj8YWT3ayy6mPsi6hlRjztI7CquhNON
scHevW7hXheupEZGGDmBlPiaor0iyCohI/fZwyL9qXvnDGSenKlKTcjA6/ov8u6Upv0x4YfTqs9h
KZFBdpQlG1EYvdErQx+rau/kwnWfxttWDF8g8v7arzpq6Cnftbab42N53hD3/2AcXLStofKo65cz
XtMBwKgs2Wz8v6ol1in3mePPyizABZ/zQloSfWmZi5cNBgQUYKPk2Lv8Z3UpeWer2KL1nomC0MS1
18HUWBVhfiQNdanFdN4sR8vpm75tu4FEk9W47P0o52CDo8FIkqfAB6bMpKP+sE3RrldOIPF2JJQf
cwHC6l3bXy8OMUu+FDrG94/tQHCX5jfoVH6EOg3oKpuOZAOUOKlwlm+gIkio70TYDouz3BEOZa71
V+KwR6zNr+LEUa7y6PDJhN/EYmLC+L0ovBtcN+tGuU49zzHzX5QmqWdx4RM+4yT63xZy7DLG1qUM
Qi6HwztiO1w7B/Q2OLs7O8KT2zXZVxsG2kacgqaTPovqFDCfi6Wi1sBMtcJPx7ayAumQ6lks5W/O
HAN6hSBdUmhhCDsvE7VJFa8en9/46U9rcprOB6Bhjwm0FgQTujFW5is3ROi3gOuxQIW3mvbzLJts
42gzKr5RPh6gZLsfC7OLghMKsM46Jvql49125zLpQJxPh67Mj62+DKZWIZKAYeLTEi9OQuknoKr8
BWoihz3BufE4fdTKcIIeRGbjRYLcbHq2dyirmGcjfrVWrGy1V4IEB8ynY14qQXRlZG1aMbvZjXyW
Zm0RyBFBZ7TRP3rYoE+zLR19IJJap5fO8X+c7c32sSLu53kjX172ixoEfzWKYjGZgU9rPfD15XfG
HwfQUmd4lNZYvzJ0k02D80I/uhRPqSXuScT0kINdDmnNnPoQVWPGXCOf0UFZoYIBwpjH7f69TS7u
H4GmpADyRXC0gNm+ZbogtSerjQwmh6LqU/r1TgxjZ26mnlAfpNHolXguj9XgFNThZEbVJU/Qhxjv
zNbaSYc9rvKOnVGS2uzdYCjbTnCJZhUo0xUS55D4h22ZYmuahwGHPpnrHzdgMZ3gbxrnXmuWeOHD
+/KPC/TEY91DW7EKk1YjOXQzMzxvrAuVN+of9xS5ZKJQlrQoCgt8C11klfhwdTUjCGo6NyIhKMVG
dJzIU3p1CcR0Yf5fS0+X7/wk74vei6cPvY9wkrzRmE2buOxJV+q+livEw1FesRao7fCWwQRvIHKQ
9rpgKiv1BBM7uE0Qil78tkJETNsMfVZjlnfXnlHGW+4aE5R8XNzsVTL+AjTw2aWOFz/qzq1PSHpm
qtXgosx5g21GmjN5pu+pG0guZTKaX0r2nUhnXrXixyQzw7Paww+F0zETDzwVz/7DfaVxN7U4gbcB
QAcwpG+HBBfvD2Sk/PGXp4bsYzZT+4WdA4AC71BlupSKIvmysfvzTLQrrX21YQ0+2xuNH22ZR1BP
a2z0o7kthf4mBHVTnRcieejVIZalg0uyZgb0lDBHszelOgyp8gJapmyOftySkvshHeNZ00S12Mev
cg8KEWgZ3vA0gnIUm2GVk3bV9jBh8grf6xy44aM4dih5rxk91dFblqYBsTDZAqmhsQLcRkdMVVmN
QPbfTJyEj9AmAvgLq6P8KEq3XNI7m5UbJ8YOATVVGfFtLYcdYIyrP5It1mRyZbUCyGgh2XkJ2JO9
dgOPLciHwJbBVYl0S8gBEV0+E/ZmVgYWGmhnAEZbEt02h5/TMOatZ7e5EPP7TWLWc3Z4pBC8pZDM
5eyvuIBo2u8BLbh6W3sU3HnJ6AhPvikuaMamoMW26falXu9Cg9kg6uP38wQf27W2KH5LRf4y9fI8
nb0fuzH8UikU3yeWp15X3hfXfA/GcpHLIq+aeO6/aHsB2TETtko55u+vkmweJayb5WSL9uVDTLOJ
bKYtWBTNYu2+FsVNUDB2bDYVbdJt/u79YZXfhpInbbqSforDwbZxEEB+t5aDE6GlezN7qDGbKVp2
OzjrA/tPYlsXcoG+WcmJT4qA/zFar5KnGttIjJvyp7txiD7Uh0+A5aIzZXs8PnwzvX6Axaqduu4N
Z1cPuFJGk3Rn4wN9qmT0cYziPeE+IH9gtKflU+YKlBBBYr9TrWEo3X35hC6OGqNGDMJOX9tOUmj8
HT+xacnvLJ+NvfFoZ5hnr7F44ZbYBvJKAer0YsBzm2nD9nCuWz7ipv3BrCqsBxzw75fMHxtDo0Q2
6JmhE8E0Frx0RBFbupIsGKvqreTuJ9sZETn7C8hsUq/UkIPD1qU/7XxR4/dpAGe5UTsZwolSqcWw
64rtfxWQGF7Z+GUM+1QpX/6EtgGl7h4OOFYZNUieD42+ZQjybJjLrkAAr70N3IIgubtqgxyNsDm6
/JE1oPEFic0LPjlsl32w3jSDKnVGo4UoWimJEcQCyc5L090/dXeKFPnUPMMhuW4s42uC2luqUnub
NsSSBuO/159Yk0yKkUC63fjNwSyQns6V6HlUMtPekyncLqyuJ0xK4+xBj3gp1NZC4cHuEtgCXmFs
CdX1Uq/+z8XBlGgQ6fUYKwI1sJbRmxBFXuYdRqtcG7orV69ZTRspKxZ29ibPxngXUC9dt4zmCENc
XgPZi+plSQUn+GQPzrc+Yn02upttB4JQS5/eP7qZrU66Rq15e9EoNqfZPQ/qsIvLFuhEkyPtAHLv
Vm51GYgFMgc28oS53V6idW30NjMSeWT6RxkUJpfkG2tRtrbKSStohNQD+WA0bO0rVh0V69Y33JPd
44R3uJ/AQ7LNLOBZTGm7yyTynpRRxUAQOjDSJ93BSYo4KD6w7d9CbN1YJiF0W70o9t94LZK6zrD4
KAB4yNCOCTHtWksRgLgMUx8BgrC1VkbSRWdiUtt8YQINi0o9+URFRZafWYtecd2319KQ0f20AjZm
8s/LsPJo1BW9Wg32+GqpmIYiY1VuELMrVk8XJO7gRlmeO9URiWKzDPIIEkmkVdyR/ojkx8STa3yl
gv6VQLBPWKutWwJI4PESzJ02MgXn36/yNm904j5xE/ZcMbitL6wqyGHfBHexmSJr1qMh6RCIqfuk
VIi7jDeHcoYtZHL42ryXdgvVc4hzuhr0Y14C6ULPkCxMWigFrBlFcO99eD0Z+9Yg2t271T5G2p29
cww1srKKbN6g+UHMlGGWOvwBf2FKXXoHqLTwy7sdjLCTMUxjQoFdPq1qw+vknI0aB0Mi/xeJ9PBV
t0QQTyC9/sSoyaBemy4iZkZbg+rhrc9wtJN3YlqHOoDJ8T+W/w441gfUEjRTfD3lsE1PwCAyk5H5
vWk3coP0H70xFqmxgvzkqMmyi2c5HCx13+u5jOo2p8pHsEAtKGZb4xjvUHrpuHczmlgf6K7EDW4b
xLQD/XFtHn2vpq3eiukvE26+frl0pdzFwkqrdTzwW8ATkzulCEFA4meezmpsHDVFPpvf0oZR8TQH
SdKoXbshdi9VimcNGl7RlblUdtnIYSepcjUisGg7O+pkxdFedDyCXpKNbp8hmv+kInxMzMK4QFkC
lneaaazVoXmfSDx6Snm4lPxS83YQxiZo8MOm6ZiaR0L0mNZAMwSFUYBnH/aUHrZmSWfXQnQ2cVJD
76NGgXp/AoVso6MDo6xWcccEnPEq4v6gqXco5Ta0EZiD/XErnb9h+nY0jY0CIxyc1OQjJJmdbKnJ
RcQv5we5gZ63S80celhcz2TyLe7wM0adcF5774m7c2tyJ0sPCdGLaw+A3GNMGrzm6/0cnArys+Am
aUAXSChjdGiuqT2KDqeyNAzTlR6vs1w7dq4XPM60sDvZP8jUMiUDYi77pJQTd/0YXt3ToKPwgM+c
SA205q85W1Uy2KzzIXW0Rp+gOfNxp2zoJ6aZ+DBzD2gy0YCv0eDTphXh2pz5UwvhMJa44Ze6r5z7
c6p+2zGR/YnOtSVUOv6gsnELv7RUNGTRrCMLUdzMQPnq88K3ptDBCfns84JHsD2ypmkRlea8KeoJ
4R61axEbrvRvzSqDpbXma1SGvGisyuE6nYhRjdAvKcoLmXl/cndHsXgRVszaF1CP7+iy2vuP/TzI
YeGhvsgClnS+f78z9ErILtPOjma4QK8ZTw0mSuxIoXSkafes2qIU7m9pUtzLeNt24ycYDMAZaKwP
wnT3WpcQ0+6xVtIR064QY2OCK/EHNe7DsPdCnXropsTAL/MGDjHexahHvlUqA1dizhqj+gapzKDu
NZQL60+wV564lRthB7DlU25JYvyAZVyqo2L6keuEXCpMGiC5PCfoJOTTxcn2mZRUwLnrMtZfh6PH
EMtwAeVO7xx1AREKMZsDZQFX04/xrayHpH82912YceNy1cKoL8ZiQPCHlakopgFsN4jw7GYmDh2Q
ZWdw093alxJjeXl8HED+BbQBoHKd5Lfyy3a//T3c4s+LySYbmli3Gcp6ssxloOXzmU1Os4TwFyVT
XtiITslElZmBALmDf5EKtSmJhxV4+djINAZidTZB53ejWDy5vBMjKKFuXe5E5iIrGZ27ieO9qHJr
A7FAHkoUNh/c5czK8Whz8yCRiWH4VhlVyifhhx8zMqLg2zAosB7Du2tzs/ujFJ/M12aWOCUwBEsp
Yz7qTjDdR49CPKhqn5AlwFFLrc8CEwYv0wcJcpyCSyTFbGqZNc0GAcB9ZZKJQXT10Y1ShWzGq9fc
44vxORtjnY0KjomFzYlcGwC3AVCv5NaYem60QRf9qh0JUXwYSEys1xeHn52WMfcxWL7Uo6B1U+Ka
4ui71rA7A9Yeb39KOeplFDxzaQTKHZa9AerF6FXJpEVkHEFh2Ky1rskkyePxTLtKysPt8G/U0Wrd
H27gFDKwEH90on07xurnNzbl1lc2LvMSMarjVKMNG0/7Rl+NXiM2/EDy049FTB8LSTOhDoRgA+zn
zLzkB/eVlC5f8VHGPqN2yEu+78mcgr3LLMQ4TmeZvTkPi6yUdBEEn5FCWIn4NLk83p/ITcMb21gP
benVOH2NesHoMAwkBykY4fzYjzVKydn5vDKvNnwk/hjkDybcSNV0oETj85+t9ohwzDgXG4T/R4wy
7ICYHWyT9st+8vazYkIWF6UtBGbModemBDZhhhs3mlQkH/aUmNMrl0m86fAbpyyg7IRj6oNLHDe6
CZdAJqAQ0XB2B7E7ilQYzpqdy0TbYfI3LoEenPOssqq+wbBE6Oa5XLJ46sTEWgz7FZVHme0YhmJ3
wtS1K5yMp5/gkQUVTMhksyei7Mm0SpOoCHXoCMhly+VR90zMmLq7O1FFRS7OxuTE7+CzbaxVQqAh
Ldlv3RmIRoh+A+DjZ8M5w4rse+nAGw1B1+SsMQOXgEg0iDGcqBaFmzZRIgEZhHBR9EL6y2suFqiH
ygy9/vBwMxIzNUcR065ICInOFNX8XMroa+fL91pqvvSo6GLSoRN1CfOj/WQc9Xx4MbM9N6JKuFs5
/hkoPmUYM3QEJfouHGB3gSj8yUsJCXRKmMOhe0m2a5EK5EmvpYLFs+pbGHtZbFQ+XFfBYO3JpZ/R
BHaPG1JQxBvM081U55uESQXPNqaZLUfVxXvhsQYb1HRlF+EDMkMpJd4rToF2Dxj8J1PLssHj2JcN
f3UnPtByBIJVnQWt7zmiGAdXpJGYpPzrZIkekfsKjszuXPugytsDwY93VdS+4a2Hv7Eod9XTF8MO
52n6sfv7INUZYMYLBJS23p8OGOeMgExOyfvsJdPHIaBYwhBQRpQrhr2SlG8wOc+yDRmRrpIC0Wd1
9OoZETlC1/txokMrP6uc+6yr8KrDGq/BN9TROS9HlafFg+CWpYO6htKfdXAmDI7aFXQueZq/Bre6
TbNwJy/bfrKc/wJVvouOkh/bQ3EC3GY7U12zHZKezLSWofvuoBn5iezX16ULFzVr4uk+CYFzNO7l
kApvMtMpr9mQC5PusX4kEn6tqqvt2R4Q5kTqYVeHXD5rQYn1kzZa+e8aD/OU8tHHnOmAOlAyFa3q
poY3ee717Amyl1Mp9urBxjRmZyzhOOque413RIG5EyLzIn/beepCRTPJVHXGifch5/dzKv1Iedw3
5RSM3kc1Kk2JoLMvlKytZnwrQQ2MCzUA1sl9nUlcRsAtt0I5IuAF/yRGGlv2Srng59T2GyD5b7Ag
koSlTeH6m90/je6lDatf/Vr0YkPtSDeRZIxcJrnbFBaP4r1fJgcHt9R9CDU7ThSOkZpBLmZarXFH
ALbIwovQV1veVtc/XYXJCgDxHjL3aBoRs8zHJChv6RijE4R85zTLzI//85zewUtT5T1Gk2d8A+cG
M8nxkIl1U+DBEwFCofDaK6YfxlUXbbV//seTsC4TSinc8DWUx6TMlTlbkczWSEin+qQmkPztdCmP
x2f4p/5g/HzMoDTekTRp3Qk47fgEQFvlEMCqWMvmK2zwFfwC1/1KS2hMFHDizlonPEEgBI6DPDFU
wBtaB7MPxxsUONEc0Mh6Uo8QtuFVwgQLs5vY5MgQbxetsnqP0nPuZ1zS2bLhyzk1994hme5iXJHY
XnlGfLVhNuP0zb9QYpUYAu5bVYoKIPjH9ztbcrST9o3UGCCKxkNlje6IE7BK476M8VIAC1D3mDNU
DEe8KX2OK+xim9NaFD1FwFbc0DuG2GqIPSlBfGriEYav0DUafgLAXRb/azrwwkblnHbiUkzI0dY+
kh5UeX2AYyncFJIEkqqs9eSW87g0rQ/0pnxzoSvWMxzFFNFBSqcdIVMomUhwJwpeUpJcQVxnVTiU
1gdOxPDZoI3V5Pfjb2Kot+46Aw7Z+jIdluH45RagaOtLaXo+fj9yYviD01sZqGMbl0SxP2UbJrxV
0cNv2Q0XSmU/TcR06743rsJiWzf7k+Qpx6g7SHZaAz+PKUBSl2WbKTrEg3gBRp1M9SFs0IarNvCy
IuD6EnB6U0kXMB/Nyv2hWaPhjHo6OzCP8VqBmvyqSVKE9K2VCYrOEgzhQLEXqx4RIJw9jh2gx8ed
OSMEx/Fzep7/6rq3XtTSgNvyVRXt74Ynd6059o1KeEnRRYMRYI5sacKkv/XXcS4crnd4nGr8pWfW
QkKfLXuSQqJ+ICCNTRwg9xNoBSdeqtJkqiGO2YFSTm7K/2JweyGNRSW8YOnlq+snpi3RODmA2vft
2Lbqagfc5NdI59L7WarDgA1YySoxdVhoEXtjA/Bri3VHX23zCiq/KYpjryui3DlKt4b6IxF0JNtP
rOfQa0wcvl+tlI0TXvD7hG4JHsk3EVyMVk+rnqXG3OeZpoRgKRCwQwvJLxm44RR2QaPfWT12ZSYd
qp6PiMQJx/5A4bOZ34QkyuSFewkYuoxXwxWNaiqZHm+iiBQBayyHy9EMYtXPFFojC5svYh04oBsA
KlCuDdb/QdBaoU6zb3zce8autXtEqttAxtyZPUh/3onvvAR7LY9OpAhFkcd7UAH7JM4lCYrvKuuQ
C4p3fmmGq6a/1KD8tgFVX+lZD4Wzsm1yB/hBXGYJo4ExHx5lJXznCFBrWhAbD8A1jTDrN7It56GW
6Oj7fmV9ziA+RsPG8qzOs3LIeZCfoPqbYVuhP2nlzgjsc2DBz8xsLR8MS82+rUYJxbaEiR37oCVo
qkTk95aO9XmO3kKS4PBOxbGGDDArKmcPVaaB0cpnu9O/9YXLtbD5svcm84RuEc4Njb3XIpt+4kRM
99sp5PIwg0hQYxxvtxAGZ28yScxsfXsala6HtVUZSUiIN2Cdh0h2vEqt1NcPzDgPA6TNnRb0Epyn
i6bCLsb44rRcVR+bO39xTWKnQZb4y70HbsZw4zJPvQ8qS0goBKtCaahuK2B+ip536D3QoWFf095V
0IHhpPul38KZTADpFH2O+Q+fPSRw9LOQZTH90Kx04njFGA+hRK7LpyLEnOWkmTfNMtzsYGEmR2uJ
3rHPgfLs87RmB+uzXSuuBtEbJrlD0b9RvfoSck2Z3bZiC5esrwkgaoDdFIai8BYe8rHlhkNn3fq1
IdSqGeOOsChjgdxCcw/nw829c/uiwwaxphdLxwzZEuUjJRzgwAs2tw522fzLwnm581DoVE7P9qcB
1GMBRLOVafyg1JOetSWSTnFM+incEeL9xVz2tlB4KN8h5XGiCpwGq0nYeu2yhoj4meCl5Coy/mWg
U3bhXjrToqjceu1l0Qx8xvJRD7VENjzHjwkSsE7UQ1xyo7Xm8/wTs8oxsZrQ77psfl++rLP9VaWP
n5ukq/XUJz78JPboOGEyqewUjyVsZk/9yOJc2MxEBleXnX0SDOms3eiffQcdI0zzhoVrx/6DOuzP
DlrzpoVXap38LpzHjDvBIo0Gx8HqAM/BTbc2nmFlLSeMzc/1Eu4Fx/vEOI5Tw5dfDi8Q+rf69kw4
bleT1FwpF0zbxtJsVa72/7F8ug3Sc+ZhpUfz86eJYtVjkL/1+ZGQ/1Ro6hR7TMWcp4PVgiKnxtMk
znXJ352gePmqx9bhzNxuHc6wYssorMukgg+8Z6QkgeT4jxL12/SITbMiZgLFMkLBTuCGa0jnLBLv
Sljz8Yi+t9gqigiSrkcFi30FI73x7tgFSiY+YwAkWsitNuq1lHJ6p8Grw0dbHp6ZtsVUz7jcQNC5
1AIdS3YTBi75Hp8qOu9zruEmWuLqRyNiEydtazP9Q4PLEy0vw8B/hOLQVMLYQf1xAz8jpkU6uDMo
5/YIH5tfvDckZS43ivoZabhh/OKFKbNJEjJKoypuTVRyGE3wAIM4XW3yiAhrNQz610fBUyHihyWL
0Os00C84alXVorn9LhJnThCJeUHnxWx8Jz4PIEmVIGtBjVAe1SwHSpMQYkHV1lF2/BHB6m31CmTd
B/Vu6ha168ZNgTmIUFS5cr2AqEnapZimRC9FM9L3QNC71fqGS4mEfG7/NbbU/LhpYRvE1CGauMWz
L6XmFhvj9RK5xMukFU/paKyDQBgkVFzNftXDa6nKzCQB0aYH0xL6H9qQ0dG4J82uDkXYE/xQQY55
AoGSFjSbNm7ugRQRpdnI/N2blBBbza9FnuXl8HB81nCeE5zz7zz2bUpl2NmGSmYePREQ2LzBSXsz
GFzWQ4WmHIau5M4c8jIrNNfF7BaGagy+UUheoJGOm/DkhOpB2GNucR+u7oPp/+X27OmJxCywr5cT
SJcCfSLX1urnE88+dzfdpf7vCPej3FZ/cYulWaihPvs6nieZBmjcYzobWE++zbwAsly2JwVbUTMo
FihXovE+snIOjAx0QXE7H1urgxdpzgFb1FYz5mVQZeyiQfMIHJHOcGqGkYiKlYZrJXr5NYgisoV+
GFB56p9i3KnCFJtKHyQfLJeqtP+JChSBnIO0I9gHisd//ianUvzPC7k64Wy2b7/3kY8nyK7dHMiq
kdfSDhskIMWHc3hyU91o9RzM7U2EBUfhYFg3/hN4Wmop5bms626eY9hjkYOikesxPr2/jWn+m0N4
APHDFnqwYaZlW8OHqTSH5RT2I0IcoEtFg7WzxCNuBo9s4baDNJXYTra4oPyEvLxlz+86RdBiLHcb
eaLsvDeDovtqYnAVjHYoUC2ZHbLmdt0vorzR0YTyw0GebxIrdB18Ss1uVlGmf/JRxYmzIxjQok5c
kRrElGXPQBoSkzaD8QqLEOm5i3s67Vekc2we3V0QYcI5uqBD1wNGzW5ML/dmjur5IVvxIMAIUWeY
mFZE2YkAwk6GyM/CY2lnxkVAWU1Xv/ErYW27vqjGlA1Ffg+heX98tG3nRI0HZWQWR7Z3fMRfgzYj
sXsgaPqScRbpIoNvTQEb/qvfZfrrnhVHbqOljrQA4eFiTUzFwl4HFtnvJJ4B6dkbzMlhTF/lsplR
h1AFBUJ7U8ng37oC9Eq78Hmy+yziHnZC+v8Xd6gwI4hRYcbVcpAKHEd9a9a5TZndLbcGZs8vuaEO
IV2zC4t7MTkDn+30Wr5p1eUmugKsz/lHGXCm+kpOclgye2LrqjnzjRziyZ8sfnR1twPOZmHsbF8i
kjGOrKtWpJ68dmy6PHsjGqL2ZrpaNQsr5bTUdS7myUaQjJrIgg/s2Z0dGh0HQchyyhKoIEbrvH8Q
fz6nO82AfSmDBNPvflPSNxI/rIgSTuZypS87aIXiMGqWrDqCWHs9nboG2IabtSKTjz5AzS/1YTbT
mEWOHnKxudInGX7YYGU8bUV8Ndkk/Wh+T1JGeAWxXIixwcD2SjhTKLXuC2QYMcUKPfprMdMdiigN
IZYbUgVX2waU4cMX9NBzbal3dq0Ual2sfaZ+PzF5BB0IRRl1ekP0KMxBIbAB5LYh9PR6MZfnJe1Y
XaVsWr5/PBAslp9FK1G1dlnMmzLSYCMoRTbH2yEXl+jDxP6p24Mrpf0GSC5U9iD6fVSqcc1urAWd
mVyr7rKWVrezkvjb8KUKqF3MZKQrqGdPlClaZ1Jhp4Thar5ExKNadO0rAwC9fC9bnoCAPLS3o/YK
IosCnkUt3GcFNZc71x2RZWGrns6QOAIL1JgYIfJHR3K9NgY1WjHxoFv3nQi3KuTSXJjb9k8SYj8M
FJb6AENNHsEWc3ltErloYpQhAyAl5ry8nbEMnZCLkmu/ePu90H//AN9l10tgRpHfPFIYY4ecuBqF
2qrTyKa72RWrowIvhPNoS6to+MM82Opit85LtwlOwDD5+G+1mH2vA2Ta1m7M6xOcwT4xs+mlUv+E
NpOp50IBX5EcU5KsOjbLlsAxOkaBNTudCnyzI1wR+4DSCkHqnAym+rn6qs1mV6q7Rtp33wVfbTRJ
e3DU8Yt6adXKKEcu6yJhA2cLwmXBgJx2gh97unuBYDKJyBV7Hc96VE7DguSHGp3YDUT78UQwVF5B
mLG6836z1A5jOF6eiTc7JhIIoPeuz7vpHu4Bg7cA6PYXAGTJTX1qvt3Imaf7vLCqu3t/frTWui6E
/h0/SmZgrjiaqO8Xk2w743C1VVVgfHMUv9l7hx2KON2hs2Jo+AdwlwjkaOVNHkMilknQcE9YMAkM
h++ix0XVffqw9QGFe8Ais/H7yrgSaf0qKOD3hCbxFKD8SMqzO1XHoPFYoNBZBY4lUueAdCp3zKQe
z+SiuV01Gu0JzyrWbUpPjh+qoyIOAt7lj/Gi0WvH6hybaJ6RiG+YA2LHQbbQKgtfyk7CiiY6DU2F
MqmHBVKJmXQM8HJxN8+6ETRIOXXZ6nz0Nuv/gNWoIoUAHCN1cV/UJBy1Bv9Gi5ePtprpscs6zRmu
s7FPuVmnI2/I81zzrKPcyDzPnr0/MJ8ENQyFbIq6NFMn5HdKBd/M+obD3sbu9ZlBLJnv0A/6GfOV
i9WHuhkQsXHzWx2HKiQtSPF45/Qn8dDf0mSUG5vm8FevR5xp6+UKOTvOONqVDB56SJQAQ02y9Ab5
cSrKbzc6fI17HgmUA2cz/d+Sb2M4KVJ63CH+L4VHhIVi1RnxH/SYB+VLmP/sKz7Ua1xhc3/hFu/D
nBICeYhmOIjpMa7XDhKjOyNctj2PS1NrMRT+nZfPEDTFQPG4wGK/3UcvkF06HQm0ls3THb7eOfEC
58g2Rq714d/iKbaZgmb+r+hqa+gWXby+SPUmIVPL/QQYyw//TqOA06lFMyS7u1R6xwChCOcsp8on
f8RHp0bkvLGR7dn3MBM/n1oc9BEGguySGNnHHq3K0ruCG47sRLdS++E1BzSpcSudFBQ8QAbZ0DGO
aBnJWYMr3pY429YIOS3vYB68eeVvDQnoOa2NyP14HC48dvPRHkd9jXQkv5k0hNBDLurfEq/g6Ncg
6KvWd4WcYXCpIW7Fp4xwYVzkBP8LgaenvGXQY2lZSTubgbKlTSwWtlKUHUZR85n9eGP7yXGbO1c1
28Uy8h+73+4hVg+2d7g1vTwebNEek1Dpa8OBSClmXOpjprtYtLP/ebL4vVpm02lNbWg/bZ0gA6E/
9l92V18kQP5Xn0uT8DucELLUMQUKMGX6XH02vO1LQwwNerxENVUVeOVDm+1PnfNBdDUFwqTVwNiz
aJf7t3eLwiyBuG93n1ij4lH7IkAsft6bFg1LZzvob6+a78s9RPgCnvugeSRJMQ5kesWxmIR0+9sQ
/bCmqchmzIkA4A/xnrDSvY9JQOZ+XXAw6/Lk1pH5GNGagyeflArH2NRFinsNAcV1Rl8XvZhA0BS9
Rf51yRvZ4cuu7Q9o60+rbsZlMKjghA0WVA/FqQkWjMUjmphQUbPBhvDpqHF4ElvBb1KmlB9YWAd0
nw5awVgeRIi6yp3gVDuwux3WXQNDwlwQ7fomGOqLl2b6I4QwP90/o1mu2J3fxNXt74b6Un6tgnFm
CJrlwb/gBiwOIq29WN5YQkKHsJ+S1hF9JUgkDYw4eUeq1LnHePQW5p94RJTSpfWtmYhkEsmE05qw
4Im+XaC0YhVrkIIddvlxtsYazQTrxNPpqT0Cw9KiV24sllHURrnbi7npeCNXCjpZgQdEkCMsmI7w
O8SD1yN5jInD1mvxGE0G5w5EhCey8Y2UPlsDVErJHWprIRNjupAz8d0yiCgxCKRJcqA5gBQ1xtz3
WPS+8yxOoep8o03cxvy+aO55kJXcMbbP3HHKWJKYO1bllBmWI19D5z9Avlx4e3xJn6BmfmGNTBxK
smTWtNyLaFIlgRGaGj3k/w6IYzqfWSUZ8Jh/BpwbYHyYGMGOgDOZyDb7xk64Wv8+yZeNMUEFZKzE
D/zrIntL0OKKisR6H2ErRga89y/USyDXbBsxAXo0X/HfZXLdr3JYXfS/pR01OtrdTZAzCt6/EVJ0
sfLz+w11NtvCTdyAvSK57TimHQVzOgvLQ6z33iBFdPf6+H2TbHxpgumW5nWxDCgICu9MpWhYf2WS
kfjBlNQ1aAabm8hPo7wGBu1InKXCRTNSd/l3Uw8Mex3bDfi5kxl02BVChGF3XVJ47TsSAQ+E5rL8
x7uq45Wg4AnLyLPh6ePfWmkGWSintSkVi/WFTBEEvoH8Tf+IF+36uybJjvidVeuztW7dBatI3X+O
8KTkKEk760Kx+uoGsMNn+zIZrPI6c0gVR8w9qJwZcO67Bu2UOpu9JuygpaGR5dPIYrqCNmyrbTBv
i9Sxh2JDYc1zhut5Ym2zZN/wLiW36azkE8HsHDrSFXIU5YcV0KYgc4zIVAPsYN0JftypsGZO6p91
pLIEB0jG1uVoFBDv0KKMS7NONn/ljJr9pVmZSZ2dMGdwI47w3pxf2820RKeLYCJ7OGmwuRtcm+5T
PTXjBj/6EAP69mbGaZnjQSX7mPoOvkLVq+KXKemyVMeQXaqZ2jAzdjsaediYldBaq+0ZiTN5yo05
vz320rCXIpH7nik4fej9kX+mIO2FQXccvpZC9YHV0beLZgtQEGjWb1y74ISA7l47UAGgHXCHn+6V
X6LFiwAbJVmvxMe/63XVe8Qe9d2LMFNXrOuEVVMyJKDy8oruMqVuQqzn30nrDKNhvs1kb3K3PTqP
7R5aFz6aM0XHXJT9cmhWjxH99U/ktwnBstb/4+mgLDeVmzPq5lJ0cXzQq+4rYBWXcoJAQiUcu33S
nNk0vPH0379q9rOfo8dY+TJP2onID5at+d3yb0Lc8NtlTVRPmaakMzyp6wUc/2vUGGZGizTLkzRs
4WnH75w59PnUhopX03plduWlenKZuiG1J7j2js07i3xcBuqAq0FJiGuOzNE7ENUMPJNvDW8zomWX
HE69bQsFINDujh+kVpG8CK5cv4reSchgeP9UbsKj/CL8GvCpP5rjsqIX/kcgk939ykyt/j+6n6YY
PEJ8M1eRzE2S8nv3Y2si3uWX/vMYMdBowesB/qM2+0KUycgAQMSSlSB7Sap3cfJt3hApPaCvHw3O
yk8Qi9q7RGw7TECGbxd8c99k6dOJFC9u8OsgQbVcDS8wz7Q5U0sP0cPBXhhp2IL0PFqTw5I1YGPT
RkSBsqCvEE5fgC3TnMTuxIxazljasndj/D2ItwhSXyD1yCZPNECFDmskpbPgQ45jghGJsQGInFuN
c9j8Ylo7upSP3CxuNpAqp6ySFK79yAHdbgd2CIBdgY8l8wmQCeb2AnJ/soFsilYX3QHJo5G6yFDj
jTdBENYtu1fPBzIXG2so7IaGGNO23YyPoyTNuk76tLgAGEns+4GR1XnvQQl9m0D3vf4VschO8UuV
cjEkdUk1nAycmqGBfiUJzU7Z5kni0o6psat2FgYtf2Letp3ezF/4LhDP9L6mILqgj8VwygIUnLpK
0QSpYuql0TTOpt/qC7FUTtoE21olL928FCcZsyIjskoUMuGfFd0E3M7CdxHxYM3rT1+8gtW/ZyyA
wkSEBjvGaj2l22qI7wB9YZ7AjsjmVOhk0FUFPgprnxYGkUbVmNFU+KIXG2A2lOKy+bX/3MD+mrIS
L7MwQmsgegxvpqjJE6Md4iiatQOS7+vsJZbCfMHEuDXEIiKu/3Ls9x1XdRNFGTPwmTkSum58UP2N
7A7Vi5zguHhD+qOxN1+HrgTEIWgQPHJhpQ85F9kP9IH/KK705UkSYNLC/TgC3j3Iw3coADwrWNCm
I5urJbpvFAMaknBRS/znRUGCW16a8DOOmTmFrYJWu5pCkTfEyemFpbSSz0QBjVLxZm/yCyyOqR+9
d6rXXmxcPqSXyo/zVTCeAtoWiH0yY59+hBrEdFm8BraVNO+xfUopJTzcthLbEHPxHil3lEK2dLW6
3on8xy6gYdIAAEimpFseLkITqfKYwmSl8ZlISuPoAEmrwpRM4AWq9WVCeRf0pc6m+iqeYU0X9051
0jcGMGQ6pMtScTk2NBTb50m2BIucJMpAeIu/nvR39JhCrfViOkM4tt14MKpCbvCPfJmWZvQ13EL+
jDf0gZ7Bxo9hkljXs7q+ZTGHyjfJnLK2uLFvitZbcU5WjBCBZUAxZZ4Kmwd5MNCXmvnkGoG6ApZ3
I37EG1rIaX2l15n1hIOq6O/Qt/jcyUK3Xjnkck9xsaZWWU8IzIZbxxPEPxn7iB41RqY9wFDYN6pX
JwWCMCsqR0BLXloX0DF7KdmPzrtcqZJaVyDC5AuTNRozH+InzSg8f8rhGrnk5GYt3Nh/zO0fqnc/
kiIkTib6BH4prplxPVwkbUCH8MzlId9NZUODpIWbWor19dFi1pHa43cqu9S+BIL2azdd/ZAeVL3y
dVGFYEGMs0SltIFCX68FFejy6OKCeYg809OFG0F7NlmDKcUVwK7sj+nHoMH1RZ3XlYNeXOTG4YFn
ODMSwQgfwviYqzfI2mxFkshcah3BmPyQ5mXT+ic2AAYlEQbFFnfs6MHm/kd4ImNFf3+hRM5PAFQB
r5xOlKOTa2rXqknNiEt1X1lXt9f/Om8QkJba6mIdADPGHNWeLBDPnpgTRtSHIrAMhgHQnUZNc7Nl
TJWxDkhbvrgWuCwXWFJ6GLXkUUokzncWhiqyWqcAG3HT3gI1zxUSO7jOI2PbIaWyYdhg4c/EsyLw
tNm/d9IW0wp+Se+tnrNwSX52MZfvEmI5bxP9oFS4i5RkAoHAbd5a9dXYYBkGtzpiqNo+k7+bqtlQ
Nhlc59NRg3RyQQGPuVE2ekJKMd39f/uguwSdfIEk8+chic71TL2TlCD0JBq0kTkuVjWrM1yCbFKJ
A09ih18C/ybeqZd7k0OG9kibhd2HEyTis49+pOFGP+DuXj4Btn1lYxJ+270Ewt36uujnBbKlRVXL
QG7tKM8gEmSv0LArrraFWXhLVbKsnai/9I0lQereRto4iSAMoFqEcA4mSo0tTHcXuo6hNi+hkuOs
s8cRm3Z9HS7/6vJi64epEs/rmYYkdaMhP6DeXLduhsAxwbR9vJ41rBsS4K+5HS73ejHqF3rjQx2L
fk6EydCvfwKvshp3YIWuUf296y4msjYu63sS1j7eY95EZ+gM+zXGunzqc54pVc0DjDK3sJAYZyIO
v8hxM792NOGrUP6gzfpyXIE56rCcmqZpS0jL85KMxYpJbW1nKZFILGlm8ThlQpHuH+XgjsmixRrw
o2L1Ns/bTUI9RjsCGulsuGNFrJBbroR7gBQu/kSuOVKjlawaYA1GXiI0cpZzoW+EgDAq5m80pOyT
C+4OeHecU9ZYurHunnR/+VcMxx0/I9L0rqYkwr9/IH4uoC2t8mynooJmiXJVwqaIN7+5Plw2+hFF
3cT9FHF1VChtR5T6BIkVpPZnZXwjKs5GQAy9VEhPojec7GbgG8hPTdV/E2eBi6sU6P8vPXsqdM1D
DV+iz00zNckRUKtHP7lH4kAX8w21OO7G+SYoTjKK+I4oUaPfQzSCOUm9PSq1BqQgI4RB5zdtY+hb
rmozZzYZXn3uBOwTjfOvvrKUJnv6Vy7ITOUFX0y03Vy3I6/N3PJjBNiVHDoL78+yrhQteWGHbBba
9PmEArfDGKewZZVn4PSL7lrdz7zcAhWSBW3sZG580azhtOmrpuq2amvTgKHF+uwYORPzcwo23fJv
p//ZY+wM7vI/RqUfgUutp60+bTcjqJcEX6Xk/PNRFwQxXWDfc0nEB3vJBNNjJs2Uy1ISfPE/+CLA
XkSEgJb5K9ThgCbwWzscGXbh0Kw0fkYp1xyYp/HqiaZsKG89XjO+FZI90VdIS1OSnL2RznhyH+3B
1JWUEhH6jUayiLtvI0usjCqIPuMv4DQzdxoxbP5NrO9Hl7iFRAKAPIAJWZCYf86T7wdOopS2vEuP
v/CbRUekZW7EasfJ2lgl2MJtuSB5Rmkgxl/A9Og0j8S+v/SFNHipTs39P2SLYyh4zwwVFZO6sFD9
681t3zfVWOHVOS8xdQUAEb9QCqDABJNpQbnVHcEKg35iEvszUURq5qEnI1p3F8MxZ7Gzb3WNWliR
CCSHcuUKMrBSo5oaMfqLw8tJ5nsd4Qz9G5BWiVNEKIND55BriwA3I7ztFunS44DZuo2x31JnC0F+
/OsTpzHYoDDXemVKAtO3LldHE8t08KMguWR71Euxv2s9m+X/OorWvZGDVZE10HItWXe9B9YIin2n
xaaprA0k6LfDJYkOshVG6E9FLAYu5N8NSvRMtDa7O5kuxnmAnqhNYkmXMbL0y+fcVmuBQIcl0OqZ
XeK4iiepLXvbmnQz9hVOrvbGwtPxOq0dPCCaKdW3WUxlR5O4PARo2Tm8bz9t7cSiSkaTtTJOUbCb
XOisgE80VeBgo6t82HrKPqLL15SAm41W82clsqu2lTGnl4EbXvl8jWbts6LSu799dAPiVFBQiW7U
/pYYVqVkgVX3ePN1982AdiCvusoNlRE/qbDxdN8mPuTAM3XZzKKTuM2O+WjAtEdG1y0Q4ek7AOev
MuaQK5Ho3WkvNXK7WCXpaOeOGwBvrpNtWk9eJCFmZalvBFYnZuxUe2Cj5S1zdzIgxqPY5fgVg2Hr
ymy8GHiauKMjdm4lqzl9iQsLxUzrVjht+JaTe0Ze2SWWbHx7ic7jVWQRn5wY9zRe5nSfPnF7YpFL
NUF0kdh0+J1HePArqYTcIUuayGzkbKYov3nYWNyLkUn90qUa9yt2um+akwSbbdC6pUvZgDTSQi7X
/13jHM57vGCawnRq5fOnWvXS3bt558Ir+Zpg7EQxHek2DGbaWXB2mXcIXFjnIvc57v8uKTXCGNJn
slTVQTgBipTp3XTk2zaJTSDGC27uI5/FzzyIcALdnFn03+L07RYFgksB5GFmJqJN4TI30B96V1Sr
s+c8trbumtqDC+UOkXqGisRsHUzwn0btFzFEzVwpSAJAXMSBSu6+Mma+ThV3Q9foUpSGMqr+vTt6
ADJRz3vBiTqHhMcAnZSklm8SuWvn8eqySbWvsr1AMtGQzrueVTSaclbGT//5MM8FaZLn/QFdTWk9
DCSUtS9yO5kjB2ddDpq4iJl7wPbzTCWiGML6bZD3kVPdJUU3CoEr4kwIl38U4UhEwcGS7SB+i71I
fWY9mAQhhazyy8W5JsSM6eSZQg8TxbKmHfwkAti+EGe4EfO6NqB6G+eZFeDkBYXKCxksMVVVYmFQ
vauz5FohB6nirqIc+VSp7/PfbMB1zcjNpSmaptLXtZQCHwuiAc5cdS4Jps1DnHFp/Y4ubopGXrZr
9SbDoswhNSrTR9PBbBqwRqN3Yj9p/+w/82ykzY1WJrgIDYKKF96CZH1o6CPGvqmnYzmsTe3253xz
CpFaTf14Tc+1mYVVoK1yvPixIFiU6odLb20kn8pa0arJ1z8onrQALBTHTylJxYgKTUv5RAIH9wGx
S3FNN4yW+R+s1UVTSgx5LS+9kVehdrYvrdgd/92uVFPJwf64qideKufHla+Y5Fzo1zpdnYBhP1Le
Z9M2+gBExEpUZzL8CSC703ntM35mZbXmqiMNs8fBG1u2hXjc9CTnGwwvxnglYH1+lUQW6wMr77p5
LwsQTjpkSMKNg24QyPBBLAtLDxmOdYe+YQgl2fVy9v5qYitmlujZ1pABglEMRCik2KccDjttgrRo
nFgoRQFg4OMEkrpSaEwRyH5cAzwx7/+W6azd+H31kdY1KYfpTQL3fHvLfUBQiYn+q8VLNv5goN+f
T/pmoM9pYs0d0eTMNQhjMJciFIy0PtZUrZ80QzltnPjCfJIfJdGveEquYPc+3DkNg0vC3MF3vpVi
aJZwPlnXpENkJ8B9r6wAK9NRxgM4bZcXCFC565sYYxZ/IbY4oKvz67uwMHH8LikXw+DxFqDqve3d
9EDoU828ck/qOTB41VYDSYSx6S0jeLZXgcebO1VYYoRo0blxilQms3+PZXoCmWw2M27ndiVmMlXy
Ykt0gbKju2RXqCUNra50ahSKq5JeNDzE7zpv6BvqJ//3vrfFv6pf0Jsg+QV6kw+KkdKrxxuwpMnD
kn99bOES4nmIcrg5RE7t0Pil8BKeR18/6dyGHL8b8n+OHal557qyhSRz1gyOLmdIcDFh/3puK9jR
ovOx0Irs4RYMhaLEKQgLHajXd/pERXGa/v+N5m1bWS1BLN5G0oPccZkfkrLV6UcFcksypPLlInU1
TRcB9LeExkZI6No3R+Y7supDaYhZ40BNrnwuFHsP2ZkHTEkL8A03njTenAc3Gq9ecYaVg8puX4/u
d1s0RnZn4gOU/f0dJEmJU3Vw5YfoaQKtYPOEIvp50ed/VrNEGiXr3NBw8bEJqxLgvRPzCUtgiXl/
LuAsvi97lviCgx4CnGan2GULBRdEmnBRHW/Gh1oHEi4DDmI5Vf3eNrUP8YIvuN6h2rk/SUjMYI7b
RygPYNdVAOEM7NVFUtOQ+7p1vXJB+GyaQDh8OmXgHaHfeukM1J4YYH7C/kuleX2dqtFfqIuAeZPl
22S+Yhag2FJi/4VAGAIZ7kqtWKr+jZMKYufVDnhV5JCS2tj+DudvgHg6KW0mOoBoNBz27NdhI5HJ
dYUFfqzLZ3JHsJfCMY5JiK65ZlLzytlYFrDw9auVE53tJ7HEW/ZnVugdo/qAP9gKyw2oSveubeLm
psGlYkAQpEpV80x8Cl1vf4PoHOkv3/R60qxXZDnpzJe3KRENLqUoKeubOEWnwM4RyXPy3EC6tV7U
O8HhZRGdbpjzvidtUJXEojemB5I4COhLsu6KkFcCzB/ZaZwBHyoGaxtxPitHfQNkHWatoQXJA4up
0w/I+I6Oe8tQibBcxruaFWHKtr2odxzJPhtUwsURaAVZbP5hsg2shu9+i8wYQoXftF3fyhu9Y2yw
dMVLB9PSh28jnOmBVvhIPogNoQbmUtwut7z3M64lcyhb5vHUT849QZEGH6U/Btgb5crGLaB1n7or
ycRv/497ra1U1vbQJXFzS7xjTBCzXly0muTqNi0Gn7FFrTo4X0jPEpeEvcUya8tKuSl6cPiQQHLc
m4z9KmPjudQlxH8h0+l6Zs6LW4Rr8+1vLKrrDLE4/a+FwKeUArNSUGQh3Lmx62GY9fBQNUq7ckI0
YZ4uiEX/p1EqQwXXzJeeGvhXJacVC+TYVpcpUyex7ooKRMtydPpocYD3pARUMq94CFNteuoSzjUc
qDCQZ1JEPNJeNhEC22yzYn6xd983k9MZ87HcqDtHwHMb+BhIqo3tbdndblkgxsP5IZyD1NfdxSIi
e6MEUbaq8BNO8uglF5otLNFJ/YXHxNLFvnl+ZNCBp0NI1fc7syQkkRAMnQiFO6HHSzlyuC7i1/5u
tvmWQzv6qHGzK4XpBinAHPaMHe+ODL1Av0Dful1uSBuM5dL/CiOZqlEN+nG0wd40+uo/yjAcDGmb
vl9S6sggP9mi4mUJYKyV33s3tmz9vmh+KZ2iLxcBOhpCJtWbxB8qVyycbL/T0gDtWF5OQL7MjBix
rb6U541R6f9PYiFYpkEYMXoAqQk2viiXlfyrpzpUsLU2LLADpFev8jNOQtNeLddZKK7cF0z1Mbu2
+XXz27DsCBX9Uwd1ZLMzjTBign57UtZOzXwPhvi00z51TcUALX7Jdjj2MyMUoRuV3JSvImP+4Ijm
dXNJ/fULq8hM87fnejO56EZCf6K5ho2ZawTvvAL3/LWCIskI6sKrwNWWAnqjM6tYVb5wiVQrTBU5
F38nx//f6bPOypunsgf8XtKWAaOC86rZ9SVzvwQ3/AQeXeFX7nI7gSZdUyMU4zF285+aJrzlfTWM
3fhw3II7b+Odjj6kO/ACI3E/5p14uEYUSXg1ybOpZ5he5e2Ac5c9PV0wEmb+coNGFYqlFC18zdmj
H4usjjRWcgs8JsU2ibvctaqP0m4SxZFF+2hsz2DpAtZpjLTY2RTn1HVK6XTSYWwdu6u5ubEXZMHH
XQQfcHflPYmc1SX/h8kLo6dq1jJnmIHg5YRhH3K4Q68YVXbEHjPvhgGHHglyEcZFpRWFBojLGHbl
aePzF9sgjHPYYfcVBildMr1beLu+cklAsM876Ky0fVdrqysnjAYXtVvVgFYumQsfBPUZu6qfBorZ
wLbhbnfURRkw89LVn1ZQN2YlVJgQ/plIWG2TXCYs0ZzTzWMlLfz1uSBcYrpmZkRQ4iCVZT1iiuBu
Rbmv4DNtXuUM2S0lB7Z8mZ5zuWtqXLo/J44fY3jGX8r3jjD7DgvJ2Dm4+9Kf2r7hUSJMIXtlSTTs
r33C88HdUwZu2MJIDPEu1fziLP9IfjpVebjd7DujAPOluA9x0s5Lfatskyw9AxQnWZDOOEuVBzSP
KbmriRfIhR0ztQMfgLWkt7fTmyXXAno6SwxBlv1ogGp4gwXKcHzfKArEs1tGzPT20F7IzEUhLIbP
zUmMmbQrgFSDmlLjwMm7ulw3MJEtZSRk04SsfthCSGXGy+q+u+CCoNVTnsE4aQD20wDcHEogEcuI
V1qpwdde7d6H9ZW8T7R02LT3CzH0UwnlOfjV9KgXYZ0MMRMmwITOkpCGjvf0PEzT+AbaSO/rkhKQ
WW3Lhbu+UfY2lXLCWaDRhtSgTOY9mOEwjDMw5Z1T29uPdFeIq/+C3uhLxutbLq5GW2Z/RhE/UtDR
hmA3W9DO1k8u6UOeMRqwBAtaNXRpvlyl3GJE8SHWCzKDLURxKZgZzRlG41PmAOiJKXtZxWTLPD6B
t1b4neulGXUE6PY5Ouls0wCr+YYjuyF+7bVDnIQT7Lza0TxKPPfIfmfIrynH57qR5kltEjbRwkYR
+wqzDEpeO/XLN1rhjY2UIzIZKvZMyQuPF4Qhp2ZI6p3+QX0II5Rw7H2vSB3w0uJdE2SPEemykpJM
3Zbpws9GqkHqX10wmGydwy03T7lMj5jAdFBwkIOJV8AQG9k24K1n1e/mkTFN2SxxcctJSIrwP6bs
XaeKoZ1U+DAg01bM8w5GOeqeJ3X7dC+cpmiAsSo/NCOvQqz3hdGIfmITLKJV87/VDMc8ZS8xXwiQ
Te/meiTC4myVNVZJyFRfW0uYFGp4cQi+VcUTt+ID0vRhmgEOsOO2QEFHUH/P55EfvGP7ovMyx3CO
edlUW4I0BswGCnuZGfCkRh9CjeB6sfKWN3LUzWIxbFCIm9+XOM0ZaUh7loL+437qCy1s5mI7mZIA
mSdEIiXcmmSmLkS9KXOVGwfLr0nKEW39DxbI6lmku7teQ64GiwBwHZWWehmLThiP4a45DX7u36gt
wp1AyoXou8b2pS/BDwBUdwE4EoGv9mBQ6KEoPU/36OnYwaRG0oivXXYCoALZFbP0AH3G34r8nYZD
PNda7MCY0uOp4PPZ6zrRQvmvnKqL6i8/ossOeAst0LrHZMPSX1YDfW34pnIX5DpZKi3IT3Qwfu6/
D70BSd0u4XS7eAKTiKAuEPp1HJSh3ACo9uWhM0lDKSOxOz4WewwsCMGmq9dHrXckfAfZvJJuQz6R
gl8Os6a+ltdsZJ3BS5Ig3pcPCi3dowOICrIAfeq3xWZO2e4u7+0qM1UqYWUgo6jzkenWEFV03naJ
iRNfjmDg9LlhzpSLTQ/6atjRSiKJwZ27e0Pma2KP4G/AQA9vhLXw7BJzJJtt1p34ViQrdP8/dAtb
YGp+bro+m2SaCc53h1yKh0mpr0+OH14WuA2oDfUE5kHA8BIuMP45x1hrD3+xbWcn4dnu/PTqeUji
hNB7YH7JbTU4GEJouqYcPxQ4FWk9+mjhdgtIwbz0sgLxHcut+y1SlbYDQqAMUsQe26iFQ5FuRBao
ubOONOxS0WZclmcri8M1s7uHpGM6RwUHSWxlIt2IuUiypz82cGFF1EGSl70mDvzHIi1LSfi2W98m
gQ+7DDps7S2kfU2IzSx97HoEJ+RTHgoyW8QedQS0L0aP59FTDBIq32XeCQmXMznacV7EQGkXGGy6
qNRaHspDBPASZ2uAh67qcb8YnoAfGn+143qh6+RrjRtOjXC7lPVMvVSFSoMdzU448REfg4zJ6VNF
yOWpxtsltCaX0YI+RJtzg+7ZNjWnJlfEXCULjJZt3ULLuzEVujf+V1peWx0MdCE5HKLKks4u4Dw1
CsvsKC6YxYWabBtOuZdizMxnuJXGUU/Ncd26/mi5JWuFN8yYRkvPEDfrAWAkZSmyDli1PBTAOJwK
mbmeH97zUlFNqjNtnUnzgOhnJfj+KHBokaowY6ClwchWLbsRozuj/n4gK/OCRWZJJa1tdwiyMaFd
3JaWfWtt+fhzGOLpKvKU7q8qhOTMp36Wt9vyzAb7vwGVrls9lPdRkcu6maLfn/i2wL8rF4vnmi32
/zqFJW8/6T8vgufgxKyMA7OXXCBIqSjKlIzxBpN5fVDVXt04n5fvy7lNInBKXhP5WtBjdhNTC1Cj
b8CGMvehTm86J44n6Fs1nFb6DQXKS9jWpSl69pp8mQTp90/1DZb1y71OBfP9lZtVsbSZ069GN3yV
gsrEWrrLoO2hVlvsP45fpDfM7jGz3v2E5XqnzMVKzcU35bvvSTNLXJbnmuTWSGorm0jObVXszO4/
jzrNBwoP7yavCXhUazoBFQqbZNMebh/iRWPJgyLCyrw2z2aWkOn3wHhdNpaivR8ytRoqcTKoWDw/
fN1RzqLd3I9WcnYFJHjpXTH/36UPK3uzTt/mIvJmRvk8y/g4GsQ6B5BRD64ZbGT/XxUnUm9SAoDj
QQoVYu+QhV3qvlnnzRxusqV+3WgMZlKZ86alnESLNvjLGzrr3ZiPBtRBjs9HXhI0DxKkVrlpXDOQ
V+U6DPrLLiN5on/HCQ7lTEkxsU8GkFQzvopX2U3JHb6mQVvnh4XuGhcJhPOrytqrLcwApk+jZdYK
mFzDigxkAfkluksjtBnqUBmwc5WIM/VcOPkV4iO//QsUdAV26ruX+f1szlNR9cheZEssaTbloT5D
NCbjAyocpCxY89jFVH94v3Tq1n1GUENWnsXt8NcaogehAkGIt6aPj+imau2k7/GVLLxh+OWDfU2j
Uzy9xNUW1xDZsvO8RnqRy2EHhp8GdiZhVdTrvW/PeHGyPXXPPelVwcwU3fntTrCZgS3QWgggKj56
SxJj1AyPPa5ZCYyd1LKjy+7TnXPSEfneUfpyhVLpHXbmQXNKsW6178ntngn8PY1bhmQZX95wG2lm
YA7Ki0IxioI5gAGNIK7pRl94SmgxHm8RLpxm3s5/JaZuj3EeuXRNuXBdIeTLgsLMXucj0gIlOKpl
Cnh6Z6O0H/xS0spyd8QfE/a/l6O9FeE+0ps7qe+uVzLNyEoSRgUw+wGI95bf/OMNb+f8J+eVevB6
gPqrVdWPtLMv3PrUkq/lDgs7cmg2ytsRY0KWsJ1ArhvXsJiB+S5U3Ng7Pmc924PLZ6GFvdE9xE1G
B2bCDzhHudclCMLMXOe5Y9cRB23s7E+IxtQUJdZOzKs2jkniRnp5oi5h+cMrRfRVWF1bQyFTb9PQ
JY2AvJ8Bxt1v2jYHjs76GJLCB+/qsMkrxeFYFCowpsVAhjxCMcIEsEaa+in72CNIk9JbKC8a21b6
qVngGswogcOMqCU5ciQ81SjyFBGaAA1blxVTD8HE3tPqHP8YRk9Xj1I19D4WUkCuNqrQFNcpA6HL
agJH7Ia36ivKgcKozlo70gsFMPL38NELzyv+iZPJAP+iAG02thULuBMEPcUOoknGMePl1DlTzsxa
eE6ChN7mPXEum+QwEa9uH5++UHmTgVgnzHlg0NwgJf6AzmeeUjD++SrrZwu2IspjjuhdqdSJhDiX
eaG2HkE2AhbIWODzLUBjosongoop0JvKQB0PwpdM0ySD9vsYrqKmvc8buW2p8w1IzB8ohBcswDm0
VEQ9wtM0i3v2URD/0ljtlRvdNihtOR7bW0XZHtdzEwDKDcxDaIKGQL4jdQRFw5HNmtMQJZu1gjzU
hSPjUtQ+Q3kT8y80+FAT0MgvaNE+blwW7WlyGYsrmvB0BiAQm/nXnU47XsrKGUjUVDUhbrLUe0Da
k/vgZ3bB8cYG0d3P2BF9YYdimNzSMMCy3JJPm+/9xEY6R0em+fRa7Vx0HXUAiELuoSqpmFNNQUsk
avnXEIEBuDyVceG9qdS/ztcNJnSF+I8Bi8+0GAEkNV0i5W3iEOGuz1qr0F6tyJo2IKmNRbebH8eq
G4Q1iIw5ECIHF99c6rCyof50W9pxyxCHq4XwiRAo5kCA/xuz77zGZoNRFxV+h/x10emJ2gIb1YCm
UYb4A5znrCDC1rzQst6noUP/smgONBgvc6wLdhSlpKiEds/NOQqG4id4bKKn6jsa8iDwTRFxTDoO
Crzgy9CDKg57DKlJ9IOiev83EDzOZTsCG74zUU6deVtNq0HcLMJ9sTg+aNp9NThV5SJZZ9Hijx6k
hg0/VnkhyKdpX30FGtviU235GW+cvd0VajBZzQAQF7PEbJpGPxA1WSVovyr+Kg6NlbHY0ZFyCggD
JJBIfkJnx7tYwpK+x1tkXRCZVSdlUaQqcVe3tht97r6A/BDLjrGXs6eo3W46/1JKxV4H9B/03lAh
VwIdm6BtxqtP0OJBjUqO92bCfDGNsPYgbcEKvIV9opUluAFVfA7MUHGezkde3AnmszOC4PJtBxgO
YfCjwz9FyDyvde3SHHRZmmtAMyA8XGHx26SBYB2kn+FxbhQ7o+aKLkyylOQuC7Y0U5a5P6s964V7
6hPvgvgAqj7T1SpCEWBX+ug1xJj1aSlYXXQsd9O6vO3x1ls+XqwxEbcXtc6x0N78Tp0GXBESc+nD
luksi+9TojXe/MrU7nl0aw+fC/PrEmnojA4HyCfDSdH3VIexyifLZRL5doIIF++7Skby7EBBM/u5
Zo19WLnPL4LL2kn5QGjFcwM5RHhzriJPwWxSdaTg7H1d4VLs4AOSoT2Bbrc9e/47Lux+4DMmWpxQ
JfevNRCj78Eqk6+hxrJuWlnQ4SZdaxjSfxnOrWCfDP2p5HtlLkjFeTs4/gbBzVmRfrF5JmRMOvcm
gkhrl3sKCUdhOcRcQZUBeIFDt9xwQUpuzQfSxIvrxiSmR707c+Fp+kGUjEcLqtfIVSSWGchOmOVH
WLOBt2veHGP99hQD1CUaIhtBLdXhUn8bwhpnDgB2WHSpfbCsx6bN4zvOzNIG1cOdC2K3/QQcbQwI
EBkk91BDdNKVEwqk6bAohMNXopa490dukviEa3T/opkFC54MF9CrAJriVFXoyMykFTeuYsoiBN7f
nFzGYz5IhhnBMpbL5pXbeuywg6wW78dioEKqDHTd6YT40tiky/0KvgfbcT5IvmqCOXRVn/YPst9O
vN4T5FgdfRO1YCx/G6PxtJzrEHG+Sx8xwqhZ4x7NMS/B96Db6pwlrY6tAU9kGlxQU9z2c+kjOSvA
BM975ubT62yTifqzERalZLZ/DzKcif/p5mP6uGgw8hr88W3sffuXTRFY5yJh2ujKNdLHuack+U/A
Ga/Xs7kvCBzsbvmROQSP+IMnz1Xmxxr3QegvSS4oPh86F7IPqf3revNch1ka3p0iYnLiscZf/f5F
KAguT/nmr3IGDzM0x8jFi5f1LyaGGw++mefdDlCcAaDadWe3PqdohEtz6hg7TKRVRzn/zkLVuIpt
AAnjx1sNC8ebYwRx/3L1ZL224W6y0FoztJUYSZtGjj8unjqzC7PmQKfl4kl3P8n7RGfj200vT2oj
kDBCt3al+3gq1v6VRyGDbAe0/H7YWeLGnJUXb2v24s2/n+zzdP/Cmb0Mj8DpchKzylQPIc71jbc+
zC/SwoOA/HJgebTTFENPqBOF26kMMNPxVCE1r7UkY48GB2HvSW0VIfhp0qwSY8wSMZsoruiSlXjg
jgPEGdPjf6PG6QfZTQ9NH2N7nMiUGWlxzSWQXbWyHmtRjkmbLbnVz2S2SSGGQGUMatJG0FgEPrhp
6oPRthI4ydWZ4JYhCYBzdgZgEFHG17sbAWRjA+DDcL7RmYLvUYy0a3LwLk7U7TCSZ7W3BXv2ugmH
Pp1f/YfHVkBISZEs+3BAKfxQfIVOdtenslGQYK2kiqe3A9mKqsxwKAxFvYa9Tq+3gcMAaWO8hIzt
pFwziRU8OpN3fAC6e6euG4QbYcOYma7sv3sTa+C8rvnd9lyXoPNWDX545zh16bkOBBnmQAAu+Oz0
YliN97JQFlv9+IkUWcFNBq3f9A7SLgSfJunY1IOEESEld5+MB2emm+NKPKhB9jYWFWp3m80wbK10
v+LoG7CihxqTFONxt6zDR05/TTWXdMf5qe18ARFTGDch97QoVQEkMLTMWxhCJ9wBz5SKtUZndvpz
EUaS0WmERbG6imPLxyr/vAF+FBCWGoBhptEFRlpR+YnFJPe8zrrnQ/nvd4Ii//2WuoQEe2qPLS6X
F7+vibR5rHuYeIXs59SmYjwZNrx0pFhqLOJnxY1ETAQe20HMGy57D20mTiqKjxGLN/H0gdKLljK1
6L6sDB21EpQLxqszi4d88v0fKGMjKylvsdsd0OoKLZRsq0+Ga20+JlKATPq+A89IUA+RcOECYEOc
SpUuNJSFs+QeL0U7Dr1eJkHNgKwT1mEkuZFIEZRoRpIouXUucVxxBDKMhMRUKiLYaJaSec1gCh3K
T9B6lrK3XrmOxuSYoULg+eWz3GTswjcLeS/yie3yVuQUYFRVMvg0JU3cfZ2/3AaA4nnT2oT/HoDE
3uLXLJtbDf9X/HOm9TaOxfhQLqLE9Mc+sFLKCocXQ23nZ2E42gWgeAtpnOaicQ+hxSsofe9by50g
JNEDxNHj5M5EbbXV3FW6gSV1Xe1rTrZT8ndsDlCWaLeO8u/rLxW0lFQE1PMrXmXHu5Y3i2DSGv+V
j2iNZ8Q2MsvtwWgkJtCIhqm6ATgXXLZc8l59sfdJdFxXK7Enh8h/htg+235+8Xa9kPbT9ZaWEuf6
004kbgU2qlGlyiGLXRCBYE6/Cw2L2RlsCLWzg17JVffc8dS2Xxykyc/9UmYIzOzm1/greDwWWt2p
xLkCQ9S3cFklacm42Zes7GTEaV+TYau59BPdSjQAV4rdb2vO1bNA/DhhFkCGC2iQvJmQqC/9Otwx
9E5dKVYOkCWSQPdcw18lyOtuipICh5X+kgNZ7Wc0Pqf1pq8bme7D+/MMu4+6uLFnb9AvBS3MdmH0
iQxYhysWLra5GF8b2ynyBeT5FXzzOx0+D/ixHkekPqjTcx0Cnozti34xosY+BwKNGtXGb5YUl0VY
JueFcdpUzuyIFSMeo5jAwKiaPXWT3kjLZxAldNFFObV2c2/X+PXjXydQoY89QyZjjEa6JZ3LUbfd
9Ck0heeAGe5Tvv6E3l5DALy3SQyJz6NzNaO3CzWESi4/oWstTMk+XDb+Bj2djVQG1sRXA1tIJXWM
Cu9GV3Zpp+Quv3JBZ3XDrAdLCysV6cQCMV7h86R12EIMa8weoahaeZDo04hr37RJ7zIiONcTZmbw
UeeyeWwCD8tnXciJ0CQkXsj8HipfjEsjnyJStDN5wkyZb8a8ErQi1895ZNSzXybuVCKka0AzjHhh
G2ujr9tDZ9jJP2YiDu0DjPhUlnY2ysYbLd9VCOrYTFmfoVZKvejMPV2DMZzeGLEuaR0Scp8WNwnA
Cj2K+GA9OsUxITVIKJJpxDKSTFKjlHozVJiqQ6aX95kX9SqHs2n+4omicf0wzXJ0Rx9RMyWXlgRZ
rIxs+BGBuFaNSa4GMKeeaKi2wXyIbdLmKh37Y9/ylgZytPERgO0QwM1K79k+596jmKpYfbBlzIWm
mtapB65BHGEMP3bCEHR5PfYwwJOw99x3x8c0vBAzC6fwLe3YQu5qXl33dFaTHH2IHvwZKiZpwryB
0DreAWpSuNYCtmAH18HQmwRCPfFgAUhTOyUMdrOGBapw3YnGCXCJXH8oApwpkQY3ksaUTW000jzH
+PGpC2LW7FYF19IKChwvy6OMz71EYFB4vHhepJYYWIxu2EPhOD1mQ5oOfan413XLRDysQIG7LsKI
3evvt7dR79FqhYl64xtBrJsqBhE46eRVomiXpaNJ3ej5VIj+LH10LhUKgI4OmvxF7ACW90st62Np
e/dddDaT/0+IlxCC8xyHKVxuLDJ2+k+wclGnrt/b518H59Ic2nQXd1bxdbsWPLyMQyXT39yt9SXy
JRkWuKjFu5QFjPdXz6kh0yAC/sK5rmZ5s4hPLED76s9+o7A6igHG8Erkm0p/fx5areeN16I0GcQY
TkTxzpGrDcq12C1e5SJ3zHSEZB0ysi3BOYeG9jHRnOQsmnGBC36vpzpU2EXTXE55p5OA8ytcetoo
EZaqCCmx52bYFuqGJ+0dKQHwBd84o9n+CbV1Q9kN0w7nBTTwORmUt2f7G2LKcV80XENXw1fnYL4L
DO2mrI6msS00lbqALnB7J+xJvlqBzDAid+hUlts4IgYaB8wcn1nusBqqRfWdCjbaZ7BOf0j4DRq5
9SLb+fexv4TjFiNbxX6DWNCyUY/ton6MqfOQoxZdzfBXtwgjJKSfx2EVGoEC1AeTtgXLqJLH9hj4
j68IVfI3OaxBkXHjKN5koBM7HveEnzDzAa6+jixVM0qhDzUZbivhaFLUtOIJ7QTYEa3Iai7vPE+K
tCmomb3bs9sEEwB6q+ztHeUL3NKLEmnoib8ZtUicX9Q4dZ65wYnhw7fR5mGYKp1r/gcURtpTCiCj
7t0GxBz1TY/+bxVvUwcAw7O1uldeApwq8qLTEzE0FaKwJLSdeSC43SaE7ocvc7/9iZIlc2lilrYx
xMr1Tn7YyJ76CS5wKvIe3zkA/ewVq8ib2zzkCFwT3SkLCEAEsIzq9Ss0KfXZuCf8SRSThCwqk0NN
km/yySiH0ao/h/Bx2dNIZ7ZKNceeZnfIxnDhNcjUfhGFjP+n3mDx3wrF192Z0XJeePzPUgNtPoQy
aPh4ha1kQIlbM5TM8Et295nWKuq/rsSo2gMWjbmSFK8l9MsDXuFuLRID9LNQdD5yuGd7Ymtho/7x
hQOL4XhNAk54HZnRCxzYpw4pc/Qdxryx3shHgloCQl2as81reJJeN2+KBtm3SWlNY3nzHn8m3btA
gtYC1giCCji/v07t+iq3UMt0dbsKRekDjIYXI0YXDpf8m98HYVEnpgLJqb2TLYAMAMRxf5IVcO58
i3znnn8R1FeB7dXS6gGk/jRx/DMkKJ1e9LZhjOreyZUvu2pk4YPH8wTgr/QGqySKAva4VWEuRfXh
0nHWmeKlFb5kUyzkk/uN0h5KduwrqvAkZL95WN/GkwqtAk2adA7XyMnaSRqMcaQYnYEUdSLv9UiJ
svgYMmblkq/anPZMYn2XusOVSmJyhT81NvXfz85bsDqtu2H5mBK2Nt81OjHqpe1quO+pQWiPQRIH
Us7X+S1MR3+bBaxTdbisEzTOkAAawOdBvo5uv34NRA7KWrwKH9VKC5SM4bH3c1wJCIBCpkjdtTv5
OWwvIfYVO8V1KsGAVHpssyP7zYrm5U24sTdMZti5myNSZ65hwW7AakdU52jHlXoPsy4dpLmjmcdm
BjlWxD9Rv9LMHDOUyEUsroWWUWG75xsF4kA7eAgLD86sHRzuNVQmR5W0FhKZQYdGzv4X/1A0sI48
R/moxIw3x4k6zI5nGzpzKuW9f8ZKY9adbVgsuvAQCtCrV1VEAMdzNxFuw9GdcrQo7uO8CfjNWfqP
W5+SjQC+Mfc78pa93LJzZyrGE0v5PrND/LlMbD5hceuhEuAdSFIlEfp3jwGs76+BNfMa1XlTELv8
Y9d8twl2E5PiYQTgF2GWCFLrjsdyJMZCYZ5CrnnsxwM0kH2msdPNOTmjmgL+/r/bu5sqcas1ursh
ONarSwolxfxC1MQZc4GjaKbfwLqYdIxe17OKZRpswVoV/EyFiIbIDmdxPqYNKjgAUBtG0nl1TQUG
M1ruJ2pMNebGk1jFq1gDLuVLdP82xAQgBLuFb+WAhDE4hz2jXl/4vi62As6WJgwsBQ0rBPkqjhi4
agciK9IZ9B7C6cKcMhzROC4qtOZprppBMdOL7am33akwx8LBSE411sVfKRqw1RBu5NAtMc+WVXa/
7hkjX64R82VE8u6s9AsjT4KDRYyhKFU8nQonm+2NAnk0GCB6v8u3ol6cPzeZwjcJ/RWRbKBnAC77
idNVvvqoYyD42iu8T+uc7Vn3C9eFOfwpo1CuGoKbw9z8MU7AlLaPcGbJcXe2WcTnaQvkVSxq69Bc
bZCJBNmqKDtV6CoHvdKkv+rP6TRPlmyekZoH0VIUKVbpGTgfhJDaEV+oW0pMjlK+oc06fWduzQqr
2WjXX2QGvy9GHtQzs28Wo5ZIlV4L2t05ky/bE6TFcvhpMvFqYvI08oUdFzyvEYAhENdOSn6t+DmX
PeVhM1K0lXpHEqhHfqT2Ge2BEdbDUI6ZWJQ2ICNGtMn2chQm0uoCk9SINtJ5CAEgJGZqPvgF+G6Z
+gzl8n5Onn0UwnUm8D/2OI8rCDj7iXx9Lw03a64G0L6+oRvlyPpCh7oORQt/PqADWJAW4P+wmqXJ
AP3W/KsRFufDoTTt9I3yukmkMZGFhuak/dUkeQeUMBLo1oiJe8/1hM4b2zGxxTcepteIrh0lA4vx
RvqR3VfMa131L6Txz/NaFKm1YaktTkKVrVn6vRUoa50Lom4BcUC7UPn+c8tQvLU+fVAT1sj9Ou49
omPXezMUikwCy1JB4x7qzIC/HqApYOivynqKk5Q/vllo1gpwPMSmVr/qgeitGc1n2UzGnm15GZie
rbQZY58zuNYR94CVxrxnvY5lbwxgcp/qySmPSQJ1L5u4DGCvk6WVZe+mKU9TGxxwhFIcp8y3udRQ
MJpEqN4YclltrmAKJ/WD/kjToiCtjagAvGLEprVd8WuJgPbORVxtnsUGilQc9n/yiBfeKS7VQxu7
aVRzkqUQcNYhQLdphmxokYxYU8o/cDKsSH/TdF5xGNBvy+SiGYbSQHKEfuWLoqNel4CwVO96OqE/
PWKbahT1/EdVMpccAnWjW3rX0vEuSprkvzVePIvqdbdA4hAztHVazhfAx1mCJKyIZUBsBug/e2CD
Xk2EmhLKtnMfS0PddA2wwagoLenUuktBpv6PmluuQrNnAgTo8QbCKYQezS7outf2bj8zWHfpcfT3
U8Eqf3VVFH0GQdzcB0n3V3kJZCfk/HSC31ty9bicLAYwmjpfGb0/DmQms9/9tbuMc7JMTqNEx8on
PW5k4mAc8n9DSvq5z0dEhyH9lzVFslP4/FySPzVPDL4o4MlgupdtGFQM3sdKgZnUMopa6UTm+R+v
wBaq7yl3eOlt2A8fkMamUi/CcdRyQ3mscLo3fC2ChO2KMkRrtlMUGTWBmimPuMPWPblqJ1jcWi1C
ydT5x8C8LRUchDthzgyeLLzO+KpSqT3K+TADkbY+8GCiDPRJQnEgb7BIRqTOTVJFUl1O9D+Shrmu
3mcJXdtINAyUtTfdaX/men+I/iBZwo72QAgjjCNAPp/9493Khw/3fRC+SGYaamkrEb+qZ7LUgkCZ
c5XDvVgBSKM0lrTGTBmcUAk+LS7FD7Pl5riPrD5CGjz27eGF1M+x8eVmQATXqrc5HxfvPDREeTnf
+8VuvAGNlbrj6Ja2MVFedSVi8Sw5H9gBCcTtoE70z5DajlNWt4B+zc4weYD50T4r8ujDn7mQ9IqC
TSjyMdiwzOpWgGj62fNoXQhs+9E49BNpRLdIApEY4Gnf0wXd36trGcIdRijoRFgqtPcxLD406lQg
6bpYJBwrIB7lBOtjtFkld7hf3d6eR9vTnBjV4QBzDPhRj+tdsavYxDFGMd4dNgLKMR5ERUUYRw/k
mxP6m9iXkyGypzw3rmzq3B8lpH+2NzsYnakP2bC4MOyJhE3HlmlPXvj+i25fAjMtTgmnAj383y0J
JDGTbanosAgtCsXYRZd1HoAfOOK+waUcGOQdHzI8dst4v/H/W+lyu14BaMZbLLldKIo+qYXdDToN
RXWV2VMcR25k3CZSP6HkulhZUK4irDmQfkzuluj/6GAIN0a/vE5B/i/FR3gD9uF+mdQ6nMrwIBK8
4fbJmzg7N47EM0U0Aboj0RqXA7lKGC7zO+6AnsjpU+9ofiCAQkPux0hexG0uJZZ5Kq1AH2WdtHLv
Xcr2k69iRDPZlocpPMpq++iyafv9q06YS6mIP2iVTFxSFR/eTGXTk2aa4LRfEnlQIAWwbqIajSDg
NQJy4X/N9zqvlVHeon9lU3d4VMZ6nfPFgs2Hn5qgBa5ahXRIKdX3Qb8bhMxuX4q8S3Olzvu6qbRg
rjdJR0pDxNNEjctHEW5+UU5OFgrvLyvrfZj1nfLEk6+s+CAL5npwyRLc6ml5cYLNBn/5wXTyu44i
C6lb6g80KcCjOcfHsCH5g7YxZrZN6Pml6ve5FIiyDRCufEQZv+qcvo3ZAMgGKx1Y59kaN1nOG38g
RxUtYh3tm0ZsQtJw0X78xUdO3eAu10H/8DKmymY9ENfuOvr7NK4knIsjgk7LJRUcA4qZ/Vg+6Wz6
x1ygPhg96Y/o8OTnvaVRKbakV4bme20EVQ6QQo5InI44kMOn3CztqQ7zDBJaRZKSeeEpKJURv2qU
bv0v910ycHYNeCkCz0cj5o1n0fii/jbjP1g4kFBXoXBnV4AqSk8n44kqt3EewQb3pauiplH7vex8
RW75UpGShPUubx/5IK8C8B40y3v4KCe5Iu38t47asftP2SUbyZvBWei9a8eH/4vrmULf/A25NvJp
4Gum9aZeJ2O3/arldGNiiiXPPIWFsHQrYYbxMmDGZfFsqTjM2ZNFsMpgEtpJL8yCTqavgScWGTla
cZLSfGcUMDeqZGU0h1UkbaZZq1DS0AyWPbva9gNxSWtejKFnaw60L6QVwIcrt6vreREcu5iBXuUq
Z2bjuyAXhnOX+fhmcQDOd5Cj5I+0GZDcDbXIVlodCpkxAE1G7DHRBbkIG+bKNtQewP1OqVAwOoKx
Os49G3/o/s7nr+jp71H9b3I+LRb4Ii6EVyy/V5+9KDkkO5TdPhwdPAtLMoVQxvYH2qHXaHgeOsZI
VT2y5m/bXPDeUnOJc6wFG6T8PVcVXKYfOnfdN3VjhmuaYKGJHG4D9LQZUMvAheeS+mgqKdcS/PSb
NZ3bSX+BtjcmihIsm22meLu7FRlf+Z4lP3ine7vI6UiIGqQwLN8jPEoHgBCH6SMAZegBTtmY8sEL
m3gA+yLDEekDcUlbIp4TNZ1QhwlLD84BwANk4Hu2i9QFs5WqAGhGCxB7w4oLfyLi6ArdhdYxt0eh
t08ulqusmn2uU9SpSPFuzqJYcA2eVi6ScZhYrNK91PoZhzEtr25xSfhoSFFPcKBsiG72Hb2iFo6R
/YJZgvN51wASdml9clGyIMHl2lOu9ZX27v1ODodDjzpDHlmz2GXZUamh8kE6K8MpTuxvcoqCaRVq
KqaWk5XiqhpmYCpl1mVE2g245Qh4gfMqLcJ8mW5hnG1L1umJATh7p0AF8qwUbSdvvGSre/s9JWzA
5Q2fiq+F2OELZK1SM1mfbvJO3OmFDwvzPpg6VlgfTChEcEJYZQw/Q/TppqhrWnR8heCGNGT2/Vp4
l3VkjjBaTg/kQbc/Ge177XsnBogDWapBNiuMmGmWlfQKGEgnvRWnk0uT4+rLSXoi1WMUoPQGmrWT
goSqDQ7E/4wAB7Ai2VfVr7Y4sHIKZQA9bDQOWcNdE4CRXjf8Dcd+6ZksBnRnI+Dqa9wqgXAAjc09
VO8UustznJDlV68NaLvqp+A0G0VJmJ+lbbemz7FC30GlVX+6iR1F59lEjpsMPp9TCZliZyilPNGU
bLOyyrVTA02TzBJsHQvupRXGX9NC4S1byjP/pfSJJiU5p1kZieuEaIz2cZUX6ZjDqG4xtpvIoM05
IkcwfX3xJRzLKyQR726qpaY5QA7nmA/tTXqAD4VgGcPuXE9LxUPXO/IAz5JJN4YWVfd/y9APPXcd
37jm3Ou9xCTYk0B5ynfx9Qzr+awSxoN2h0//BSmmGk2yXMYYdUC+6zIlks/kCIBKADOPMzNSKtrm
MvLBvMgorODXRATJg098qTJ9sXUbVUhjSFoqsaK9koTfyXMCM4+UMCwHoHmPEADTUitF461OpN90
3sJZygw57H6JeHsZu7aA3DQXk1202FVnRXamlW0bKnsioaXLLBQO2S+iCmEEX5B8gzI7ek0UN0GF
CYIchQAuRd2Qp/d8M1Vk2v3Wz/Rlw8PZ4WYNgfgQGL+G8x21xyuRAvHG4JwpaK2X3tHHlsd4npPq
Fh9nnafx2tz2f0h7xC6O5hjNSLAarYwjfb/8K3esux1zsyqoyeyOmmrnPWaPIchhxTngIeqz+lYp
tF02gN5Oq+SCRUz4TfCDFsdhnDiZ1SQOu3Y9MjGodvIVHMnNz47WuUXLPJGJMOBWl1AYVlyDt/Us
Y5+QhDa9GiEGeT7qwn4xeQHFVXSOIRQPONIyh5vNVDqJ1yuZeClkqM11MMQ4EA7kP0Yc4DAOo3i5
hqccfam2RbQKGLGKr0ZkMq9BYqM0iMMjtzNJa4GTMQ7kuDfp+bqATLNK8O8MJWwGC+lgEJ1zNm+Q
s5Xf61SocjAAEtNctjfIZc7oFaU0EFczCfahTR2tZVAYAUPoXxrifp7+nV7p9LbQJCZM1mdhdhXZ
DyROodtK4CU7X/nvfXO1GS5kIC7Ew4V5mcrGd8qXGMSCcfM6/RbaPqyaFBaCDHF/84qTi7LjX8bg
uU8/xnRR0q3U36HL923zj7NDh9dg1hfuhmqX92PbDD0zh3dw+mgzoWCh3q64n43h9ZXAQCGfBRls
6UbxQIxvmueAuvBrQTg5J7KpYBNAK4LlIjSkUSKEOvWJdm86ROp18Mui21w4uooFkNU+rMAFUnde
pWixtwwYS5sEiW5qCJ+LA9IUGeXG6pUACPAQABlZIMYOqkiNuiJIvvWxpKMYRe+YmDB8E0SwAXgQ
Xb8VljiJ5LxybVFC/e0DyteaxLvr/8WB3hzzW8BKKYTLTsSDYrsrXu2HRAQbkrqV+cYwQZmIYDLE
py/fxdc1KjSICFJa4xFHE21sIQJ4S6WRzYYkr4VDaIREqxeM8zBNNcw8coosfLslh+rJ8pG2ibpR
Ubhkl4wM4GgQALo8ma4UbwLYqC8c9yLPjYkDepIy6T+NHPMs4yLKecHKE2hQbl9vgmI80FRvLGiG
XvV5ongJcS4oY+buY6dshazAzmnnasrr1T8mxRU9UbC3NKvj1JNNZAx55dObQgko7YTx5h9rB5qf
KUQH8MfX0a6ymiaBEa69Bm8rDEcbLPETSUphTcOfMLF49OIzQAzG8QFEc9fnllqJDDKNzfDimk6a
InaH8H4u8ePzIfQhS6WVgsxRRvAD8ra3RKNsPj1wzQG24lRslhUwAi4ebDfdsIXbtnnbKSZPeTFr
Ijs89on9cZ9jhF5hlS4sswJdsQuXh/TWPck9h/Wqq5z03p/4jMZyheb/ArV9fK/wvb77Sbfs9RW9
7WnszOw5J3gV2tt9ORzstZZvHp9N3J+svLUOPXjEOGC+2npzt0E6CRErQzBqm2/HrX62LCVvThUX
hNXFOm9G/j+i/EIlluKikV+HKwOStjlTf4ZkcyVnmMUdGMq22gIX3GLfKbuD/HPRTm99vMX12w/x
KheLx6nYCennan3GnoGJbYKUvhj3GjEZtOunHAR7UUsU7ZjCqv01PrRHc0EixW1wMmIgsfkxg3ur
yYGTm2pvHg0nWZ1rk2exXCjdcuXOEYsc5+dPnlKVOognjQPSgmv9QRWb31OtS39eoIyxipBqIX8v
nL4lwZqNUS+GJjS6m9bqVN0NGDnuf8pcUCOx7yrn9MlTE66z/3kVsgcRZVD00Bk1UOqU4buDAQ1j
gMkWjuDt6q+f3nAvJdpzLArgFbuIVRQMJdl6acSEIwB2KRRdX0L2BCOzRdhaTiutVHsHyMYfrc4K
hoigLQlthOdeqjO8HogHknB3KK11dc6EoY7LjjJVl0slyz5/dyPTsPpegBl/fhFJu35jYgnFz7R5
Rv6EzywTloohQw6iiEPhaj/YEYRRMjlqs948P8MymtZspboHdVU9fTyVVg5d1a7mU6y0fwjZj1Uw
9826eFBnFTIymc1ML1umfJ5E0t08U5RF6fRIr8IbFNIVYEz2tVEhN+zArdqgSkqzoiZic6CPC/lI
WlRl5m5HXmElJq4mM2hvk18B1YduqE+wBuIZaaMFs9srMIREEXIhL8ZLFLiPiy35RKhmwqcjmgyn
xTB6QCFpRRyYO/WzYT/iWRVJHaF8hlUse2XFyWRMqJ7xrvm3sVSLSjn5HVpUq77UOw7X+t42EKfX
jUlWNJQLS+0BkMGp8JgOt4+JaikqH5fw9Mom7nvSNUwLCySHat4wZFk/aTQKRwGKvOIsf4Cgnawo
svKorzq+LEHu56/tH6Fe4NpVRtB2Ry4IWedW0OuaNUFWX8jiRJ+L5CXt3AbPYf/tikBsH/4Wt85z
PaZFJYo7fs0Eygo+5WlSY9Q9rajCMmhJ4jJuitlAYgdCA6Wvzg7TyQ8xM+I3Ly/YjelquuVNaM5c
7n6jALbIfXnfcCmSk+DvdVFym8dKno1W0ZXZpDoq9wGAvsZIpMVkPEHtvOQmzYjr+v4NHehEehmJ
2xQ6xCnVCq8jEKrrR7y78Shbc5JCSD2bxmu8mR7FUyA3t7tkrcGQNlbdLBZnilPoyRLpxF0+qf+g
XEsanuebPdd6V3fGLSVbeKSTFsWXQe2L6FTYu0SHAtc74MxufUT6rFV7omM5ewkNS4W17MofNW0g
5WUuAqBwGxMNAq+WJBMLBUUo8YmQoC3G3y3CyPKTk/GuMUYZLpr8JcIB38kA8c9z0jPDNmuF2GGD
KdnqZtLyWb8841REevSFChp8ldQYUik+EL61MZWOeif+AfhEjic2h0DdTCZn7Ybr/EJWSeDA4WNU
K5E0zpSr1oRWj6zNIz9s/rEo6ShL40dZEpgq3qKx1O8oGkkkfiy2AWRxXhgHTgFb+E50PE4VsXyB
huRSA64FDT9Dtzk9/wfrbyXjxoneyTeFL8179eEMF9mwsUUAAMKcUcu4XpDN2PFeiHedARhc6foj
3jIDNrUR+HSF56ya3DCM+vmd3sAf0pe7u05GmgwoOKXh16UZOZQ5sPiaWJX84HdmMWLglQl03MDy
FXtjsq4V78cOqd2e8ggNWlVIdZgh30fUt5Ead1gMIgzpaWrgvRGqkPDW/RrmL+lL3pmrRvTVwRDr
/GnX5bbYIBZXRccPxSgogVhXBM7u50JVDMMYDokYHcj4WIFDI2PuX1obZnq8qoFQ1XJlZeC7AkWK
9WZ3KQf/cmq3StNh/ubOchANG4SU+DtVsOQlMZoAnyBRfGxtTRN5AqSxWPuPyb9ZRKjWn90oLdDL
nX9TcoAhp2HABZaEbrae37G6KjNaHC5L5UCf3F5akXs0oycBarrEl6yoJcE/mXsWlnC0AVJK08AU
NV2YADa9cYzqGbjA/YJPIE7RAfdkcE0blIzbZ3t8Rn/G3ELhGiDac8f7APua8rj0yeEV5gFZshL2
YxCj1Qnrsspn3mRkEnyI7+73RL8uy/JR7bR07NRrkrrYIVBg4Vy+JiD5K04lMX8rJdo+a86HRFvq
LeTDbprYo/FsCi3l44LOGaPWluMWOiRuOgiB5lgZIz2l05/btmYnYqpri6xJteSPOmXUziPxe7Kw
MdGRSGgKt2gqxShQ82JzwxaD777rdaNBHFWUPAh+tnkFr5Llm7wBqcZ8Ecrhbd+j+V44VLcBI5Va
t4+wACIDk5wdpmuFTbUc8kdsL5cCJ1RTZ1Jsw29/g/30TKDKW61iZbzmHlpSqG0zGprVedn4/fFd
EJghWW3S97Pih7WvaLSKyFKmiFSpWCGPMVxQcTOjpoz6rCYKEKubpvKipBI9qGVys3XLnGnmlEah
NpwbcQ0fPmz7Msfz/U6ThmWeKjIqWPQC2z5ryUvrs8U0fS8POJzvg1HX/cyvZEW7e3I543ljhNWg
Ql3VaO0iaGHeMUOYTJR87P7fmIg8CJYNrRzAAhw/qoRBoIJw2L+wQb/YrpNhLioYncXODbV8jhzX
zTAbhe7mRXzCoKtj3/6mhpIMtemT8cB5F67Gv9VuXW8mVroiuwZH107uslgRaJdzVJ3VVABNcyI5
hnx3bkui46r3yoUgMRisF/7JoSuTQL785qHpoveOeOQq6VlTHXPbfPR8QDaLjIF0qY496d4Z0VkU
3AGLjDJWNsr3/XcuaRNpCOquoec/TJsq1+ggRNJbOTvLI39w+Xf2H8RtJy4t8GgetV7aAm8+MJUk
Nbg1qcYAh6CiCAbfBL9WCqjKH4U9/8J8IHHfAEXF+LdESS7hIZs5vvYfyd0NUGcXS1UuptkbcVKG
B2iLYlY+0dHm5RKbcQwKk2SfkvFpjxC9X6eJX9JpireKAayR2CvKC+YaGVr0zcHvpT1T4UIOWDYl
UHzNNtQw8caVCJ3R0bW/6eGiOZc1wtXzMSGqKYOyWwcY1tntBrWaXBK2RjE13jK+rH4XADGl9bB9
b+ENk3VeJdOzcFyi0B+sx5ZhFojOOchlPKznWST5sWmEjnKVpHe7URWCsoaAOVTcqvZEJpT8Cd/3
O3Z7Q0rNUnsBSlVF5m5IrrjwG6ogFHBUgDqarXg0MiXmSIwbDWcZV9ZaJEa0WuCkRF/lwE0Fpfg+
vJLikAk/AuIVZKAwKoS6b7teeWRkJQXEPgwvV3mJl3P458mg7SQKCIbUlNWXfldwRqHjkG1KbUdo
z8cPxAvulFvzONxSO9i+wv8+Id8Dwv49N5RcORkDbcuupv8JoqkRqLuXjUPqR5YwCh1LDoeX2PJR
IzTM6FnPFt/mmEZUBY1tma5YTzT7iVCx+SiWYTwScG407rZpWBIWUxV/D5deKcXbTogPAfILLWl6
+laADmDncGQHctXslUMQyOKX7GYQcZAbzUwh7lYTxwLBa0kvpG+Oq537JgHUP7sgwiPhIuQOzqk5
UD6XmpeZMevHSNwnBPsMqM+2z/7cL1ux4Awj49Kx9Q23cdd7Z1ksfSfV+L1M/D7BRXHTAFTE9Zog
i9vCmJl/fuI3tuoFQcxHV0N266SxVzdVwdq7GOXV+iN1mtBmurKl4gQKCWvOGVGDqzDbOCRTOhHr
OjuqyYA3R8iqVBInBx8pF0/Vrxz6CiCS1pS/E0IpJlYCBCKL/BO0P470Zl5h2kqArlbgx4pfIrkO
HQ3aOrsoeywDKze5gb5Byi8kasIgpdb759afl7cughQJgmascK65K5xpG0a3rPRVXN3XpvpoYvwv
xLmkPnlHqRvneh5C8th1jV6Qhfhg2E9iYo6hl06pSWDNo2aQXp0oFDvbZgjm2zug1Ba/ven5lU4o
uvSf9nOqnJE/U2SFC+0IEQD9mE3X5aItqwUIfSjSiqYPObUOCo2zx5dmEb5LcgH/e/W86DMR/rX/
PW+OzHYhys9nLnBdFI8IrkHVRrpA7gUKL9sd3ydt4HtqQZHdw6VqVV/BNw+Kpj7iYTIGeqyFQObR
jd1zDWm+VFm/Bw191a0DHQxAu0SJiawg/FjRKyh1T39ZFItbfDiONR+cDqCKJrvSdlTkbkuyeL0F
6IDRhC8HTcvYycNCQDXivmjp+1zb6yTj5K5YL8jJcKr5vnoQBj9Tku5zmrkdbVefmwSv4ocJdtg0
E3vB+8WDtb4PlDz713tg2QpidB3k1tVUynkoSPFDUt0dOU1KMxxpR3iQu5xhjX1rL8KJ/NWOeB9o
ASh2DewYiDmBm67uS75HBFWCWE3isLlawxlR60mezXaD7ut8WQXXAAF3GrhbZ5CNt3cBat+fTffo
pnQHFNawpGIPbXkCgKCHNGAkn7SdeefBH3bsGGNJf2lFuTpKm+ncd6tuizyK1aLX3zgUxU+Cwrus
Pp6fNYfp9oB7KqIZuR8NRCAhp/eZ8y0eMKpDoHiiVHa5gIFPZkuJ+5g5Wue0LWLy0+wGQJjloOZc
jU94yvI5GTokgX7a81kYFAKigKQGyEzshix+AuCoPUFkv2NYlmQgCefmWCALRRoJ3O1lQCgATWKu
F+l8SMK5AAQTrNZq8L3a+z3yXjKzj5sHBgPRMS2HgOwbL8SUcupxadRPeBuGwdRvuE+Ye5Nk6RqR
CSGUlyUynRgZj3Z6Hyup0/kjPK2yQpxhnIrVvL97zxq/Q7hg0NDCiBKMIQ1Kq6ocd/T+u46HRcHQ
ssIfk3fImwLpC/jSmWr7cGx2vAhO36GnXgk7DmFBf8JIULT9OyeBXEwhp1xYfpZExeEWI4ZU1JAX
PCP+qp1uEZNc3O8xo4lSCRP28R2xIkETscLHdmLSDBuz6soH2qeGtIZMjNFQ1T1a8KVCBmhqZIjp
3sXG7x8LK6ynsv+S6Ln3wzuta2+g/TIGq52I8AQXhMOnX29zXciBknXIOzQhhtgkLNxbvmR7crGK
skF10oSrprdXjFQzNoGh1imjrALHMzWuJOWy4HWx9rPiRMfr0wA4SuKbsANVtJYsYMi/HB7MS+Pm
ZcDgIi/uX/nlv/OPDiUNllAHv8ShtmP/CSPkibaguTCFerWuS9zkoMwZsAey12Bx1aRxIX+3RicV
SXuyvd83pA3sLV+V+3eUminZEiBWcPAtZ9i15FH3ADGbhkt9araae9soegkZQ61obSZZWYPW0xRs
b9T1J3erfRWr6fAZnKa7Yd4ydvHPVLCew/iN8A7M/2auC1Li5UI6Q82gvGIcf2c+4ISBSSKsJGtb
bcGoRt0WLHhs70P3HeKDX5jSBSX1TejJmpu2KMLigUsP3Ara5lSx4AsGhN+PsUwSKemYxM88EeC5
xkNnLbI5KsZ9Tq1NIyDJaAs1ds3ZjdAIUdPgXVdGyGB6K5Q4ZgRdCCkIJs/KigSRT9WRJEpEqpIT
y679TW5HeJ4rW7aDOmtYTB9rtU5CfYMgBCU7o5rnIo97Mxv9oBNgcsy9CDQgC3Ic+YPaDqszGo0i
lETyN8JgQ5b7vuA1gA1GP1HGLZ8IfPTpuK1JDENOCEKLJPSUiTlG/XunedlnGf78Vs3W5kVFVvo1
/8PLOG5wiZUZLs2Dhh8p3b08p9PxlMgSrpb0ZqLSQsRarbsaNotg37dcGD62nGDJ04mivFPPDaeT
yUcFXYmT2wt4coBooYNtlg69vFTnIpohi0CXdAvbVNAeuxPKWn+W2E+4GtWLWwxC31WF/10AerY4
v1tkH9JqO/cYW8H3anjomjfuoqwKIZQ0AgJFzABoq2loTmLXlZdpJhExyZKUIvL+lVrQciCdzK+s
Ua6i3Q9uSs6Abqt1sn2fHBFveC83pYUtFFJTIdszx3pBb+V0jGzRo4ShPiCi+WadAAOK1VZBw5pl
7LpX3oBB7WnpHnlCsfyPXJvAOt528FJNHVqgOs0qydlcTKr5YrFBYFwLjA6KAXkmDlS4tyLchJkC
lBdopuqC9NFE2N9xGqmempPcG0jtP6JY4OA306i2x1eCCdWgD6E/DxzAfHDqC+frfQ2gwTvSvKPR
eV0nyMk+kUhdF53ZySuYXnbbSynnhhPB0pgbfWeqsil5zjuYDvzhkr8PrWAEdhDRCx8G/6nNYQao
K5EF5q+Mr/BRginD/L4YxgeThq3lmvX/aZOMRdN6hYfaNrKgeDaMLEchKfzwVat6j4iRMMsE2guH
DKLjmvqT1HpaXpVKlrcFkIvNot8yCuGpIhAnFvIlIGDgP3BHIgqMqVI4pwm3JJ+cc5SiKUrmu1Sw
ecrkFckm9BQ7Kz7emlyiGktMJaLpqOK/7NYOPezZ5Olqy7f0rBUwuM760qCjmBwZS5FLJ99cw1RZ
BkV1PCqGkncpQZhX2NI8IKiFSjdQ0hKfZru7CCs/32oTIB+OElVi97/OUjQnIeaUZFQdzEJgHnDl
teWESkDbptX3wyMPz2KrI2vFi7/CPsELsR6rqbPXfUdDvc0x9Ql2rKbSX0+tSG7iF+JD0DBsy5mn
VFQhnCx0D7iBYEfSsZRA6mz5qtufJ6VgMCfyDemaFV/+rdSzjCMWA5RKMc2k3DpTikHta5VOARAi
w3aRPMVfvFNClps49SBWTwGTj7V785qAF+Kx8AV0NZi4eLveFtFQjv7dHpTwCqOGyeTlSI4bCdLn
6zKQgM1Kxz1aTX+NwDkCBs1TnKK1oTezc7iwZtg4zSvSggX7QL9Bmykp08y5qeh+1Zh6i+pKDMvl
zQ7V3u0Tq1T8iAYYDZoaGWbRANVvqcL5qM4f7ZZCX4M+vCafZt6JP2UcvlazXU6/Nq8HWWeEtpGN
gIKr/Lo+0aHA3AgrWUcOlBuP3NJFGNp94igc7HPotUcrEQKdpqxp8kkgISC+2qrYC5wwPxj3Yy8o
spUi50awRZVjLvmBjlviR+90r3OZKr8Dijwx3IRdVtqIqha7Y7no1om1oyEEofOQdQxs8kVviGGJ
UcckKnOKZqpPCvMGzOxHeRhSNHIMRJEznAmETe991/jWGp0IphJtp/QCngzjCjtrhlGaF7cUoOaI
IkmDE9CAm4e9+crNTFLT9PuCQM2AcQfw/3zi2Cqu4yugjcHKiGsnktZcGmOC0vq2IPZR8MgIex6u
0/CMx28IbLzunriqcuJ7tNdO346BqklWhfWh5YVwzceOaRTDlyfcSvFLBCCDmbCfVDw52iuw/NXk
TkpTudaeas7/LukRkrx8o9eNYsRvaBl9S2CaMPoSYIp00OIgVnFdabLwqlE5vo7E2QOIZhvQxibf
oMxLEEC371fwiaSA3YmtLCKf5QbtRQhNH4fvyZN0hpyjZsvVv2KtVN+mXuVZY01m9DC9mvcbd4xy
cBOicI5YP3IFCzUZH6N0vvymDzrZDVemLcP8T8PzY31HNML8lSx8hpIJYM9YKzu7zAufrdlUoUAX
vNqWHjluQzgNZfl5RuQPRXQn3JZFDDLSnys7k8HL4O6X+AK9TN/UMdVFJHlrQ+i34KY/hzaJhoCn
GIdAOQoHyiUk2z89wmVGsdX4p9UXOpBCJs5l7RHKU8Cc+ShSK7INOVYfn/40U3bHk8e4ONwflLMo
4eAJPyrEnOI/odKM02y7aja+8tPLDYkWyXk/x4eEpfOOD5UfBV67Z4IyLt2AziwKdVSrrymjNy+0
ljOZOub/kqXXnBEMnJVhkUuXRSfmZqAbDf9tET2qaX5RZwIwrHmzNPO09V3LrfiMnLXdbofDISsT
9mnC5XV5s26LkSLBwnGCc7Y/Y8JFuptjUdZKNkJNat9/Lrth/0h05qiR7Q3f8f+0O7NA0a3HWeOQ
2+0WqFGdu0n31yGXxBQ+vTsZGrMxHIIyHG3m5kqET7mwh9CVRNxDc8L4hC/6s90wN37I/WSCShlh
X99aBlLj6bHBJFwDQR2JL85N097n1b8YHEAHG3zYaIli9WVTEW9wG67b0YDDxA8nQCZH3rgqYOzA
fHaItiVhmNUP2Dvk2zdYcdrCAQgBDBUfJ2hAOfWbdQwtw0PZVx4kS4vKOnC49bqcqxqtSfk6JB7k
PMAlfTmS5HksHXj0CMzYhPeIyP0LmXtNb2i6TKGRsN0vC9KpE84P6NHPGCqwcCFA/q2r9J8ZCzRv
4rokZ7MzE+fo0ZP+3QznzBOaPNYIf+TQc+N+9wLycaL6SDT/4Vsjz/jA3Qs1woUwEX4YHL8UFciA
627IYv8e+YdfAXfOpp0Hr7RXaOsNLXYUcDFP04Ko0me/4y2c4/J+/Arc6Cbi5AhdAff9qBgW8SNj
OIV1dG5q0MssjUdHkrjt4QLifYdvSvsVoaqixhuSqn+Z1d9ZDKFlGiDwZeB19bz4HOAIXWDW5MFn
zeMsUiY9aB8S427gD7eOOtMrvMCCeQXjtjIAy2KkcH15NNth1/ewjFZnoYvSgJgKKScvPm02N92u
4YHkSsIL5Cq4C0KCMsaUqs5ZY5EfX5wr4falNP3TvSSbeoa8CBogjSI1Ore0LsQny+CYcMppdb6q
9ty4Zizff2REp7POyOCH2UL+r5lSHHApq+5604pvKPZSJHU5uAHkjc/lPgIafTtT3uNv8sJrpLrh
rWjx5NVhLDGYIKGSLRGriUucWaRihdNVq81DI+I4VjP3aEliWCU5ZNzqhVZIdGYsTHa6/mIc/Wek
GXJfH8sykahQ++MStOTV361voOWJAiDcYPVgWMQkvC6uo1rregyzRbTKVg2orWmSpD2xBKAVehdQ
RBfzJnTjIvZF9PI5QOxROaTIh7WaIZv2XTBVZN1ErnNjHb/73WjR9rDO2Or5ImuBgIp4TmO/W6dK
g8izS0gpWXKxAZvf5ZCVRqdD6lX0lBEfE9xu++OOPKSitydAmlutrbqvcVZr9i4OI/ZW4vWVRM+P
IIRCZqNT2Vqqtz6t6hk6JH/cZzgqIKdBPjvyWECa5XdCP5XjCca/X6wahiDjJAebtiZ+IGdzmd6F
5cGIJd0+lGpKeSIM/Damrc1aqxZN4SnVPMxP/XN+bSdSHg9h2DtiR2MFH4BB93ljfTgxi71c8P66
tktTzV7bN1eg5nq0cmpTocNXM6z4AT5XrQrXbdFiZ8qNoixY2/3ZdnClyN6KU/USRIMjumeqXYvl
3o3F7Hwd8zli1wN9TI64yvfifWV4iDFifYZdhVm09tjdXST338156ueekp1Y36NIGaFSEARxpi3U
y9dJrJCF+35n378Ya0vk/eGo5k4rO/ucq6UgavBVruxS1jfncEydCFdJOxF7XYipSUL3YGwbu7I2
QBvHpBsX61QJRa7wR/Zirv/iUhGyP88xxNFDt288gLvyI52oy4UPq8nZOtZ2wGvb5HRlGL3A+xYd
h48K70L8JLrzCERhPRmv6rBjsGfiWctqZdsYMx8n7wC15JXq1xMW+VEQ7ra7E52imMa8CxHYgt/6
Juvs5N1dqrFUwwtZtmCrlwIR35KZmuMfAaT54rTg3wGv4Q16lJkXjKPXsiSoRiI+wHMgg6vkarGX
N+KcYPl/59tNrB7FRUtLrgRnR1q4D8Yb6qjW5wpLyMFY66j0bMMrcX/UZ1eEn7fEvkMhF6r48BgN
aNGSncdv6DJO0kvVaL0eXkyR53BCEGxp4ZGeQLypt2iWnn1nL3NCL2X4rHphGeV0WKeIWET7qPbn
hkdCBntE5bTZNARgGGMmycKYB0BxclqgyrNR1tph9gMC/o1nCtXOIcwKmiQsX3twR0GHRjS4dZLt
xyOoVfh2XJtXtWOEt/MmrtHjcSKT5jEFEtGQF9JEDV2Ytjz1NTErHrNotTpRoXor56g3k3NSYWqv
RouNhAKyLfr8g8nwYo8W/Z0O6h1CEx3Hx4JcOhoANtayGZLvdYgfP8219cMec0o7j/7DXP+FC8Iz
/zo++M5jT2K7WoSRL/xcDJ7kKFkORKTPMzWfrEqW0EyxabEb29CkFchuByII9011JSfHDOkwot4I
t4x82/GwaxwxZeA660iM8bEXFHLqiVpqJbuhwnZdUMpyWdSv8aXZGsrYCbwKoVmUzLWB22leWjJu
GkJ/2r/Edk6x3rXmbKsiGgu43oAv40kEdwKwHjD8fHTNqSjfLIMwwuYDMbQEqpdHjZgMTuYHK266
kmIYrzJe6gMryUZ1+urWDu13PZDgCLAzbsWq6dNss5ZbGHLnKzc0jYGFhQFwp1VKLUEsJthUCvjq
jX5A+9FCLAWD73qgqAxtQ1puYYogN47TmkS3NluGO7UordnUuGnD3nuOyBR4x8FPoZLIlzlrVLrR
H40QIXK+4DgwQ74jnIME1rr2TKoDp85M2iFcWZGDzSQA7lo13+5NkNN3nqhkZ/XvTd50DP0JuYa1
L+Stv2tYrfwppJq53f1+6+ms0d3pdiqHshllBv3adB8FXNWIwq0yNG+wdkFmSsLf0Ag34RMSUljL
WMq+Jtz6KZjxxHYxjiU9sm0MR9DYR8pGumgjloOPUz95ULRnzzgM+Iu9xsgTSY5n5m48VccjZl72
eOpjMLD4E35E+OoFhAuChkgSx4BnnpTEWLDudrr6LOm16KsqMXl2bpZFW6lkI4SPq34abGQrux/q
Ywfrag0f1nX8K+amxHeRoVt7wFo9XN9yWdXlBz9eMpvSjby4Ody9pX31RUrFatkJC017CkvgNy47
kesbqVM2aYWMFqsGDhYofBNfZBM7t3cW4CP69/TyWyohK7FWNF90YF/JOo5EPyrYs4+Z9Gc1mvrN
4dg88ydOCYeb1L+6VhO8SlNwvQK4RejfVQyXl2rBk0kyZ1CN4QDwY+3J4xmiC6H3jURddeJadgdA
Rcu4Ug9m1po7pXAUTpjYpW0expYZEX5kG9iQMCHLAJj/Ck52NbZsrU81WuveUFAzUs/3AZybEB3g
CmETWZaX+0vqZy8KzZtjevNnIiS1BYKQmlJTfC0GzM4X+m5KDApLBHlAwnyaJ0MFY9DVsS9/YXRa
u/pW/XOzMn2TpJ2NW3dY+r30105gD8VS1A2UzwP62knU1yNVX4aYqJSErzjrvQlBJOT0nb+osZRK
b+9JgyXwH8/51nXIw5CRb/itB83y5L3DCw1xZCzurD7uVBf8DrMaettgo5Z4UOK4D7D/RfIb04cU
GSR5uURMDTf0KC5TSyWFHW8BfO7v26810cQb7T97dzcH7so2vt+JGdXA7X7FtH3H3YVK2zUORZ3x
5qPguJcocY8t4U8QW44NWlvsKohNRlxggYd2tMUW8t5pGTjPWSwSpnEpNHYh/2RWQbAWClWtrO0T
fUzS2E9oKBYC1Z6SCHslKRLyU6PAp+XlVNVT5QgeHLeHd64Mq+f2cpEtfVjl8tpXn3KxY1gYxmUH
04BuTDKd0lhxe6ZbRNFceMIzli95hjldIHzH/LOlD93Eyd3bKkuqBzbebMEirWdTAOb5fI+PMMCM
bywm7ONTglULpKipkkVOTlewwUq5IL1c5GWuTjovFQuel54LY1sOnQb98YKX/00Vze2ANzPjcg+d
4EJyYEc3TZRDFWEtT+OKemFCSo/+GGO/PVIQ/8nWqoG9xTilR4CbDNixmM3xJkUpeValwX/cRFQE
20PPT5kjoTfgPRLPlpRkUWAoyOJBX2jm23Z1ckd4n03bcZAhh9Yx7RpeidWpoxe5C6YR2R6yUAgP
aFgBm/9CaOxc62d4sT45imOMf4fuc2CpQGgrRyVmT/O4wo7n+pNdUC0vAXng9EJ5Ci3ugbY4rJnT
xJJHPxOhHAiwgzFLThU1SnKAvwPWZSGtraQo0Gx03xNkLXgFU4231X0QpjNsWfZqojt2RqzPXcq7
c/+9djQV9qYOnc9qKbmHs+5COgJSJ5TGXIK8pM/q6Ssi5O16QePqWwrgOs0tTZc2w0xqYRa7V3bx
prX879vCoV2SFKzic2fWb4SpjxOlPhbnXpyu6iF16PqoYqGm6HQ7sH7dPeoB7TUvfPZaqhC/qxEl
c7JAT2Q+ig602pdVYPY/X61jXtO1BV1OXODREbqRxOUM9GZ3TKsa3KqhMq6FZHIFVOA0PzRq5nY5
Sqj0bnNjmkFufRZ9KOmfYdvUV5qLIIg0FZnFfw/60F7wXJe1lHDir+Vw/FaQKYJ/alR9ZpYvF5vL
6Xd59F20GswIdUYrJKF3+c8yeKme7lALcWqsi3V0ZuDTjoDkBPztzVXgHDKvONZ/+yJDmRFHz8dz
yb+YVJxywaLJehuf7IMG3E4RkcRgSObmgZuPA4XmLrbPBU+rMmEDsv2Zu9c42OSu4BeewtG82jx8
mEP6bgKROlWhFrLWWm+As2ObgelIpN0j8FQoZdlzABc4M5kUmE1B2JJQr/5tVbOMUUAdrbqZPmnv
NlAidd+WxPxu9dXr/+KUd38ukEPWLbdLkmYi2gAhffpVjxbFyFngR0ast47GQ0LcvXY/1HRpF1Ts
Jfck/YgMX7DylV7V4fJU09GIeVr2z88w+KtcaSQpW+lnJAraLArpY9UOqPCDXJNDMMiuzCcl0/x7
+H/VC1ApY6yrB5qshjOFW45KnURd5BnrZwXp286kcWl4KpPsb0VDfex692n+6+OE5Dbm9DsyN3Oj
nkFxBv69wMa0H4bQlNGabtm8zOIekqRSNfNlJVQu88ubzTdnQNgyQTdtGo3FXpp00x90kAdggPzb
jCiFJiEJ8sWtM0RrZIWKpSU5rars3/0aG3PvD2xeQQOjyDWKeOjp8YANDiL5WOM58SnIqGINlOwt
DM6C1qujnS3xaoG73mIMvHrLGXzOjxpfKNC2axrp37TgGqgIwpEuRM2WqkaQNiaiE3N1hOMOV5wC
Kus/jcm0o47yFHGfsxCvosnINZwCN0B2Y4ChFYID5/0fA8JrkjBQds2AHOnKm+ACs69+a12sgZyT
IvBLVP8bPB77sxD2nuQLR9QPMj9Nb2nyzONG5zG8iy70xO+YjVOjHA382T0hB/VA+8I8XQ/u7f2W
qc9iu3fHlH0d0H9w1TosKo6B5TeyENLR9HaXzkstosaTZ037fM1HvKGtpcqohGRmtqjAwgQttHpT
JTx9GV6jCh8asizU+dAQogMvKz71K3Jh//aon2w+qTJ+/3YwOCmICcV1AND4Nqrwk7i2l9VtKDSh
pwnzOgwg7/nQT9dzthzx+lDaxU24gGpy/tlCyxQL0SzyOLL4yi+mYexS0S7EiT3bUesv0HjZD65F
DkErOi/0KlMNCx5hvLwjFbaPBLvxw+yif8Fc99rWyDR5HSNVDXN7GiIfQGl8xlP2JjXmlR+qcJql
vMEyhda1h++qS3luHMLlAFszY332Pa0ajZnUbnWopIuO0j+zSjFsogJ4IrHPckQ7SwN84/YDO5JO
jykgSROF5gkdtpFw/of4qJ3wI7Oaj3QodgLuAMIFbsibjctAZrcuM/9vkLSiE8cTk8xKzUvXoaBz
MZUIvbGD68C0oGjzoURf3Hi/srZQpS54jW5aHtrV7HZ1j0PWLW1fcTfMUZwY6Tmuifx0BnezSZoL
KCWAxdOopHlXNQ/bfSDaIsFYtNYhHjL5oPsUogdQ3LGOUmSfYUTmu4vv52WjyYUJFY/wIpTNK+sn
bqBQvpEiGwALRTrxXb9QqWkHzotiaPfbL3RDmLA06SrTWpb8Oxv5vTXhFHk4fJVMGiFsJorRwe17
JGGvti9YkGdPfugzrXbvysWt+hyjI7VsDS1b0z6MRCUktmrPnSdS4CQilyG8+Mrdcp+5wY2qN4Qx
eq8jXkHsMdpL4rDqHL5vpSRr6zWi2FEVBhDeg2vcc3iTQMPZQJJqUo1E+H8JxycI32xXDa5jyhCN
Q3zFvViRtMcBKrxwDetEhIW276U3I3EIDJQkGAGYT0TcRaX6efPEUn1slyrE7u8MpK3TfDlQI7/O
PN4/C9q34URKIeSN0tLoxfV+U1L3gqweWmksczsaxoKmIyY+7wdBP7CCH8dkf9g752rbRA9gYAKJ
DUUE2pP/Qs8pQm66i1z7qXx4unFelbgR725RFqOiqEusScrfBisHsE/dmVX/CvvQ6rGaG33LtyQd
+28OJX4BfDx7ygah/w9/CVYnjoihcs8U8x3Xa+Y2WmrjxvcgCJzjshMLkW4OoEZk1xiuggpUgMBc
ZvPqMn0B70KHlleB2uL3Avk7nUVRtM8AhqLHOyyzc4lx7Szmlx/Mhq5OY0GVlIw5/aLc6SzmhCBK
oR2QqEvW/NwDaIHh6Dn+EmbxbsH57kYtYgWvD+nXbx9IeykyMWeD7kjuBg0GH/EG80Jf23AkCYNm
iZUclXJMIcmpA6ExdxOR7w9omMv5KZl9sXPjW48KK06GKfzLoqdaWIup/QwQ32RGOfTOr82lzG1B
eLEpu/NdqnBQfrmhcgIwTzf1277JQVFEDBO/3XQpmAWIk6IWyekhqJLpF8rSlNQ3PaA1GQNMWoyO
hU1gLQh6KEzPJqMmd/vu5xHGq2hpc2uMZbO+VqStom+sTBtOL4cNpMpXo+aeunmMZg8E8FcEbEMH
MLVofziBuX0YgBfEmtHjTCclb2XvM8qeLHLjs0mnSttGLzLBnGfu+kGx55/T4d79I2sZCRsz6zCE
j9UViiVKhHwts1aICeo5vs8NyLjZPeSkjJs74ejI0qSObeuLjDX4WOJspkf/Y0Y3/qBad9VfOw1b
lBLTCmIg8iBAWMCkT6FszZ3KYooDRjyfLa9KaUwoqsbCJv0tp0P/uSJh9/FTQInjeFcpRxl1MDEY
pcXCK4QmZIHhGvjlUwCou3e3EdrIufPN3R06DUW7/bixeFGxA93P20lmC3hUyEJWhUFFXTUOuIhm
3f3Q1qSJAsgy5aCa21lgUoB3an7t/TePW5jR8vWx+rJ/hXzFWoVkUEiz4rbpUmS/uGBImbAqwud8
R0E0UaAUO1RWKNazrZpE3tw+iULNrH9GeX+k/02h1DQBZosKC8kUIm+FBSr2UJ17Z63jW7qY0rWI
sTEhum/i4j/NKUtLlUXpGVbLGwNPKwYKCOEgGtIhg2+McUWA8Tcy33dN8obL+aIiLg5T5S+/I0sX
oHoSvX48Hwv9UjiDbXUc8/eFg0pvp/pgX3hT6JK4bXpI4PLmbBdBu64Tk99wHHRwuFit1gA17ITN
Yp67eQc5veYiUn7CNekuV3tXPrHBgpYVHF9jQSusM6XHx2IraV8yUEIgZVe/53jmyHFLZPyiiA94
Ir3/f7n0OTHagYgqZsjWk05mck7bMC3FQeLkmsDVBmJv3kpSwzQz4gpXJvE420DhQYkPOX1TCEZY
q/CZgldw4vJkSzfU5JIXaksD95Dj1ddOvwmBvTqdNQ/8kZvM1vwBs03e73aTOOn88JlTNi8hxsG+
kxu8wyBiZD1cfdM0zosNH0Gz/f+2YHjwiJ69g/C0m02vhcMyDkM81IiDa2GyHvt8l6gL38P7huKv
0Qme5LkMMO3Q4ZXp20Ke1OZS1VECq2b880GfZ/SgfAEwfr34PpvclvQhAJgSvCB4TAFekV2AOpru
W10T48IBRJcGE4+Of9qBibRwEazZOKCMn+nq2czOdDVpwcDTjZukN/uQ18BoGeSRAsgNa4IIKLiz
V9TP3rtBk3sGao8GSW9Pj/a2VoYDAlYawWXUZKV5kQ5l2ZSvs+vJwoo+E3S8Mp7fm6AOKuCgyJ6i
ebuz1axmyCq+J3pKmsYaxToMatINkG4vskK15VywEm+1YEuVF3HCTtNho06F7dM+cN6t13/CSvXS
65+iuAG8Wmo6pnYoDGRGLHYxeJo8YjFweAx/p3i5fLYTrpc4EMnE/0xpKHgNzxua6K0tE3fWgdjR
a0Jp+pwD8F2N32WUqZfOQd14GGTbxm43QRclW/002Xl/odsvGYHm5G1qQdaJmMqiWeKu2xjR0USV
DoQ8tWeYZ5I52ZFkrQtl6Gg+L98FMmzsZ/xUDDEGFZO1W+Ze55vIbBvzrOit3gWN0Ps3VMMiBuu2
s30VHuSmOIxMqiS7nF1n7tdjosBuU8/r1QxCDHwbgIhQGP/0wbX/nAXAH2b+edzgon0uHwgNFEdm
nbK1+o654elWqyjr+LX7o17wXSMCPqAX1BJTgEub7R9drLbjdx0rV0zrzMdEljT8+qRyZpp2Azq1
p1WmyZelRxgkT7rh+yrkUKe3x+sYsqkDJS8RofRbagfENmP4GSBQ0HVL1zjrS1ibI2AGMYGe3iN9
JEYgqAXtt6Xo99Pnhs9JTiiVscMyETn9hmXYHYczt/auukyw1YKnIMzz7xGt+Ce1fqBmRfnxE3Kp
JeXkct4FIU+lKAFTpb1fiAxnsGOM+bX2L4VhJDsN9PkENUpCAqU/wAaWfKUzq/A9Q0FF7q8/Cu6o
OuYSgFQpBhWqeNlCuGHZ3q+s9KN0uOog1omBkpOG9VCM/ZKSNt5CDvRGbL2/zWmZj7E1pekXOdY1
tdqNqbJSv60bpy/bD687iXM4kvzSeYNEpQ44q0bqI2DwRb9MPeOGwDDg3d5/wBZESsnDQ9Y+hmsi
Cqdk6Tc66UIzGcTiP9fiy155iZR8qQkmlWCBogNmsJKFn61MG8sjXu7Neb9XaHoX6J9ze1Q1Tt4u
gauTrcmIg/50TlJ9oGsF8MgxskQt6iAEDxcBl3ouPwMfJkukmURIT2yWuACkv8fkqLPNqbGd7QMf
1AaRgsydJu5B/xDGatk+jnFu5dE5Wg6AUIIwlsRXCFBRCQH4Dj0OG8N/pB3A/moFVx9S5NGfo87r
IwRo4LlH8AWp2Fg6lBbpo3Pyh5Bv1KktvD6D2GriksNFAtFb6t+M27j8dHdVK+lVQGNjDo6YPibu
K/KCtE5p3vCdFClk9gspIMxkwZc1TTLlT9DVOiAhupj1wYOZx/XcGNVvffa/l5oFb8JN+qUxLT0H
xC0zyXc97krJLfemZsIWXgCUOFgpFiXQCKezyIOCOytVhmeMHW04rOaTNlR4ZycjZu8bCGjk/0Yd
zX7hJUx7AlOtZwHZvc42UEIwQ/7ydTA9td7SSS0Lw6cHp/1rTseHRXx33XmF8rFVLlXMignQE6MU
p6rKJKAVFo1DyN5lF1MN0eIGXfRmHdE0UQFJb9jAbjc8VOoc4CHCYQk0FPh8N0BuWdDNjYzKaM0g
Rs2vWHLANd8lvQKWiPdrgiAQIA6YmIXZjMg+tDiAYEPvlQT0Ruut/t7PElP+0YaNN0x9tsfi92DH
bhOSd7uPX9RZDfnZGkAL32zJDMmeLURDoWPNy3TXx/fI09p1LDociWqETXsctAdZ8e/tCowX3Asi
W6X+3a9yqtQnfkBHHRc8vJd3gUk/+qmRVdGY3eWt4HRJJgqCzlxL4u3Ewun4rcGoAmZTEWwdZxy1
MnD/V/wHo3PkKXzO0dkrqsOiogS8kCq7aXOO2zJS7N8bhOGrQ4T9j4kMuwGWQu2onrXn4QXgJEb0
bFBfuX8QgwUZRWlMkPe5YG56o8qy3+79id7mBaTr5CwEp+weuwNXfZ7Ur/Zut/lLCk7xG9SEBisl
V4iLdgT9OWplGgL1UdNshole6NOjRNFS6MoPNyruRLqVNNS4ooJTcrDLyjfrlXLYvH0fFnMV70cA
oCA3TpFrSaQy/YGaEz2Det+Y51qdYHuxCK2hN+59SDk+Heu+260AQBxaI1qJ7zGG8Z2bSYw6rhxN
fpZvFn3OybKQoKCiDy38K3SHeSv2Y0YM9nkbuuxXzePiG3xzdotf/U3XF0Isgei3d+EPXhGEzhyc
+g/dFeuezAWzJJIKvmSddWgsgfjaUHyf3t7g3LnDhfeJlS7BXqkxaMh54U29GegwLUEnmMp6JOzX
WtjRanLOhgx4GsZ4jR5wO9IWFN5MvoNf8pxpTyD2rr6AAjLZp3HI+BPgKTMTbEN8AqU8z7KngtWz
+EGEb0JDaN2lng61d66RiwZ3w1gJtzr2keeourlRQKROoXtkIqjBXcpji4+5mEU/WqezUHNd3GCE
7H158t/FmMJWv6mBdZVbB0HKR4QduDnVFPalyB4ErtIkUP5QeNa7jUaNhVi5Et+pU5ekIKfaTA/q
OCKsR5FYppC1cUXK6eqi0UGKuyOT690LGWdJ5ZcjqD5N6iENA2W3Kkf1jFhnaglrxVq5hrFfUYZv
Tqgav9K/mhmJnjamu3Q3mWIwlmUeTCTPCbXdlcjd784W3CRkjPVpCHWZ52oZC/OF+LF/Zf1BN0tF
a8zm5ZNM4uocV6RHyVRFHRzaxYN9DDxTc+cEQrzcWu5XTdQVZlP2G9awu2pUl93CSSplkZnrrUFS
n26yfqz4l/jldi+e/YsWRlICoMMaKh20vwkwxRbCev8ezXexTLQK9GfhJbgipvAl0ANy7aWFt5FJ
2fhjNVKDhWyFch9aHQURJJf7QeReKttCXvRDaHyTSw4u2g3tFwHtQ3BRh/FgWdrpP9nMVAcU9dI4
nbpHC5CksBEaJ5zPQxC5IanQ/5H2F3aF6xrihUsqgkOiGU7koSH4Jned9Vob1s4WoRS1caGSxi6j
Q+rJdfcyMfkZgoZ7X9pU2ehLVRljhosqOh6KoZyvsQLwvSWGqTaC4Yo03mXy+sk4JCLlEGle2plM
4WiSW2A02JWcoBZtpF8TsDbM7p8JSjfrRhwY8h6cJp0S0JS3T+RxmYu5KO6NWbh2kUTLY0Ou4qtl
C3YriVa/MFLiSiRDpnnzo60I1VM7yTL2sQCbSyk9bQBPALX5688X318Hn9R5i9RsGk0QsBqSQQMa
q4opMqVFt07h8EDA0+sf0W6FFXiDiz4eTkdAI4uHbIh5RZxtfubirT4euO7rJtRva6aGfZSWanMB
fSglIuQS8yclDM9Sffj0PQdvHFPRdMa/DwPaTv4JvrqDIubMMqid2AKEc5lD3awOMjsFLoFJdcXY
nO/VwolYm8QQjukyRKg+R2n7Dz//5mmekGnWeF5HpsgPTFJNlxrPumwZ7r8vzVph96xVXFr601A3
mvRdrTf0yP4Tdg903mdRvpeP03MWWL2nODqPRfdEqBjm/K7aUmiUfGuATy+5jaYRAaZfxZDevkqC
Uj8xCZesG874+6nxfE2xfRdFmVCDvzFbj33xL6x/nBBzrkSwr/vrcPxeKC+JR5JgvrVHtEZbR0QR
thK/tXltuhG5bG6CdUOVQcl6XjfKU+J+enZiLCpnR0tbeBhsV0z+KJPgs2WaDaOw/cAt3paX1vYH
Dn0nvc8dwSAH4W7M2pUWWz8txHjtDosawQsXYk2O6kblusuAO+n6Apcc+DUmXyOMTZIIRWzsf8U3
VRtBBMgTvd7v6FLLHWeCmf18Vzsr9tJabioxYYU2ecSqhcTWDxsmp2oAtiFViLorJQBKVBOokr+N
4zO2BpssGIWShahlorUnA+n6hHpHIvXCBbBJR3lj3XgnOWeDl4rEePKiC+9/lzZmhFmD6G1Al4T/
DkEdqzi9bkJdIsVe0wK3eOjFqJFr+nVIG0QRsIzzAaTmmyyhjcb22cvlnjRGa1gBEC5WxoRHxbpy
LeCcwgBRXS6O1VI7JeMbfU+t321cluk+rjbngiPnxY9kPVbAEkL+70B2ITQvPGK4nk857oUnwrZ7
3CfVWEINKsLSaHxxpKeK/zLmhlE/spsVq1Hz41yjyvQL5iHfsX7CiXsp7c6v/pl+zTQe90IGGPOe
l7QM/jlIJ74rHKrC26+246eeRjbusR0V9BXWT4mjrht7klrVpRioUdGe2ApcyFvNY6esA1QSfR1H
pdnJdD0toJun8i02w+JVDkAXByhk7MunFJ43k/1f3n2crygDBgdEwclNcFA6zu/+0557DM8873IW
lKdV3vRLqK8OIG7NE5+CA1br3g19UDVTin5oy0CHl/BJpjXQFs54vrO/5uonsefj30nvnyHeJ0LJ
diCyHykXGe/gfxBiJm25tIr5f3chk0woYah9gtiEA2vU4pwtRpuVl68HXrSsvqKHXZeHQmO8sTrj
W7YzMLplPUJEu7JRLQ92nA0IehmF+9/TnSehseG3HUxVQvmBrZUOm2j1bMcEEUzu+rnqUdL7vHGQ
QqkUXg80ksSGatbw6Ra7LTGOsRgTzZeKj073GqvUV1Bjt0ZnwPF5W4+KJBh1D3wnnZ9hlqlBRfh8
y/yp6OWiHkuuNCjZeghQU/f31TszBZDfhrqjjpro+8I4/iIpBsd2W5sZoLCvuUt5Kpvh54D+7sbb
XQnfE87DFPxMCPSMvvHClSoyIpQEHleMWTMpKPjQ9bPW6G5N+jMRfzUuCW8er9b1NPxho0orZHWl
4mggNKwm9+XDeHxsYypWwZWK8jLXDYOtMBcLilaxNj6f66grezVWj4R8Zrwg7JGgRjLwBnqVOorO
sYG1EEoyAZz2ppRGf5sMEaR5DzSr65r1G0ggYKZB7GcQmh4JwcQAaDgOSENS09WYH6zRkBsRfFmJ
wKvTqK9j62mQIsnUf/zlKw0IXAhMUYyLShkZQzFb7cHdCMzUvpVDlt3PbRfY91HwfiFCsdsb0S/9
W8uAcrOSIJbAwYZWAXcFHJ74nkuywCnf9iPUG0jjKt+c3z9SiQOOP2J3AeiRW8HHh3TftwF6QCSK
uhEAJWEVyu8/GLf8evgEyMWMojm8usKwhH+xt2d9y+ffcOt11O4et87gswScDy4b6bD8hzWUUF4w
PyfuOcQYwwzNv7eJts5C3xJqd3dlGtNuIEYqL5S91KDhdf+QWi45h9oQorfOl/2X5e8w6x9ysmLP
lus7f6naFTcUAJ37H9pNdELGZSsmIEAwAEqLmrtONRvxkn5/p6PVlBYTjF+Nu0N9V8LLtq1FP3Zn
hFf2hThxG8Mdj6/lb7RSWkMv8DGcun4uZ9mfmrtzhxJTBPtoLLWFET1r4NTg0eRfHHcsIBEUM7Sy
claWHlwWcpxkVoy4a8/5k5vxnqWj4GbGclcqN8JnCxJ3P2Y8e6CSqGOo274/gYxyVSb9yG2IMet9
nordsaLtP0ZA+NCJTxkGum32yG2M081nj4hj5VL52hzUFImQc4lrWGt1ELrwNMr3Up35bxlqdtW2
Y2ZGj8xIPHZwMyuNUrAyyHsYqlJf3T1dMPvGWG2Ms3N8JY9EHMgcckejEdRcL1aWkZENb+cQ4OGR
j27WEElePJyGsEuB5Kqwgyg60bVOmhrjHlMV2OGp1U8ZaojkOJUkGsKGABvC9mxTXysSUqSIbd8l
iGUe3khknQFdjmIYh9u6WecnG6O00dj4dgyy+hyHhlllbR+f0RgHPlht+2YM4zVz4iH+BsslQ3pC
uv7HudJv5OnGe0lptQZllbmk5FBRRF4wpxoBXxnCmmnvr6Ab/6QkzcT0n80zQfxie389dOCKS7s0
fIrFk82/v1+w2VE93wU/0clm+LVA3RTYu2cwnbtihROpl4S7V+DQqo6F7E4zrWXsW0UkGLRE9vFw
5gPhkWCz2PY82/e/86kd0TQ23ryPbivNeyrOmH7i/phWgJ+0S6HXtDa7qSOmqbQK4qpdqP2Gpv65
dG/lGFxJoTgxNEhl2tS9KpEb8WtdO94SYqYIj0Ra3SVIdAo6Do7WKN+MHwi84oqPC+8TCA8naE1x
8vLPumGoEhDyFyF6eYgFQa/bJ4s5J0+SCz2yyYx2o7Y0wSp+2Ypq3LcNf9D81m53i0PLn+NAgN99
//TpEmldfLA2d4MybeRP+ss7fbcKSh1hBtidjsTxopUWKWoqmXguNskYKgbKzENwVIsOa/Wtlk9r
ktpBluiKsKnf4qf67BvO/xv1pNacIY/7wxTXcWYaJy4t9JgcB2OxYlSekocrbAUNZKy1zWSX9WjR
anC+RIcgCJ8D3ecGSuk0d2lxXBUI1VwrhEu3OuMmza9f058pxl6pEajgBchX0ugqHZTk3hSAKPg+
0VK9cYDNd7mgcqxxT0rlnav8XLeh2dpaGyJ6IzLr1nNup1ZhSmD7MoyaHDd8pzEtvNH2IjYTNeJo
GtCE4esmk66ZUw542n6bHG9wgjUGv1g4S9z3y8JzSZLB1dHYKwTnh3MC4NszICAcm+HYGxHkzI/T
YSdhr3nA2vOOTEsk1LZsDGvB+5FASpXjXGuAfC3z0YlUyzBj+y9JYZWH9S+14eWBFYhTFDZt9wXn
MMvALERdSVc/LMaIZHMyq1mM/Y/fdgNJBAcgCqbUsAOYzP/7G+td507JjpZpzCleBWoaJuUAFuwU
ZoXxJl0e5VB7Q1yqgut7aS1TyVPLzzC4lkjYnRdM0OSvJDItA/kCwfOObYCoxdSw18TdyjrTBCud
GwPkzFJV+oETkNmBvhwxwvN2fms/7TFNd897DVWP53nYpOSArdgQTIcu02c7Xvr3aVAHxyDdpAYe
bl45nhUeCFTHeI/R8aB46OTzL1ot/XqgxWVozNEzlhNPrwo1g9Kjw/gb80TzltvdQrhUl9OfxpC7
dX3wmF90Oni4hru3ub5pvRW2hkiercRX00R0XvQdI24gIQLVna+nrsTvZaYI6hnOt6sUfxpQA+XZ
HT3sQaX5dQglydn1f+EoVA7HOX5J6wIDwntSta4B7k5/eN6GVTKHuz6qDAui7EOBKK4ODysJsJKB
3SZ26AAP7mkGewF/HDMfYpIrqq4b7/VQJcAEw2K2aBfgEOk0ZMZU3XwnnXnF8qfKgMSv/0+Dkcrm
UUXZHeD4HLcFUyNkKClc8F7knhChTwj+4DhSH53VV3RszLk0f1x63bwpeKmnqB3cxu7GEurJGyxj
CNp0zBUheZBSWDGZbnLQQcYIimppycZMTDLxCqMlU0Aq/HuaG6+a9zrZHt3saALYAaiu0xNhNbkT
kV1pr1AJVXJOTaVeGDle1xsofj1QQyExkis+pJcNVXFRYd1+tKkYJFsX2Y/+t7dJh+BZq4qN6YXn
wpMpWjgqhxWb1/cKZZdyoiTXAoDnU1LQeBP1sZUtbzalueaYoxI9pc9wsiGhnEXq0LiaGfM5wrCL
KlWWIU5Z0PIxxvOIxunPXCDbenPkJu/0x3zBpfVkVag4DXgEYkRb7y052C8ZeiIGEX3hOuJIUFXN
gzkBe4Kb5DN73d9T/x4pP4f2mTvQ+t3CRfHXJ33GZIB6mMm+s2h0FylrJPYbz0s3UArYqIe4aSXg
uydIxz/z4fYbbEFFQdnifYnRON0WdEXBybx/YfucAp/PZFbmD+bLk65MrUv8gfau+UbwWcTYlWQ7
kRIEQAMkv1fzGPdypqHOnNWxrreDucPzzK0BuH806O6rQZ2sVnXBbhXfUFefZ4/tun8U8R2m/bnJ
d436xbzTdecLCbKFS6Vlxun8I0X+0X8Jr9NN47LJztrOPizmtrTN/8I/JXPg4k7b5T9kQVxa8w9J
rcLE3NH5DiYukEVab/SNtScBl51j7OGCH9Fl380p2EecWqYjOF2k9lVift7pUldTgoIKQJvFBmKh
NUJ6RiozQt/V9fHRUndANbpGb1ypn1fS76F4qRBJ65GfiHywWaehVYOfoFKsVJaoHYvcO34ClcGb
WdUFuufsJUkn9h8cLvodCKLbrqhPy6oIzZPqCzaAiTZRNvemikSn4Uj0iAzUsagCaLvdRjpXQA3a
hrWXXNHLMvFtlAR2yOJmaseKmiZO++4Le1BLAcTB+SiZOTAhvS3DfFoi+HQjAWen5yK6TJ9MNmjZ
qdHPnXlIXSZBoxKcTZz5D5sdv0TgEzld9BzwCTldSEhHw2tdrZkmbpzhLMIIDJu/EFjGiChxsmW9
J+9NwN6gGGJcK0py1XypDoQMuF77bUf83ARgykLw3IjQv7hhX/cuZWVb24kEBcuZxmGybrebjuV9
5yIQyXTiDSLrlbuAxoCCrdVuJ+fufw61wda8hAIVtTCGtYgCikYo8w8QHCI/FzEI4UZUwGv9ddin
GItjn3pa6fBNg8twpojwSfNf4sgkaSNrj0uhmO7a6gm7X1OACuo0l6kWA3cyTnwR3RUD2GPBknhO
Fmnm4rJgJoQ/StG0IPGsnZsgQ93/lND/+tketusyBj5SMrb9bz9i863opSEXFG7XZT2HMwoX8cxH
9qrygpiLbYNOkxtz+19n+WWpRzcSGuRRaL3JE8jp6EwDUrNStd0gzMwyq45O8jp336kczREdlRxi
qgMNp0pD4/w7yyhQF8/Hp4iFFhlVe4aiatkxsVttIoBF/rI+PuwTvwBHK8MeqW9avonJJ4baACkX
6WH45oIwjgbXj6b3yEsCmC0oRT3OUKLUS3iCKmf09X7TaXjvsyjkHib7TjFXql1xveuPqSlk33wQ
/uzrIC4LX+n4XUO4mDH5NGgxXOfSWznA4vYERF0VutknQuy7tAigA59UpHoYQ4qm9u2PGcvOJWCK
TMEStLL/KVEVSQVBHwXgXqwayplbepnP/6BFmrcYv0ngFv+DjWTfCGBXu68Wn7c7acm8rExa11t8
lGKy1cPkyV+IGx0oHavvhD1HtLmkiq2VwsimpUKAD9nHwb9OkTmNw24v/pXn7S3jw5JTg2qmhHCv
GBuMBie7ZpKSKJ7W8zrtkyN2mZzNPhhIObza0x43AyRDxPTHat9MltlA6YYHOkIka3TvRNExOe9p
8F+ta+fHe/qadV8dg7oDVXjIw/w1Me+ts6+LZWECPWmo+1LuWhwBtMS+qbOJE3i0f0BNG+3PsP5k
2UPYmtYwRaxSYdUWuE3vx2bPkop/R4jVsCi1sg/1z9ckj05ADCwGQmT7s0QBTzWe5z08wK2wq6zj
Qtqbundh2slz8xRic5gJRpycCEDhv0XIFgjwWfDp53m3TvhNY3ooXnUlPliAFVQk8AC2BE9F7934
PDCxAjae75EdDfKit2i/3YYmJfhtY5xU2ZiP+m5pc8/PLGuiQHXLJrB4vh+fSLR+hCyw/EDh33xP
5LjLzS9BoHuNE4opuApaTKAbv95DYzVCgRu42mpIHt7gzOUIKi9oBo1OeTxNJPwnuKQrbM2v7tTL
TXb355WdKv/AJyqnyxrSpP6mS1PKFk2wBwLvkFXTtYWsit8n9fA/MNm1HnvLHM7/FvLztwYwvYHz
oLrinZJmpiB+2IBdzOgzq7HRn/WFw9c7h8IeJTg4mnojUP/mbk6aAEiy25rnnNOEYmKg5OMW2yFW
/LOvL296MzsuZJPVYSNgZeAQ3Eoio9fn99VMIFHp/NYPFMKIW0qAtYRtzvt2a+Z5K+SX6ZBb4It2
RFM9z2yVPZlq4Fv64RhSx676oU5GFvJk/Q9mteFJNGf+akKCMyZA79QWywDJa7pov3yaSieCM/WI
91AqVHAsEWGh4aEnYkgGNx4MpiBulgGblrwAC8wGqCoT5WS6USGwIMYF5rwBnHqT+gy5ZpOT8I2P
94XvQoOnCXtelBmbtq0CtIsNyKHkQFX58bskUfEpASlfEsncQXso7ekmJO321P9Fy/qyVeq5SFie
G6Ob31LjSPZdPQB5KjRgartVqvYHK+xTSm/1Jfgf+7kALw+7r7/3wAcZCs9oTXRZRKkUN3RY/sVt
mqVGBxImsMm+Ej7en3U6DOlNkPpwj1pmAENUPE6TlRzdARO+pizND3xGDzB8ZWyH3MKST3dJsFLZ
qBsGMTRaEr6Zxx+7JZJSOU9RS1mlkSDKDkvLuRIWjbzEDDwB+cn0SRHNaIGxGzguuu8FUn3BOqOm
FUFsgdhkV5jiHJ7XRpbHD32CjX8QeQmgvT0dDVrexWuXqcM2ULUM0bF7pjd6d+Yj/g+ab6OfJf7p
A/KmnMCFOYDdWuBFjtWkGlLJuXuUJj7foOxD6naEV0qqPc6gIPDX8PBPLfMcckZEMRDQ5B1LFMsx
FMGeyUrvkvVu107qbLC5aUK6/9w1D1ArKcK5mf2qEHY8y54XhPWgKQfyK3nkkb5fVApqEEvQLlMW
ZzR364mDvF8DW37VVAOO3OlzlH9TPVBwzaVpvGyFduCKCiYh9GEWfNLihIAC9OkD2wb+vRNlJ5pk
URNzk4zlRU1BLagunWOM97+I/kvd43I/BSfVyrPvQsoZIxQikUnrkC0wMUdShFaXcjZGd9KnEvw6
VR7AeLxtl1yjLH6GnNxSu+kgV/FCi86/5XMfhKrF6GQVRCOCwza+s9qb7ALWenGsBxEfRLSFzqLD
QJSbisAB9ZtViGJ9Qf6Qfxmy5/xS0Z/VUSIxj/jjo1wtY0EXLIIGilSko5ZSfvOlgdeTYe96pnDX
cJyvzd2luk6Z267vmpK8U1sccYv/X3xEgd41LMaa9rQLRtArdH0kQrpaNqHhqKoZpaBIsEqrnD7Y
MPktOlx7nRK7ya2W/rtY1jc/OCKCcGzmpyotQgSCFvyosqt6FzMYH+5ThX/31TuTgaMYY1Tt7/nJ
Kd/nFXnUfYCqaFKSio0pXmoSKDEu2OG95EEFzV3hXe9zFsz5+fLyBwFaMzuVlpkU/Zxvb8kcyPMi
KBwcKdc5kgI+BQCbakSh3WKCVVsxHCcSfUrWFXkQUoMx3I2htFscs8/9/WsYoEhLn+HYA9vI6T7X
afa6ocE90GXNrE1iCDJ0NGqI7yzLz4ZX78Qgo3NE8x29RmQnSvd2pO/wlwjFyqhMuqsUjxPJzQ/X
fGYqXnKDHTIeDjvkvQ4bmdtZKdOCUBeFX3KZmvfg0WPWkvuATrJGNEFUizYe0xvPF/uU2/ApqkiX
GszkbF3bqpEd1RDgNUrmdaGMRdQH5faMK0UwZmcz/Zp8v3US5ZsEjKB3Qr3r8JhCOWuzyU+1MUnD
1PMsuOm5K/PBO/gtiVGzQWPsoR9ZqEEyZ3bZOkjLe2dROpacnWk6joNYSrjW23ICAb7XVpFTS5ft
B5EwgLlL7RQT0GjHeslBgTovXpGomu8iEz0qDqH/lmdA1YgQK9TlyRxwXfauzwfiVDEAkidKYC+k
qiOgsG2wvtKSgLl+ANiVTtD6A2VczwKZII6ZMDuyaRTN2aldQDASGhRvjfcXBoe4o/XxCBmkCa8K
7xJbNJUlUJMH7LlUhrXR6ATaHCv2uA6I/i30vuYTuxcqXe6iW/B30ktpHHrXrtXGOixRtrMAZLJJ
eTRY1j+a09FUnypYhO5rh/jBqjZRe7QzNT981Q/aJAO8cO0Vo5rEFP2DNiBld8B3MshxxIy4N2Hi
+qnG2cFvTJyRxCPFv7OTUJe1cdd4NNSUBR+4rqCvLKMTvH/ElI/AnQrCRRMKuFD3I+LAOjP6ex7F
s0XYhKTDq2cgn+EU9CVtThPdNoSABQlewsyEQ6diZl8xdx8M9j4Q4X2vl2MS55DAMluubFjqDdMU
egnzaO1btE7zrLnXS72Y/QmDA880ltZr+sYt/13+UscrksgyESIg9Sf94Y0gvE4oFv9KtDeMhd3a
4Xp7NvWqTCa9YUnqZZy+qeO43+je9zJG4ml0fyu81BaYyqt6guQz55/By8ThRe4vKu6ynJJLIW3M
ZQFcKwQIp0xIZ6QOy+CurStbH8ufJaV57F8l9TWs/WdEq+KXBhoCDSjIacBwiaaEe8qd56yreMGJ
mCec3MR/Yne7k0DyzPPIdy1mO8h2KBzKTHREMil3G7Y6b1jvVZfkKpmNbC1Cv5naOERuArUAQbeL
578Q8LTxwJKE5wFmVxJ+IVCEbVBjju7vGC/p5lz62lzLUojArNfR9yhgxmKolMprGTMaqgm2xMR9
318RpjK64UtfKxyKMb6rBdmiGUWmXDESm5BgMPH79ry54gq2g7UtAaI78n19DMM+Wk57SuVJk8Lg
q54J3HD9AcMZClJE+zZ3vC4BlC+qtXh+l1VX9P+EPIL6LDICNXiMfqyHX5GNcC8aclUoaV4VCb/Z
t9js6q29DdKjo3sEoIMKTSshygGsFezqBjwG7JdjBUBG/HKl9gBKDyOjr1GPxGZw6gb7f8HisS0F
+xwjnKg+k4b0Act8HXeHbtBLLw5V0xDWYfgXps+rcUMw9gtGNRl1o8xlqmoGKJZTfC0NwmsjdVo/
CkAdiMti9ifvvCKEUkLO6mE68/RApF99MR1ua/jtmzq9ZUfy2sI6TGUuWoHRcGx5aLjDrTNti5ad
w2KCFHZNCw3tdMORYwvHEbgjKqJ7nFNQDITYVMz+urykU/gWRVg4oAwavqzqm1bycj12eNKcBv0i
toTC1HiVSsx+wnePY9RtKHKuAks38qFIavV6uD5pIIbytzrXrURglz5DceiKWX65Y5TSCAu4jSqD
JwYMXf8wGH4DIMD1CsaIi0b7Hoizl7LwRlJiiCZ9ZRBKV5z03MPJPMzpcm9vEcDpQ5Gd4opQrGwD
QbvKPzrilQ5qOTSzyXaOB8H7kE52qANA4VS6yEL4PVszbSPQO5QIr/TC6IclS/bkXyPTSHQvBg+I
kp3couO7kHUpZmxPogbvy6uf92nNe5P/fNdXucuQiGWjMUOsTczAAm5NoY7K8ABaEWIRP7+v53PL
EYlHEkPVorYX4QenQWNAohhrkcnFviS3rx99Bw2y/k7JIiUIHaKtK+6F6rtE7ooPQqBVl1kU3gRX
ABN3/J5Y8UVe/Cptdc8CoYto1XaAHvycvrfaTArL+NBhMFJ3jvL+XgwQyv1Gr65AncK7g9mc/4F+
lgwJQytadwPRse5IYrlfQhkXr92y6lXFh16eadA8ZhEIydyjJ+9T9FFZryYDm7txZekacsh99TTX
7oVieuA7lsukEBdNR1feqXGjqaDeJTWoipsagexghLOxKd6T78M1BBUsYklr/mTJzLw6kYdIGm9T
CKZHqOerfONskhuvCrvsys7AR1+cSLc4QPkrrGOQ+3Z90qRgu6loRivvmucNdGByeaCiWygy54JD
ORXZsGwgz+6vkUeuJ4efybMKWAtcm40EdFdI+KRchH5DFvaRjmufFl0FH7MfVsbYKYHObxYUHeSF
8eGCJpXv2aBSbKiK4vOD2/k/bU1PNwGp0ij8fSQG6wZueg9Llqx3HVgGRTcROiTRLpPHv5cRLb1w
7J1ks9ig7V/8Pvx3WseSciwSPA+M++n/j5d/HVn+tfcxl2IzBTRUs7dDyV8Jy7obvJ2I+Resv4c0
mo5Q3rq0o8rxS7L53W/ZiBFma1M1Cw9aydOwDCtceLoDKMIBZV91Qb3QXShe9y5IrBWWj1O7KaRD
RX5ODCfifwArTkw7sXo7o7Tfog84cJLzjkHAWE0gjbiZWCI+LZnbGOUT+90HZT3QvQImyHXCYw97
edm4nAUBdpU6S1ODP1+kwjqhlSPUliCtuRe3Fb6r5qOAZ9Rx/XJZcCnB33pJ7HBlX5+z2sP8n1bX
7vdlOCfiz6n0J/uh1TT0z40tip1tfNfbTqI15/FytUWerfaGal3EIM3h/d9LyPPKRdqKpkARAMD1
p5xA7o1pGQMxW7ej1mvIPP7mLvEpVct98r/AtdWB+nh1+nd2s0Oglo8eLTp9Txte/WcslQWxdMYg
ZFzNsvouAhgpayiX+9dRfX2dAEwOaau17TI1NobbMyHArM7hk+0vpJKiBPALYE4QPO8zBK8q0w+E
P1haG+8jYTElS9tKnCiSzFPh4qwnzatRuOWZbWx1tE7O2lmzU7M0907ft+LPPmebnb0CIGbxAJfW
xKHFGqg/DXTqkO3uIJ04KFLy4uGXUhUAa2KCD0w1eim8OQsb+fXrec9EBnmGiXu/FXFpNDRlvaYa
0ilr6HYmNS+Kdsl2dVgfEeMacUb3GUiNGg/FEcBfD2CCpLo5/mA0xcKauMqE8b6ZCqKooMRRK7Ui
3FZoTDZ+WoWTYlSH+GL8/9WZ7zw2+Kr1Z3kWIdsE7Izko3WapimKDXWeAauyJRX/xA7NPevrL+gA
1uavPTlNi80Z+NO6XYQg4q2rEIB2fCf7Jc/3mr5UDO34T5BNFC6KR2tYWRaNLlx5wxaYtiqBcVSl
82qiz+sFxqANhlHle8JoOtxifM/oHH6Kr5DKEm5YTe49RV9sveeNYqWPxTzIXpN+3DJsfPi9JmAo
8XmkqSyFYf1BE48jk/PJYrF3PlFNnOx4KojRcofs0kumRlY67cAmp9Zt39cuB1wVTTTSOSnwekxj
uj9bi/zlQjZ5Omh/dXhrE0UzsWaOIu4oqQ6gOL0UCmnPmRTIWNxFxgh98KzxZWvvOh1eBt461Ijo
fh9dFPI/OIuCnintG7/Bvi0Ge9tAcM30PzZ65eX3FP4hytOh4whNcqzB0oFYeflhWonkPusC/QDn
2QMvutDsiJSExZYYs7TOwIszpmNukRNcl3hi3FMenj/mnOPuL6pew1gfnUxH6g6xANL8BI2XhUS1
2vLudfy+7+s02O8OdSqQo8LhjIlu5eI5XcQaN9FtItJhA1OeE7g/tKZlRmavXo8o620mhOGPHNJs
QKYXky8lG/G8DFS4dlZnsfqOkrjlKIBANhy2iPfZfgsf0BTLAgHsfbUjgDFHMpL6HWsZEYE/xo/g
joVxE9jsbLQUCuknX1ElfKX+CTwE8lYJ+x0a15ZkhZyVxaqDZ1KpTKQtdxit82TtmZDPU2HhTZ9P
bwPPMPT0RirexhLhzjSv4zOfmst1welok7vBecv+ukVgDLazrzlZiRAXRPlysgGWxnFoSL4YUu9e
m8+3R9O2bSVuVL2FvpxAfBZSDljbwYT+jqi47WmKeK+RDqmou+la+p8TrgSd6ceILmo0EbOhQzxi
WEDzvLxHI2V2NRkm0OonCfmGRfqYGpynW3sLiR0IWgFxPk2ubvqklYzsW+PkUgsnZ4TFAxmmEH5h
KTu29bAwjB33mFp5DB/6SeAp+IIKsLjYZndCiFgnELmryN10v4OHGJna0nB8HyjRHtZgfETxYvic
Ecvfdml3Tjdq1kHdle2fIU9PwDPX7ijUtdRdgRaBNxTxZZYCXWPqQVEeYXYxKl3hg81pq5BTN3dW
hDu/Px20zzVYHu+FBCD0zW55aQbk6UQmjYpGAhUjIyM66wfB4J3QD/B9zL7orza1g/OyF2iBizoX
Vce4tlNj3QNnfOc+FyLflunFNyS11nLvNEeSHcwEgoAOx/f7wxh35TBkhbl/gf10QkDGrAAu+7jM
0n+fPyA0b9ERpoE//US1DUms0sSq0DMGHEQiPj3T24qgwAV7oQVf4jUpkbwgakNlx5CWPs5JHu3B
q2HW4B4TjJ3bCAEiztNz4eSxqJ9slMjhGGXEH8+eQ9apG28Td2LF/z2YSA4EDuGosRxlm0AzqENa
qp09PRCgSLo+Ov9RM4vWtVBx6aWCZUOCVE5yOt6aOTO8NJ4Dg4pB15vaV+01P+iVZ351ZGDepGJZ
zN42PJcAGVec8P52wD79hilycLUjI0wlVmFLv/kMzI5eWHcsAQ+PAQN7bCJWap01wLOvzsPcvMIU
i2SU5qIRwOb652QQ7suhgEICg/O6KalnkRvaNYrDZy0lyhhVZcJMDMkfMBfExE+Ck9My3C884Iq1
TLAcQFjG2RWRA6aKirCkqK8lLtmB5WjIdcoS0angR9cJExzWlN2Gz2NqAN8drzirBHTIQzVlWh9u
BcRaVJ6A46mr6DcYHPhltXvq02ac0khA0TrvAPL8IswI1NDW73zJxpa0h8Kf43X9c4n1JMvaxnhJ
T0Ii1riK05IaPxlU9wRVcZ+jCDVZ9FnAd8jbUrz0fDSXGzYHOxtpxEgLQVUG4IZSaQVcAVn2c0Az
7Wg3iORZeMuOJDiIcMPPhM2EA3oJ4pGd3TY/3lD83sMkXuNiUxaZb/708sIuwclvj/NB+PigBVdi
EDyduU9ta9y71OmATPVDAa8/wdKEiOOwGqM/pe8TpYZ9YegcqeDVQkUAUKZ19zthN5t+xiiLIkub
T9FF52SJ7DVMaqPK5r7uRb6GGF31Uqm4O0HIAxy0w0f5S/2SfCV7VYyeTWwlD+oFUSJCzZtPgb5j
NilMnbAPi7DaUpDfsbYamiVHlwFHvjckAr3z+mn6VWWhkczobTmdSuDCNY7nZa8ClMa84BqZslPC
o6p4QehBDYhjLgEyGIWV2wsCJWdoo56PNrqq8wqOeeVhesqpLtqG+Wng3gSBj35iIQNDGsIA+3AX
I3CMgDswLAFZ8vhe+OcUM+RqDmL67nRN4fWo7/U0vv8B9kb5N99MTzCo5OinYpXQtZKZu530MW+i
IKhmKOs0sQsfl0vLmhrKCa01IML75xb9e8Y9TUXrjrPZc8oT40xpeVG6SR6jqKLU8SwOzZCT6iod
LUD7lV8l0a8Rx3WjRkaA5ktTvKTG13Qv3hYQfRz+8vL/k3CA/VX6SMSTWFbySWN04LFbcbmxpRLg
1bQiAoQS6wf0GXTk8DkXx2vVPLp5ZMl4ikI8f4C7LFnmHy5TWf5bQa+CB3wzD+MStHCcy6IymBso
4LIPDTEF8itm2d3VJ/TeRNqnV+KONZjmuWFNg6fsbVPJz+GkxGxNo8qKQWKzi9K3DRMfDYOX9601
vGnV9OVaDBLMgCnRs9JwFaxtLkF8VVC+/v6fOF4XKT2gxvnaTGYbJES6k86lReu/QUJS424Qqe/L
HAJ7PtQMAD+UiMLNuOJv4yalP7I2GOGjI32H2FDKtQnYuhdzmmwFzZX2bI2X2LTj00freHaoFS9h
gxhH+YzB0gBYRm1gv4j5Xai64Z58yA8S2way3wlu8L1NDjFcOyios2XQy/T4c3MO7oVvmr2e9kDj
oGZQ/XIpHEcxIvYHzn+sjhS7oBlTxqafdU66Ao8kgcJzVfTobFzwTGGq7FQov9sUiU89fz3xadXO
LnMgCX+Y6L8BiyLtNQzoBkKmAsEWNphP2kid8nfyaxBf5Sv6RsFBkzrJ0OoVpQEMFaZjihx1nisw
/uyx49GteXpMY3TxP69BgUPW4F06TllrPls//WlUfUHcKszHIIbEG/HT1o+bVB2RuglASIQ3j4DL
IrLZiJddSaBL+Gn0EhkDCiLEsIc8r1IlEPtbH+Pbcd/cwh5gDZ66+VpppMRgCI+e12L3HOx/KzM0
VbMlrXODwgZ+HOOaecIe6GqiTAxVdO4JGalFfP5Sjkkakdvb40DnAWquKjllJvi1tauVFZSV9gWj
Po6YruqFL21cSpmqn2XvhQ3BbCmLkRh6scRCEcywp/nfbLl2C2nbifhjK3VECElAAk8yOtvgIGVx
OIL2E9sMJhogREuoR8VnK6/LZOs/lBUF/5BjH3ntm4xajKWvQXwP2spN9CIftTa8Ehgft98zdBHA
4Bp+HYzgX9v2OufDANVLB2cnaeLUxvLB7zaGqJZZQcTUDVxJpcZffGfhgJSd3tsRTEl5D3YulaQq
NaUNr904y9qeUVYBxNskQ9dO/VKAStTqNXVdq7SUmTBJbtLQ88XJLzR68DbVR7Z0pXUQZlqrgbtH
DtDYKrZ/jE82XKhHXAZr2L1Kc0VQELOVkPU/8szsbbfyGsta6MTwRBsbQSsftlkIQtqTWoARgmbg
kcmGVVnmRbO0LHsVdNDC+97vYHW+8V+ZUcYGxxGEfeZ2xzxu98rR5u8xkaLUUZ3EOw1VB59nou7X
5KtJ+mkTM62d7XgWz/MlnPqv0RvSRHcWYeKxUHBE31o+HK24Q6Hs+oMHn4CnXcxWtsDq+lZE/pAX
LP7MkDxEcV6RaJnIS36ft1sVVWuUNABVPQU3FF3muOt1R3pyeOASVlyo/ggg5/xGeBG3OrshkPZR
dBPlS/2UeuBn8w9UCtdX42PY1gFBluQtg6V6wSM+Jm+GtWwwGSxpzAbZvoAFBw4KbIb7qu5Z8ch8
W3KBga5WmWP5b/4v6K6LQwqsLFkboba5wZz6wYG5vGve3D0kPrGMjlsjwXsLpBUwvEQeGv4/fCsR
w6C80fNoaTYbz3JWn2N3T8auBPNsxsm1Rpx3DMRo/OYq4WDDOIFkrFtAw0qmCAASWzLrE4ZXd8Wr
I9q+pPs3sS1XVAUIaVKXkkpN+WFjH3wAYgW0PBKe6CvL5epQ2XENACJAOdIkV/Tpss4hMnVs9Qzm
rPknkCGndWVbRkUQVTrocqGMQP7B/kMK8HT3LEDik6C9OA1oX7oAa9o4qEEiL3Yfh7e9+HU1iirf
MI2OZUWU+AGTmuZ1otmrdqrRDC7nqvoDXnwnYxMTUIgMIBrlx6h8ye8f7otHuTn+NWFxKCLEnmUc
rMd9q3iQhKsjsPxI+Y8I+gPiIsjT9o2sJA3zpCL+rFA2sFOmLWrSkPUwucEVRRx6lEbkT9X8/TuF
MYeMzAbPmc6BhK/IoWTbylByHglBUghXl5lTpOVHbNJgltwi1A8heV22RQWgweyMu4vm1s6vC9pE
0jjlsqtIR06xm7DEZCmfumdIUref2QRXU5YvwXaXHRNymBNkpo3we5licHZct4SFj4C9ArzJdkkk
WRAt+wFbGfCxxcnZD3+32TUIXVWMhlMrRDhMYH9zR3NJXwqaRbBup4bgk7MdOAT8XxrYksYkw73j
h6u2kZaGlUda+9Z3kMs/OgIjW2rql6oLAS6ZVRkbbNeulKn6IVM/nhuCtXDpG076VZK2B3TmItMg
Dou+/QnpzXHfWSPpwHCx0+eSUIPDlQAQsg0vp43pT4LmrYtFpUb6nQIkgQ66DHm3T/xhGfacvRCW
DL2080aU8TS12EMr9I7ImGGHi+R/JKxXNQFfzjMsJBgh25lImI0LHlFzr+EGYqOeDP5kZvpyI2mT
bBxw5Qot+pJjsBFJz0Z3595orZUlkbxKZhjpukUIbGfACmkLIdsBIFvx9OVYhA9ys0b9S27Zo3w3
+e8dqZ21rZ30Z04HPLJMFxiPLEsUGk/Omm/4EZn/71ErmL4Y7hAHJy9rAgJDml+BhWz90P+atCqb
mBrI/+AkBEOPhoTgbmEpYQSn2Fb7K7Xud4ZQvaUFGztVGsYOEzjkkbnQmKh/byJV0Xx7B8Df2hh0
bq19GCyuvItyw5HoO8XbujdjWyO37GpjN13v03SCwZKokNgZ5raK6m9QCaLIJVwM433B7cdmZfs/
5StfphqD1THIof08y6B3wd0oVW/yjaeG+oEvqtCpN9RYltmdSMcced6hAa8h6Gbt2uE+msJz9bij
z8SjolXdAfcPlxeu3GjWABHBtdMynrlx/8W4ZXIImgLPNARhXAE+chYD6TMz3oan+l1k8XZPMFFb
vbMYATEyp4/GBZRKtfuAauxmyx0D4UGykMXdbqs/bP+HDe0QpqLitNJhJr4fFGGra0k/VXQtEODL
zhosib7qil/rElLDOwQ5mc4GtAEJuMRFPcoFy/6zMP2FRFserZKVVVxVEJWIaQ61CDx09D1NR+J7
Qswnk+LBoEB7Vs+eQ9XP8Ytefe5t+sOIaLTDC4GgIsAVvXrcOHJfx22Y4Tc8Rzz6jgvAFCqvnW98
p7HaANHP03u1ayET9wX/mbJY/0wd77sLRdxhm5Y5GW8bbd0ilnV1PHaWzhRfBlVwff98X5t7mIUS
jvpTebH+AnG2pcEnuUr2UojQFFN03EQghvz2dGOCTRrtzoLGLYTAwmF9myVblJbeMI/gwjMJgQpk
9S1X2+3E9ksebkEbkJHJwfbd6uJw0rkG36iqTRaLzT3gg3jPf+L0sErdT3wuMRUB4jWa+zIbvMEn
oFTHelMgJhDsanHVmKjW4f6aJ6BYFx8HSh9iJXjWsuPMVHMUjn75fxXHBbnzVUqLHni0fwO12VeA
BOtIxCfnqfInpgoZW93Sv59NME+rYiIHO7Eo0PkWsjpVUe/HhVJ7PDVKpoicROAdvtxM2Ud41jtw
QfXiemlUVFmwYIBmS+mGqb5tBawkgpHNt0OuYOmeyBdjdHDF8Re35oJ9sopxCbCC94X31oo7rbb6
5suWDeVfXR60+z+tMMMLXvOjVrPMSfQBXnPpcuNUlxsEMN+yennBGtWHdlzlF8Yr8wsAup1tE+om
8GuewsbgUlgUCXrjAXkDMCdFjRJh7QLKPLeQYZNJZcieN2AmHRO/5pugTY80W81N7CUtGsB2dxEv
aoljeEh3cu6hlfDvg2jPyR7rTFATa0Ox3cgBiwIcM7HFaDO5MSvw3mg/lyWHSRc36bhmrIOQ5qL2
H1Bb3mUEJ1LtLEzA9yH2za3kGHyygU20UrrSdzZu9rBlPK6EcKAf7BVFWffRunGbMKpyT5MSH9CN
ZSio20Jdw/DQTieEnjcPBW//ytJumiAL2wcmmbQMioP4Wqg6UhdfZP/Gvc2vKiWJYmoHsNpK9Sd0
MFUOjjKYLdWJrnS6Pc3TNJrBbvJLp5U0JcS5QplLkJPOt32ElP8gUCYZZEOLZ7nT/UAvmULEjTZi
pAQObos4VMsH1znTm8V1JSnRdQMLljYRPWBP6Sr4Iri1Cg8om0RdEwZjgQn9mvxfkRVtyXNx2yOe
pHU4EdhQ2NLPqZRstsVCJnFUhaVNuriPCueJCMpy9Pe+t93/GotxmOg5LwRbePynes45kuA0KmgD
iU6UHr2g6Ln5apAsOfy0kRlzD/JSrRkhlRHrvZZAS7FA4rzHel73zh3pdKvgI3AshafED1ijy7Ph
7Uw1soCa+VF1ySQx8Ic1aM8b94XxFO8AUeVbcHVAuQhaj9omsPOXpINwdJHHO85d/EY23ltfMWBf
IyfgKV6GyBe/a2ZjstwzSAYsRY4+wkUqveKExNRaLXP1pOrCkd0K9bhkJpX0fS+xGF3O32SCn+xQ
lCw/Ys12qOlpfdPbIRj+zkrRk/X58kXmQp7D3Zf3iRVbMNVoAZOV+WQDQUwPwGzNE9iaicxQgRYO
dwdD8AvptSWiavB/jbOk8Q1MbTWUlgfqpBl2GUA//vWudKezq/PpNoMzvaO0bOJv2Qky6MfTOYv+
4qOhQUNy1+3zutBKukJ1wAzT6gq9gihEKmMDsmzUp/WkISe5rRg/KS4CG1zsZ6S4bpSVaDrfI/4+
77cDZV/pxGU9KZ5DBBNT//Dh831RtAbCfNCOoU3SBssrOsCvmduAy+/qWKFByF63rY+FCKAtvyuD
FcnWUxgONmvqM8GjT16k6z2TbZn8QTr03Kk8Hphzpbjq968N8+MIRNexm7MPVBBmSllT44kcs1pM
XMm9CZWl9Xvmgsvx52uQXDLDhvU8SvadpzMsFslq4ROwRnTUXHcLE7rYbHWy2WTPP7S59Lr8dEg3
vf03Wxvu4kZFr+YcfI0a2mE1bL1hn+ygVkMIBujvlCjVoqDgbZ+mZ05RV4VlIvleuUtq7J7NxgtV
1mwmTF6atnSh8MUVfIBdpP4IGf/gnsvJ8UupTWXEUyohAl1tvMR0fVRLGv7rD3ryfXGAnfi6eXBk
wGCiICETEuUD866NyzFxTm/tk7a9U3XxQBK2CBpiKGpDNut87RtAjYFOA12t/5hmmhu2QkspnWXY
wtTxT/oiDV2mdinhjPSa/P99v6jlSmYKep2BXuFTWcENl55Eq8/JskgZJzjYO6CRPZTEMLXWfZdX
BiYIO6thyyyMMk9kzlpvpjr2Dvz+YX883d20JqB/bVMsXdjMh2FtoZDY16Ez6pI/13Ezd+mMGA07
ok1WdJrB6Jy8csJQzQ6PLN0inhhQdhh9op7t5UTED9vQzayprc0+sZlvR3VyUyB4KSecXPBZtgi7
dv9DpNNW3s6zFPX9KHLHMILR4uUitZEVA8mYmlVzG4lVmqEYiHboOT/awrCzM1Sd1g+uGn20zEEa
j4/CY4e/uJdEkxMM99WqXGDgafhNUQuayVnO9Z7NC6dtlxSq6ow8yF8xGoQa7QLho7rw97gbhnsa
R6K6VpbFE9TiLqWKcIfwmfAf8epL65bo0idoaIFh8NSSavxiosNcOWKuWoGhR14zQswuCFZZq+6u
3jG6Do8wTBdhKQJ1Le2rCUsffm9tOUHGbmuVwc/5cssQltBA6SypPykO2t5l4/+lO4nti+Mpg4p3
/UaIE+U7oEqNImsIjCbWGZd/xf9dkOzg6+m7ppBaIELpv2XH1XgL+Npyd6eQ9s33YCE4ol3b3Hyo
ZwqpCq0afW382/9axerGBvZ1/Y9p2HHwRD5odadfc2/3ljjm1WbEZleufHWe4/AmoaEqBhjCKPIS
EL8ZYQU0wZNEW+ieL7Y8fxWd2KruemWGTsS/4vOPVWl7oEtzzgShmQysbMriSp2zVnIZ20IwKV77
VL8Bn7Tp98JC8eFuylzSu5NjEtL1uKnnXuHELyF3+VshbSIkn8iVHa7ZItttPG19429nmrRdCN2k
lqZuxOjsI3p4qIXv4V59RwhODxzwx9Qh+xQkJR+567aXmNGxYiMnpV4Xb+i8GC2QnWN9AiC8mHcv
NxhuhGfDgtsp5usvkIqpAUZc743irQvwkGxSR9aqSrFWtP9hQ1w+6x4Ch+0FcfPeFrYy45IR4yJo
grL+ebUobe7iN67WqyAbqYnp3fHuY9uf5Z3ntu4cJbDn8HU6uQIt37vh9GDeGKGtTa9cKdY6f3J5
rZzSQhnw9GOmVGRoI+i+dzD38N28zWUzqP+kQPx/laK3rnbYvmmIJitF1YUuAebyk61VSnPKW6xv
ImdOWJ/UI0SikpuRanD22Rh3IyZizQrxgwNu8gdRA6kYGt6nMrQIz5vZmc47ePez2RktBstCdiqJ
BYVi/jCU/Pz0YHPkePxVaBr4hPTBs3aCIpSOfGrVKqNeVq+qMVI6ksBDmwSjYV5Qt1gI7DydIduV
pthFXsMtW6ZcWAqiAqF+0JLzoskuwrJ1VZBGbXzUWjQjoi4PjzqD8YRcZyBi88KYFgSPZKGvzuaC
E89liN/l54VOY1RQZpAg5t8TCzNaYM8K7fqiZaUTTZpucxSX9mW0X5bkzfKfNqvL306FSmgTmN+3
FvKFUPYCJW+NNpC5hhcEijoMfEzbLzWMgr1nvge4xz9Vexci3jGagMUPmr7h3T5zbbUyo/mdfC2P
NzDFIFIV7qV1nbuUXJNMfoqHkjeZHaNraR0ZMedp5xZfxvFKKbNllYOm0RzFEsygNpElUojgXm65
wqp70HAFYlm25ORZTrQup0xjmJODRNiy41NB/Qo9sdavxbyB9lxc76vjKEYpgVwSuXalBvapI1Wu
rNqJKlOLCGWdiLRV/qWnH7d/vg3ksrbgFwhStePiiTOo4FKmDRLMqvEVlFhOoJcDhM+Ur5pqFbPR
/Cvn1td0l6JWhw7FBmQvj6lb0cXmA0AmQQdaUlQKW59BlvuP5Ly3Hw/bXf3wSmxn1e76vX2waizS
U2VsVPuJSRszXOE2SYB9ZFP26ioP9zEOi+m+n1DDvreYlWDzAztx/Nki1HVFoT7MDMrUWXVy8YFG
dvvijwlobkq9jOZToBaLYfnrGFPyMb1GB2bmkn2IqDWNZQebXiJYRMyKmv6MxYT4aj4348vwr5zV
j9nv64/FLgSB+LqRl7ySoZxBWeE7H1xkI2JNIJE4hmM8LRVpDK+vPutRqaGeYAkVUi68QjdfZ9iL
D2lxAFnZ4oHCtPaUuS5SqQAzMk1D3V9XS+TfjzEGvglLWnnz+5nMU8d0VLVS2MlWIbPTY9PRjs6C
ockDQlZt6i0l3NkML4nfic/r96JgDCfZKkPAvYwqHEQ1m9yCxDhBM3TUvNgCh44l+fHenQozFztI
9YVvMD6fZg67UovfyKBFttWmNyNNnucvModBHR59wgOZb6xrGCYKUUH04IRq+NX18BbSVvfxjwKZ
b1lX/HtYCKahdFiAJ0H3XeK/Pxq6EYSxVlt71EKbskbujjOAL53+LUiQsfrET+YFtBfXgUBWk1mY
1tdoZPFhgRLHoVtx7JAK6SLCQUcTq4z5qVY8muoMtpfwmpUrSHaSMw3PUPMLttb1IUXwHxTbPl4x
F7T9puHUUfqxGUlAT1dllxB+3iJgcLtXYaQ341D+S99EKq7VJyV9zUvByc/ci97iN9hnBo/910SN
dZiJ/DxSeuwh4C+m9sxPacna33xB+vUIUXZUsujHGNzoFwSQyQxL6bfvDPw0bdMdAkWVB1ftNDyj
JqupT/NuOTmTa5W5CMk/f1VV1hz/fMXc/A1CzMfIudtWlkb1yXloU0ODA2l7YDQ64dsptpDaiz7T
/sN9vKJWLBp73VFlHNi+dWFFpsuJtxatDYaA9Z65b7WZUdT6G81HtC9KeiMr8j/1McG6I+pvxaFU
UUByoRnrzhioAtQGMwcJuWyn8cWP1fHezLNn22ZSHshy2SpLkeivpUgtClsracCmIK2ttigKtmTj
E5MP94i2u2j9Bcl+vhqnr7Rqumtcz9La9BaO7xVSmWkMYkY+30AjIVrxo4zC+a4RlAK03qfON4SA
LYzSkudu5fgIBG+J8f9kewTvfcaPx4fWCMNQndd98+gBjef4gV4FnPC7xUADZ8uKTD8VobcVT6ds
5rdoVoAHbI/RdxPgkBvdDYFvQIyuvd8kPuuVWe4YPI+DKLFo8uSy0FQneWs50qcN6aUJ6Wh6V3vx
35egpqPPChwTRq+rfnNz5eqjpfHeB5fpCZQBCX/i9xUHZXAQCg9C+R3blAKk2biJ9AEuGdam3bHy
ePmiIpo/DBTBYZPbZVD+DEbBBDEBXKp1mSzUjNAwc5reQH52pv2hWTvUnm9vFzsBqp/myek/31HK
0sYD5zuo2gAl7yYl6LFwvZDyx5ZuAFTKwdsj5ASCV2ib451lbh8J+i4Z1UwshBoGvtcNZJj6FcCe
9wgqY+rlGpm/nKNIY9re4ltdcvF9kWJHyRQKF/lw9yFgipWfWFe9qVgFh7iQuyWXsQEOZlVluerP
n66y1pvzoo3czCqft0zXPqJPBq+D6/ajmdXj8PimiuhFVpObQbH0ClCSiNCeS6OZTPIJw4VvKipa
08Ye1vhrwPot36DSkS9SdL/eRzXuRZm5vr+H5TVy1A9/ijoUJ5KwtDs20XhncbwPBjoLUb9ZwFd6
tFl/iHa/lFuYVVgP/w/CjyOU0r4sw4fl934a3ChwwiRlG/zPlFyLqRBjYdNwFVf+Q+ZjRtcDCRSa
MGZ7NivUf2vfQ6LPahHfRCJyGwu4dSLv5PmpDEOIgZKZWe8H97M2oWv4B5KafcKlXq4Lf6vjELhv
eK93MtZypenpMobFdfNrySBoEPJo2ttwvJs4U9iAFWxiUc6UplsPZ+lUEIPk50SAgLx39jFtWROO
sWwiLqshhIgfdsgQoR1lqcc/2ieYLteTn20SWtXvCB/jku0UMcazRGm2iVn9ufFDGcVmk+LcvV2w
SYnE5y0cGgMjvfZw269Nlb2gCAVu2pIg6s0D8Jswz4vunBfKL1qUixGhRvk8N2+a+LHfZEQnwAxA
zRsPcu1uvwPnceWHRplahdElsMfddi/BqlXduHmPvRg2NJsRKLkBP4avA71YZzfEojSzBvUHOU3Y
RIG+6l5z50Ub4Td4159HcLLMREtlAB1lqMQNJhqj6/N4RfCSlgGWNkDtafsRbC+YE8nsZRx5+a+5
xP4U4qcDxw7U4/DUfuFjA+XUpdiBwRycnzk/Pc6A0AivLPgob6Zr3ujBy/IxU9YWdushAbzqOf2x
K3zR+7mqp6LagFMhlmy/5U7Md6teTrSTrxu1igFiV+UgyRG2uRPxO8f9wtchjH+tlzmwY014t0ye
2VMXrPzE+/sOMjqZwqsV25khWgFaXz9ST4bFRbrvmYqKDCKKP+qnh1oSsBPVa1efdUzuzRTV1lKv
N9HfK4gS2WSHggd2t5ptaeslnM/Kxd/47JLzx08QpR8Nog+xzlzrslLYbvzNe2vUjhDMAfi+BGw0
LtiOvj/bKsZNwzt1fcb3H7iCUjF/p/QGf6eJ04MRoTwL2mesjIE8P3V2OtD9UCb0SwGrZcmfLH99
kj1vc6x/muab//wo/LScgOJFB9Rf8Cs4J8PJxDUrlUx6iCgtEAIjH3ffrH72ACTpKbPWFXf/lYvy
OGHD6kRt18i+J9iHwTn0v6zdpMHr2jGO+43oke/0L3phoMfvwttQrzp3JnEgUEn+N+Z7xKaR63Eu
zP3EnDVEiRJ/EqBtMf1ifaViEobNeQtSmLSgIyNMkcuSJA7Z1G4K9oTBWu6LdIgBCxJLTVmBw+0V
YjNeo3Lm6CYfNsgG92FUV5CdGaTgXdyZN+X6w9yq1/lWYvHIsGpYHTY8eyz6FHXwrCp+1x+jjsqe
04k/8TMWcdE2hHgD0tLvk7G85adJSb5UkrP/zzQwpbmXWIjKcHcTjHceAUpMPriIbd1lO3xNoGD2
7q5OFQQuf+jYtcczSv8ix4T3m2SR0HFc3XoqkCaj9htw3/bcTSMSJsa6mYhrQJd1sYX+3TXMpSIU
ggWgRQ4Ke90YWBxwoDLiiXywMQmNgapw/TWbsw+gagz7QSxeGY+AqqQr7B9uvlUhIsD9BkJZuXZH
u0uUJoo7WkcnohdxXvGhlSArxfa7LqVNQwW6wAU4XNyspVhGfcOfU7NcKVgxUkj8Qd3swEfNPwdJ
sw/aG1NM3i7AlrJss/qgGqtrF+NXMHPkRErx3YMqAKcyR6MaYJQM4mgKNM7fH8RXWh/X98XfldEz
iJGIXUeMMOzGXFo7g655NVSCZwKmicwqenjLEmGKKpF6zUnV1ksLGPChjes/U1WITvHmvcjGaG7D
2DJJixw6IxUutUWq5oDvw7N6WZ0wGKkLBKIAMpFL4+45eaynGtsu0bPgOJslww0v7kWzoNIkue8S
6TjIudGnRFXVTIExYLMDxUwg5EqKXb7eJtRCQ3J6SVKr/hBXklX55ugomILqtIvpbD5MRKyhJERv
lOftCDJbGSRKntplZU52nBorGk1u/yS7b0B+Mudv4MM/9LMhSQxeK0iF6q8UkgA7Dt5wr9gJXYpj
5k6pmKPtIs0ln03Oa5udtWFbo2jcSTHrz/m2aLW1vVBaTRRbyWh5c04MPMB5MIPW934OfDwSoKyw
/kBrSiumS10EsqD0b6QPEsqpTN4gB9X5HUi14TQaODNFQtp3YvMLSE4u9RwFcZo83o3ICxYb0QaN
9IU+g6p/y8wt+g8foxqtFstiZcwKRfqp/UQXNa0cz8d0NkEvcToQRLSmSaBY+BHfnxW5wqzjikvu
fUIDmVbU8xG3eQI0x0FCU+xJX9YFmWt0DCp12LWW+h/4AHLmYC75IGYZUYT636rPrm2iHIRCeYT2
3+qJmILk1l3alvAs0jsUy1dkyMJ1e2UCgewBTOUBz1CZbrE4keU10oFUqruU0YsQ9wVdc+YBUFuq
LyBxzr84V+tGL+Scm1dQeq9a8qUZ9t0E7xjbyHzjy0zZWR9R48QcsD/d8r6QkjzOIkDye0QDp8ev
H4LvKLnXKG7W0iNDsx2SreZCFoI/POXyFuQswDODTrp9Lp/j8bm/rZO43j6S6gpFqWNJ1UT81dKU
iZnxp2ltTDXYGJprO0XPqb6nQtqo+fixPnZBA+Y1UOVxFDDZy/p+erLVH0r9Of5KL7GPQDbdYJNT
CH6qqTxXaT6htEDUixpVy5TU5a0mzXRFSzGPRNSGPYFJ7RRTUJ+lc8i47YjzRL+Z3ZZEMlBEen8u
xljGGc3nctaWG9wXIz7qTXoTvLHI83oRA9PpbfDIk9kYBTJ49I7X0kFucY8YXygPV0Jkvl6/6fYk
pt4UnvzOQvz+a0TA0ri+HaqPR/r1mokN5YEGk1PjnTLGqPt3nsPuudYx+aJG5r7wHwWa/v/dbzbf
XZssQZK5LGR1A5uzGAb2+epXTMXzZFmI5eR/AcKWiaucItkH8Vz9Ks0FceGjxWpZoxGziA+64uhZ
nCQiYy4UINqFQ7UkfGJozL2dIoqYmbiXZNZO+EOxThtrT3eRR9Ci+j1v+jfDOcIMckCQBLPYVBou
L1sKqCLAB9GSK/cJPfbs50AmYyrom77s34tRt7ctruU4gobMnWeHbi/nELTPod8EfEYSGxQT2lpJ
YCuO8uuFn2nop5qft5WZUU3naRXo+j8Ejn99u1bsdoiZR8aMAgu3/1/GIMC8iBetqFOA08fhMNwO
SQUchkRvIKW/c7qVaQ148WfjVp6ztd9uaXjG4qGLnuHhadTSND510n5wC7LK2xMgo6PonUvSTmjQ
WS/inp7Jvd8yZmDsTqhGkocR6F2XH80PsJuUDFbqOQRw9CTQ0pgyRqVdFaA8cyq14rvar3xofVwT
2+ZXbcm7HH0TiiIwfKPJ8EpsvY2NafAc08DpFpVm1nFTrc3Mgsw4bkMAAC2eXT4Amkq2KEuD75FW
Rb/vbdx3lSCEzNOiCRrkdcr0FsiUyH1ofVyIDopoR5Oc7Da7RyOh+Xh15jf+us9Wdd4rTDEO7gaJ
pNpVWNqF7ksv7X7Na5tLkr1IzlI9Lrq6SVP6c3Ht3gvs8pMRSWUYRVcudHbnKWuYBgf5N1zvHq3v
uF1+fhRDXjS+pD9sMmTt+R8KyI7CknheL7lzC/m1K4GF0aF6b8VbP35mtQgUUFkztH+tqYy4jRLK
Rxrx9M5eSBKqSSlOLDUe7nFypanZnVC7GsJUJVypI7vbOezi2h4DSqrFqkNi1xI6Jrqm0HauRBMl
1BKuJRcvjnNNwZ9I87dUTB3gwqrDLCtj8e+rw5HKYqzlNo2UYPHm5Y2bN+TofGC0d4QU46d2mH5o
9L0wTv/xu+7asla8J4Nf9xT8cNfYPH/Md6P/QjP31QSEmCVWy2UA6K0nA7NtpVi9MzQvuHqP8Xjk
6RlikCIjkXR1fO34GG4+vldFg12sL9js7ZZEilOu0VLc1Jddo3zdXqDX3V5Gv0+d1dK6HB+B1WY9
wlx9eHIWXM4Ccm8zOZQYZrCFNrb80y6iOMFFpJ3Hq8Q9NETQ2+hZW4aTrLrC10hiiScrFPZCNNoj
4VE1dIludM8tJRle0CqCtfskZb9Gk79tsu1nOXpGPMQ8NAiQGNtPMu1tyB2FPztyopQFb2k06OkV
dPQ0TXwWiHAe7A0ERYFniFuZZWuX8ubJ2cG3zLKQD8vMmRM3UUJNmluu19LJEIFmFMvqItCY6P20
4xkWQrvobinq/OQthYCov8+XES7eQJY3ftdEG8Du0ABLjJnQhFZE55wb386Me+iVxycteoc5V7IY
xZ9OYTWnSkaf8DXJO5eifXQM08J6KBWG6Wy8Ku1cwQSSSE8AZ+HkOowxQQKLzXEgdIumIjVjl3gt
W6PsvvEBzQtW2nKqT7953q5cCSXT2HM+82YAYa1MKT4T8MTSFhdy+Aqg64Fsi8Rown2mZGdYBsLE
XHvvf97G6g9CUICDIM/Yfy57F7nxAsujaTesgx5ZUhmu0S+eHCS2BZLyZvTVefpG2RsR3Sc9icXr
I7C97VGwENK4Ip8ndXFCUo0Fqwt/TBgm3fM6P9cGxOMhLgUX6YAKE6ACO81AdeiucaWCr7wrNVNP
uLC1ie1d/5FTwvZVGHsA+aH+98VqTNZt0yNsnBvXCcjOsU2l8xJlFXKvGDtB23+ZjIIWrJA7F8Lp
cxAP9T4kew2fLgtcn9RFoazE+J2VCxcI1Kmyqb/oCOke70rLEe/6CGVo+Vls2P/jv/1OHcyiHGHI
kRj+R2MMK51JCAlVSmTX6u/H8qBMaInbe1H4zdRx50Vji7BiQWTxyME5nMOpamcqC+hGDJ5kdJHW
8hgaDzFifZQQ8epMMWJc34E2sC/f6q7RC+vY8+eXWD4+oWx5HSyTynwXaQBVeGbBbs4Z5RtMXoSL
3S5V/l61WTRyY2/bEdPloqaQMKigM6Lcy7n1oIhFBvYVW8FSHYAgiWmT3xnQ4UPE8afgCu7kbRfp
6dg6Aj2zgwkFhx6n1i9Z2CA//hdQm57gjEo9NkDsVYIrJ8utWPngsH+x25ITVaAOeFcyAQ4GcEry
dDq62hrav9mjdAg6XPqp3k/soEW0itAv7mZHv6fObtrzLaF1AIP96eKTvCwAAc6mVhAjevXbWMei
Z4Pga+vrPYsILcSsvj0OCJIred5hyZlhAhklWR8EVLhvKfHr0GVNZ85gxEZpDso0gG3AzI4wNHgm
23LBuujr2Qda5/uGpk+V82e06ByHX0OB3mEUti1b6o/ibeBw9UPzWpDBHmUCKg/Mq8SZa/Pn9+33
1iSgEWFsOH3dwBnwI3yZ/OFm0DJpz8mmP0xvc98mjMLA0trhvhsxm8CtNPE5O+IgkLQW/wJ+KrdB
0yXRoKWNjCT4TRQZ8LF0fv7gdr39Rp6sM71WZh56gXR7m5dsjbWRyS05qdeDc+Pc0PXfj8rSN2ur
nkQrZ7JUTIZ893jamNNjwm1InU/Wb/h3ZcVEBdR6UL9Dtv4rt7nQgc4YSc/cm0kQt1l+gIYgHuQi
adTEin/8fxJP8kDvsfsQT6FlT2xERvUSu1FlfX3FogHZxSmm1+QxlBB6BUizYKwtwFCC15w1oJBm
bF0CgkhLGaFC/vmzkXf8P5cbq+Xh83sebausjpHmAf0B63MdJtZ1fyMULWCQEPsnOLJhjuQIIfIb
A0HWnVUOJL9/crNjFULFThFyOrFN13OpH9d0qC5lQKy0iJ4x4HiBj58z/Tw3aYeoYjcY4r1Jx2rp
8cMjaSqGfYezlnd6whYgYOIrgU+mFaIX7mj3iXv4HohzSg88A8sx+/CFw30sw1rnpiSOYN+DGP3V
edS4B3sLKYSKcM9GsVwnbDnmyBc3tTAMjY5TC1ZnOuajgu49eAn4MZSu25VatxqQv0I/Ua9Jp+84
znSr2cbYX9FAe69ow9olTrq8f4yx04hAOPfYpSiTtprIephMRzMOH3PEK53fGqLh3JDoR8o+svnr
VkkuaqOOzrkIoe4UPWO7aT6652FZTYzs1YuX7+P1Tg9k5NSb+RVtmKFIT93iStliXJiw5i+UX/Pp
N8Tvochlr1IUrBtvDh1qvWPH7FCfU5dQvJjFRVljtXHfu+KVM3Z7HtlKfioXwTzXCSMJLtziygAM
1q+n0gRrDY/uOPCzUbB9izpwlwlh2iDcWVRbwgRkcWFhkg1l96+gBDHPyq1yd0KGlc/lee4oxDOP
f3R/l70iNpyrFbgW+F32fgLENA/dYJr/cblNXKVd04Jwr/1imo0DEsHtcheRSx5E47wRUXnTMSmN
DpJR+ylsM8QeXFm5SJCjxTaeY0mvaos5yrmsJPriwoN9aubKzZRyqjVCiaEIi6seeG2MZSG3QKlG
KcONaX0AEGe/66aD0g0KhB/RmVKg4EwWV62K4odowdD5hwMCfjMqa1BB1AUYUwoRbXBxGXm3TWUp
U0N8OYwg/1jC4dT7FAA7ge1fkpCAr9wAmDIBJ9J2yTCVGPa1/pCXqidpLoVrm61103cDa3tstTMA
WTNo//9QNXm1ZbnQLcWEo5kGrhBNy//enP8hP7++wVkBGXzlb9q7vhlZVXJr2JY+h26EpthCAt3y
xmeT241RFJOkbsvxlm5KaFmv3u5afugHRj6qcpIDoPgbl92PUeFijh2arWjE1NbcE2lNEDInBOlS
p/aefwWe03b3DrB/6/LOqenQHCKXcbGFVeTU2bkPtIg7f7vIsu4L9hKOPN72pvR7HxnGKDuTEdHf
zoZLa5g7UKCKPK1NvrEkgfdosA71ETr/FXgnmTgdLZ73D3aTS/yZVwSx51PO2sdzlu/6mDPjLK7a
MOpEQVVuWv4u3iunierrin0b+Ku4yjj7KjlDeCFUlJNPsegLgtQVrRdDggxfntKoj853iJE04c46
sfhVnRE9O0I+Jgq7z23xblcUOevHzQO8AJuU3YcvNYagfvg44n0e9Fe4TtnRvohBCkGvkbVfNfxU
PgOLx05NmZmk/pHNq3JBj3OjbS7zhJD1aDB8jyHvdnWx5hLULVdggaVOCgaKHT0vdEZ3uIQOLl10
SE6nG9flbBm5mfMuMXiyG7RHF75rAY3uuQpBwQU6KPkXHu56xvJguwltitzabmcEp5XMBgwBGYJ5
Y7xxC+T2mBEn/e8ReHV1+FdWJVI9GO/5/W2B5e1WxhbB+odnDgrrrJGi+I+lu4keSHu170lHGs2D
zbMcF/XWrcY6SjThqoJ/1DN9a0V3Lvcff4AyRB4XMqvAB2ryzlocQ3uFrxg5YuDaF2em0CsN7TWN
o7e5di6uVKdZt/S4oe9KMqjdt5a85iaDmxU76Pkma9MnizsvhHxjCEF6+8TPvybpW3r6JWew6tcx
lMzv+ltFkDz/ZOC+0DY9Q14Sp7+olMwYRLonYs7QcOiyIViLOSHH7PeLunBJVG7UcuUL8bH5weaW
/DAjc9G4UoQUc9Cg4mfv7IQfZbPhNOzZpw3O8ryJ22ghjPciyLK7LE2fikdCeHXuSJ5wwBxBI+XO
UeiAQLxa6txEfZnMILsgC0nOC7/ghGIMelk/Z7bzfF+BCkGfpg0SUNUSPmNimA/fE95Pjqu33zpD
DsneBJZwNWgk8cpxxX3ANRO8nS91oIQNbo5PQjxWghN5BqpyCvZe34PSflQpukx9duwcnvm9mOvP
x5oT0Wiqac3v+/2ptzFdl4ncmsAy3RLURXRTQup7al5syx9DgI9FZOWQHsPouqWTC0GQ24RF7OV0
I34AtATwbvnooysYrFJE4utmXG2Ec2xTxI3oqBoceIj8NAP+ikeyJXxG52pgSTGqWd+N0tBwSWWS
iqb9EprjXa34teahQ9jnu+bRWRKt/zgYKggOUFuYMm3OEcy6FKIeLHUVaXzzZxSiUHUqadga3NRa
MSR8Wy4LmH4rbFvwqSODgHRxQMG0vmpDLVZAoVHD2DTruq7qUJVlB/qbrp7J+2FwnJsjow6XJQk3
fcfzf6T7bNdhGle+N0QyEVABryBLG9dwaFxVOGTm4lKb2gTIr9hJ+wtoQf7rh8CRyfO+Vb6UDB9J
vghzxyYUYwOucz1f3K+R8KUIvI2zcoOhNUkPIomvs+APqAUuqx3owzpWSDO4D/EJsUjdUvBglTcg
rI852txBjsRg/ekMib86yZYo4Nc5GaVTjkXf+m1h7bjLZZM7nWp5gP3Qi/dVHQyZxKR7qChTDf+r
GAN+sLYN/rbqFtLWaUOUZp/uDFkySTITm90lqYgbIyP+WgsgJW/UiLApVsGTb0mEbSFNzE+K6Xh/
PYqH10w0TcPlh7VfuU9FN3gYvwpA8tzmXfrddw0J9eOCdnR5hAu/Pvt9yWpqikIhzlttu4hgCCxR
dKRtcBK2dPdz3og9K1zNRSCS3+wQ8sdxRMnmp0kQqSKuR8cKfvfppniSiUKsFzA2T/rKwIoU62d/
v+TELw6ofG4EhWMM9umWbBEq6KWfcnW+eokLM/JoF/6BEc/HCIis7M+sSe2tRWgynGRRkGICD2Ff
xfiQy+T5zVrm+VnUizog6ZX9n7+yygxjTOBFEy3Rr/daDKrxWjJ5EKHfoGHKpMJoKVEh6wDwIjD2
k5rhAFC4BV7J5X5ViriuBUz+H78KhAG5cuvPLlSC7lE/sjz1bZL0xxZSxiGxOKxHxE5+H4Z02R9C
OwmMaOznrnFgFoAvg83GdJB+3M5EBb8eGoRjuaykCcUJaLDfrtXeE6ELOZykNoy37A+muIF4nq/V
TxCO3d11kGsBiDN3u5oVuyZfhAaquU1BK33fmTP3yWcBhZ7iUxmxgc5DqqmTFRMonbRU4Nu9Jkom
LXCB79W6v3YYNZT/N7leSRoV6vDtTo0dS5QAfCjBLexg1ju1/vSKUtJlxrFOyYz1+f4u6HBeNbVy
hhEcbfAlGLVQXEtgapNhZcfeK1Ecr+MToCUuLumcHjEY8kPJEUomrPXycDivOlMi5rSJc07oUU0j
zx8Y85WGtICAFPghcNvhXnuv0nZFjombi45gvSHmTkihGrdWGtUp4sk0cNSMx2ShPQ9hpZhJ4/zq
6ZjIvmBU+l1MciUNpblDd3ks/QvGkQrxRS10ZRLr2SE0fZJjjpv9BAWX8j1ggt9qvzrf57Zn3a7j
ZHq4zInqfnYSWe9KN8oMxX8XtFsgD/qHizmFfEp1/uHTUiWJmcYjVBf0MKTKPa79/1THhzvyKNXH
vkkW91ElWXdvtp0dFlPCOCbVgyJR4dlDe+wuFruXMYRsPKP5uynMjK1TKn4KrSckfWNPB1db+uwh
UasiFXRdpOGc0Grc6xnT3PS2oG16NBPSfEp+sYC1trqVFDk1jYrEE98FqCEH0xjfbYpbBa5Ok3xC
Z7Ra74oIj7CMcD4w48JVHH74hlKf+nLefBmjuu7yRSoXns0JYlS5B8mVFvKYeks+ceLfSpZZW6RX
5vfJQ9hmZuZwmycDZneyRO9kcAcQHSTn0EDku8RQwyJGoDIN3xoPXpb31cd0weZQaPi76VMDsn1O
Ro9IMnDePzJy1NkRRTFuUO/wti4ikrE2ommKmEf+lFIPQnwj/BHqT3JH+gH/E0GY+jk0gwi0PvsK
4MYfJZZ5T5MriXRPSAJIU4CBX9GaW5LZVKk/sN+eZchcIEZMwAOSYtiboT4PCz01yGpwMFYmkTqb
Ak5XBpW2zywReNMraz3S/1BGpJv7UsTRvGFo+C+M2vRURpynSvwOYjx/5RpWP8M3rrjx4UX3YTC7
qGmeMMHhOcLNuEXXWlxq8rbMulGW3lAJwjf3K0R5xb687XlOn11nS6Nsz5o9hLCKQ/UbW4laYM/N
solFRgF6KGAp/HCkWARYuapybY1UUpuVqal1uzICSdTD4laDJeA797N2YjAqp2K+zeIl2TIepJap
0qmMHO5AgnF5VtwYczXDIcbgk4DkKn0k/b6O4Syub3AGLpmaKFB5X8y6T7dw8nhRFjsZRckJPFzl
hQg/P8BU8aJYEDqV7Mbh6NQ3iV7qciAQv4TeqKGmKAu0aPcepxMpCdcbvzJzrURfTmTcz5Kmouuk
vWTX9CRRFBoynGYc0IvyBJp5top6JzLssckiK7u0KhNFRIqHkQwRcbXosbzp6RKmxVvL5Tc3zl+3
4Ybf1A/Dy8XpAflSsTIOSpXQuJxcxxBkDgYSfx430GnsQMrTQIB4eOG7UFPl+JRgt1KYvegqY1nC
2bvpglt320rvpdruEz6hjfUGkJ1E1bR0yr6l9/GsYYUTHDZiYMlkpZJmvTnAkuLpJT2+K/8gdn3h
3/fN6s87dk2t01+XnC/v0pyOBHWjS9q8feYAZvZL0fsbNUX/0c/qofPQDEjxNjG4IcmUwsn5kwZ1
vn93nSTh57H2KSaE3uhYWvb5d+OXJrqBtZlO3kMVzWrbUqW/38Fd115FoB0Y6WaeBWgT3Gwz/Cmo
ud/Q2yjFFlYoGKl28ZilYaUlnp+xCTQswrMYtZG5mwiCLzgHdIjWpBZrDS+8N+Q4SL6FkC1NZ/lC
NfVGtJmfpE5a0mPtkSdWneAnm6w2T5zu45D9fQF5pWXPGZ54KETELiw2v4f74dib4uODeJ87pvxl
7y9eAOpwYKgnIctzLkzzteKnvYCiKflORxsA8ELfk5Us4As/Ojk6n3juhouE0dtd0qU6yioyp1ZD
Wrd2nzdgI7i7QyO+zJ7Y0jgDl0lvxU/lpZW3hQyeOmpxahxrVmyGr+UxGamHPPDcb48LXXVXi8Je
SK7/97hki4tETyJzD7DM/HL3i0vt5mNTotprHxAUqLOG3h5XvSUCl6uCleKg+3iiqxjslNHZ3n+b
nKKoseci/wQg1nLxr4ET00YKzDSF/pitO1UyewbHHl0hCRuInOnH1sboqF2zSb+O6kh5rYtP/8G7
jhHozvXZXgEOLdmSEkVOQttWR8COAEeuWFkRnNg3LAkvP7cYooES6ZeNxDF9c6nJxDfpSkC6C9XY
TQBCbX3o3LRM0Ct3cbBuOFfG60wNZSNmxwGTJf/llh9DFoehnO6t//PR0xES7mNfoLV01n7UT7Fb
iOhTG3adOf22sd2gaDttoAC8J2Xrx/7qGfSYbBF1QX28s47xzrHv4lwOQ1HIrhdkoLplUoWiI9L4
TgOxMfQfKumFuKNtzyQbuMlKY/j7W7Hlhq0YRQDSx6EVLKbFZLHsb5Lxdn5VG90lYis8agxHbWtK
12/8JqkSyKZCvbQSDyB9bPAT5tAYS30iO5X7SSKSS9f1v5RTSSAlfHaaAPGxIkqlFLKMx6UzrgCt
ZC7BbnVi5OCVsD6VKf4/hbpiq7+KH0mY+vgHwB7xFuK1QKqamYDfLTMBNQ9BhFiIDo/otZCLf0iI
CTCVDYKpm4bjp6cgn2fjtMm2kR6m3dYCvMzNgQRLc1kKmnj9leBT3o7kGQ+YbjXX40j0+ePt1ROB
3fD35VnasAcmW4YOyHrr9KDuSwX/IfJern/rkrgzvOYDLO2i7m0h1U4iU70MSUAunsML7k3Io1Nm
Bid49Ywqf8Tdo1c8Gpzx/MhikzKfidYic4sXVfIeF7tjvdUI/J6FMtsgNg7zrN1Fi0Sl+FmaR6bZ
G6AYPB4XUs1kChL4gv8MYSzSr074REdRAwvHhArOJPfqaohiunvo92H3FtZ0w4XlT9SOyAO+J8uO
gp2SxObSNz9yoddRnY/AAok3nQ4Tl7z90Pp0aEUZ10P0GK1Vfq+aUJVOOvCxqu9H8qg4Vc2Q7u/r
PwH8l3pwsBZN6Vf/XhpT/1jxOT0p5VvM0/q2XPwuiXJu3Xhk7Jif5/5/aoE8BXzhV+DNJ0ooYVD8
YyIn8CpJw/4NYz0YWEHQcK5GcEawelmGQzuZh/VBH3RiTEQBAsXF3xls+HA4t2HM8lMXJ2h0jFHg
45UegqYVaXV1wmddR7klWxjHVt1MSfUoP8oZRaz8Z0fUpKywOqzUixHtCW3IuDaj2E2/lnP51vDJ
Z3G87bZ8ZctFVl8mlBsOk+HuZiu0V6LYvYLt6zd1sF2QiU+VMh7jUMrQ9Fr4PbTckk+RjkWT+lm5
7vprNqmyu+i1Npv0l6zAhs98fSBkuVPFirzdbqte1iTVkEr4wd+K0MuZWHefTb/QQzNGSWOFUe4Q
WfuvVLvXbOs3FwmpVP4YU+R/Mt+ClkkWUekM6P1XCBmTXsW7Ycg3rhTKe66FCkERIpvmn6YoV/Yr
EB7ufNoI+2CP+lF14SIjat2HsGrN1aRA+XvAQ93XWF+BaCqXGTS9gcsujWHnpdCEE6kQVLnEViGn
zbaSe8eRYLX34wHWZOMQ62KGvzFj/Ms2g9lzjgaNCYIxx6ABENaJImIa0SXLFIoVJ8WFkZGUokeq
HA1MR0OYHZs6uGV9HGI6a0jtFALJKbuCi8i7Idz6msZW3grZYerjXgIs2NNongCTe/i0QzC96FhP
sEp+fQhf+VAdoLrxIyBQ4cKfAvW3vZ4F4AqtPxNXNGWm6fK1YrBruKRntZHf/wO/DfG9S03BvPK0
/nOPgoBgetCwQbEY+Lar8Lg1cDzeoSzGfBMq9/rPzv/oo9kjIaYXWyrC+jOJsYyAg9+HUWevdMDt
NxoQlCbMHMOdudMIuxCjZEwn/W28tldl4ymDgshwnC+7FA/oaEXFg+JU7J/zbvrIgb9Y2cWXv8O5
NZgbbNvqflKSQzAerJE5rf5pyIFxp9VCZDw//WJ7mpUL1apu3gh/JXJ7Sahtjqt75mrkP0MjBuaC
c36bv6SVO+QEttHRIDQAg44/jHim9Xb8UzhgrPbkazV1eX528rJrCe7Anoq3yPnn14LBAvYE1eE1
CbE1ec4UEJBsaMTen3nMaDX8iiz0tjAdCh+xX/TtArjXn+CGAiAw0AAmcYMK39VWwWgyD8qKiTxH
mE5i0YlMNM6FKMbYqXiqI7wjulsDCU18OxdaLAJdSWU0lb0qWLYNDdp7NVWPe5TseFdOD7ShZodb
QY+0bD1DSkb65jMtFQLKAGQpDeKuNlGM6mmuGAeBPAtE2ma3VsEQBG5IJyPKaO2T5AXuEu5yys74
GCw93MOtYCCh8G1p9I/5lRW8idosrB0cfb0sr28O1z4mKo2G9eoVhWs//dt+R9OS3taoYQ4EZFL0
g/psGkoY8MFGci5NWTn8ejQmViz+6ZmAPUZP+w1Qp7Bm7LA3CWKdCWFmZD5PbzwaQw+Tx/rZTP1f
WPHLLPcQYsFdM+Q26hFH1AiU9XKLIcF2lzmbdEAHQ2WuYti3d0Ten2f8+FuDg4WFt/gJF9032AP4
iSg8D2o8Fn9HUjCAUdw4b8NWKtDdxst6SFAMIe2Z1CKr1htCkGM8Qu9updCqTwX/JUqk/lVUSacO
3TkqshaneUGv/1zCI5tOAMhypQqJV9NVqzu7PjZdC8z3rfVulHTFf4pp+j+KyFlrO23vBEcUeJWN
jgAUvOyfAtgKJMixRlNSM50NvBszOncinHGarRkVpwlfa7B4gpGTjWZjmmR09tnLmQu204pu/6fC
n7xbKeMSgqDlK4gGgMZE96fN3SEtT6bG+DU7r+5vwoYo1jWyrhXdIjyPIc3gc1NcFYuqdKNB8dGL
VyluA74LmXsQYreupai2ejKjEae96AynJti8B+j/3dz8YrjimZblgK3DQoMVpddoiClZI0jwEPvi
ifl2PxNvzUyccZS0RCt1G8naSPssgdeASoKcIELGszBSLzGZT4jT68GZz20UcjMs/RBPX02kagTC
s24QALJ/s5jM6wFL/x2MbCTSuhxYCbVuy1yf21uKNJrXEXTCqPJXjlhP+Pg9S1ZvbwhWqhNzsdFA
BXLmAHO3B4tC2wv770L7gLWraROd3LAmPgLGeJn9E7wLaQpXQ9gIINkWZCXf5mARNyK03JHYAxVg
S36zKrak/7CHhczQjxXMt0NelOeGnjfEiFMX3uksh9N/U+Eo0BDIGTcSZ3+krjT7GW6mulFwmKmT
NTVL/TXNzzidEj/yD16zh3VV66qZdxK1TW0+eKTGW4DL3+7DNGRsd5hN+tHRqKoC/KaML4eQDb/0
/sjsJtXYrIYNNEtQN6MLv4OUlynSCXJzuM89PqzhVu4rncqtHORko1zXipKMkcncVa5UjNxaqpM0
oXUC65acHqm8ArlS3z+cIWHyrqIKamErWDQ7y+uIn4v0PpNmICLJRLpTdV2kJAu5jiuyPCo0d85E
5Y2+wD38r1wY4uE7lXPvQlWjevH/wvAxA0A0yP5WMfaDb4cRwVNoM5kwTzHFv84wKEYSPcFMl7Bv
UVzVizQW5ZvlCZW5MGtToDN283hTZgCR/y7lY5cQ79/MPyFVfRTtDCxpcU4gLelYGozfpC8PKOdp
ScBDHnWpQbgKU8bu7y2juCKZxCMJdFRSf/8FwzIr2DLxwYukdXB4/xCGGRqBNEBbHp2sMCKY51lu
jkyyHI6w/qjFFowPulPfeBBgrLo+hjLB1Q+3Sdw9r2gNo3Iy+xLzz+UcabPbvaKOl2kW7pq8NSyx
/G9mwEGltgKNTtB+65tJD4m7hocf8i/3vZH1kQyeiif47mb2fRiCRPXouoaKp3b+zlKy3cxBQB+z
zxZPrf1MR0lvIDG1XGUQzaOLIV7B//jCUol/By0j5xs1SKMm0G/i9/XkCY5TZe3oqgVVAX03GiZP
RbP3ZTMmvsswMHLRtYnHZsl6IQB3cAjjnztgeQa1BYATE+rOIRufdkhM5QuUDlvi+P0aMhoEcpQ/
61LrWlw6FgIcaDIvyOlarfRl4/L25qRAZ7J5g4k5PcQBvhmKWVrhvY7CeHgQ2WUlrL7DUdqlkN93
OpxFF47Ioia7FrHAlSCZVMh4FkudxO5qgoObfro0XX2SELYCHF7C7YE/RXA7MAdv+Mg6pyb3Yo4T
DqbTkoGbEZXIglsT2R4cTIk0yHaHtG2/LEHCW2OpAtp70vjHNy8r4KENahBdFF37Pa3G1QAJ6krx
gt02CFF0mfErz90jILk7NjZulFzkV8IFvx82OAxQjVupBTc3rpEbNwQbJbowLjB+RWZm1SLI+iIk
xO8tmNGKZo3+sndiFY85bVuw54trF61t2oha8NaPKsPv3Du8ETpsD36gUgTn6X3qHT3mVezmVcLP
ghUCv/0bihyqWXouDlgQUjDG9VTeXY1PMOBwqBnaG0M0uqnfmcIgEH7HHO7m25jGtKVsMFFyuvJo
+ibkdkZFaD6YOoWglvjufjB2T07xH2w2czfsKKkMPt/pqFTQDIwZ9OJq5mXqUGF81EjlynJ6SaVu
j66eqdODi4hh+4xNn1bAVEGQuYob7Zi3I/xCYso6C96yWBF7dFNEXtVvVSfsTSIsVpxJILudFsO7
jMCKAUf+LQzFYhU5+y55rc7Z4skwr9gkWdtlZoQ200YJJu8AblsTl9vI6ZorfDMuUA8+jm5Y3Dye
loDlCnp9fN/pR2GmDs+/pdPStcKnZ+nzT9GOoJJwUGy4nX3Z+K7aABYdR/kJ2babGC5osQpBdnY7
w0JfD9/uB6Xr3CvmxjfhSPb/Dn8gLDhpO+5laikzoRY7U3IwyXe4qL/FzCiPtbh28HwNxaxhDnq9
nZnpODCGMi3o2CzcVKC1q+0G1261nr6zzof+16OJFuVIw8lGx7sYAvwLgPTU3QO0KvSnxTeAWz2I
iH9al/5slu/3Bjuat/wZKfoQd96wV498o3LB0VJCCoyNvY9ah11nGXJHPV5sAbZkuT+CsS0simhU
DlNB/EtJxITgT1yJ4NMi9Ffx7/P6GWFk9X+mGcV9DzWTWXoc2KD2P5sOXVkkOf63OELCG0XGx9/S
VYtPx5NfAcZbghuDzr3ITqzmW3N6OacfgIv+O9ldBtvA51pjT+4zybYJDclmmcs+siIkjSGd1EJ9
5MmUVIIY6Bh4HDXqvIvdD0loZ8KTGeerYnowrluQFa4JjibIDnn+jPHsYeu4pnzqnN3HauAGiJFh
MRVHNa7BwqaAhoaCNkSVJIXaj1DO8VPgmb6AXaf2wMA8k113b0RvvUn6uS9V0bMUzGYDLP5lvfAK
ICA/qeG3Zc0EOAw+mni7DQYwgPSOl6piHyCf4zQ4AtL+g7fdnrngnfm1FqoBNEmRq8jTcAvN0S/J
kW7/npmJxwcgTo0xhDR8N8qDSXdiX1N9Dml84xEZDbOI9rLWucYBplfCFO9e8g3zCIzj+kLnxrNa
3MgSoep0x+TPdX1lyLQSUf903wEYJEf4sKUA9mSHtIyGncamZUxngIHK6HWtIgf3F+la+FDuk15q
p5B+EYXAil+W2dsSZvDaBJahYFXqM60CeLAUKQdAAvBtR7AiXJEefPday+ED+uYlEVSER7hAomCx
uue7+cQlxiwKuADMXEWPBcdHuPGJUb2Cd98cfCR21Pv+C4MhqErXRpj9rH2rWqtA9L692lDJj92A
9zKnY+TxCI2n2rjKDBe6Zy89xnURD/3FPQqo56oQg6VwWI+kDL3416IyPRQdfF2B69JqmieX+1W+
JjCGCcf703s1Rg5dkC3n1lKDDfjWz33XexEMCat4yyL6wO1p0/4uRr1DTE98wvADjaAcfQrfcr5c
KsoP7VDyDY+bmR+5YvYJ3rQ4Ay2bbzGzMgUuO0Y9aRDlLYHylfb0H5IMccAvlka/mJm8GOjtz0f0
xrV4N+WGdnYrVRJodhvZTVvqzG4FFxxt8i+FZj26GPz1xQEK6kQbTo0GZV/rQByzkWcoXRI7IhwG
Dxn3naTotWjQQqo+Z8anRPQYhXDYcGFv30W2tGPDACyL/T/nsqjU+w4E9UqmyYb8UPTkQc/Elylr
7pFne8me2a5h13lafu0VhBGpSe5bqw9G2W2kPqiMQST2mVB8uqpg3fcYIeIssk+tOhadqgOXuEym
vlcQSgQsTBbArXQ1IvzrMl4TDV/OB61TCTQMTaK2c5gDh94q7Kkvky9QNL2UX4msrN251joUiz7v
heZd7Wp2bJIYH/iK1mbzj0iLPcsedUuTm5XWv7KZm3OwO6Ys/gxJxJqlF+j500RULdr2OY1mCCvu
nKLf1MeAwMV2oks+nyfCUNLXKJ7A5ax8ic7FwIMoiyAvaLmLstzdDznw5ssjDKaUo2nVqpkj57xT
+xNZw+aEyaZIyydPGEieJHFflrOYWQfTWLGmIxwS9f17NVW+/y8M8TumonwvreDEuttY9CeOf4Cq
Kf8GRXihbQNIyVb56cWOo4l6DNnU6pp2R2hxux83iYVAWPISnLQoJ8OxvmJY4iXhho90o+K6t9Jh
fUq44JQO950JpWtRFZlnlbTNgIgUgTbNfRpnsgEYUepYZxnIXiArceP6fHudcLHJ3sIWz9yZLjzG
XFSXQwhWCHpc8/M+C+AM7gpv5T1al94VSDZLjmsUpx2lytFW64lX7MGa3I5+RLABcbwm+A6N9dkd
sNORf2AhL6buEe3BWuNV8DbwwohoxcDQIuGURtWcSOXOgb+u7S25PeDvby2yAYDEoMN6Dg+h27Gr
Euw8kSgeZYrMq0zriW6JqM0mVHRMKKSTXMiSSVyDm7pQMWjN6rmAP1+shrwSHjQmcYcLhwQtDmd6
xHqMV9ascannUFKp+V64BTPpn5o1F8W2gxVNlInda8UDvFISQtwjg7Nli1Ax0pd4c45ML3UMQlkL
t/8I+dG3YlbVq4u9sw6MhL/DCSO/pqDEphPC/8oy/AFujcjzhuddUH7rHKNZD9XEtQL3GhIr0Nii
R/JMYEvf0tED2cD59oYz2IrD+uvP1QYgiAAiwx6SnmN3njvbMw5+ZtIpkqrK4FSAOtkyzRspeJ9r
kynT8M7xAdM9Zj4VA+ItJ3Id+KJzWt1Y4tSnXNwK2iiFO6Scpyl2NvQkhKVzGyX7kBm004P5f7e4
n3f2izsAuQHjZxYBYqHdgsxZUIKgeIkGI2GhS1qpiNY4q0H0YZobtgOQ6qq02CH9R/Ee5d3xaty9
H+0K4uEc+3LpZTdR6arLVLa8QYAlDqz3Be/yyteC3qD9FM86hGvwfwSsCaguRPD9lyT3l1HLwoD0
918E8uNWSzDNvMU4zI0rhilMCRd/X9CFwu/fAAMWBlBSwsZjYTja5myly/P7bD2fIwUJfZ0ewc0x
IaPuyQmuYaiyNDM0cds0e6x1LfYTWoHUDDEA3Zg+uyLcR35a5xlbDTFNDSxsaBo9xKiWoomGEi29
izaPWe9F05lWhfNRJZ3H4Np1quGdJtnY6g46jmn1JX/6wS5nldmRkyfYpBVlAVhvu2JggoHi1snL
ouUYfT2nWSXJYiZvf/2JnqHu0x71y/ZzYristyunlUTI0Y76mTOdFr9c49upZB21mICUdSEZQ8Q1
2OLljMv5gZU5Bk9WxgMu6+kt/RDr05VvvpNhSLc5RQ8Pz4yfMXaByh/iDDNl33nc0cDs22wx7Ns5
0G4u/uIcJZLY2bXHFSBKjqA1R3Ep+3gZqc6gY4W5C004Qw+veF6kwwb3Eks908fSIMSoDv8EVc+l
A5iM5yXGsKTh+tjx4CBkddwFh+4M1csPuFr5+DmGJKfr7pLQhmT+nymwy5aWJC3Dbx0XovixhKsx
IcdDtJ738NUyu5cKYsEvvRtvxGwTYgF7gE2tirqA1qcPuLnYmIyEp1D09IsTbA9T2DDmzKJz+QRS
KLKYFA6VwuGkFde2L7XpP6cdGYSI29How01HvNjJVjCRlsEalc+bcG2WsW2cNeWXxq30vLxilKr6
Gxsr9YWDjCdo8IvJIcVyh/oRgc+UASKxPvukGmfJNi7zVu/w0JEHgOw7ryyqdaceXx4YbQQpFq50
yQo3blQ/ryQvOZt/5WuQm+3ukgLTb5SKPUQlG2DsWTVwZ+lz3JIy8kLmHNcG2vhxdOLUfqgL4z9W
BhPwGEZNwBT6bLNtHMtcgoBkmHJG2dtDv0WhqGz0kbYcYsjY6xg7kvaiP7HYfNtMg9trOiFDCqKf
gYsrbvdDyn7C6VAp1zS2GzcngiBScelAr3l2Jt6OLgpercALJFE+TqJmwrLx6gQYqGnLNGAK9Eai
iKNAATC7KXU4ilu9SD8wVYSYVHPhtD4a2W7LQTOclfu8kpDqpdvAN83XD2JKkjB3Inrhexkl93Rh
V/uykNyEN0XhsbDFLsg36oDN0PwKc3ztqMd9nrmVyFG+DR7H5I/7N/K7WKbeLCkIsUOgJbS8H7cL
P8pyt2eyjJ1Nou0R/mlm9B425TFBW+7yGnwy+4EIWKMOLvnfQcTV1h3WPSObi3tv/N59UhAKM7Nu
CLtIUP6a7z5m2XK2dvxBvwhMiZrPmXZmaAKcxTY5PkY1u5Zey0VaY7Bc5VOC1V9snw+2xfQ2ESQy
PbXUOj7dtgtwatYL+LaafjqF20ol2rkHR7DPmQb6wB45cKSF34XPNg+EjMGz6q+FpraBrqcKQq9G
LSR/3GKI3a1jNuaCl/V8JJVnUuD3CMYYUGga8agyrYy0BZ/Wl1D2++p0LVcnPFt+P4xBPLK6OMO+
+C7MWSFlaTQssOgJLyeBxp/l2SlqNU18kiHp/u4i6bHrJa/xqgMhdUEKH2kD2ra6CHS7nzcOLnfF
2LQENgHN/Tij9Ot+zBydGLTh2I0g52oO+8AP4aBrGX9miCgaZtc/9w73xtZ24qhgNw5aLPWoUmG+
wV+wlhOJXvL0fltHzZPt1dTeYPPao7UZhzLny/8wqjdmLDY8il+MJV1csmyKofhtZS00JhfWQzgh
M+NdkI02kw9js+xDfGIR6cR0M+E2Fq0pDmHCZaJdEQegxcag3UQQDTH1qoc1WOeNHVDMWifqaJdF
wQXnBWsAROBGoEcwz1KlgXnhKAhUyJxH9kbLE9EO6BmbnQbIHlRESJUbCpH5Jb+EUM6dK2luJ1g5
ZI7Mcf8R/3RGwDWFjdDhFnchNY51emVdwODAl/Po/l+eQCZSdbh3XORz+L7ke9RPwlr07CQ5ODYN
b86GLfOVohQNciW4r3T3fSxuVggwz1pbLZfBueBHS5JsU7NSKm48EUQkj686F5aj8sBo9rw02NLb
hDA27BfB7pjy+SqeIjFUxwD5wAx6fq1nH6V8W0YkhuJQvjyaS9f7xP3NvNvlQuYvLe5fyhqW1+Xl
bNyWjnnlmGaTrpLz/te4bajoeOD4VuDOn2bdIdXGF83P1ODf3YNI+yevEXyxnmgLxTeSB7bAWrwx
t2bxmXbUCFbDl31AjTYDEPhldK1JFccfQ59hMTMVx9yPEAMtq0T4OzhJIGff8RP1mfvNXXJki/7L
XmEvzVnU8mzmxyHtPlNww8F+VEvM10+lsW5ZrXe0XTrC5dTM3gGcgfH3ChSVdjj6moo15/9AR8UK
5TNi/ngJ66yLbzqhZe5V3b7B8UWS+6fyLDgTK4bo32P3sSE+taVy4B5jvSZA9Lais6GfmHhBvrYY
81s4cP+UAvO0vANPG87mMHHy4UtJn5ifcZABRQMTzXZTVp3xIR4lWjf5YEIa4ttcsWuFIn+1Yfx2
qcEXxk+OOP6ey0C4FI76ZQxdNw+GKD0+fakmwFa5IbR1QYOKP9mIsgx3/G5gW9TXPyjJ1nhHVNkJ
ZMHTdcV/c+kjvPkIk0NOtPOfhVa//eGORqVVlnfpnGVwvnxL3jv4njw5iQ3F6oMcQ6nduPT7xLL3
gCOBkgudv+V2Eno4nagc/x9hGfaDY4hj/ts5YS0MyTMe4BdxK5rDbDi6Bm4TBJe792MzMYpTpPNS
Y6cqhGsFQMXkExMBOcVk9tNOrKs9fbL4ynIpremRytAoXNZXILHh5Ivuu1+N619J/re5AJEW477o
m89m/OFDtDCQ2KHhqdE71P3W6R2MVr7FaMw2Wh+gG7t7l9HlikRnDg1sFOvF+TAdyc3nM0hhZ9uY
v39uP3faSPSLGzAvZIa9ilVcACbC9PYm+zyOKQChV8b6iqHx/4W7eEyU2ymWYIdXWrZkOhsd73zB
afKajQnDdrZijYQoqQ8WvMkbqMO+vi902AWD7m6Pxo7e3Ak1U0c9Py2bl/lxMgFTU6aCJSJtgxYo
fct7MtxPbOjEbE9Xzopm68Ems8dy74EIte/Z5aPbi1K6gOxhIhuZ9yQt9fExlDVyTY8i00N08mt6
qc0g9puC0wcT6gBTgExAGIsQiPi0LENyEJ2DWM5uvq8uu951Zooc1VGOl+SEnb/gIFkF2JAVKQ+1
Ezziba9Bgr7kRvMvuFx0NUpGxLHjZdMgOZM1V29HeG1UA20woKXkNEhw7NgPHbctlW2o/vXnKTk1
tgDzzXfOJdAl0MNK0WTriQwIAiIApJ/H1ByrrgV/xlnBoroKr9/JV2CTZ8GUqZm3z/miGIcaZTW6
yYjEGxtIchnNpvwh8OoGW0nV8TciWLppv4q+FWuh2PGu7tiFMX1Tdi5m9OA9ZaPS2jzcwyd0NL9t
CHR8x+15cKoFu+/82PrYX0XTTr4pob4Y3cuSjkLGN+/xAlQfLvr+Vm9AewA+owGL0/rXYWvRhCVS
Nm6Jc8knUw3IM1JoekMIl/93CqbgY8t7VViOLI3cXGnPCaPrmhB+2xy6z6ayVn6/3B8Q6p5qJQhT
GgE6u+3kDrUIsulArq5HZQS+gDcJ4AhKunTp6IL72zuzQ6PhFG36wAHYswMqs19PEWUk6cYVCDvg
2uW7L9BVDAwySF4KEPdtDADXHduTSasDhm53KxQ2qxRw3Y26c3B/FmtQhtdAY71jarrPKxAgzX0S
69mgKYXvQrfnMY/ts4RVPF/E8ItoDY+83AGtkv9F6+TTu7CkrhBYYDBo2F+eLXBOHyLU+Ijed/X4
NC+6TKvsvjiCHJaNmKqKQdfPYnvOCJy7xSVD/fCQu8bhd+4RSMkODO0v5tcdf3z93vjLLGfeE2QD
FnBqE0Eq41TSgtmsuuWbiJRiRKJCIX52ATDKj1zIC4RlfZpvMj8zfaEr2Rmg6fbHV9mw9kTr9R5t
U0KnZdiqNTf615ha3B8yCKcS+MKSRC73jptNL89/zuv8Qs46VKTTeYB6FJK56Jl+h6NCa0etRUtD
DizoOfEYANYE/qELb6cRwdJF0HVm5l7yBpIN58YGQxqvnduyycgufnXNbFgRv67pNQMcTRDnXkrh
q+bXYxScxKyfBI7aExEVeZFBhLkyBWFHCmAgxVuTcLXbXmcbPD+/j0/gph2qDVY9jHpIDLRwkOsR
P9b5oLmOO7QOjPNn+a0sk0efmsxVORQj78WP1NCVw+eytrJrsTprDIZNU4aBTFWLEePCRmoMLFV1
nwfL2Q+Jdxz/pHHUCQmfEBkSUob5tUcr4/XQFHvS6MFAHFKvFdd2IC/DxMpWFvpEchrtT9r9TqwX
fT/+An9xWgLIGmMgzpl6HVvphS5seajqOPBX8SYFLjtm91v6KJcNsM5XH4az8JFFUtes9ub1UHoC
K9FVx3t2j/1j8BoY4AnILYM2zt1xd/316ZozndA7N3Q9axsuN/heHa9GOnfLVWfECIkVv+0ijLjd
+EROh+UmJg05NlQ83TDpWVol1gmnkKOZK5CpV2rl8KRT6OCMdZ9P9UhmF2pzoI1KgpuTlaOpijrJ
m9BW39QfDjT0J7e4yKiJZqNghCNYFAexow0IaCf18uoRf97qPjF6p3z4sq+cyMEmrGrrUHAolHAj
1rja1gt49LQfp3vvSZuyYstN3JRqo0mc63t4iZ3fZ07qER1l661oBYWJ20tKANx20UnwnFFtq7jP
yJzUPbL8iKlvKae/7Iob2k5jAV7/kKwxIQ4/lmAkQ7mW/stWu7+ZiFXrkwMNv6HJmD2DeUz7pUR0
r640I6BOQhim7mODIftiSrzGd7DeGs/Ou9Krzclz5B81x1E6M5omTiez/8uDnRWOY5r066aEpZEI
YPo1shyiBRg42L3OCOfG4PLcq/cNOci90b8rZASMijpEOqJb+7pOCqOgEC9rrdVPMu63YRGrfsh5
pNREgaWFr/+8N7lyvUPazDNf3STu3toleEzVLFjOj8iiKiqAllJKU5wYkktYsN78hBkd2m7/9/3o
FnLvYBOdqLjQFwjjJmg/vjfqzHaihumdsa6zQXQadUjp1xvYPdn4lLSrA4Rh7xhU8H9JDoTyZFVa
MqFwUbdMkPvRjdm5Jr235Z8nl3gYd/JMZver6L7lyrMK1uwyovM1iry48WUsFedHtd526Ep7brk9
4H9K/TJ/0jSKDlbgKNZTgShdpvlyqtJbKdVtIp9K2ommItdSgHZvsjp3UB0fRaLQaYygFb45rBhE
TTSyHBukyJDIBTHMwPmnR+PFz2eJtZM5oYvH95oEhpDmfWhnYMfbZuISBLRPzugCxWKXy4v/Xqhw
+0B/L10ZNpxfK9n+ggJPxrs14SpBY0QPlxdf8eIxI484jASQmnDTrsT76QQLLLfoRtiSAoQ/bhpl
ur2kIxZS8ye5JKRSzHDwtPRS1jEL64Hiedtly96iZo37VAZqj3MEvEHSkE6EJhhuH9OFCtaAaz/7
9qyadRN7cSLMS5pMqtFnqVeX8Ypnv3quQnOfrI64SfiUyd7VXWBcV9AloEpFOXgCPFZwXGa++VgT
XQ9K/b5Ko7nE4Offd3V2AoEhSe6mUuZ1W3ss07HnsFZ3cn5qc1WOk+r7UWnCgkmumQ7byQqhfYYK
mBpjZG6TsYdSzKiTxnOla54BeeXnBkHx7Rp8shBV8tMRW+nRXs5yIiUcc8NhC3nnUqm7kkjSqrtf
45T7osf8849exM6IC9fKyhPHm2C40rpUD6eFlXDpR6Ukbu8coIeSNfrXWKEMcGYQWhmjpLx7o0Kp
zNRPxw7WDSIX/2jXLV5KBlTM59AAIEKxEuEW6wvBwufuh24+mDhWUqLXcDriZhiCcLNx1pKkweqU
G2XUOrnH8bviQImQ2winH6of3KxbSsdeuh4XPv6lQUmd3YNeBTVklTisKueluAnUkiRCyMEQNTV/
Y2rqCiFLGfw2kySXWjY4WDXcyZXeXP/CnwwzZqb+VTpqPZF7V+a6BP+CWpz2QHuTLDRjmVk5+C4F
k+lrwify/Qsd9dNPV5R+GCZ31QDzCMYkCtRhgoON055chcaHyfB50aQaivpjarVV8h+9f2gxlBQy
NWq6XT0lnBWu/e1n4+MJ+3TBL0aUeOtmZoga8rUY5QlE3e946AtdsjWxKRE27dlGYYfdno/Jh8uL
iWW5hLUeMoIK+f3ZnrEVxEInEBNZ8/56OjJGTr77vDkNVmyipnCwyfP/YfjBtoFCJnTuE4pbOafj
rHlXTuU6BLVEF/oXFSj5RHI5f93Mp5Egc/w7nvc+wry8JWhc7KGRFl2sC08SK81lFX/D1jUatdaH
83D/GtHWbrUyTBi1tWNac49w++EKqbcfBb8ZyG8YJptTb4NTGzMIE/puuSYbqDcUxBfH+G1QW5f0
yUYUoUfaigAEc5Rxf85gzZQcuW3hzkNSijIHnOPUiFJnP5XW7ok8u4oG0+LtW0UO0gCqMpi5jasX
AfMas2R9lh8f01F0/la9aiexiBZmgHOF2ORJR0iEgyOnfF6PiQiVCKOul1sqmZRIFl6ESk8kUTCP
MXr5bxDOjVd7yzAfzxJgjDQzTUAP4lboj7BfIKQuQGmAH345c/zzkseSWHyy0ekfEEHeVu6iQoTc
wgNq+KK+kRZD154Byi7eZJ3TQaqFc8rSC5zdWE/01NXnDfOydY/UDIgR3FImmgIC9+FKihpsLOHR
RyIezU2g90cHXCR/cnD9M6OsYHi2FwRryZ0PhEtHTD0RC1FWlCS6O9aQho7o6b3LdassHJXPf7Lp
o+rFK3Hy2AxTXShFTS4KnyNvbjwtu2+VEUDjYH2RyCuI6ev66GOWJFLJtfN/dT05jEXx2UAmpnPV
oWbzjgw13SDCtJSRLb++JlHAhs3FLNoNtTe+V3/7s7hC+RZfBd8p8r1X+36UgoIWHBHb6oprI2DE
trOeG/F18tYy+V9KFGJKnaQJE8bsFn6FHu3++7zoqDmcqsqY6r8+fP5D4WkVyQHa3+rW4dVV2ua5
DMljnWDIzezDOqjqomSmKJmaOCKdHJUGxXUOk1JckVdrfatCSR3UsK7Eq6/0/XrKedXalcVY9y2V
3Y8jFzfsYC+JhEmI5ejbJADOYnlUyBPd54CvB9VNhnXr6C26M8bhhRABx4A1PYAW3w/Bl2PKVVDR
i091jKHanevMJQgpJve2S0bS+VaeZV1HsVcyHz2gJI3ICCaAB0lPce8HISbYwPZplx+eSwOrfz94
G3kLYNgxPQCp8pxry9j61BSf0AgiCbTSYlrho24OgR9tzCU76R+TpauHgrsw4zbDTspQ+CDWlmyV
bkUluB8l+Eu4XROFQh8EygMI7ZiYsp27vz6AS8TKKnzGZ/zQNFqMo+TPk+xCspdUrAGHt3/ji3vT
lNgLIVRRZCPz+YKs9myVwv7v7ahEV0CPlag+lfvDastfRu3FN3YApxmS5DigmiQbSpI/6I7aGZrh
ex2B8CYL6A/h17AihXNEag2mxv/LmuZWwKSdlG5KliUzG/WFsx7fSoYxW9YcgJulvt2JE2YRm1TQ
Ogq9xtgRXs3BISb30VHfJnjuaYrVeLQ1y85ehs4xhE9E8RmZx7Tvn3nLF7t4sQcgKyg0XCbIqVID
H5fj9sJEdiISh1z/hx/mA1cRYli1evRTHTm7nGzDqvxg8e2y+l0kcMe6OjBi3W80l0V68XUrnYIP
XCnB87AkxEAta/uc1s2+E3LX+YmVNgp49eZk24RN15mTPQCx33/RY1cGBStsI3K0A7GdDRzKR6au
qs5AfHH0vKqR6qBRMspeFx2KQxYG4qOMK+oRp3DpV7eT8VVyyqjkK64Kol0E7qYoBXX6+vgGAUt5
RiNBfeN2v/Fe9yKr2dkoa+m+dSitK3nyUVGkFMgZFsX1g/lTfWvKDlwhDdAMwkuIWDVIKPn1vIiX
i4c0uJqcgHoUiC/YgDpV0zK2Ju2zxP9TJ649VYEK+2bpLHt4UsYgos2R6U0b93RFvELPnckXPmQA
fs3NKX2HSOMxEBN828ivn+S0cF7GCGYFyB38CXKul6UdjnzcgjT65gww+3fQcWIq/ckrEaQ/9edx
JCu8XAUE0oJ1gTZA6Vd6kYO4AAPG8TXh9/oDVuEnkp8WFqqxHWmhmIs3UOQQpi5aCRA/gNKu45F2
f2v34X8HKwLkyk7brautCKVRjq2Uhi86SYH1GUV8Kj4zEqzxMCHmJr6GcJM+3BSFbJIJoQOWVPmx
JxYuUjff+cZdRZGYM8XyYD7V5K/H8JDmkr/ayLBDNA16tPjbaRwCiiYPZI7YIyv7jt4DshSgqpT3
UAOABrwBpMUO5SLhrbNWPO89uUd5p9YAtFm+/DbWA2gXW7ZgNszAS2ANr9Meoeq4pxIH1HhKBNcq
oIETnkkP32uBZq8E9JTj5x1Yxq7d22s3DyvwPbAxFNNJon8ArZjU9c3h2McPM+hIG4W+g6InKs2/
nwKCa4x3nmugD7DfXbQp99slRbvYxTVzcuZyRgCvj+kCdJyYYsWz64ZwIGYO/AcC5oPZ/wvOgpr+
xLoKjz3U5RaItxaD5xjfJDwFu42ue/SL6SfFrvvv5t2MFnQIHXa+E1M/HONTSM+9HGtYkyAtViTl
ql925mqSVJOpsQziRvMrOBi+UG6YvFZtFWBzv7gvc/EW5zHagDxCsdSrIzeubv8ZIvBiC7z6kQjp
ljz+NyiooPInnn38FqqEpl18OV/yM2nqLl5tBQfNSpNGBgSUm1beMB1UAnM/JJJE9j+1rBSFxCqG
wSZBizmQxJkpcztLUcHeElgZELGZRPEEkci/+0MKiN3gS8o9zBoIxAJtQlZiXFdzWOGzbA9PC1AY
zjIVT8qk9ydl5iSgtwzwyfkNSVXbGjEQUpMJUUrpucUiu8ZDkyhn7huenO3DSGQ5Euk4kjQXtpn3
vcPTdy5kaEMyK87taQ8oTsSWix2WfHkgKgcOZ2g2Bf6/j03wrATdzUXowVIgONDERWXPiza9LXqP
tMVyvkWlJDu2J8q/6772PkSBkMYPniccU4ukFb+/S1r5a19iNB4vP0wG2YHN+Rabk8YosDZcQ9eq
uFdweitltwNROP3SdTl6m35P1y7qgW1qONe8CFduLcwjboCGJ5+bgSlVdjf/qtUUCepACY0sZIQC
g+1YP/CatNWqP51OVSRpT/vYSh2m91JnSX4MCUEu/Z4nF2KxbElTsgyWpSFzS58DbD76050qCrFv
8zFFu/HKFHrS3vbDCBegHKq35m98uXDxjbdEzpMGoECPvNFry1EuBXoF0IKZ/hGl+89UzejaYYj2
PYiWZo9Hy1rD0BMr/zBhL9H3r4KtP+j4y/2eZPRaPtUmkC59KvyOzpaWlu+31McoeeYHPOdSlBvn
9+52aBFREcTxDQ/KoSlIxweEq7EdqTfNnMkkJXxH5vkPQcK/Nf5REEfTtjnA2XfYX94Efmtukse4
WiuD0qaZjoUfC0aC0JMcFbU7F422MEz1zPnu44kIl7kETGhkFcDfFNh3I2N/KHvLUGbmJ5SczRZu
LUeZyMiThtjtlBMKUTHabblwLZjpRmJuWorWcxOdYngIqlb4BluCdUU8A5UBWq2ivk1cxx7Q1hgJ
RkgyGX2lFqnYBVLNq1v3a9rVrypDaAC8A2EcDOgnkjdAx+3Rfw4OVQZWO5G2s9dxBEOb4aao8UJ9
cNgcdoQ8ItmdQg8Z+MZw9F2lgjaTv7ST3rMOeW4wJXE+nj/VknfPKgOAD/Ygjb7Q0d42hYLTslbr
IkUxg9jtte9pvF286adre4BrVhxJlYsXxWtSphSxaNUydUwug0lrdLgV/LvRGRwkYd6RDlPhtnQd
LjY+smGmqTgQcrzDD6ln/M6jogxi0klTloH9AGPqJDGN+bjRII2wRPO1XpvcBIjNg05xX0wLQRkM
550f8RgI6h3JAxRMOqJE1MmkO4K5W3nUSJvNeBRRrrwzio67QRJqx0Z7wLBvldyp7ikqK6354hne
rivRUmDvdt0o5K2PZkqggaF0BD15W/JBGsMkHabEOgJEXQ4cq018adWgLArRoJrxn4syVSLqB0b1
lDWzV1Ic//wsrNSVw2+E5BqQjHpzhryp5iIhfNYTB1qDPqzWWlJSbbEStWl8ytsD2vmzAWaaMZKU
1Y15qgqDxjxrt3cvt1SzvLlIMUJnJlPYBHQTlzWpSkdlBDdVHHpN39dVVTKIsNhz0QR80RSVv+51
9LfMt67mlkDz8P648I8yw+Q4/Hbf9A7DURHg3rklQtuFy056Sw7CZXVtGyFp7E1M6NcGldPVfwYs
v7M7j/HQS4iW/7vOwd35L9H4VLcF79dzgA0xytcSHYGJiHN9G1863eB++SMbOeIS9Wl9/vzXkVC1
YUILLJuNQU2UvgFvzFlG36e5sUyzLG0rIKdabCSdQse4ud46OpxDMq/6TQX/MxLlTKOyOjKJm25a
xv4+wx8IahHvw6IkVxvf8T0ahlxVvcMH9k8gDwH5yHEXltQ7VKeZ8/pmB5WMfdWoGE1nFQQPjj/S
z4WG3IZnbQ6YdYMyJ2mBzeM0KENiXgkR32ee+FgfjDYAo/Zwl7tw8FNiWXL8//DXqoULvDwE1wTl
QD8qrC9JuTj+OGoUAow8EzZGxDCd3/R2UEvYO3294WAyDzdhtFKs6ueCM4gqub5EbCS+SHefTbMI
hJ30hbS/ySIhvrXsnYGRpBrBqfnsoY/JXKyxGJZyAL9xb1Jek5ud6aOGFpotcr/nQWIXGeYt1o7W
PX9RecGU0dw/gLvXQ0NGUl1dYJIfhYS8Ans042msC/hoZgZGaJ2O33X2zGKOHA0Bp3zrez+V9+hX
iR9+ILmkswLw7MujBLwthqYV6YdRThrFQR3kjyePAszRhTDJ3iSDK7KDtv1FD3HBHC1SQPFLwNSI
qPhW+hXKourmH4RmHr6EB+kkuOp8BI/ssVDE5SWZHTKBtlfiJhcQPgD2joDpgV5GoTcR9TuYPkv8
KbIFIAwtYPclwo31E2nFMFbNuC+UtXJBKl38nnneEGJVjcOgCh0MZYrL3Pz8bnowBtyiWmgx8gwx
x+K1OobG7/+KhizFoqxAaV/kz+IiRCyN5o0ISeM4b3UPsT/JWVgpHTDJFbaQHTLlOTSCCzEOdgjF
6sF3AkjLvPDUZO/lBWSbTJ+XmZjPy71ZRo1uuBqwjq+50JWOCuwgB8iHgkej2xMuZeFsdEDRyWSz
71R0AYZlYuFRg8sQfylaHU8yAhTLhCcVTRzEesvLIO32urZjgUNaH0wuq/3pvZMI2HIlpYwvPpsq
alTdJSsuN+cPnxIssoD2lqWoRHSMhyvkvGmQheK7FRG7IrOxYHd8P5b3dpfEdZCyCM74TIlGAng+
Bk9UTRAVeb81bmO0dmRptVIAHp7ZDrm2qoXYARPHItPgmDzGVHEE5ncgKcic730gB1mW1BtfFuw3
h7WncSt0aM7gp+bJ8PXFtHL0LaaCOHs3lBciTdYowd5dxjktHcAW/1gvraweKU092sW9GBZtqeLF
qILaA4pA9qOu6U3IRhCXM5/7mzNY1I7uXY1wvfTKzQWErHbmCz/FpGvSPyOpxPqCpjOBxLJbfQCQ
xKlLehqWZ2fJDSbAQV8jTiC6BO/szHi2HHXADuzWc8NXOT1ga0DFWEP+dM3AA0yLO/inJP33BKx9
oME/fLDqwq2ea4xlky9gcj4qBmurTjAu84SMqs9/xsdtVSPiV6/KRGJ4NJIGP056CzBQx1hhCOIG
kz51i9vUj5RTTY7MyOpV4MJDGFoXdAjEfS9ZLsDBF0F2af5iNnBCGBqPiJRd4ta4aG4OD6ioPAML
EGn+ACZOktSnQLvDRtc0bsA0P5BL9Iqpbqsa+3gA/c39PSXAO9DCPMaIJuohvnG1m/SKEexq7ptO
g6cNeydJBEyqhm3EpODIgvtRHyI1Wogi2Xl9CABttlryekFvBd3KnvoG8776EfE3Zlc7o+ZU4sXs
I5x9hh392Z7/GDcb1+sgVSeX1f/ewh/3lEp/69VGIkTFzZXtiAkGbIcTvCOus3+bX74boooqo/po
S3kvrQxiDkFLz5Vq5pMdEqZcBKCLy0GEfCstMawczzf2L7huV0T04JmA9ll/QOT51/2FjIaL/mAj
hgyFQzRzjJ2h6SJJdxcX8fOLkKZeJardQCaFTNbpeqnb72edmrx+BLZnOej+EErQ5Ag7u7fiAg5C
Jx6HUajFl6Iu5uwYS/a6257NThLWigXdSb7lD06xoU8SsjTrMY7f2xsRDtMyIH2cEFaW/Mlm+k7P
djcFl+CVgWbTmwfUNhnMU4aIEAnANgSoldoZ/TLdO4Bt96Spo+M0fPLh9IvE1wlhj/HVfkzA9YX2
PTZVBNm2HO4IAcpmpiFfH+VD0SwQESixviFUFIrx8Tq0BBX8MKKKlnnHnIWRgIYNOgXo2vE0VL6Q
B01yLNUq/ublOAQBxtm6qR42lx1S6gQczmGg6q4eCZBOA6d+hD3GRMT5FqCdlieG3i9eX/8MNzhY
kVwDTNExwSg1aXnS0EnFhFkvxLUVly9C3of8kzELhXSQ6WOZxhVqrXJtsq6XWnsDaWBk7S7kTnmd
Lk75xKrHD3QmZTAMuGH6fAqEyh+YGGI0X6tAiz9SV5y4z8CGW5DeIzs9F4Mg3FTxc4kMXFcFvo38
Zy+FwRJyUwmCUjzW36rUcWfa8/8fjKKB1RHCuMaOCtir1Mz5UPrIHGkry4IvT5es9OXu5vJ7Gd9j
z9boRqwAGevEVfkzwM0A34nG7PItPCOhR1S5V2fNdZNZ5tLthFlw3Ql5hbnAicYVv7Q2VTkFJsS1
Ke3hqNnnQYomcGEQY5UaxutJ1DkEs9wIeDVhKBwJLpMo5WIWFI+8SKkdGCLrFSSiy5jjJNWN7eL8
4eftPfZd6XNnIy+cp//K7exxuo+AjfSquC5CeOuI8MBR06EH+9+TcId465JvlVz5GOHa1NpDnv6A
nLNsKsJZCSkGLnbKD80l2q+o5CxUjU9nGfiuzq2xkgJx0NXCa3Rzb+ZnvUt9EoQzqSg5G/VJAZBl
KQT0wkKibJAyDnWmlpeSznrSwUlGBgzQiHwd9rCVm217RnbXhVKATsTdMaHKv4kRU6f7YzDkWkcF
U2nSVZRofy/bmmgtovG2QegkNoMC3uLqythm1jcVcG/jG9wakPFME+SadBYYVVzr2LmS+SCDXfNR
Y5OLPJc52VlGMH1Ptv1pRFthwZaa8Erl/AbptJObbxUXryT9z6feJqchPHnsQNexyl/Q1rMNZoKS
rJcBg4ts88qgEUOHexsbY471MgRmOJeK3EjXiBrp6sShDyyuJ7xiXodb8bNQtT+ZsSI4+y+NMqyt
EnGhrOhVihL0Wnh1xkwcDfb9/r8OM0i05qHcHhMWsGg665hMYzZX0V/ZlMQZHWvIwk/aLUtBCeh8
QKl5MiojmMtTqYCupuvYjymzanb4pD01upoisugve7W0xi36yMxNUlTPufoLFyKQeu5XJTvmyB4U
PLjzAhUUDVuK0gSANT8PdvhEODQmGAXIeqxydCCFDP0e2hlwU4sxUbMN3efSg7k3jIMVE3wQAN/d
nKQN6eo3HHdH7Mwk4TSh9P/XzGtzOdVOl2cj2Ny6pGRCBVzIKwZISQZQpxAwRRu/mCmacQFmp7PP
o2kyoA8UWewZ0L58q1d7EQ7YdGzKxPDKSRf4/qXvLD792ht0ftgr6QgY99bcT6GA9on/ce7H/z5U
7Ye9DHK8YGuBj+X4aBbhMpZAJO6kUI8x1lULFLkZfoyzblJY+IaGQ2OelCpVEt2ipCZvFgmNz8KE
c1i9TvvUuzjxOJ2ZtROwEYciwsbN1huETVAdpA2/0tERSGwOuM7OOuaw5j43uFmx0g2vCnJWKsyC
89nBRvh8JRzHf//nj0Ue7Csk/d6gzzFea3LkuxavY0ZPRdZvM/CQzw4lpCJvW9ykt/RACtV7PmKG
xVMCDa77Z1+sPOwK09AKDHI4ke6p8tXYmc2fhzhTh0fNf2Aio/2ctN5dmdXO6nUVJVG131+symlR
NWMETcKanN30HUHOIjDPo2D2YxcZSZyUDRwj9bpDLxC9Ccbeexd3TIQu2S4zG8weE4gfvPn0+787
hl4wXhQz8zr0AljPZmPCEPtRwFwxogvvXMdu9UEQBMLb+1rPSRmzOL53UZxRHJcpgCBJNgJT5/dA
9VDsoOihn7CLBz5qlzDjO5pv4FujX5uf0SYfK2iDxpaWMEDBaM/FVY8c+D4ZsHzKB/RotKEDy/cJ
v84oyULCbBxYGGMa6KlieigdoxcACjjMu2ioE66fdbS/InWzOF33f0fP6C0t5N0jJnK7F1n/uJJc
jYSm+DuMOqy14xYSUO1DUoq2fMJe2uOdRzEA4RfrSQtU0CoiCUDB++kjl/PWBROrkB7cWORCNIRG
nDKKfDf1qjX1/bwbYVIMHiJYO7sTn3hDu3/B+KDFjeLWYiFy2ssyoXtLDXRXnpSv8KDFjoQ0PQHG
UzaMD8sL9VVK1aezdaJqtD9i2bpmV4ILT+kOjZpEUuwsrIOQrGCSqcObJ0/myc9NB6MgJ8dwFwxD
G1ahbvzxH5G2hSvMpPOon8IE9IlxtcFj+xQlm0dWTCPVOnOwYzz4JuF5WqFMZkkTl8cCaq2dCAQS
Kb5C9pEvC4EAUmUN0HcfsYij4r6K6KIUGuxto3jxXHacl5LDncuKs839+SL3ri6l/BMLue9EW2tH
XSsTi13Eeac1ccS+OJyTDaSrEet1FKeepOh+Xhf8zDHFh44xGoW2RKG3yz+UXHUn9s6L0qZD2ejY
sQsOYhb0KqFVtNU4QiHJdN/68oSpLbbFqY20YXLztmskmP1twQYfNmXqBOnpjxqfHDHeTj48OUTd
IluzjftelL6uVYqoHjd6SH5tyAiLYsJacNDF6MPDUm3QFS1hjOiTB1J2uN20JW/O07n81iZtasQK
oyPa+BGnOFT0ECZuEth2WJXDF7lQaPkiRPbexohHjyYslvGcnBUEYpk0uVMD6iDmVvLGNQapfwEm
wHUnbKjSiE2tXhT8PQ6vGF8fhj4HSB+OEBMfRYYrc1g4L5seG9aZtJ/H6eepjEzjHTwyL7j6GFEU
G8WW9cqzPx161MfuYzAoPSeSwcSKRsQ/Wk2tk7lNJpSjVpP+WwfWaTQ/gxbY9H42ZGsUTZ8HZi3y
uUGkFz4LYQ86VkSnZv//riCrvquVkrxxUcAGVGkeWeschnQDoKqhi8pOMefF9RddD/+iEaXnYdSC
z9t+RFJoAypJZIaBMqQ+7O70lx6N+Ey3wH7GCmSUUahenXC70+R2PLmHlHUckElOb3wZgRxn3Ypo
01Eoun4LUeu11BXyyVTCbER+BUlz4zgwQl9jc/cmMZnbcA7OE5005ecRegn3c0EijO+joEhkuNfn
ACelRF+3w3nK42Z+7RvdxM7IiYIlaizONv2z3+gJYkDEBJ07epEzgLnPebalgsK7WbbuUE8Xa/eW
pKoE5xVL9WR258yWUU5pVhEHfr44xPfaboU2cC7nrKa/pUdTfdESbjtjubMx+kZTfeEldgGBRA9n
I77FRlgYiUgCLq4iO7ut6a6nraRKtGPtqifmMh8QvGmoa8ctLKatigYNzuiiAI//qULR/TLwZTUA
HGpoBoUJ9zGDonaVn/Av2RFvBxdhERap2QmPFpWbDfdWr1YomeH+Oys4YssniSVp8Sg0hER763Fs
M3BN3fumfZx7qJ6ROsid9dZY1Vt5YpHapAttPU5P801PD6cSEVJs8jjx3+bPDEyYjaaT+Ik3k5Gt
e0xh5dfzm+hP1VeNWiGtvWhB+4Hhoj+J2b/t2x+4yur9y1vt2ZyraNgSqMb1vn8MrGj9qQ8if5vC
WYstGz3nYqc5bU2ImuPprIYX2rhDDhZ0p6UnH8RU6yax7tx8Ypz0k8sfYWjjefQ8cpxjspFo36ZO
1NYpmP/o07S4QoMKB1VmkFayNQyroLhTLrTbUoDWwfasXARQzqRjgUcOQUmYnJgJuiTfCNajSlsu
mbB2rLfV6vvs+wUT+bkGKnPGxTnZoVVvrDgTAp+z60vj0BvYxgLZdtxEzS5b6+8T8mhJ2Vu6VuMa
aUdJ07aaHLywx/WqB/r98PY+j7Co2yHsUGMsP1ZyUg7VLBAl79mOzgmoCVwJrXq+qEZk6wNVp5cp
/pMOZQg+3M+71cSqgjfCnTMJXH2vArvpcYNMfdARhFnYotmCzbIKt4iZgpPPMrOKlsaNLcabjWVE
PaNP8V56x1M+LM4fUFQKNhyPN1XjBBpATGaWPkvcPcysntHVvjLdpKieTYEvcG7U9eVQczcfwHAs
0ZlixYeX7078W3vsuPE314xXjQUuEBjREBWrl9rwA/X28EQJ9TBrSq6yfree7gSYQxosbSP5VtfL
YxZwfyVqCJD91LIXhStb0P6AxyP0O4wUYYDe+z5sWYE8d7wnVaZvSYRHxKkcsjItJsTdEX3nuLhM
0hoZYM5BWE5tmnd5cUEdTD/9nFsc41/sEzeHak/zLRbtz4MLNGXqnIYskyfxhTyvg1IXkKXUs2sd
f0QOp4AHJ9XDKHLxu519OYOxglToU25igOEQjrBGoDHVdHU65AlfSHhz/otw0+Sukt3k1L6Oxy/s
Pb2QExKY9iupAvrbLpXVZVu4/W/0HFi3aqyp3h5GepxAzJ2tXLdgs3TtA/Zx6zmr1XIkGqUWQU0C
Ey9bWRlCLJjFMpt2omJuRWldqPqpjiqbT/VuymPuZd/kvZeXiiEDmYoTVKeFC8JyVcGA2NFg84d6
/WfS7j1RNIqsjWwMSV3kjwWwuB0FE73UFCIpA/oCIsG9jDhlJFFBBKco0mfGnG0oGDGrDQiTqBZ0
KeMtrwC1wM3WXoCsJMSkkmLVmrnm1/byATjrqCT+9WZh6XWNKJvw4FjTOhuKPWudL9SmQx5IU7sG
dJNkir+oVbKxhOp0YMk+p/oNPCGqtHeu6gb6h1roWzfm8f0J8svTkh3Dj3PbaeqPl0GuI05kIqRg
8ditgDa8ePyZxBDLH5/5/K6cRDjo8tFv+UHlOEBJfy9lQhCi3WF7zbYN2Nam8AtTTkfqByG0dq8C
0m58HG3OKQs2Y6//KBjM2JWd3IG+4Gb4tFWyUJ/KHR4Iu7UqesQCYLxjcA1wug1EnyOKjIHKh6z7
J4k5It1ibbm8KF2ybOh7Q8Q1MqgwEznc/ch0C3h41n85l+xzgybn2rTI1mINo6o7ZDm96wiM8PmG
o4sJFiqrXDJlRctQyKjcBRZ6KHnaR+HwVUhcTQHZMZeye2aNca7E2ywE/Y3YJZXMBwM0wN2K+flQ
CLN7Djm/5W64QktYGSKW1J22zc/QolMv2X1Pz6Gv4HCTsGXvfJPua4/osmzQDySGbnyh33gJjF27
ehUjDLYcGtvSBYsqKyHh0qAR/MAQh8VWmW8lyS/mPGlZmKrAWGZDDDUlUiONk3LpFLmFfSxTLUH0
7sFZBNewpwywHFRelAC0ZsM3iPIv7bQk5k+z90INy87/KB8wzPfvg4pFXu0oSl4yNnvZlMbKKfZT
PTtgBFU1Fbm/n9pDdBefp/pErcumLRhp2vtVSOO0pDT3YENDSBzQWKPWBUbBif17hFY5KY6yBKlh
OCkSiXN/y3bh9RD+u6ahq2pXJJfuq7qfELVG8YDd98IGjbCFIp4EhfQSGBti0ETJQZ8Qqy6kzDSf
9OYC1PVzNOJds/MBrwY5sgnIOrwtR3V0VMm9sunmON04GvWSu7cAIGyi0+DhTe99qiWwZhB//f2q
Gal++BNbK2LB1hSaoBRaWarvau0Ruht/fRAKvMHfQ+95Sn3Hwe+7GI7V15dJm/WO/naBDizMRDnK
jn3Zrr3djnC8Ek5ZW3gliT/DN4peCOM0rVoFW8VMOD6HcM11Cbomp2x+Ufv0d435CQpX4XmVRCe0
S1YHG4GlXrnyeAgDCK2CZjkS9/WZsR/D75VZDUaq0KCyiCqqKeHEOnR0bL6vRziQkfV5lr3r/FgQ
BwtUX3S08yfPyebOCDKcSlWlFuPA1GOBdQgt5PkRpFJ3CE+PE6Jw9wVmYpvc7geUr9ymTC/QMyt1
FE7IaH8RjwDmXpehKihz31kcoeHShAfmLHMFXJsVaYiCOdHtEhnm+cEbOgwE6qkUoLAeUUTHODp7
LECvh8lg6wpvsMjFbgu+S/5/Dte72fT7xnzkIzRXUl/zZoXhxwb5wea5CfQAWrx+4n/TikhJwpvK
Z4gpR57Uuaw3cfY1WcJBqTciSiX9uMPSg7pImYLD0frocB3gHQrgjE6ayfekQL9kyO5Cgk2nm+zk
CTmXz2G0caFedrN7nCQ0aAESvasuWLXwRaJdrPJcy5G2YuaDCbxV7AcsBp+Cib1khU8Z27p7sa7p
CIf6JyHMszmeTegVOBQ1d3NMwdi5HjjpVE+k6ljhOrqzK81xWtxIl4QeZEvRCpz2SbuSuzd1qJCT
ORyn0Ew2fmM82S5WqcObdFypbDVEDerR4s5oFO4UZazBxRuxUyyR+MDs7/1CnzFqfqD5rsmuz2lx
Ryfn7ZvJH6a1mEdV0vipqaesxO6X1LmbId5vmP+/UU9mzKHwBeKs5+LYS+8MacMIDzWHCLzwnsKF
UTbPiULBxYCsdBanxOapZhZ8xhyFzpji5blV0SW6BjZHpaBsew93KgbmSBSNWXjCKT/ij77Cy7XB
MIsG+8ERUykb0ovcddrY8Rnh+uZJjrHSItLSfXzWRbxSgfgbyyVJC0WzIqJgnXbY/lptk8b3G7Lx
xOCje/RDvzyZIacobAi1qc07tU+mKKVnbb+NEOeUVAlw1o//U7xuTShfjfXTeRZg/qS/4EAsiEtC
pORQ4kchlMoSt7I8JsYkECV29gAMNpqiaFuKvIZWZPIDqmn5bNXfXJAPjWctsuaxchRFnIle5wix
DntS3AG/ywUtPJ8f8O1908gw6ckcqA/FJKZRmE4oqyphFV6nqGDjHUWiAM6b9GRdwCFrw+Px5nQ8
JRulqM2UJsF67YG/CtPSfSrDEwsrZLcUKYGjda1nYoCHu6Q2SZbDQPZJwZ4ba3tNKJdh/hjgqaV3
EvGKiVSRuZqBeaxrKIXLmlgZy0akbUWgSvnaL7sBEpUljohTDBUGLK/fjsBNC/bu3X22je56PvwJ
WPpX+B4mOS9+Zl+gUIEtjzUXn6ZbVaXZ0pY5ePoS97WMbXXIiEO4nrghrkGq10czcUfUyd/1MiYa
x0klgI5S2DdNn8xaU2tXFrPwhiI6bNpWdTRgIjYXDLBPxV+MoCUMEeE+dZkk52zQSI1Mg71PA4jS
ik56Gv/Bs/JPO1WeUFX1jhRaZPwP3mAhdD4nYPQ/3piMIG10plCscffYO0ZEVWZt3uLI7ayJGB0e
gkXPIacYgyrgWIMTrPkUHyDbKCmuApe2zkxpzo2cBuATgjWVMTNDua2SFVy9tor21rurjmRtOGji
N2H3c0pQdiVFArrei0eCS/uWjCz1zJBVJcyleqZDrNBrZ9P5gqIwjXhQSjkjW7LnxUCFWHZ7ixPm
xBpL77chBYNVzZ3bEBf9M3nfdQl1C+LzFMTeCxjacoooVhY2Ue7n+jfTbkqHZLGOXXzlVy041pwf
TCmugr8EpNpAjW/Rrqh0BV9n4VXhksoYzSURh3SQ6X8PjEPpc4yAarLN/2iqxs7hfowMiDRyx938
ddJlb8gXmdGAJ6j9lbT719lfsl35cTeyOjZHQbKNvsnb+/onUtbP+HS/wAoWM7AWnqJdJdKfnNT4
FpJN2kUIdmyuZmzZ0ZH+Ptmz0xlKd8TYnUnmn8d0XaAQXKu991hXCPqM9xKImA2XJrc8ape2dKCu
T7DAMzzsOAZXdOYGbkBPP75HP6Pi8c4mD3V0PJykL1KZn7iF2pdUo/HmLGtXxx1AErBovhSdNo4C
KovWcNUz/r+S2C+ta2IcUopeQv3yDutYQV+zBiWTfmgzzRv9DUZdc1d94CkQGw2leFKd14qdgQ3v
43YKzLBLPj4NUcEN5VybZc24pBNupGPH/8avPT9YDaGZ5wNsNqfGDKIWmjArLrEmbGrQ36Yda+mX
NJOy3u4hB/RX2vFjF0x6shIQcBXwnSN0Lp8wrfKyEa/oNUik4EOjoUEOdC0xL66+AabBJUMZ09Cb
p479V6fNm2jAEMDVBvSPnHvAwYQqUDqacsrSF3EJmzi95F8+Ng9QPk72UQ2gRj6etJ+Nqz5YK3py
sGllNlpt4AQQFr8AvGLxbIrNRpeNS27Kaa32AvMmETe6aabgcxbzA4jGhUKJg8gtEcaflrEc0jTZ
10eqVySaNiaystZt+xqiKwV+IUZtHWczOsWSM6EB4+EBtg2jzt7E7FvhJ7xdZrQ60ttrDWpQJgZy
7ej/LMP7CLtO6Wuzh0ElgfDJwuEuzS8XfNfkd4HzbYCgylJCRz/MOlTCFstQNybFrMnSyp89srll
yQZFYskWzvICHgvAvJzS+8i3gk2JcGIMiWnJOFRsuojFtzoA+OXalmSbh7ZQNQpENXvQkxQczlRB
TTHEuf3ZyiYfEvCe9w7Rdxk4p9P0UumijAWiTTrOOz9l5kRX/mN/k3VH/VYowodNDcZv1eRyPft6
Fvlny7AH1O1tYs/SWQVos9Q/JE6GfQoQwdnLW1oZBdeVDFQkHt+s+Gc6abc9DnZCzyhBCL7DY5lo
OxgBEa8x5gVEUHmlT49VrjylWHaBEtgstfM/Wvz9i1k7uG44Jg4ACgvaZoqh8elZjXpsqUCEkYUf
V5Ttz6cHkYTiYvZ6UYUV5X60YDZ6aeociH0VY5LWt+xrDoatgPlhnfuYsXncqBR1JsSkYYtJNVk5
n5JV/Hy251ARnFF38Xf1ez9WvWuDoiqupyLbyDlsjwSTTTxzJCyCRM0+rEzxVl4h1Dn4pOM4lWCb
EbMkmlYF0haEg24a1tMMW4JH5+vWM4mXZ9UHvWR1942oWeXkoCMnJf4lQpE5rAwSs5Go0lFgG9KG
Zi9h+Xme7DNq48oREubDPLqdEgQzpgN1G764OViYXVqpOIs5vqIFL1l+y5YHyg8XdkYg7AxrSvlL
10/y4XbQ5c5peo8bB+Ifdu31BPi3RuX0yMfF8+aK/J9/pKAeYDWXDzW8M9WB6wOkFuEIfA3IscFV
U1XuJiHu9spUtR5utLnQixKCD/UYOnxxtL8cBstnlnGEnwdsUkmEk7igPVgo1MNLuzAHNCHPdtOD
fq+ya0q/oKk9fjbwIAnY1f+L+dKmm69xSG5oL3AwBDuQXTbavKqDFgLiYhbbj17Gxr9wPaet7kRf
07/OiK49RCuYY1pmlkw5Rxg5HGG4GriKBSIRe1wmD9Wa+HnNGg4cEGHuof3hPYbZHLAa6WGIKaB/
Vj4FAFjKQKRbqw5JblgZqJ8mfavO3PlhFrK+3Mjaqk9yHiwcIf6/YqszgWTZlr3POIcavoCQiXeN
CSdfxyl7rQ9XFCoHW/m3RZKn6GGD54JGkqFDBxLDcv469wg4RwBRmmMbWH7ZoZAA31EPFXkX9dTx
/zjeIEygkAhA+upgdJ8Md2QlRwh3SVt6H3WPw3qTUQEQDjzoA5Y2DxMZpi4OKF+JqqwyTDPqxnfe
WhLuh2BSbNIAs6IoEZBhtQm9WePUhUsyRZCwYDfYw7GuwxAPj1PvS9yx6c2l5anIKOWuxZXD9tV2
6C1N1nxwWTr6A2pbwqfwnxkWM4WTXtbIyE/kij/B8oWpiK01+KMFDr00/86A2jFdyoJc21IbvJxT
l+WpN/tCsIeWOP61Y/AOaG3qTP9exX8DfAxl2P5FAeSjMqrRwIEBcTaCXoyoNsmgfV7XvLY3iIAu
JZQ1fIp9L9znRHiwxjm7UdkjJFK5f8pyf5bJiDpRV1ejRR2iFh7RlkZm/JtNb3QL1aB3epusqjo4
x11G51XrO8beuKW/Ljox5Y/3/7kwhGHvkYCMLGSBLmXQFq4dh6cIDM9mb6lu567+R0cw7kCPkQJ6
55SIOBlXsttILmIjR2xWZYRw1lgZhJjOSZ3ACl1rePpbzQP1ZePL2peb5aC5L3RHXsBF9WVXCI/X
WFT445XGHDN2bZUZNOLu9pqcXb12NAiYcJghAjQpeMmGHimv7brp5EOEfOwsmA3riZtxThDmo3jM
6agEFoTyyUvB7I3b2FVUzTs0OMtCVlmrc4TGHOrTCsuFza5JiI7cJjLcAo30zVk6/vz9EzD62Als
UN0ghlxXrsOAu07kM+DJx8RF3z+hBVCLJUfvynaMZ0oohwo/yYEYi6DMcUEGFH60iSOguA0oNsEZ
Ukmxkd19n1dUu9cxHwoJu0MSk/ot7brAfREMWHT5G5o7lruSu9Amx0YwQAYuxg8623dLNe5aIYUm
L+3ZJfhT/5KrwbEiyNPh3OQ/ckPCxoqPwL7PmwfLyIapNUVBSfYJz8fLu716xXdu4H0TPeejDE6Q
ko5Tgz/ElYJHixDPb/DqKy5mmRINIcdit8A9Re85LjxPvmyQdaAnAahZl9KVqfplqmos59vkH05D
C6S0Rlyu781UFP/1hXpLmK39elFRwrlew2wZePCPbT+oPYMtIw3gE+afFMCT47f9LG/J3nvg2Fvr
JyZBDbJDeuIEEpNkJhTBOWJx50iLZd0RgE8hPnVvxk01y9aRlRGqK5yzimaFf9G5+vVlJmJs/IiJ
DYsTB5e0SnUc+0VDcMvmrrJ/FtFzQKYlrrA3QMYfhFsESPjK2XMfiEzlnScEnAPwK2nbUdAKbE9y
s7+i5bDw+fd8AQq4el+pc4iWkdjuATOeXbx6F8uqAfo1zURzIZ2c9VHp4RdETgTIjMYwX/DrguEL
GCRM4OeJaXF8jqGOY4mOs/E+nbNz2skrN7v51Xb401Y/+erOTXs9LavCb5EXg3VAyS23Rotwx+sc
vH2LzslR4GjtNYlhbLwNGfl4og7JQ6Icb6Kc7SvoQRvcKcpqYEgo4NPy4rRk8vDRoeAvH6WvVPRH
s8nuQWTgfOI7iM7sHwS53w95vx3u4dGiyz/f+OprQdPkx0KORUvZwRARkNIUwhorP9iH1RVVDa5l
qbapFo+NUc3nnUkIpIpoLX9FbAwgp80YbW2owJm930KIGyzmSoZXqijpQraDb6xbNm7neHIOMtYh
OLI5kMld/lJSBO/7P7MWAOcTdaqGgOgm5FlcW77H1/KkHzzWBRfZ5vJfnz9b1sxG2y1Mx03wXhIm
qQBa0m9KYu0+KOiDO7xmBy17QGZSbCvgZgyZND7ILL5hYevuHI4gy6wAfXSuKu+hC8I3R5x7b/jP
I0KmfEseelnlLrsbvHfLon5ll0p8fNZlVYHs7jeuHJvjNGzzaQ40szCPEtHyoJ9sEvSQUoHpQ5cA
UlqO38M0NvLIHv5VRBTEygMZ1yiE1ym2p2oMoTjmqe1rig6rOPBHHSOyiMbtQEm0bXBp8dhOUboQ
SHFRTHUkahZ0s7cH2FLZol1J5iodpzW7cF1lZT2LDEi8+K7AXlnZF4T0v5I1MYiyvYUYW16emj6+
knmWNgCA/L0IxQmkIZ6vi+JCymGHtUuJ6Tna9OXUOYFJ+oU6Ba/QcRM9AeLT1B2+8yB2PiNmlaDW
ZtTCnpH7VRufeFsUFnrwCysjlw1+aaQHDisZq2ENuddqbeqMrVGZpVnY6ZjOGkVfpe7muXngOzk7
fTYHXwXIqiUkFgs0yVNiUC9TuK13tuwMx2f7XW+AQKxqOmfHSCTPsw4l0AKW0un7vZbaOx0qSGhM
+iOq5xVnwdcvxVvcXC1cjcFXRWRcLBAdHfD6tAD1HuYWFwduPzG4+vXRkgbG+ULvD8NeN96XsNg4
DpvbKezvzMtx8uPdIusxZiezwgZZkOGUE55+mG0FLjYpBoAQN8gMkBGQ0UW6UG2lhb7Ue0lX3xGD
sXWAP7oluGk2ImY/N3+KeIaMC9WNhcOSbi7fh/EFtZM1/E4VWwiAv97c/m3KNlnVRWe5GXmezvpJ
XVolZ+ctBv29kDSWSp/gLyccOgHEzkOWmqYm5AW3QWtZcdFsk74q1LQV7RnXJ3vbfhJsqOP5uUVO
mUcPezGD7g97pkREB9iQlDm79CwCn6EQDPljbPVShp6Ndfv8k+nIybzDJnJzWivBtT/v6PZmAGrP
oXyLk1GVfc8C2wDsG4aeNA8B5QigAp1SV8tjSzgPZ1wZ/pAuzTRboNN2/sLcNKrmKrE7Oz7+buTi
KDaOOeGT7PtRVOhHumJ+FP7b2ZDq1hIDhdjB/AeE5jD+cE53a5heK0jOM8gxsx4Ha9U18q5YmNY6
C2yOIDRNBQEmncx/iDDUAiqDwPzTYdNPmDW6hw56bIFYcYB2tJqsX3qXtxqqVV/aMjvOTkp307ph
jXio2t1FbEgmCD7nVoBHPhTIVYLeasz9XDu47Hv3JCifHLfoGolxwrWLTmSkKncguzqTLnMBYgnT
QMq6N/FB8ohzYvzlqgLML+epIB0nEjOa4Q4+OHCa/gFD0j1A7iUH5oSfAdH9DLrn98DiEOEKUbsD
RYdnSaAXzu7g2dHDhXZ5GIWQZSkNl03cDaNywqe7X+LugNPP7gt+JlRmDtYMW0FyyGswm01pYa4u
s6Q0Bt4B6+X6c+28q9kP9zBgHL2mOtqvKP3TK3KJl7DYImgOrxl1RMbASPmT6l9OnwZLMAjjHVlU
Fzm0/FNavpwtL8T/RCv1tsGPZDQ4jhUi11DrSJ3VZDjKokSVoTc07Anht2TUGl+3tPjXmE6fN9v3
kokuJfvanj/gRGILnoQDeNHos2klF1rHkNgU7In8UX56iWtWj/2Hmy65HJ+HWJD0X/nmZbjaJPmd
IPuYJ5ygRhki9E6yFIoBWJ2MxCJ1s8wL9uHVxyX8V0I2xFoVzgwh1v67tjE484J6YYfhmKdqBz2f
iRqAhCCopryz/rpvBvJ4pf7igdHneZKf7W6FcR9aIjf3RiHXdPsOXyvKx3ntgPKkxI5atmlZxPr9
hmXnKKidNb0tCQEZLDVOMquIZvADeaciykZsXw77W//W6/eXJRjIbnRrDVsROnGAn3k4Hykfj6aF
YDhkclhkvaJNTJ5wIdvHi0UBma3cHWMFfpO51BCjsiNVNvwB6gr3ux3NKxeLyWQlQylRDc3SfnD+
DAzhv0EpXiDSFkfox9CDXZOGUEOqXlWbaSYuFkqIGDvW8xWPi07MsxEcYkSN/tophL5ryuD2VYUx
2zNNC9TA9Ixk6+JDGiQIr5lomq+yHj+THnhvGzsdU03ESylmRQCpkyPIxIhHBMHlV5TH7RW2S/V+
x25VKG/InSYP/COBpGcim4yeWZUAcSTyzk6XxGZBZ2eRR2ywa5e73Ze0hGikCLZwV8kKKyDQZ8ZW
wB1hkc899eY21czD/gL2ba90U46U8qkpDgNMr7QKapprVUufUMlSjEv60Mqs/n6tbWLCyn/iwiYX
KHOZXpLt08/sCRf8ZnZ9CfrPCgc8URCcJrPyjft3Kh+eIrFsfKx07XOY3UhXlpS+eQN/W2ie8I+m
50qdxPpsf8yACRdvyLC/wB0VnhdfMfYRBLIP/GBS7yQZ2eBPMUfrTBTCYi0ZlpRX9diNCKcYHoZU
63dnIilcV8iwghNa0BniNQn43LeSoQCuIuPKV4Nw1k8b7vLOHxADKWYL/izwzPYA3tLU8Wc/yAH/
l/bMP3+k8mq5XerpqSbq4r8t5OAT44t35jYkxVTScJzDIQoL/XdGDMEz0cuVTZZgNAUv8Sgbx3MB
KBuNnlNA4LbCRBNcaGTg4CnZIFxAsxpDeWYMh0euwZAxkf8QDdciT9pb1/8F07/LADvEOLrgbVkp
eLVvb/O4vOCxGwwRDOENFl2qnNQd0BZRH9mwx6QKs8mq+Uv7rjH7ojmJ+DqJeSJG4/HP6NhYbuvz
5jDZMiy+e2o0u+balshkt6oM0eYyM8DfiIEBxof9YKlreXeraOShwxQ1lC/Ywauon08DLurvybMO
ip63hhAHd5F/DPaepU57KH1YKZOsMK2gEh/0I0NvVa6WmK0ySpvDOzx+SYZC05IgkJEx8ozXhRu6
e2596IJV1G9WzpeIozrNWVskzx97cQcWG6rqMS0NRvRHwp35RUUCKCrirNGpDftLGAEiH1Q+jLnh
utSuIK8UqqWSLDOlsxTokXYUNLf9uyJsubj3iHOlvr8pwsOMrigcepjBsTXP6Oe4iy93J6mCeq9C
n44kNyPXdPjzLhtTKAdvSsu+7G1whZTPmacnw8tCzFqBLbT7G6ivGyCBAvrqc7xqHNoEqT+0Z2+/
UBgmGB2z5paxvVWLTIvIQ7+FtwPdVk608vOr6od+iHd/heJ78+EOkllTQybknbGfVUNY+0uLdZEm
V/W3Okr/ntO1olQ2Il6NvpE09yLfxu7EGZ4KuGveb9JQJiBgdx4iGhPyWSxH9ZTlF4hYfFkbp8bB
x8HALRSbNoDwIZg0ODeAPFAqKmWzDmokqQ0eytscA45c2QH13htWjOGHCLzemFSgiXXK5GTFN7/G
/auT0dHgCWAKcg1iky/GLbiMOGJ7N8g4N2gl6JchYSjHEoSmoJIAfIx75T4oyXuWmiefYf95+TkU
cjJeYXh0K7kT9/SQCUMMG9Uzy46VxJ8ePrWPLrwWu8YRQciq/wBwoP79UKO5+gvhuqVR8qHtHaEg
9nyL3myQDsFMRLooqJgWbIqYMNIwNncKl472hNuYDlKu7dXiXB9xGf/0xOhHuG5/Z6d0HpNbTkaU
8J4G/MykVEU7Fz35wF1XGRZOebhv17P6EVEUgmZy7j4qXkVjVwpeEkJIgSC4PHPH9iItaTDgWUm2
veybuVBcWIuV4sLVynOpq1m4ECSkFLAGlL4mkCr3cfMeb4v48xxVHhiRrkVKLI4QERo9h/PoV51X
S01XtjcZ35KTrCncT8c4m9l+a+kc7JPrPznyDD96Alqs/jpFMsPSDi6hVy61dcVthFIuT9hqt9I2
X8J+L2mUE032negzDS7FNIDj3u8oRsOeZYilEyGUovIjcvyoBJLoZFSkQ3xMM8FASizCDt9+EhK2
1CxWV3rXrw3AqkTM6p2r5R5PmWg9j0prV3RKjx5/8Is4x3K6wcr7jkfXyHs4uYDrM/LyWR0eBiFr
w5WoC3+BqJtj7P0vOYpM4nc0ZDN5HkWfXsCsGzfLVF3NjEZq1OgmCXVllpn60XAjZS777iTpdwZQ
yzixC+/fWuDMY7vTwB1D8E3cpJlsAhHKo96Eb9Y6oriaiJUq6lbi8o5q2L7uTJUqCmk8k60ZIJc4
AMPu0V4wUKEtRq0i7SPjKf0Iqv0RovkxgXEcegf+NAKQs+zNYyhoQ4AnOYyTFilp5XLucOKeFVmq
7Pu7VkrW3L3OZ3XrwgE1vnAuNAG4DahOTkxQdcR86AX8kgRogaKezHYuSUTdvRLHGyQ82Lgh+qpc
hDmXgqgLAS+WUuvZ2kr87hPx+R+ZoLjvYoTydWASnzFFsgLlqguXXEO8k1jKdcA+SQ7+q6A9pXg2
TI8+cZfYP67PXyPT6h9uTxj4JsDPRrscybRmQ96pW1grLdyu5NfSjK4hGVmE7p3N3wa6wNdF7FCx
9kNKFiWekUi4vVNt6PLQjuAYuhNJ6zuKWslpHsHEUeFDR2V8OVk/yOphfPcb6fdToWnzo6cQ+Bqr
oPdVu2RwfRRtGrp5KPg5ygd+3mz3px9v1zMNbn1N8G4CFLCawjtNIcrcnVIGl3xPwwTbkN/HeKGv
LVK/bnIVxCqCvpDvGFkqqpOj7L/wDqua5mIXrDyXV4CWm53TVUcovgLKC21h4ac11FTNLteZrdpb
K81dkoXqGSz15EL9G2aIpcNSmaSwFTZf+XGe8EsSiL4slTJ6aGvXg0aBnEsGKeTseAsVu0PiblqC
AXIcQbJulfgW1+UTS7ZL257y8Hstxn18e2Vq7rsCMXGYFevb544pZpAmJbXvg6akXrX3hBuYAXNQ
zbiHomxWbuLUwTzlFPTMfUQ/pk0QE5zbVTnj3CkY0+IXNOFJqvJsx4fJ/5Z/O0/nTIppqxd02kUS
KCPqk9mCy25QiqSPLk6DMusmi3NgeoC68IOHN2W2I9vEMpqnmt4oOltFb4BoDjtaYEJFQO3Vm1t+
rH3eFAKD2aGoNeW4XiRpBoFFxyLOrOrPj0uGqMd9qQfPkQsaVaESqV/Oau1yN9nPAAT4yIL50sv9
s/WNKQn/l1+QG8NIXkn4apL0o6nQFvw4vbo/8ntaOLhQeBzRKR/XTkZrsoUtvm9PAsUy7AHX6D4W
Te9UsdIgY+ETqeDYwIu/waikIkpRpPjts9COfV+Mkzac9o9DWTS8yVqgG0Ixv03GCYMa1Dbpm4PT
tRI69+PCwq5ewTexoASoc8PWqTFFJx7ESg11G570ANU1DE42rIvd3SHZL1OiPekXpqqeBz3W8O1M
RPoFabXeIOfmNqsRKt93n9kcVAv4URpdCvPFvfpDFsK6GYulbKxbJyqMADI195fUa4ehV0T9/EMR
WjLZerVm87vbDnvCW9zwqkaQFjGbnpQh4ZhawEa8IFwMsdfm9gntptqePAeeLeL1sKJsp4TkOJPd
t2DEbH5Kgy8xbewAKJDhrefzFuFm9NHns3tAudOPDaU/LDgNqwcH+eZ0WHlxu1nVT3a9oVTiRv4u
xcxroCRUkjo79JZzzQlCAACjpsuSM6b2+gV85Y0tY4ZqgUmdYN6j9GJJvzDQMogtzX+lHvEJI2j8
kGGZA+KRIEH8JL4VaF5Xqnx9c6Tuq8HNi2DQ86cvdWelehHU63dou+T3G/TOuS4eP5uNBk+CCMbi
Jvtn087AwbStit8gzKRTx23oWRYhsMbBkgo0rcAhK6+B4VO0srQ8qNB0V/d3HLR42PBLr5ByMNjg
UA18HUyadRq+34ZXbcv/kFyDH82estZm4//P7a3J/np+LGeeAhHDr2Y+BmkOK2elPGOrOb+HMrRw
teYDSApCY0Nlx6SFmvyv5+DnsSj84WDt9Mu6MrVRkSDor1kzVcTViJ+TsllGomIUgvwMpAC3K3rt
DaQKykeD56k0fp/U+mrkzAJgFDldtvB44UmOyUK5UUBIuif6kPn+4RBVoHhDKT9pq/xX85KHUaX9
WGTXl5V06VnNTJTgzkciQKpM/HDRrhwhQ+8sKIR7Msxd3RvPZQodV8ffoJZ2XDhuDpEZd1IDs59v
k6pSPblO3z2Nl41EM7NZhbQje2UMy9GtdWsocVDVmBgW5vJrwJhFNZJKTvhILVdA1p9Snr8elmbM
dt68DVKLgjpbh2XE7HvSP3Z2AH6JWVFP1HxWBe5Ul3EA5nbhRgFshvwuhT8olNaBfSm+QMMJsVY8
GHD9LPCj/OxKBXalISMlIfzNRmd/1rSnT+lgAekndHLc/0cQ+FKwo9oY4US7l4HAW8rD1XOf98L4
wCWis2AU0pkWorWQRjzAosGLDgwxT9Z7g7+DkCNSHF41gzYKRD7PJL+uIsmUaTa6ZgWPiUx5ePFJ
0IFS1ZAuxo8zjjvA4JEpjFgIrjJRTppEjRaKlkP3ylVCfVncTiB094v+JNvyGF3z1mcQ4Bhu3lss
Q9+MrlCdsIREPGgORv/+ea6xrQVsldjvcqaWIalQhC4t/zPNc8+7ot+Xqj/AXz2wh8qCJacRZ8Cl
sdUUE3zVSWCQoE+ilmNZfzhqTnB/H/qaVZWAfumOpD5PJg5sBSwkl5sHo0cfH2jje1qmbcSdcKz7
Ub4zz97Fb5GvrNM7BEcAHZiUNHi2mluDiMX+5t5wsl+Tm8op/PbPx+7VW9OVNxdQ2W7IgSnEFQdX
xOhasp5noZcY8re2WUmRpwGRuMUkwGAiXv/ZnUR1kNqkIqfLQE5cofTqw99SJ9KYIE5KDkt1vLQB
lL3AXk8Qu3UCDxkp9UBqzgmETfoqNPG0XrT8mqPbxPTFamIVjfGst5Bn7Keri5/IVK/I1MK95di2
otl1rsBx8tIvzn8lssgNeuic2WZGSRiVtEKLlT2qgsgD6PSNXUj+SdJeVH/QrQENZg4XCyeR5Tt5
CYbr1TeuUB5jkTe12L48bM4CB3re8KoMoEY748Q1KnKLOY+kT9bxsPL0gWFYHmWnxayCL+23PbVt
WbL5sBnz04lduhKL2Qu6d9nOSBJoxlosNbtzNWRMmfPfQORxKFSgmceevF7iFbtOXD79h4tOquOi
PremviynbKeNE0JdfxUubkBPjpijS1rcgPjPz989TZEZTUyV0KGcdTkF8+WIe8KVZ1XOIdac8VXN
aY8rMlsZrGM1tYFd3JUZy4qcavNJTKpTH+AD0qR6zC1omMLF5luQj4rfAo2ZjZGapUNFneYUSfQD
EGi+NwUOy58t22V5v6xC9oCdyEicXi0OJCt6CydlL2gno6IuRDgFdMc6hohQwIxVUcbV+uub4Lru
dQ413v2f1a6P48pLvB+jhVNPzxvAjCF9E4g6Lbd59m3ecMMYocUXKkO9qXCTmcI1pLeJao7ioViA
GQmgsvcwB3dBjWDrmdRWdtrZBBbSdPlW0g0gJNTWaEAKLjPHAMMFC7gksdqzBnF3H3Bi310Byedk
uX8/CeeO55TwjE3woAtHUoOwqYqYPEy8hcM7VkNOox4z9ip6p+lHRtPl3rkiHQHfINVS8g+6U8O/
8FFtp/cHzNDRPGe3OEN4fJLoNCXwsjJbjyep/PopEm3kCNrl6xmPXgu6/XaYtmwmp/C/4QWai2G4
JXupxQt5X4gp/Bu4ogBNgvguayCClyK7dNeHHiDlXnrDnyV2jyBYBbcfjo7sDZj2AmOIUR+gFdVk
EpMAlT3EARHcahvdcjJeY7G/a1Zxb6ot2dgbq6RXF8kD/156R3cNOipJFL5P0rpLxq2pPuFbx+rx
2daV5on+HLtclqOxMkreX/1wKKnSFsr+najC58DzBPX18JszBBX3coQK6qe+EHrOANAFA2a9mXj3
cC8DlSDVylSHgqMauldpznNAK8W0zfQ5naji2U7xcce9p4D512WXD4EcEpDhXV/Ufu4CNBFl2qrQ
C9dEMQ5Cu0YtH9iZL2HnHXf/ibeYZ5N4CpkKSWgev9SjvMiTdPh6O+lgTkCVSuAuXvM9ZSxfeV2P
GEMHhgLzNpoYHF7EgtJCXwO021xrcG+RqfOwZIy3OTNzCgYRVYA2fjgkY99wD3kl6jfvKQ64gv0b
U8evIgzlZcuO7Q0qtyR2y02DDWAX0FkMea+kf8CPvZlY72Mv6gMcu6nvyPH5hu9vSQPo81/S4CoM
hCOUDApK48mK3eheHvwHtoKk173nxac1Lq9uQRik7ZA1lrKN4bUcoK70TwkGyiT1lgaZolkry8Rf
UBqwnbAHcq/p3Lo/EyTieXKzQcE8NiAkn99vb9zx+pPWGNFpdiCTUS2f9X5Yn6TNsujOyN3DCal+
s1yr3OaQijtjg3UZ2l1guuAJlirAHkJJZlm1NI8SVYYcrrXs2o6zHEL7XO9w4/Qeec4ghnCaCfBJ
2jz3elsp/auj6wum9nQW3vdkAcG+1q0SR1q2XUyevca7pEONWvvf3QaujGA+6oU93HK1Rgmm0JWU
rg6fJWXeIrgPKfRtoEWcJSenvKrzVQ8gIukiGv9Q7svIxrYbjKZBsqxam289FKgdsun6Hvhegon8
TQ45rtjVIEQYZDMREy014AtIywQ4j5wWTMRhTHf/h6V+T02U6HtoQLK/6tIDsjFB9LKRmaNZsVKz
UHywdaZf3dxq+DdklXm5g5Tkk1w3Mnt0JegfibZDtLlXuGmJxaP29VgUnuhcNmrMkgjRVdVjMm5j
CDAKP56Msh8quDG7nlMINoBWGWsKgC3YjCC+Np1V0nC3W+O5Zl04cmEc4GEZZE1LC0nEBqiklMBR
9WploHJuP9h1nYxaJCeBrAIAW6mVa/HKWmlse6TODs331FC3c6/zWjbigXdT6U57COoUWSM1R1we
pcOEmwC0SqSB5xw2/tYoLzM1Q0Pm670FLiZXWs8T0tMHFKwlMIEUsRGDSIYN2MtptJfYgJEnHTpT
KfB+Xzmjmc7yY2Z3cv1ynQTcxeGsfdTCsctUgbkHuYYReLPNH17/Mx+n50EqrivXC73HKycngKt2
xEm7MK3UL1wsln3M11x16HclFx2jVHOAl0U3tebaHksq3+XEIqYYyNtZ8Pxw1SxxRcmdIdOVwxNl
k0XiTH317U+8A2fuMcXfvSS58n0lnWrYaDszymjyYfdE9Iqe8sNPUZuatGpbaODHUYlU680AKhIv
druRamSEgnigd1Vo+L73ndzLCvBpzYTHpAORpbYGofwJkpFCDVl81OeRDLzxq5bwrlQKQRRdtedS
AI8YX77PwV5D597ebJeRqByTW4bOVvDwLwTHh728iAjUrXeMMuBx88+lrMRvPbQr70jYCU//Q88O
7XiSt0bndXHTS6qLrZJUHe8RWgJU5NawzQl70MVLSriE5cJykGjTv9UyszDk3wOq5KMsC/SeVKLz
KZe2hVjh2d3Xd3rQS5bUu0cHBsULQUCWF0B2nIXGZfUe3C9V1Kb2LptE80tN1NCu60dUtYWlVWBc
9c90u8RO0UAGXQyeE9DOA4YIpxcVEZrEquLUpdxLhBefqu1DxH51k22qVrRkpBBfOG1dRowG+RpO
X5gdBNENoIz2vD8Q5UtHuInW13/h/5f+4ULy+fg1W1Pss0ma5oavtYm4SUB4e2ytFrhMk1KOwfDO
U+9fcHUsKgJo1rv1oWVl1cTucKK5FPxlRo2Up2EjQJbc5jqrMD+fYwS+pybHMXblkGPxbz/YYarL
NBB6v25qLYMsiOLxgEfh/Ml9Ito8lXqytodZlUoX7SlWufverXs8gizgRj0sN3TzJIbIMULiLXpU
iOVA8VPOcKVIT7E7Nn4zu1BKPNN1ZCWDi9E+JxMKJIJpl1zkHOlMD3Wiss8zS/gqVjKY/2ZDrkOm
hdU/4yNkwvlnPEyftArpwykY0ev4zXW9kMxlRTJTIoQ0SVoGve9RC550TJieKqZWyXWoRqXJWSwu
p303ALIlOxELOeFwJ4/hCCNpB+J11/Z73T1vcHs6hgTkoNe2K7juFgl9psgBkWr+Sjf0F3yI3EPE
hlDFPcfLh0grMO/Dd8dLC0g7LUiNrQfbx347NvdY7+ydi0Z31KMvn2U+Q3SeUgCCw0Yeg+Z34f4p
/gU+vVRXzp2exox3FygqowBF5g2OlXUS1Oy5bGRxVIn1JXeq1XNzSo7kWhn8QgnS56HN1LA7nc7l
BuxWJ9+un5QqqnV0L3LUo7XS+tFWfq15LFVlyyWNZRWPt4U3rEKX8A4Ixbp2xjHlqoS6ZiGhYGDz
Kk0blp/1xTyEHEXGfplMYVAt+tqduqMrlWlp/OsYVMbDbMjyiEddk47Uhq6GDCV37jMJj22pon1u
gyLTGcqGJC/4K7UxlErR0znU+hC0nvdTurNTO6IHIfECqRdMzMbvwR5dT6rdvxbIBJAaJMLPK0A+
iIULnK1LZ5OVEUlenZpM9c35JiJgAKvpXTkkvgVDRqCmd0d8s95jpW6fb8g1LgBI005vluuVOgb7
IIL1uX5Z+0H5dEKMRRLGT9+xM+RPDE62+ruOfBFX1FW5OkGJWqsKM6AI/W8fE8tunXBFFEAWZnOm
63ZeXer2pDFEA0jJtTI3+aMGabvdFrVG5qeyvLRSE5ofahn5p4y74KMc/Fu4NAptHnqXGR+0vpHO
O3AERYh2JneWlzcdwN/UAhRQuFTZp1QhaYHgjDE/7Wk1CP5YiTNq/qPZGgiJ9x3z4bs378G/gUCR
ntgdNHsWPOUVYf1PusNucAVXVfUyRgjbFXJsgRdTHY3znYbx9XGmF7Y3IIN2gzvcRFV4ztOI2iHR
7rvWR10P1QdErL0VvewPSnLRHNVMEApFE5U3jJXmZ4rSm+pItR8Yj49/cBmBCvgXqf8vbsg7ZgyP
z//kllLkoCeiKRcpveS/pBmGzdXIz6TmD9DHO0XaWvUVMiMIXoKlDBD09V8I6SuRBBrZPs+FiATA
lt2qnhbEdB9GJQEf8OtjuzMsXGy+ZBlHYjXy5NI7WGohAKJBdL/21nIpvqAuupecIA58Q+5Z00Y6
/yov125psB0UwE2AZ+KAu5xxMPhycmDvaWFIEZNmd9QzrijXS5EH9gJFo6/saMOpDlD3hLa1uhI4
e9wfZ2QGVU6al5El8uQcFILjGwtOaIw1vNvVrCsLc6oxvxqZY3wDaPqiIenXPAXajSwR6fyJHGxY
NwezrIpJG8kEDYXYPCFzrxjy725xRmt/QSNjAwqhfTY7Et8Rr550uFM+dqj/BHrpQS4Q+ZqHdFZ1
Fj99D2KdqcjlqpRhvb0O6ccwOZxKo+EO7Q5rjTe02RzqE4pBJqWwhmDPXWZDlmZaoNnV5xFUDaN0
dcl8u3DPlbAJEZqJCzQaaJi/UugeHd/v26jbTmMomSlqKD4GwO154sQhDzerwWG16aEPEV10xdjQ
iSsc4kuuALmw5r1mqagCynbkplnmYEGhCc6v1t01/Z3ASJ7F5z00xOmSzNXe+CLuHL1vsnsuzTOa
Lgg/1IPcPOxEvr7wBzxk7zA65SGHjEwUK19btqCbVqPoaYH3AWx9Cw90OnCir310LFq9Ox1vzeOE
H/kgWFsMV33jPMP+uDGaDe9cYE69jJImW4wikHK+EMdNDRmY8V0+uYgrd8jInR37kMJL/ul+V1Xn
EKIU04hengYgJDb22bKp5YVzM3eLT8z7HmmEQ9aQWszBqJfZsT6gZ4BmnaLw8tCZudC6aVIxkQY9
qhsTbOJf6vfiIQv0N+Y8RJU5Y3HBdnOCaLq2ExBhZB2ZqgBEYTjKJ58t+d/E315SX3t2SgeyKgvN
WBH35Syfr8LsF/B1YK7212JUco/HXBmw3VvF+EaKzAt2nqFCkKDrclp9tID6Kw8wfLh77c3X4yZd
etTc4OTU4sXuC1IOKyevcKXoKfOqn+sQxgLgAmnwbVj1Rl9xB5npUciXVl/DXlARNl96hk5X8cBw
OcWFnbp8ke3Fozse8rykaQQA72tv/A2L7Zg1OwfCZUiyx5BsQVjhzP0Znm6979xX83SKrI5byf6+
r9jeOyFgaGFYd1aWXpy7ilJDcZij2nkvE5DhIR1aaL3rF1UcOy9blCl1huTDPdtJk7x52be4MWuu
cpGxKlc+2B9OhnrEDCyhtiYqCnYU8hET1Lqbhln8bNZe1OpxFG3pxWWLvJjIYkUTVQSM8nNqDOh1
Z4hShfe7RJmxdEToyiJF7DYm0lx66MEWg3zC/I/3AX62EnwGB/17woC36DZergVVG/yyUOC/QUkh
JCvmu/2fz0Z41dk4gfYEkE/TtsHhAemXPu5/xjjjUabIl924lTuxaerZrr6wCSdCnvrmKUdt0aai
23Y6EmdS+bUBriwKzvPolLNHRlQW6XwUU0loQ5qXBEOt2Fu6yfNnYb8ZyWudePCrbQZLi8sDZkEO
0hZp4FYLlD5ukapjh3TTGCia+7fd6wkJZUA39sqvylfH3B8XqrT2Iklw1o132j86FriziLo+Grp7
3mIFMPcWvd4UA1gR6akEWtoO0C/gOvEqb5Bdx8IuAMWL3x8i7nNL6ZYZUUn1XTZOQWapM7g2bjEb
mZf3W6SSHUUDNMp5QmO/qVoKc4jtL3P39uOg6naHK9KiI+9afTGlHS4B3jzpybj0reLlX8R+aNV/
bcK37julm7+43Iilwpsh2T3EbthNnHtSZK8Mj+4xuQYupoLmS4euW7hCqD2Jy7KWhecgMLu9P5+A
PJz1KqAM9BYudp+ps3T5obZq4bA7QZgq3tEfXN1OibI/6/ce2iMMV/q1JEINk+gZEN8fDJcNBioV
ZmjaNrw6UoLDalPr48BfUt5sQkfZHZBQk/8iATBzOw9IHqSdFRTYEGTiGgUwz7Gz+NXk/tSsLAQO
vwtRb0i3W0aGfFBMnSxyqs05r5Zn60W+AFpMzEpiUt6SWXcAiZQ4bU4Vq7BbjpL78dbshEFXWjSY
p6/jLIm2sFLd8ipNM6VZ1wWFjB/0uL7szFK4hfN09xVpI2Y2gK87PoHfYeZZB9T7dGkzNDnSEg2A
k6t6OW9PYusACdtQNmmGEO/0UuKqneKZ9VIU4yL99S0YylkJ3iYULDOwm0bg79zfSmo1luokrgCg
XiNhn8nJ8ooXD+UtCvtCsHpy/CmE0pSw0oxNthfRXhTQJ2t6Miohb1NWjDdbkh+rpcdzTknjbrle
n3HwVJbw0bLCD3whfI0irg0djZMVC5RHtlc1XBC0o3ZzABYGGfaYl/c6xquZuECCt/OPbUMbAwMl
9g1lOFCjNN019V3o0LxH+9+j6qPX3NqHDr0FkeCVZnBxO7252fJAclYO22XPST7GLGg/5uQ4UVZp
xyj37wTaw/kORy9g315kRNcP3PrgogEVew+qEX18iAALu6h0E2uuUlMVE2XllNYnDMKwsG458Jmh
MIoMt64tcgPCv7f9QJd0qi4Zp8yUq2D/W52cfUPqU3MZLdP0yeUL2aH3R5c8zsM5F2yiBuFjnd1V
GzY3Cz/k5rUvU9jlmNyybueNvckhV8s9a2VDrSR431uFU3E3wkfMy9x4mV6L2A5xq7kaWyUagp9C
+ZhKfwhsQlXkb7c75B45RxtxXu8B+qdzSunxXZcczeolrcFSJbbAINGCUdNgPQOxusPkcFUhQuKp
2MX5xAFYSAIAY0yjlXjbtYOvRvbyh9cq9VYk3ld3Yw3endG4D+k9djo/wrDetXC5TVpQ/+rw9A8b
EXsa7CJSetRAa7TEbMuqnecV3SBxLUHiTRsdrGkEOMHaR+FHimB4g3x0+K3TAh/KGft7aU0Q1Qec
VZ+86RnarcvW+Fgg/Yh6ZLXPL7jhwPtwMJNbUIVhEDYsg//ZjAS1Phe3zRGWKtdU58M3rhReXlPY
aL1/MY0FWJqZmP/0lkwk3EMqUFB4pDNj8N9gfTel9C2JIV9zJm5j+BveFCLUbgJ11ZRyrYU3GcMl
V7A0NPxNmbAZy4o51T2vrFg1iU89KNA2a4Qog4XYmOS3fnu0d6y6Uo3t8Vu8qY0vwE3LZMxBetyJ
OB/IjMfOeRHIj0ze3/QWcQbFFHKMNPQ8VkABVZJBfVyFnMH0VNwXAbFJmnTOwd0yKq3+lBQBj9Og
5ovrTNK6xf5Bu8CpnsIgMttzxmb+LC1iowZ5rihZYq/LpCkwBVukdWpiHaNvlUz9GaBbf/XA75/7
nHK+HVXqv69n6W9y/++nOpztil/dwqQU0KEF9P+dTPSAuLc9GXnNBqasnkvASXRfuMYDRBp53rDk
Aa9akNQKchARHpkpTfQuBYNwn+ET6KWwfUtMvZsW8+rlqhduQYTsan/SWe874HteOy17cH8+KKxs
thnjN5O0JJQoC3ZLfJuyARaDVT6l1jwzGPClgpyxutrA1HbeGv6wDuGX/TsEXWB3Yuc4c+mZufNs
NJdFFmR13TTaBAUXWIoqauDPEFrOjK9FgBoDgbAgnk2O4C8WDIPsXgXMjSxzAqWbx6wJk61Dctgu
wG84b7ge9MJhz/vIACi1VRBIQVaiqcK3HutgoEOKpIlh3DdSOfpFm1R7EPKgrgyd7oqh5zpA6JhT
7kGlGiOMJar1dlfzxh/LIWLVGf95asB8PbhI9nobJA5ez5f5kAI6Ow6C4ejI+kDdNNyaQjRypdgS
vQjpxLYaC+Z/WWx73TjUvmcJd5aiE230kV5EjPgbjpJ7rjf0u2G+bSR/EG5u+HM0wHGWZea25co9
Cx4kyIaO6zOV3qobmw16MUQc/IgbZCjDBFfvaHwmb7lW1i2Z3hoEDl7CK4YYtI0axpKYhnuyQv3v
23H3LldXXOtOma2zx66IPgLmOwgC8rSTumpSi0Bi4bQIUCBsda3MOeygFpKsyvP8mQuXkrvh1UP/
UKh99CWNEcb3xpeDtn0CkJC/2SYAULT3LiXg9GtfI9sfz2ogr/T6xDD8Bo5RraDUfk/m8N1K/ik5
iqCq/A/teTUgmJpXqyxnCGC/s02+zNL2xRRo+J6A0X0qHsH1xxHrg+hQlLANA/igeCWFNKoQDWuX
qpRD98ojSyny33ipNdBLLd/QbJ0ZFQ/q1zIzEHHs40bUZ07gmDYsiAgP1cmQbQldE3JMK+tvU4pb
ffUUqrBLqUyl19A/mEtUi8axGsuhRH8gWMOgymqGbOONMpqsKIoVzvc3QIcntVLMwXyrOhCtoTqm
yMoW/O73AAYoTlOW3Sr82G+8yhouXTsCi2Uj5ES3FODQmBznjtFDqVDRQ66N5X274LCGXEEi5irG
UTsdLLOFOn5Y1bystq/L4gLghofV7lSuoa0Ovpw/c1fJMzYoeSYLyvD7Nr7+EjgmB1j3szk+Ntyo
wIjorgjYIgdWwfVXfWhKV+s6hSAfU43AlomKTNKiGigB9pF/mT9g0NL0StumOdvNSI6fXeI7VFnC
Mudz9pgoPfkOMvpp+BKx4QBsn26Vz2fWmk2WFzw5lHUwyYKtUMcV4njODJ1wKs5hfmBIubA9VpFl
A2D3VUCT7I1y/xdtTdYjs2RsHQ6c3VgXiaT+7a650eoYx/lpDY/4FGFzNg5nBdzdnudXpA8r80Tt
DgZKjHjAiS66OwPoKIySkCRb568vq0ZRtJyEGn2zHoI6UMExMfmlPX8NLjh5F/Ph7ueFcwawReqz
qR3lqA5K7fksztaUIM73X2lzWTdg/Fr19s0pMDa3g/8aMZL2qxKcV20Zr84yfkVO1lQREGQOxTiF
yzVgSqeDupBo3uBW4O6NKUpcQufP31W9leZqPI3gOeXdwOqapXLYH/gVKUujz9HYmIrrgWu0XxkS
2HFgZT55nfa3nhG4PtklQpxGA6m+Tons3uSo7coLArf7psNRSl1ScxH6aOdvy2q2OdB0oHpVbCx3
cb3noUlzyAhX4/MbJsBuygYcg30CVEvRQX9h/iw9gWo2MLhdE0iL9duZxDGsPKowF5xGruoSrUok
G13u7/GmVuhn8+/LZeE4oi0R8uagfP+SfJxgCTEn88xwNfw03Blz6wHz07A71ujAAVqxeEQrALJg
O2nPSjdKw8CmQrcAtZ3+xbC8my9OI9n0TECYn5yEQoemfYGJElOXhWdpC+TurQLccTc/cETkBWU3
Mz459EpLxA+o3gafqdyVNVRQo+ARkGIdinFfD03blfWlM/Kq1c/hE7Txc0hJ2cZ3Nb+Uy/YDMWW3
KJMpNC1B+cb6M7mL0BBuGnOFS0eO9GHnKjUtX8+DI330CIEgVQSCHLDttFCGg014oq49EdYK/Nfz
XXoF5YSzQoC9vXGHNL4VXqUDoqMgrHu5Gd8hBwQ8VhtTTW/PeHM3gU3xsqyQDIkz5LJ3bxfTeKbP
W20ZxNc5qenPPWiF7IEPeSOah8fhhsF3IyELyEtHmcE/hHBsQaY6Po5s6RBxGOABLVNL2lgVjRk6
dQEB0oJhZA0uDQO2hAovB/I0fhfiAupy4mLwVC+cax55rUTqcgNWBch1mxZK2NE3NDjnoo6h5Tor
EJBAtQ5DYwXclbabJGUHoySnEfr1PQX71bQCI7BxJ0okKzwJKOAFNEqSG2yZO9l+JK2ic2a2XdVK
YlkMONK1IJuKQxEj20uGOrk4egL6jkbvTt4hpq9h4i1DB8TjNwCllK88kjc3Xmco+XzbX6xKkIAz
TMr+gT//SoE5OKT16L3GFEUKts+2LpR1uYKHmwzs2fi0APgFvIbyHkf6JmxhYCNNc0V9LHJbj4oI
TAg/TkCQCleBDYgiRcxwA0wY+oOriG/qGBYlIg1zi6hCa9NVb7bMMsypYavjqQjaU50FsEilIFfh
ATja79JKUukRcYpU4sX4+CjrwDHXmfs6Y4k5zhiF69KnF9mluv+kjxvPgE9XInMCM/+WLvDGd3zT
j/NjpCtQCFBMOtNdehErIu337CFcAsVi7KBDRFMwkvntJhREED8hehkY4Or88AZX3uV6nB8A+1fR
D/lg6P4A3VLgNGHsfJ8TRIQ8raIEGUDZGR1b4q5xibbmP8Gd5stElNghp5SU4pL4kXK0L97UaJz2
OtYSGBL9VM13XRfh+P7NVMbn6TqqcIHn5+FiT0YT60PkDLd3oCcpP6YvoULmRh06wc8vZo7nbenN
YxpV+yxhAiMaUPwzY0xMxrREswW3bQ/bKrUd3HllPm4JfxP9vwAdMovOu4HlE8/aKEDI+2EdRDT8
adDB0clZHUmI5JyN72+w3qfufoX+XX+VBIIyZLj9nBmJ56L2jDLTK3/ezMibHRLUUvzUCt2MIVgZ
xYhJVt51Ju4qFcmZ0xM3VxirAqGb8VCQRkKqEQ0UHRicxfblxBbCwmd8MCnAjS1hVQIkXhawFYLJ
dpcaE+LJaRfQXf/OE1Mgw+RsZgTfXUEm0k0LOOIDHRJZDrcmE5pmKzpNBVlwvdx1VSexn88pr6CY
DmXD8GaZKZ2xJA1xvYCM7BuY7ELBDpY9Do15kZWDAZicidAZAs8kkHQQ5Y7btZUPRWpmww2i8U6T
9/ojX2osRFtLdlT71e16i47DmC/QGy0fGAyGRu7yRoqB2C6O2E2wGdij/gAe9x+BztebvXFt+tFu
Ltzs4vCVUCa9HnnUge2uNxHco/UVOdFs6jGJIrLCyfh3mch8/+xkrFSC7QW4lcwA81pFMnPcRUlX
TKA57rOd3bcXA85gqYWTDzjq7pY+xpUcFEMIAknPUYcoGCn14cPj/YcXtjAGGi6jU6eBvha30yvF
DkA3pmt3WN2Z4RKdSRn/QMyEZcUbVuDnupuTjgY4HvSVQQBNX42sqtrHPB7x7y6viHfbvOx7RtgA
cA4Xqt0+zrpeLTm+bwFidXQt9BumxZD8bXBwl04s83HdSTFhcV8l3XFsuQm/+Da0s5BiG9WERyNW
NlJEFylXzAIeXYtJzIYVA/wf6/oCul8UNrMJHFb3kOKGcl4Nl3WI5GVWaJXB8ZIeGVNWsXWSxOll
Y3ifnDZbXBDm2c+CeZYt0gsoMyQ5MHhmiTkYE+yoCIrvnR5nWLd8nOnApdmOgsuyUeISgLJIpSzG
HZjf3Cz6YlItWcoxQzPbEBOXFBONDSuoV6CKl0/gWFcVpqUKR+fWkBlrP5Dbs/h+ZTnyAcZ1+cb8
KqII1/vrcHNwC3hqpWQMuNEa2G3qmsQKIFmSHt5ufteNrubAknaBV5Uw6viNloN2L7Uszczuyage
ezftTm7Fi26aBGCeS3PTyLb9icLKpGcloSFIomVdVinHcfmrk5z89tU1MrwCELfPFA7FDxTRHuXV
EfZMCNfUGhObFZQPLAUeWpyZxCmLimFSrGFDs2BCkAoCMLsxSVyrSNQi/LMDbDZ/VwzPPnleT2zp
x522QvZOwfbvQ6zV4lbgys2s/YvLHVRHgHBdZWp6TZ+YdbD6EkOqizyBc4okB+lFBiWSIn+WJ3XV
/msQ3mhx3GDK1dodSVXBHF8vd9Zrr8obXQk4gNVZJXM+kXDMyjZ5ZjJvwml0qJOns11ClOTyEPF3
gzSPny/PqEYon4iSB3YqMZQKM8tUmwx4ksw6YsjdSgzGYVvdfsX9UAuVDVIazaeCBgKEGPkG0SZb
yVg1y7EU9V238zkqDrgf5POFeaAR8XxQRyUJQrNRJwwsids7pcqCHgeUJBLHbZDCpjf6IG4MCtrH
J88vqBhxnAcaO2JdAYad9+QifHGGnrKSn6eUVBq5hc11RqxxYVpbmBfC64Fwx1wTEzVHTw1w2gXG
dXfq9BkgGPWooKLHKcH7tebToZRy6wv/7zOP0/25kOwS5ULsA7LeGm/HcZGnCkW594p4cLmplEUL
GBiEoWE0UBLPmAYvUBtwKuMLhOIqubqdGVcwWyhDdRzF1yE7zJQ4JjBsVk+4D+6NGQc3ruwN5YGR
hokkCeCUhYcMA8ZJsCJHCo/Mnz72WYMZMGdawvCiHX5S0GZRx5PLqMAqHDFU0I7xiklEtxd19D8b
P7u6cgoxAyEypzhuww2wMPwjzoxOyOr1GULKzoS/zxeNszhk5dE+3/7VrcURV3H/PYL6CGbAldTT
yXx1tEGHf3RsP3rCY5thHeDKUyTIRulmGc6U3lY1wc6M27TQd2Azm6nZhYMk0HeDks5EUDN5y7vi
AN1kopy29PcXThVrGhbv9QXq6K6ocJM/n5DpFETWn4cfyCNGajCJ25B4JnCdtF8KdF0WiM9aO4Hx
LO2em00NlF0aYswF6gPQR0VKDY9Q8aRG8wNa1b62t6zBBpSUtwpJG2BXUkhNhf2hGJwmcsFgdrHy
LnysP/3VJCbqy+JhsphNPhBeGTlArlXnNyewyFR7K9u5jYOT+yyebkJM7grJg17lnM4RrFd038Sm
Y4ZHZZMBmoXo/Kr+wzY9DQLMtO8hx65jk6EamFgSjPReAvGy9YV516kAQwk2+FGqrOOh0RE8FtJU
L1cTO4hdmFKBovhuJk6fAMJGBLIG7ilfGwJFM4++33dJlQ83wSPmVzcc/GkPIcmJ+z617cZ+bamU
UBlY/7VvN1NzywaXCJFFnPXBIwUaS+u9vzKYZTqdlxplBrT/VrlZVW1PtaarkHcI9l86DL3gEqQx
Fb2PTOZa8EmLjg+AkwsQMQ9FbiiPZT6Sahheo9qsKrY2zvY3iDRCDz95Z2iBcoSe7AeLcFHR4Z+P
j3eE8jBoFUkSxUK860rXDzXngLPBPQk+iLqUDNfof0X3kEZGyp5twB8uxbM+UCf9T4EkIkP7BNUu
5t0eMz9aQ+/XHo1oY37tAGSuNMuUz12ZbNOcFf4dAaSjJAFi8kiEi5bLKRU424KYpuecwJ4wEqKf
TM/42G58LsE8mPhZkZPar43s7GoPyiF8qdidcKhjr+6kogu3ULO4OIRl6MXK+EmUyYNGdosW5YKb
MAKCoE8e2/BlX7kXtjoQhlhqESe7fXrazi62C+xVxZR1/VHBwBVFoRNhxQcyerDzDEgg4e8CB3ss
PmZKQcdWH3JBBoNuJI9Rw5YGUutEZ7Gss+ESIB7Ebr3PutfgO8B+jFA2S/j/lGNEwauF3b7KtL0D
VHsMV9UIz9CmhvMEv+221ezHJTX6/yatoI6ssJrqHZldisygnVG8lxkD34GYkjVTWMRj5mmmqcFl
p2Q3Ayqeth20fA53GWvA+lMOnW+PwP6cR2PjZzAhJEFh3gk+Z7A2r9dx5vOYNdNU0mKraPR3Kob0
PN1Bns74tUWE7qUctlN1s9LQKqTf58ViNZXxWbzMG97pFJglxPiq4JF5HXHYLtQZFAqjko5SgDGK
UxagueSlLHVD2D3CkHVQwS0hgABPnflPWf/+i9MWVnWsHpo7o9RRe/Q0TtQA/ZLLo19uSQvi6Pwz
Avs7r9w421gY/90tv7b/nnR9Cp0pcUYvaJAQ5ficcbehs4Oqpk5GggUeC3V1Lhy2SVKCHPTIqzS1
Obik57IfswpIDSKXeRvDAjRPWFaUIlCCbrZh9KwmsxGgvDZCL8ALCwjr+Bm9DuEFWgNVNg2iodHb
1HBy5F8vvwxBGBzBLfGr9KPpT6Eh6jpTzCsFzKaPCuiXeM/htzNCa6/DYOy55+w9EwxaX/3cEHug
Si7yipspL0H8mlnq3n3mxK3zys4yNxzYwWtPI4oFcF9Bnl911/mUVY3ieKCzeC4Co8xRu39xioju
s/hTDJKZrTtvZxorrWlHQ0PNi8Z7XCmOUS7WfbYXR1RjiqIc3IUTq74fQmFpIIX2R6QTTbbm2NS0
APklwIYE/ZHHvF8L6Vw5Fw+KuMeIeWZKrSZZjpXDFptAnnbUBISXSmD4VIrAUAdRbSwxucNLb/5P
Mslv1nW8FNitTuiJ0cUQcDhYk2YIDiFZb0iKiTp6ezU16ZHH70SIWmCoAPhapnoHRf+VSO9i81yL
+828nhfu7wU0N5Ghp6jJaApri+YfVArwxGmnHy0b/QEWq1a6BUn/aWuNYSbJET4U+8Lb24Y4NcbJ
NLmfhpROYogFWtnLelVmDgGQct6nCfFEcpnL2bJ+5JcrZssyToU88XM+uw7qB6ANOkOXB1iYBmCJ
jnyZygg57wHxphsIfJCxxY2RXxnUJnNu0pOWufy0WnPLwpPP6NkKwbTulaNtDHnPSrBnxsMLaBX3
FNmt9iEJXJDuQcRRennkn/LKy4/7sYylAuhZFXR+ULROlD36YuUsWE64lnKTZJh0I2cXpZGIRZFZ
7GqXfAWyG87qNNF/2usGGe2V5tEVg2WAKzxY11JiD5GWzXr6SZoYxdJuBkzN5+cxRmeSznDl+7D4
ehHfuD/bRUgYNlVTRjG9/yW8aA404xG5RjzKJVXR44qDzzYzPLlbMV5IGLwAANyB1DD87cG14mxV
c2aQUOp+juEln6M4qbjBZtcoBcGQ/jPqRLfRhvLJEFYDjhGdszLy8e++WSRVyeM2LcQ6jHL9FgM1
wvkhB+GeD9kwY7eNWm7N2RVfb0ch4e3ZtrXHTob7foEupqNP3VmbwU4bPzB1/0d9BRiomaBf7ftJ
JQu41OJW2AH9hzu7vhVzkaHS6H1qO3JCltUA7jDIQDO1wguGPY2rKLIKNfr3hmXTmdrDVDNMfIfl
Qzn+ttbnk0gBOZUyd+Uik1/HG2D+jXqMccFjWAOwBgw4zNF5w8ObSbTsXurMRUbVxeHGTRoe6Wjr
mMrc1Ex05gc2qBa40tbDXUg0h4O3lrxcHX8dx9qe7UzfzFNscIwJ+NeAtHltyw3w2POZCoMOz2K4
qgdeg4ZVJQ/QhlTQl84zcEOwArf5ttbQ0/fQw7Vqh5T0vvir8qd+9mFckL3Vqdi3seAhF00r5gSE
8TqYTNNsJWpXqi5vLu3k14x8eRVBu862pYTiGiaonwyAfUp0g8P3eIlWjnAdnHdEnTl3N284gH45
i78ky+cW4QLiGSzqmYW0SU+UQrN3lzKxcrE/e7qy/G7KTtU+IPwAwdX4XGRCs2XQDEcqCPHt02RR
kzFhMkq5j+mU5eMLMo6QdouDWFYmbEdm0pmFTIq1v60ZB6BhuHM1+Af8moYeBNCMsfvMkpnKNBbh
BEYKSUnwvOXwPXf5I0L6xstj9BhS+0Jz2nMdMdntMXNpiJ9pErzJ4nsL/MHhtLutuzBP7EmUPkN8
C4U7YCt8KvRnldaNNImiNUTxaYGFUDus4/4hGfmDJg4d4U6Tfx03gvYrtwnapYp36n0NuVxxhwZp
CpihGG3Gapkoag8XLMewFScTSCOIFQG/jNevplY2LMRD7CoEuqWzWb8jdIaxPI49PC3++gMmqbnq
/xCBOD2agmVaGsDF2JW4ijDFfnvuQoRonGhb2xGMCthxcmsultLi998MhF+XyY7v4jJURzki+LaE
fVtInt/VA2odqmI20dbSa6T49Sxt1KReu3OTJeRxSp5Tu3ZDkcEkDJDRak438wmvh0Osg6I/iE5Q
3QzJPahHfcCLg/GERjNctO1T1+867ylTZ5FdVFd41j79eZg5Of7/cMl+GFN/a2UMcI40ZcA1tvSH
qjDQKXWHihNEU/LCb57QliIHR+3jTifAQ6MhY2kYcMjyZe0EL5JfZehpxBnp7O9C705LJx3VjUuS
YfSEw4mDY1iJc9WgqZLj6TM+3obmf8PYJDmthS4/mNBHcHViGwVGJ24idHQtSGNcXQqd2wNl2FAk
GOiZgQOTiGx5MlBlPATQnZ3eupPDr+9kX2oGn68YJ6AJWxY2E5THe/dZ8dQqWxKj9H+9KpmPZWIH
v167hH1iYpp1vzT988Hk6jQYQnxv7IUii79NzTm0mMl8Dwwb0yWfytL/sR2db2a+5nACWXxCu0aF
s9hAPRRiRFE3wpusBROMoUF0sFlvPON4bAshbylrpoedOCZVZhV2MvjrJaTuuHF+cPKAltXp6a4A
VSnP36mFO0oDfMQoBPdySe2Qq7sP1U8ohUUkcgNmLhTVt5hHtVXkEmPBk78EUYfexcfjk1QjvXOf
YIyQsd+TgmTap6SPZXEIoknGw/IPIGlCEbCPIAtYza4LzmCZUNe9CODr92u+TKilb4itQ4aJbWVT
7j5NtZl2o2FR9T1yToHnFG2NxyCNeVDIi+qvHRyH4egGaUW5jna089TIORRcGwfoEmySpxPhD+gs
aKkaV7BPrFA4kLM/2XeytGtk1Xl3IcoN+E55Pt/AiotkAtFEA+pNsmyCzT1O0Ti9t1o9+mQMgAEr
aZ5B/8eVICFH6NM/iYZOa4yCTjHcq5WCps4zWSC+gzNXgaH4A6gyq3oSXBAmPl7TKJ9ju/Jx8fVF
NIhKAfYkXCsc10f7LPoS32b8uId3ak816pqR9Mh8dw8KotiVSQX4YJthktKVuXbBgl3K9FssnZ/s
Rdhv5b4KiVJx0hMbCrGrrI+w5TxyDQ4eyoO7OKc4UcPhVqvPwn7rhVTnD8bE7esS+8WdQHutvdL4
NHSOSYVDJcMJ+X0wYOFKbRqLaUDIxUhsqREV42hAPmDz2tAuD+5PvXpC2vUheMZsCey+7upCb7X0
MIaqJzNuRUUj+pBjZipsSOSmekk8QIlSLEvl4d1c93L2BS7TTP8B/r/zIyjmHkaG9G2oBDVyiVfR
0cNBbA4xD8chE+b2KGBdD/GmdjJTcoLxf/mSgXgHezCbLBRV/glvJeXtJayeZ0n7HkykCQhYphGQ
QBrSVEe0PB90AHP1UxFykvXGmDRjc2q7K01PFeptXyXqs4pyzVCPCGfRsAyacsp/V8V7PzPIqBlx
+UEc1USokVphZkCZ4KtOZ9YxyhgDmmkk4qvLAcO77EAA31+S7+etf/XDSryUF1qeAO9GDhJkEnL3
ROyfai5w1cFdWGdQPdAxaEC2IpqG2Q0JDeUpGA7F0jsHr7F+lqckcJPcPUiqWIrdegx54L+U+cUo
sWGsKrU0o2hUak+UadQ0shWSaf1PYA7fo96Mov8AUKJ2FE/UPT9/E6srIMuPT+0iA5uSRpW9qjaw
NxsA/OQ0PiZjitjDNLesae5LKOrsu4m2RXIw5Lua3t5sIiHHF5XCLqYX7VFJz6fvwgke6S2zLYNU
lIC7PU1zhzhoJ83OaPU2/TBJfxjQ4yE8P1WrBzIOyDp63pdMVvykE0XjXajCi3MCKY/REi5Z5147
OalGYiFs6kmRVm54DDtFoEriqkyBsR4F6mAabHfosaJ1BQCm0JKPpTI7axr3+Ebu1pUIqrxrcuiB
Jtm3odXtjLpmtfvYdKHL9DAfx1U0h3QiZCIH7NfG/DIVJKB0AXAcNm+EbtGgtWfVBMUBnQmPw7SB
CbeJ1adlxHxDx7fjkYT+kdoSdfs4M8iCLzJkp+IlQr1owl4SO0nCtZ6ypGdyFVJNR+Zzfv4z6Qk6
YVl1APw6Swn5V4sZgokWW+dy5PQT0EY3x2kQhwI20FpZEbXT7Va5hDHbqIseNDzHCqhMWFYqcrXt
MVDW2WQmUR/7BWggmbiHANfgwuUIFPsOgvI134zOgXx0iJ4v8orE6E3cb4Vb0jVLPBCgnBSHHuFK
sG2V4XDHOPPFbNNO9vF04b9r8a0nxumoYCk13+CzxBHQe9DW0D1GjPnCAg6pLC2wO/MTF703dof9
8mx4gPL3JNbb4UntqOlBCPztFCZqHO/Sc8TuvuL+JaxvbINd9UTCfnoN6B2IVgWVNnn165haJqt/
2ziYElE5F8XZWaYhk5j6kG4D9h/mjTcwfVVwClKyFUMZXH70EIfAKkwaRT0E/fuBZUECi7eW4nmT
Lz7EzAQ8fWGQ8bPen0h13NR1st9kYGOR1cR6ac50WqfaqE01gVSvVMGAMp+Q8nIa3GonMMqHfACK
61GKPniKhOD5AEhtTRNJz4S6d2Ofwk42RL6LcTL1pVaYZK+HZB+A3cwzZVIy/Mh77zelrnlfOGnn
BsgcFzDhuRUBsOXgYAcpAgIQ8L+GP8LgwvKjXdrImNzpJPjfeFEElM2pmM99AMyID/gEVKJen25h
ZouMtZz1g+KrYFAPk8nFExEfM1m3YK9jc1U/h7WU1geDMt6F4GY5frlwyMvISEpA3f5joxiYuHqT
Y5p96MPN2/je0TKTEcKjCQe6iTdyH3wEDvxxzx+tTNWFDb1A7Arkpw3rBJVM2QH7WLYZwN1LpmAF
1zsqj6GWMYAnowF9PZeo+VXwC+I+3MQ0Y9lSfJMfhFu0+eosu5txA07O1mKqq+/yljnFGLjGQmg/
PhShLVCT1pXyDH+G1baxNutyP9gCU8orWtskTF+cgFVP6vHQudmMkX2PRnPM+MDK73i4hbqj5Koi
gpGgC6k5xEPznaR1GQ+6OWx6v85SVbs1gK1dbrJqZqppFESDUvNJxBUp0O60IY/D3Y5ecredoSgP
Nfg0CyR1TJozWAqU20c+bS8N3qP8KgKbTH3ToWXBZ+4La12XPPRwpjWiBwfHP9J8uym2fdJHeYEx
vEkahR1IAi/B22AEbD7s7EXuEs9J0ZEW5H7CBM7e1WyJtgF0hDRORkkdAhQcaDnxTYvEx6oIZuM7
DTumT0MQ+PDZEZezJuGaRFYdJKRQJahGI/8JDs2xHV9lhAlZh7zR8gS+yvBupDph1Rf90MmwyzCy
Gc2dVInM3K02dbFIW6XzzmZkhG3vsRzaY8Bvj+4axuJzM4sQAY9UQRtvkrP50UynTTNumGdATYRM
HTwyiEKgTEK4TYRllstOHbhNbXs2eHZqgZr4tYRwgUjwtLbOtodJeHN/ZDZyjxumbnft6XHLORHL
857n+sLjVWrcsZyiTf7e0cYuYxBKTeSnjfvQROnZx44o5Q1RrrCEhNNFH0E6+iK5kGQzywA8An5/
Q5Hu5tYKRm6wqGWugJEfQRKGXnluf3f+b+GqAnl6N8XeGgkXa0kKeVhH8AyPFDKLVxL6QgMKa3Tr
0Fwz5V2svKB2dFToTBstYFA0wukVbjQCvu8n8b0gqx+chy+nPD/Lphbq7xIyPqZU/qvlBgl9XaXm
M/N337kx6vAxW7HoxTcRALWfyt0tIlhsI2AYSMNCtEUbi4LHE7iixw6LZkAcjcUQeTYScuAQ65as
Gtj5POZfAZXnwTPNEvVdc9MRPwKq8LaL1gp5RHd3VGPqMeVCCUhWmE10j6p7i60qAeRixr5w8Gyc
n7gNpyA+oN72C8ZpVBja856GaYy9mnV5Nxd8OCpdvOeKbp8W2LJopEn8MUf5R7WBqcOfdH0WdlCf
Ugq9vn1SqrjuNfBb+aPBj+yad6Wvk0Wh5/TBjP8hl31qFKj59jvkLwJvJmoBivFT0lI8+sGFnb9/
GLL3AdkCb87kSCQZQlgKHeGXeh5D+QvaX2ZLiqLEL/7lyZLzY5qf2bJToG0ATJ5T3hDpvP/sJ7bp
dd93bF8YnslRxh1Gw0q1WrBJpcgZv0rqUOTyzSV7DSehg5tNjMwcDQxR5ugzFd7x5CWVpRB4Pe6z
7ucudR/mY++HdsBk0kl4CMc6m5yJ4lOC/W3s84a3+Xp4vLm/hOxGY6CwtcKMjTfWPuag2NaN/oQW
I6G5TPFKEjsKyPlNM5AifSDqCxed9sH+RTqfWM3YhQ9eBwiwVZDnWQ/hxqGGrVD0vVWlcFwxzaYQ
hvF+hxA8Ot3puNLCzzmPpIrfFmnAUpHlo64tU9FvtEXa7IL4oGqyeBxjxTI/C5bMSyH+C5G1oFV6
QdGblSIzVcNOW5bCSPmJ2nsgJBL1nYd/H7uKxBbtz9xVP6zPG4XDoWYq4+0auW6b2jyj5JgXgSDp
Fqnw/uEquY6ze5EqnWx5KxbAJxzJjMTiKbY6wouoUPE1X6BDBGSoFVUumybn42rQZPU+kLIlG62T
FcyXho2A9R5eZCz2js+eOiOpFp3UbBuToJiVzEZUZ5jmJbvGmE4VYdt6TgHEcKnVhoI1NAHDNBxe
UT5dDtITwpqhY1hSzJoQkIBCvnZAHgGJFGVVTuXsX9uzzq+QXuBD7CZnrWyoU1nyjB9GSwBQf51S
bHFuEMzBy78vBqDb+X55NJDdoLN2vKZlZZSLU9UGTVJ8OkEOD3gfu0UAsYRaWpYVqTIzxMayot3b
xgD8Ibip4JN/oeeYm3lCqYHJy3YcYWgn8PerSAXxH69YBzg64tIqngxNeLj3HKzie1GOg0tXwPY2
kwi1q2SgB7httJR+cpa4YwqWfs+4JvN7q40fgL36fHE3u3NLeAnqwFnnwBfQdOgtnUf5WV6jMmhJ
P5oBNNtpMuHePT5Ok+foAFs5/zAwx6en1CNhAsheqBDpgboiPEUJbXnN4PCOlBiJp/Ei1nn6OLFl
la9qm1xfRg38bAnE6cHoHce8AP6X9HEYl/q9kJJUACdWlnWq1+JzFIEblYhgp9x+dC3so3++Hmeo
756jBGmzqoBOjWqLAH32hezU1nBeKYjMVNBDz3W9hfIMH6QRxAJHSwl6FwjZ2RFOEZqf9Ov4Oekz
3DldtpwpBCQ80hdDCg652Nu2yUx5C47Pdlw4tt6BNK9Swyg8DorIPSPy9C2JaVu1mDbvwgBkMYmE
Y9p2Xh1wDa5VNRsXyWwhF354V2cLZJWNfGiSMWjU3AFTfdeE5JR4ji5rTm/2UdjgH5KK/5zhGw4Y
67BsBhhAUyt0a+RWdDy4GMGtJTcap9zarRK85z/jYfJhLrhR8agx2Q3phcV9FaDhhzX7zQiyQ070
8LXGyhIvk8+d69k5sXgAz7St1O9b8tZ2+j4mTOv77w5345B2N0tZC0TkWV//Qrvcz1LWZDeP8G6I
oC4eG4O/uiSRotqE6MqvBPhNDHxB34bP8JufhpNNxH+X2LQ2VYZ+XVIawCqn+8xStscKOZAja6b6
N2/lQ8X7TIWqONzyr/w8KWxEVO7Yq9pmIi8juBTcUEnudp2eU2L8pH6h6ehWf5ozbjlDDbse78/9
Ij0sj4EdFuAPKzL43lHAF+AI0Rmqrkv8lvoF4PcweT0Ufq2lRV93NV3V85WmihT2rH8N2RpT4uJN
tTQrcuRa0EzcYKaHh+KhAXQ83wJfbvnYiP5Tf0ElBSeS+gKTzeH+W3BMURWZ59iCSvcGOUqwr+tV
PJcuUspAQ6xU4SbN9yg8v0uJrLd8ThkD4Nc5Z6vd2YeUx66oJ+HH9m1Nl5ZdlLt9m19teaCepbXu
UivJRvCr3ZN5EJSU53yZUFfGQouBpGr4P5FZILV/WRNt27BNPKZfoXufAz6JjSyyknL4YPRfbLuq
I1KY/OXXNRMn/XLUVzyEaHaDR6Ez6IPyMBSC/B6kHdJyiF+n1oXJ41E+WGHbxgMYKPAGCanUpJSN
ojr4pQzkhqN6P/ISFdrZoMse/lh19A/TKs+wHe39npkg9a7aglArzn/sUEcThhp9tF6Fh2IPUUL+
HuTvShwRhM8lDLPk2RumVO8ntOClnnirxCtP1dA2R7TKqYpNs5oyXQqCIesWENkZHC6XxkoTr1YV
60cTUL0OCApeKg3D5TMp7NGZTvkRAqg14D05F3VqW1k6p9wG0mt86InLJMdTGmUMHslF4uYoObs9
3fSaDsUODX2nhoTk0/N0HdWiqppYP25q4azAEOttoBO738kLJanWFy+ka7Q30oJAmaBYigFJzWAn
LtXvUK1dL7h6gUdTcH77EbeAdlSyUjWDS8ycIi+0YrlGwGa+VbuCQN4MHFSlF9vduDdZ16rH2IJi
ZVSmp8ZicmemtAd001NJKCOKTeazHHdYP9xnMesTHuOWBeUzfnRyP9VIYnqWZGbqjsCDdl5xnOW4
NIntPv0waRXU22uLdErZw8MDDrTqMnYWdjjcRYpcIMiblOuiOrZFxYdRVU1UPcaHDSCN+gmLxl9k
vZRlm5HKC5x4dfdPoh4xl0aWUwsEboQpfOjOYbPEt0THHExCHg5n4gycICyGrBI1zN+jij5G4cCY
xN1LoGL5+A3h1w6fK2OycaDr0kRYNrBzOI5n6pUCfSiuKVOfCaXKwUkJcRmhSVfhW5315hSH6feC
avd9PyJ6TNgbLweLBHvOqZFAF2/OAKWPn+5NeCRcxmxHk85mozYbiw2tWCKdWjfqnR8wkP25CX3L
iRdPNcHqkuoBCLd0BQRptHTqzDPij6q44Y4QVcIeT+y50dsyjdSnndVKZ5BA79f/MpUApjemUj3+
GBvwQEgakymkKr8UN+gFFNE3s0ZO66yBbSsWbiMppo8eB5ciSCnC5z199AX2pDOXxsedfExHI47G
bwB6Wm0mOtScnIIkitPx4bDbKfmXzS5QYaLdPZE7GedDpxINVIhoJEuI8aZYS61CxAvAjrXMkN6t
9JheDEcloJTj25Zun432/5PPPAg/5BuriYQ5YLa/VbGEcssS1/2fSCvheZ/IOKlWO7UmRYGibOaJ
Qec84IQIRRs3nyx7SpzuEkd83j/V86FDwFdRKGrcZ204Z4CcxSuInxPMrXtrfzeDwhDSWgReyW9B
aNM3XwzqEToe9NTUMoknYHGFsNcvXDBdEzokVHw585W00xV9EYj5M7t2ENOyh02Y2+QthXyr0G51
6U9TryiF27BRV0CpPUp94zBG2KmC3qUTJJzKsqMNFjrq78ycNsioz0WNedBW2/4WHBMMP1fgRwX2
7B4WxLXphFhTC4Vb5wfTGCEHqEG90saGxLAa8Dj4MiVk7ZYh6SD2GJr+gK7kKe4x4lDBhE20oHQs
dbsRKK69EfPdQJD9We8l5wY4dLPZEJVIJdRpOWlZuSK46pMhkkva13jWc06aNJ26ngjY7ItwfIX4
/Z6EBd1ExSLzn41yf9PuYhYaNduk280iBVGUsbd3Q8JLKYgA4vTYdCnGqdcDerYVyY+Zgv2ro45X
Zzmf7xLzklsgQzEfoQqd2ahusfoyHdpsqV/Mk45GzHgu7QVkHOJ6rkhGe/gFn+z3G4xHslzbxqZu
JBA+6x0tpRs+feu3oOKrsFaDS9zR0GcaxxV6Oau5J3JBDM9+VoHcAQN06rwaHrvm4NkWEsGtoLPS
3xNKjDjCEtJ5UZOqObI5WxavLle9/XcPrxid1MQ9duh1sxxHOIyV/iaxR1QZ7WSgwooGqTQfZFqM
uxaOV9iCojVdVpxxqyEZ5fImI6SozlXvxkjZbTJj+091FN5h91pkAU8bBED2B/axoXc37UnXFOcS
Ig8NIrTNFl8Noj33k3mxbe5XnUT9MF6MrGOuEpkwwL4GS2bSsIB9PYmCWIFSL8QItELNlv1GJznR
PYDTSrwAbp+F9ccHZuXtS8tndQRkuH+i3Ibvn+bu5LUSoZmP1oTpnCNufVwyHGyX27W4sYiyOqPY
RbGbYLBwKH/Xzll+E14HQiGUzEW2KgmZ3t0rfF8aE+rY6Vmv0/slU3/aAPVkOIQ6TcBJLkNRXP97
pKC8WAnITgynmUZE3E2lzsKQ27Q5XoR5Fc3KSFFZI2r7cgX3sl9ipHMon53YRvsFhQ6x5aMRwBhu
NyriSNlvE9ehG78rK97Q50zzdVS03HaAQlP0HZNgQzlbAnCSnbeu8J3biddA6Zy3N4UlPKRZIcGc
V/mQUoSE/Qr06Q8FJ+AKZAgZDIlcsgPsrwzziZSiEgQm7eb+n871XueDiewPNOACKHDI7ADBuI9/
F2+niTAbCqUI+HbNKeyB5iPMa88mN1LgnlLQOzX6LrYW7DbYOLq2Y04BuoNVLve1TrcdcQo9CSJv
8kjRo5qukUOiqQ06XVuH8sBHm/Vty0QhwMI8ZAaJPnPo5hWWwVHTYuL+0seG/7V3Iwn3DbkKGU7N
g6/h1KJpwffN1SoBoAdLkLXYcIv99sDwvviPfEqQdIObBsdI7rHSBDzrNfOu/+oncfHrBAigW2GC
j5R36hMuAf2d4KuYy83dqNDVc83rrJu5ySBB/YgP5VHJw1wSAfpdMR5T3UPPpzPgdSCNwnwoP5Nc
xD80CS5WtehvCGxxviJrCPg08RZR5KxfHb+nvp1+7ut1/pCMhw1iiCWiZGJeUQQS6zsWiA7ka55E
H0GK1rLHJ8WKua+JHEeKMeJrRV52H4SjjT049xIyET82xz4F8vJdvo+DYuT+UCkEivVLPTYMiyin
93U9SeBTWBQcJQ6vVrimWCb44ou+XUZ1nFcPao2Vex+N36UrvzMzAZv6GNe26mMv32v9/GCoE5a7
3bOLNzhanzagcPJaoy2MHPuyMwEN5o3F0eQ8yEClPv/Ls8RO5UVn4ABIDVJXh7Sq0mfUtmyeAdaT
0lrTsnXuSq032Bm6AzpCUZVf41lMIdcBQZrle8JDCG1/pVdY53vfT5mUgEkLI7gugwZgCA2I67aS
Wsu/TSjTP569SoMm7p2oBKQKQ7hNEBHiJIOjmx5Xb5RvEQ1dIEBgXSfn/1wa1Bgizk+vCX3LxUB9
rNwF+sU13GHnq+tlh6qsJZaV5XA2CMCfyPbRUmBwFkzj4cUEWXyNtzE6uhtB41O5eAN5k0vdCoCc
UCxICYl3xDaxeXDTZImYxQQT9wuwdX5KDF3MdXdOhlRNdjQxjQ6K3Pza9f6bx9AsWRXUZYI2p7sO
K405kCgy4qXwvqqxKiiS3rI9pN+9y1ZY47RyAP2v5a3shoZhW2uWqs6R4IyECHrARZ+ZOo+ErK5/
3HHJ+MHswZMNjQgxImWJgIbzAhrJVyPI9Cy1LBC9//qliH0NclRmvKU9VHiB/BOaCS8amwnEl6fO
9ACphR4tUsme1Y/mRWRlcbyVhhhpPpW8SgbEfeDtMYqKwIzrnHnhzdz8UGuA+TVf9UcvTbgqhPr3
P4YQc1Nx6P7gvY9CxYRdQY+VdzHcT+ZCO4isSbYcfWbYcV4IYnyyd3oXhpinJ/2hlsWSNpf3mJB5
TWMA6p3fBKg81BI0Ft2Msh/QXXxCRyRrmwDsBMMEbwepOF2ewWNVlUCkgIrXH2Fh3zFyCzS2ymCV
LHI2fhnM/3/mUfKnPH2HWyNCb1zqYpIvsR0Q9qWG5ABWE4RDYDWkjCnSrMMVgBvlYhQCF12Ff5DR
TZlzeeQdEooyil54oLWnNxEOBZLQD7l6ZazvrmxlLhOPFrsYfrX2jBjDyL8g+1VRf1Hc/4nbD5zE
VKc6CguYl+SUbjQxVk5/wUIu+UULo7fqhCq5TE4aU9VZXfAdhfwZdwymGy/Y3zFs+AgxYZDabyut
CZpm7EiA76tj/vcZo3/xtNri9OY7jIYUXQqSiqfBjgs7euu/xkYgIiU/TVPsRP4c2TmMdVAm7rgJ
GpdOP4UwwtW/JcssaV66KCbL+lafmZ/mHu94Fc08xiXOTZdVJCK7ShjmAb9BXXZYVwVWTdWbB4KI
ZROzYfPGVLQ3mt1eBNdUwnwhYRRObgUHbrxiKSsADIsN+xPqg6qa1dE5RX06aYe52wHB6o026AEL
FEVb8i4M/QKriYP5t/NZDnIIKaVsLt+1roCcpQOZV47u3/o8FyWDn+k5tklqzBKlrEvcsD2Jg5DW
5eN5B7XNhTWiu3TEAQx8q8sqQf9IyOyKz5wbn2nY+ggFFA7ggofxRuG5Hfe5qEO9oiFgykrmdkul
JPyl4/HNVMrqAcIlctHK52Zbt2T0lRo6DuyYbwo32TtPy6+oLyJt+2izF6TNSUTiczTIdBJHcXRd
xzns7ZyeEt5cAg9zg2GaUMhPJ/gqFaR+Mi7Qb6DecK/UXvPD8MBpnibqMubIIrhXzLBnmVlxIrHb
80NIrDLrC2zKumlJ60g+yzQR31/Rs/1rGs2/9SzrL6oG2Ze7upNMBLbBwXabGqnr1XqM7bRCH/rz
RJIZiXjshTgPxWAfpDPj/BoLWtKlb8CeKsrQEX7qpqMkwpofYtMisJCAOHY2rx3Z0LES26eWZ30Z
pyxQtyJOPJNrlETuyUILXu+vTVRrYWB8ygZu/Ht4Sh/ej6F7fzMjMTa5cuBR79IxZmeipRLlMuCU
ToPvPkCoh06kQj9z859jQbjpjbW5a2CJiqqwYkIZpavWovvGNrboVsWRahjqSYbpmumidQzXlCYp
Dxsl7naT30qacPN8O/p24mwkBeBWO/E75/+rodc5632BKfD+20iObm7o4TZ+hUGe8Ns44a91xf/h
ZoyNHkLPoYyg6EZwlP94nxi+GGS8SnFC4W6TXg1FMO0xzLOECmmS4Uq4H1Jptrs0CrumQ1AT9iK8
lpeOBG4wByZE8JoEAir7fFmw0c0p+shDC+KsPrrp4J2gzXtiHMMrPnFXjSqZQMHk6Rwb3iK95OWX
2lL3gr5F1FIPV9HHf6PvmohGfKHCNSmDO1gkPBaCNpOW7goQcTbahaCtfOR+3B/5HpUUu0BgXQSF
VBv+LGrrPpCy4xoblRvrz4+cknB/BPk7PG5aBG4UVnH8XYblqePcTfdUQpP2amSyo8ZFK33LyLrU
dvCD2Qi1gXJ4gAiNZZ+vxdoF5ZfaVXCIR+NQyN/9A7aZnEJ+kjvn/6YRTt7XG/xD2ZSXzBl9XNxw
cqPzAbGamsBldvMRSQuZqtoYOTYtrGDioa3n9XvxEkDb/xf6yoshdQyRW57VmLrdIbXwbyNiATiG
dKZKDi82FkWmEwar8++5PDeWekqCA+lMohjE7zo01rcrywERSc7z1dV+2+oGEjPlc/D0Ha/MW1CT
jY8DEbkSmAQZ2eEh8eJharw78TD508IobKqCiBWOKk9oNFIuY33y4NvNAxtLfqXXWPy7th6uNCjd
UlTBZz4KDdau9ZwEjPCH+4XFM+I0E8QLDQDCHLhFmMzJZVA4Wch2PaehIWKsAASK9JDZhfla0vEP
NvBu1Wmubv/qt2VKWvsebUKz9azumaAuz++4AU6yJ7mdVOhZp9An9r3XpeOcOcapqd0AMSXWe65U
ldpzhdvL0ac29f0EJJbPsGsBnRn1wQzaKEKtgfGKzSUjKinY1cNkMEyn07Yi5XkaM3MBflVDHZi/
1f3OgBHTXpaeJ0MATWZLZqB+nF82C/WP+/2cdBEZuLIP7Xk+utK0sXJGxfOCF9dIJch2/H5KD0B5
oquD5GwXMTXD3dZ2G7sf99eaHEsK7pKz1Tq/ja9NTBgRYyD7j1LRC9diHSi8iefl5q/BCWplPaTr
qus/LA1AuEcAZk53OTaNtR/1fHcs8NntDsZi3nE1OF401o4nORM1qMCEkary8xA70HuyJymYYOQh
r15VyHSyJ7AGa8e+C5QzmiATNuwSbVxT9KSJWwltXPhSQdnNXE/kHnm+1+66v7OErmRdcYBE+GNP
miGpBhxquLwqmhYIH46ncWeIRsXGnEB3R7llcMDT7zEGpEbwKf8KNStVxMAEEUwBzB5FWKUSQmXJ
39iBPy0/Sqv3b1CaGgv6ZLccj4O+B+q7AugP3FL9kStBvIFG7QfMGEUp1gpsIO/1/XPrFLCbd1zL
5UjIpp56th3OdgiA3GG9kk2f2Rw+09EPX2xRYHq8jk0yJBhttsR1uz8hTosYBO1MwKNEN8ccWMaF
0ljQTj07GGnNpefMSr2Y9RvxGDtmW94qSrr3iZ1AynLRa8bdvAIqbtSHQ/xpb7kqdva3AZCvW7ZU
4SmvL1hYkNT2Md0Z9LD2scqsXz0I4NJOt/t0Z1P2Bcul0+wWtlcjisOqAAv5bna/Xw4U0/87DM6G
67OeIHoZCe0MS/gOQ4cUiRWlFtSJp31J6G3jFA4+mDutpF1PumvRi4xP5vdYjtEE61Hh+MjPSQjl
y3QkS2XuN9w/PUfJZAUenI5f5p9B+GqsBJC0WvMjDTFwHSelxAD/vMKt/skE/Pk1QxaqcAcredoK
RgFjyTDPwGdfJPxiDy7wpoMpC5i5xBd2W6TdsLw8pZ3GYEkpeZPzxpeAqoAuuq/QXYt+uaUiZHmc
ZxVs0M4nF3Z+oyEA5thLyAfpWaFlrg9lXmZekyMwtLqQ8vvRv66U48NskfJy6pSMHan5lJm8YEsT
PVV0TQVkb49f3JA7JKDZqWuj4dyrQM0o7Ss0U+bbvCd9u+NRVNJOWvRu4FIadb6NIdbirlmH0Qmx
9VzS5bUTyUYXpDfZYmGybOms0VYzQUvFwmr9WtO3FMdY4Z/PEsXympnwV4GEpVLJyiIOVnc42Rd3
xYMvJTDgruzlf8nuI3r9a4lYTnntQpPfNykd5V5mIfikQBWcLYmjXIh3riVLHYQr+wLtyKY4i8j9
RDmegV+pe6PsH52Gv01qjM2tDt49SGO85zxCXpfDJFN7z92YH0loSRtrWPv+RlxkxvRIYD/WmusP
/Zh6GuFLZD2rN/uzTIu45Xt2S/RUvazJpEpgVXk/Px6OPnKH5tfFcMQJ+2PhgoUcanF326f+tJAc
40Ihf1MvGDRUOxBMFp5OWSR6jHgrMG/jRh3Os8VlLe5Y4uvqTG7raVvdZm7YuASKG+ftK4iCUiO4
FbuE/RSklzgfW7NdmGwE9IZBDAZvgoogUIC8r5I75ROohNfPAfHudMR6D+XdyLR54whHkfSeICD8
SAYOGZNadwutQg7E6B8XfXftk4/ISbS9160zwhjyhjcTC+0ZVT8d8Bf0dRtnuT4XIftBw4m/IxEh
YYGuph9jL53PjoqFfaNBgGX93ZliBUfkq0eR9Dcgz2RFW9IaDK53fSvjSno2r1vhidXdK6HXxBtU
C1HOOuiVOR5Rrgc73jpLMtkUm77LGg2UH9h9/yRxOZZ/7hAj/ZkXl0eyzeB5AsiLW7Rw9jb8Ywl3
7syOgYeghsTxTQOy//nR6b+02IDUnRbusMS9IpDWjct0GNDi2XjnLzwy0EVsigLoJLf+Moc0ED6A
qTQqlhy2EXfJAVZDlrwiBmd6pwlasrIzQQRiMkxyGbHUFvLVjwrskngnZ7JB+q7yOlC/Jc3WRgeV
KrOOGn5aNmKWny34PWZ7eza+4mUBsSmXhqCHX27IOqdOgBNScZCMdV3tnmIHWfbaD1m8OSPOwko1
LDR3Ec8Qa0I7cFXXq7yJs5kAqwJaKE+9hOayfBIDCd4iXlFpumX8UQ4HOVQhh6NYe8kLwIMyEQAl
3DMYplIH+/BRQ1OXNBRL1cdpEIfycjQ8Ne7reyOyzE6ulgkEqy5Pza8cZYkPus+P95sIynsYS2Wz
0ZmddAYTJy8hODCwT6q62/a16k9wK/s6e1KuomtBBKgHww4nIs32fkKbId5rpLg5mNzwXwW8Q4MV
KRJyFLUi4fnfDnWO7VoaqMdZksTJbHsrk9PFp40KehYwV6dUObG7SJMFvuwQeTWh6DBSNw+WMG+N
f68Zq/TZjsZOsWJFgmA4YNTjCVm0NkSDf2XyAg/NokE80iZ3+0q43hwYTmj9bFC/SlpV1NfehONf
+MBrP8oeWGZ8jT5V7E5LkvYsPpsvuQUvoK1bNFXrK6DshLhYNyqjjk59oDsXhqiQvNMYhgGKp5Lu
jHw7tKQVi6Aosshx8dRjHBhgHCICzEQQ5GE/BqOVNXR/QMunf0e5q86uApaH4UNc4qfIZhafYZu7
wlnZLtT9pv7mgCYIcUsD/VeeW2256MFtvYkbEgkpYRwW+G0EkWGW7174F4k/nO6Vc+6QNXEnvnmX
qFAWknVPC8/K+rufC7SZQnLStvwaC8wXGY1Rt+b2yiIJLFFzVtNaCQF3zmQAV9MMFNXvtW3796ZG
KY0fo3EAzuRzjJO/73K6lKxqFC31GAdqtnkA/J4C/s/cN0orcj8KYhteBN3fRcQyokLkJptM8Z1J
EZ5HQ2fa6VIn0hDQILcRWS29Q4Hv1Qe0Fa76Vx9cglADeOvTQWUgxMStNKoWM4D4sPCnU2hTt10g
RYrtPJhWDkg6ou/QBT/di7IaFFuXSFrSEN0Y5vV+G3eloW4/QLV837zWvcAQoLCmPEOfTW5HEvWC
ehMzcdvxFztYHtEA1wwCZO0bMKeilqVWoMRLUmVYRp6PuCpITG3Bii6aYAOCf8IlyqsEzg6IiGIi
HR4mXuEGsSS1Y7YFo/g/hWixE/E54HsId/fTDVNtavBtQtPGl8c4NWezZQwthb8Ei96WhpvclEbB
pN1japbTw1Xh7zdibz3O+g/y319XtD32zkLm2y+PE/DRdaJ27piDpF4KzCYKBn+VCE/L6dlBM4z8
YOIa0O1PWsxPSgbW1Pz6U8illoui+74TLiTXbKKgDhU0GaspOZEr1AdVzViBotz34eDSGPTbXesh
WTFy9YKy55DM7FpNlfKWLfMhPfiGScFPKT20BZ0cpz6/A0Xc+hi4fNGg7yhU1P6suEnh6Hn2hlNz
hEj5VJ80VmMkT1wnUY2soloxU9froWa6dZgZ8NijmSjapXqGsDRjBRMS81Yt89oDm+Q+kBJ0PFB7
pjTumLe3qk6XzXaDqd+95FpR9J5Cwi2UUXGCvhWGm5sjrTLb37oEIb+NydE002m+UXYfyHKDMfBy
rBPPgICjZtF3DbvRA+O34WgsZq5zyj1hoaWSwcuSQ1xlm4qaeM6xPY3mgOCiX7ZfzmVcpBk05LyZ
6EdGuZMT0OEvlpL3X0zY88SMTVKZflq0vmz+SEybeQ4sawJ1pnrFxamxlYBrjOD05xfBxMU+3+rK
odvIWD2oMeNftAzelS+xG8Yq5ubKjsjKCnpSmX/6fbpOY/uH/+IUjppneFAJ34bCKSzYQCHcHadb
Kyjy4YOjiYhUWbgZoQy3xbei2f0Vc1mja5Vxa+y4X32G4pAYg6v8yaLCnz27Ueh6n6UA4/m0UqCT
hs16R2lBmE8L0AAjA6TZCdaZ5d+7heHcTBwMSDuzIMlymVmZDhUCnGAWq1HsAtn0ZKBR0Lydyhv8
2LXC7BkMX/nvKKKq0O2SZMd6WT0RpUV5/nAuIIVfpS4AvIUDsFk6xZLeovRCoWJxofqGuyiDziMd
nHoEH1BkWlIgKg2Aa75zL3WBeRfLez3xhDNqE5DJ0tT0jH9QLkxt39UX5XjGAjFbwQJGX9GoNA9k
Yr1AhMieIarNtqlw+GJRDgNgEP0FFm1hKw07FUIlHWKijdxIHU0EjIM0DQleRSVVL2UUVbGY1a7+
3x9Shm2fwFb8LmjU6bXtdXuXWNRURql9Os0xviDLzydZb8ggrEs3f+rcEsnAzB0eeBcAF9iFa4lX
jreElo5Z+Zmrvy6Uxz/PAOkwsF0NTmEI++OZCR6RkJq0/lqD4tlyLCR4Y9SybuwTUomWhGEk/7Wg
Gtf7TGFKdSv5BgaEQL8P89FfxMQlRHML0Mw05oaB+zJnsYgaUZY1XTRwvxoJ9jjK+0ax9m3JwgFk
fKx70ggR08XOHQWCtc3nDqOtrMlzBEh0Hz38cpLst5emP/l3XBM+VJiYNsH8kFcsjxY5Ei+IaM/r
OZUdclyiXD8wdZanD+IJ6Ct6hMka24NV3HshJs0GGgAxid9BPgLURY3Y+XRmhTa2Q1LXrFLGN1E0
SI1HWX3CUiuQHd9ws0H8dbq5xGvh+BE79AjCjEmldTKcHG9jGiIbtYP9tq93ycdBNkeexnWi5lpU
Y94uZcepTrWpL3sYuGZ0CIHnoxZ4tbyd5Hc0bY5O1cbD+8uwRXXJ8s4Ca++88iBYI6YmtUA+h5Fe
aeC6/trs06dzvrIeP3JXHmond7Oh0m4Rgd+icQHi6YeeLGtOLJOMthzKscLntvwpiywAlHNANyR3
og8wS/m5E2caIlDlBdd/qZwaORDHjA4LP4Wc/q2lX76Pf2CuiQCrSvLpD65itmnreB9PRo+yBn97
pdcw3WVh+j/Zd/IcdwetTQtGWbqvUa/SLHfwzNWCmBCxlLvlxsWIjNiVUwMp3UtgIRjlDhYS6MqP
8y4WjDCwVXCSbmbOKGbzyIYGzq+Vm1E4y3eKOCauZ6VeWrfLKuT4UcWU38hJ0DdsoBH6eGU1XmlL
YWuHXYR64v2Tu4SVwujdhKYUWJ5EW4vpErhcVj0AW0IQZAP+h9Qj7YjHP+I5iuqFJL9HpXnJ/hEu
tmHaqhFB1Wb68O38O5RnJ4ZU0fT4ptHoDHEkOMoqeyxFKAjL9BjdcvLnXvF9RqenNkRct2ne9UE0
bJOQLqjMSGZ6rTkB09sEtDGx0ggGt4+jVtJTpV0XHBiXkQQhmYR7Tfd+nzZ6OosUF0pM9Qs/IsFw
DYPFBmnfPHYkFE3tg1UR3cn/zvLe9stJb2dAlBvu8FJSZsNEFxFXnDwW6gYcetVAQMQNl0/mcO4q
N4n6ahuMYSIoXm4/vls1SOMMALIZPCMVwG0VWwbDhnj+xBJHl/JzZQ9OHj1DKroyFuFbJHOmcei3
GcFy+Uqn97heYjVfKyiWxQ/Zkoz5af0m848nYHmWaH46LI0eYzCYVF09TPgowENS516n0c6ddckb
7T0AjcSoKWWItkA0T76Q1VLpR6X9ABp1N8b4p4LdkY3DyQNksgG68r76T8oq41fTHSg7dKiA3ora
J7hKOJZOkgg+q/SbqvgNYghQ8HSUdiV/+E4GlECr0UT1YsZ51wsD6NYEZeDmIQ86YDpbA6oAZcZq
nz9/gnVMnhVT+NhNcQXqyX+He6aW6T4WwHyA/s8HvEuPzvT/7ZGqmuXC+vWRU1xpUaZJ2OuRiFd8
grxryv+C3LZJ8ukOcWRWG/3odztY3Ys8e6NS/FZz9yW39pH2A4RQbwYTtNsfPa95pYqqgsaWudeJ
Qz9J5uTO3vtJtHiKAGHAbX9rSCwuqmrf0CVZjNCi6pkpIDxE9j2mB6A+1uiNd/OZ2WOJK0y9xVsS
OU+4VpGqDogYWwpnoQbLiRQwNE/VKorkVSpwmFExE2O9OGGFOwDgE6TPTlm66YclmMB50CRCQZT6
aoF78ZguDxLCGtEqBzfiTy3kLZJS9E2//qP5EvMMqR4pgBtA0FDzSrmNBndwzHnQ3VQ4tih9gXrH
wTk51dwGMx0xYCygIjgR+1zkeZcHgKcGU+xYwgBIERO13uWjyRLn8oQNVidq//2qmEtQjkruLWSK
lPJA/GqY9GCVgXMte+IfqMcAu5j+/hF3ihn4CrjooaYi0ar4iVQCyR+QmM6hr4m0Z7a4AizPqs8O
IFGHD9QhB90szc71uPzxYZjZX4pmkEUAqvLFP+VRpOGdNme3/BzYtNToD3ukH9rskd8Q3MEl0GQR
4w1K9o7okbDOQLsHJt/OfWyglikf7gHWzbg2pfCCEBWico9GRh+GZHDcVd4PnclcRzkxKCqq6/ao
qM7bT1o7pYAu8ndCcNT+KM7EsWxt8H9D6Q6ET5UWr3Qr0mHeVeoD5krlsSa9nkR+1wtVz3oLuFBQ
Bh9KfWmtdhCviMZkocacL+Epj7Yl5ZVcfvjos6EnuqQxohEAyaAMlsyghSoopxTCZyyObywXWVVJ
leRM0gy47ASQnXz6AH/CYlNSQYoUGj27LVXmjG9zlQla6NiNeR5Hzo1JnrIGtbKGtvYEWhplUCKb
21N6rYbYduOELql810Gu2ZnJ5gR4rXv6AmLeiCcz0BJIsSX+qCMKpNDGVHWU9J5g2hTnIB4iCAqG
9wRdjVKbGvLLTHqvyBFRkqDcAf3T5kHxU3r5HZ3Xnhp80FACVnCwx+dr/jWHfXumfDKbR81mhP+7
eWX30Pf/IR+7MEKAmzeBJk4NJcao6sXnIJbK/Lbwby6HBgyda63ujAesn0Rz8+8+VSiEbc9SrxoC
NC1SvQC1bZk8SF9Hsklhookmyik32kCciMafTMhIMo31H8881S39Oj0ijqnJ8h803aCbMjN2+grH
pl5E2ml/rKPk7Iy1ERcmoHsC2GO0euszHsEyupEwzZKhNvx/Eh2KsAmyRgpZtl/JyjoDbPQ5DHPD
HXi/0GAYKaVHCYL/zqcUalDzycGPDccuGnrXuLzawy725VHFBYKQW60x360Y/6tNdXDkEAPutiM4
cFQ1OsiFPAPsOjaw+MQWwB6uc+IdnpAnp7nFrFwiZlY/6cYarjOidh66nfBEMWad2l5U+jehcLRM
FfEMk01HihWV0FZ052+o7s39FLJ5oGZZkCC42S09XhI3xocf4TqNEiQ+/nk5DEiNGi+aRFdSK1FF
3rUgHbtLmgMsaJo6jKpSFSWgzAVuePxyIZC2IiSjFTjT2GVyYOujqw7jsf8E1tlXKlL4muG5HbkY
kofCi6xpEDZdYvY+2KG+xsUiX/ybOsKKP48Q+zj4WtzyYn6+0NRrWDiXv6aVtao9DlFqw2vqlY7b
P8iWMn/j5ylNSc3b55fD/hucGUGVraCTSnQ96unDAT8xraOvkppQ+tUajSEzOJT2wzKBMkcT9Iz/
y/HC02/gzJDWLT2+1yC9VoS1KHalI4ktNCW43QBrK6SnNQEGLAl3kcbM7HK1SoYJ9NPc6VydwjvI
LsEULWYk38uMkgCBg7GQX7dNgQGkAAc339qbrlyg5vLVwMxNWdSyv+Z9EbYhhzbHlVChvLs1lEfv
INZF8jdvkh2T+FEF/zVcqkZgCvKDbuJfDJ7x7FtyyBuffosa+sSmnNND8l6wzJbeaihTY5WPjiel
7SEksTyfCQ8jvAhRExnmsdA9kQtn0+B5de2CYDIPX6aCAuQuTGM1IQ46x3YPizMHtXfPEZkT3nnC
2ySc+K+uJeWmYX0DgXcA5Xzd2f374rr9n54LnsBnLZUkjRokop3Z6Pigun4C3XYqulpY2hHj5oZo
/vb8Lu8qu/xGQY7WBG/039TGWdbaIf8S24ZMGPT4C1488uDinUySkeyBwAg9bESXuvrYVCXbVOM3
gxPEu+Ej8dvGaVTgyuLL0H/uhLcmJOTgWDeQRJaxnk7I2NTrVCLCF/5MS2Dw1q8Eyn3xe2f5TBTH
Lkv5tZPhV/Gny65GzTaHaN3Fm9m8/Ud3kwoU/PZ7TZ6JORcb8fYrY8z+B5jvLK8RbsRsVgJqULm9
o4o0cbuMxmtlULYsD6ZEZzgf1ABlxAoKIWL+NIocO0IuX9Bi0pMW+f4swERcadUThBW6dpMUrU/D
Gf/4RsdHA4GOpzHjf9JVyLm5ObfgRERoy75zTBpkSzuNnsCTmN6NNvNTQrPbtT9GcWiUlwtrhl+/
CD541Rstg0ZPGrfeK6QVLl1/paMpmH7RqxayI0lv+k1Djwj+ggRAi/Cr3f5eswWIwK7aA+D41hms
X0LWXlA9Xtk2mCRcxKX2VNgFEW0/oFhqyi8XoqiZBBjFAXKnDQ+sSjcPiV4ilzWdgoq2HRz+PP4+
6VRDg6qlkhzQgTA4+8kaWDNvo3BoNASPqdv/tYwDCgX2Fn6TeSBBJ/h+8ThOrozikonRobkOZOhr
QOos7jQG/nnBuaRZg0RtxYIWWQjiVRuGB66eih4dD1Gpc02ixE9X0OZyD6wd2rop1EBSfg1XcciG
1PUYqEsprpACF+yASeQubBSaFIBu/Je13dIcynzdaip+9NYLYx1QwM0PH7bL6KkulK1xTJRK3exl
Qqsbi9g06U+e8hodir+bBMPNxZQRYIfQMvGNrexxN0zZVANEItWnB5Zq4OnniTD5QEh4xC8QUaCc
9J7L2zz2f9gDZkA1mDdFlWM98NnUzSDh6wyo+4Ru07sjhCivD4Po942x9NEGGy5T0tqDxWxZ3WeF
R/81p46/SKK/xUUP8GIkJKkDqO5fkzj2Q7tsk2U75YzqESxiy9ricLoO4wF86K9r67sReOgIpgi0
7LngTioNN7K7xnqFSx2M8UkmU092UFfiao97OEz35BItZp2UG37YujKWpLOB/zAjUaqYgZBaLrWE
qYGMg0trIwrgz82mKAViJE5LpNjH+MpdoMsZJ0Ne511OmrjAiM0Upl0Hu1TWOxC+hOWRe9OEBUMI
EvEx1J+V2Cv+mNq+Viyu2VDHBNxsEqJmbHC8x2Ck2nY9LhD9TsjhwX4uVq5Nelzh+wOLV6ClMjlr
McB/o/YyN4W85+cCCImaoNX28MV3QoIUJ8zPGu4/t+zcyKPN70grmpWB5OEWf2zrVr4/mrMlW/YW
sCMayuFCu70ftCSmyWPBHMd8LClyUwQUw3McuoG1TdvpYQpjw/JVRAlyeuqy7okVbH3eFF90B7fI
H6ns3QCtA7ntIw/PgVlz/nju2HK35YpA7HVk+vYFhfdeYQ2at+iFY2DjVr+EbgugX4H1vIqCf0xY
DdnCVheLqYtREihD+7jkMXbPKPvIkFt46SbHsssfRZVWJaTtAqJLak5nz8WkmS4HxKPcC7MdNQaY
A9AJKv1Kqw/aKbCaJP+Xl/IrdKuiA1KQoqzSw+DYR+OdBA7y7354uxjQ4MTqKn1tGVNZfN5cw1yC
jIiHYK7IA9OfZUZHY3b5tcwvDUQZ59lHfj38AE6mu9HHsVknla84cCWz7jsgvlmyvsVghw/8WLoE
k0qwsoTJyqfXt5mIAsl525CbR4oG3i8O0qaQkX5EoEvTXhsocNePppyw5gTPAsToOYbjPx2jrg9T
okEoIQ6oqbApH2ew71mytetgCe4e1a+6KSPDuwUHYPZ1/dAOskHOLyUjySlipCmXdvBWovMEYSe9
g6NmFcxFLwjxPn7x4bzWTRBe10+lBxux6ttIj4LKRcpLxBEe1oN5kVyCroW9N2/I7inUfpVWf6lf
lfvbajsIz15DKx0wM+kihhMWT/ND0ThIGaYDywMvZ1fTtH7DVUjxu8dkxq2CevE6PJCT15859LnT
GRk4n7naJ2sL9dMfo0lc74kqHJq//UaMKjbJejNOHRo3UWzcthf8Cq1kI1uPdWyfi1axpvY/iCPl
PmqC2lYfMmz831nhCaHL8uVvgy4q9ixsVQ4OMzZQIjOyLBHv+fDMvblxGZpMTal/Zhw8Xts6ZhaI
woYI2AQfEYlNJtTAVMoi0P1aX+422iWp3B8Pphs64I4v1wyyHox6UlVdh2XGXeWOZSqeai8y95SF
T0bQjLVXE+UoPgO2V2XzpWc/Uu8CXKaIoOfOtRTZ8Tg0lx8qO8q7ihLB9wwBfyx8ifnrqW5FhEM+
pzRtiiCAWz2gSZmG58gHOzNs4BKpYSfX9Fcpj49JnJcCOCRi/KI0DTAbmPxCmGl5Xj3gOBy8df+5
jqijteooCKLMyCATtmK3Or0IS3mYBsJJrf3EpHL20sguJryrXx3eMpoCB8ti5mykXiofAbWbU8cX
yavChk51UjS0P2KPg9mrXo1TVdkF/d7gvxMLv0k/LdYN1NWDDDvmh2FxO5lr5PAGO5rDg4yRAGPW
OmC5wzOLAeZhIrA0RkkipbOtRpwJOnWMYsjZLjXvOVcz04Kkt9pQ54sQa/OyknDQTvB+6xc6s1Wx
LdUhPSoqdnNpgCRxkX/oci5j29uhEyRIh5zxnOWsSwlbCV4AN7G1kMlyyogpsJXl2PRnzIOZsqma
ZmvZbp2nGLNhPW/ESysTzSyb36FfXuvVvY7SzQk4GU8F6IaiQ+ehl2Yy3aEQ29UMe3Tu2exyhori
vizZTEK1fhcVv6yRooyV+zdGzRzk+tGWX3Xk1KaSTH2zQBlskn0qTFE5Ac7IGoZ9aUcXAbh0XrSa
sCmGjC7At7ZIObWI514fwwDMoW9dDKO43MkSvbchyFT1tD6oM9BDZ3xeUMULD6bCSB+9P8XjGzjS
Tk0DEjKGRKkNG7pjqTYw4JOEv6bwVGWJ3QxuDiy/pPTKcnOa8PYI5KPWqTYOdIy71oUqJ/LIT4Iy
4zfW346djogScC2TbiVdM6aHBsl88fvt+IDgfLR/bXSIohZihT2tHCYRFc28AfZh12Jvw0Th3crk
YVrAKaB3WFD+GkmBqBajcj93mn+Bo37GS+l8jc+oYx5uIv2niqp+mZ+DcURa41lEOnwSI/eapB9V
QvqX2wo3AgmCddN8j8kVBOb4cWkcqQadsXg09vBhJlZCesZtdd3M2JGjQ9Sm9Qu4UwDK+W9GFAkN
m8HCpPIQ8scs6N3Hw1rOkbR2nrAJJB3tWWUs2b87kWY1Ns+5cMXMBFfOT7n8wYnYn/2E0zUjUvv0
XNw1dcYzi8sv7pQn0kmfe98mjh3WjVsyEWeJgxRxCS0F8UIam4eHQXxgbTEOPWzI9OxYZqPVt4SA
vJc5pi8GbUnqKPriMpuWjGW+G0ZchXjwSbE/BjqSD940myHe7G6YjSu8a3zZyXv+OGUc70OMBTnq
EajU9nlEhQMMV1WWJh1ZrlUOxIQudB0+8YsS34clZBC9+lAUIWkcRaj5hr4ULq4NNF+HtuI63+4b
UrRtfFHdAdUkw/2ztHIznDiAvI+ElRGTzJisHqx2iiJzPQhhfTj2lYgh+KJ/xdvHXDSxE9xt/hex
Du+lKCE0u33XaJ4xUjYY1fgXKBZHNzD//dZnXX5jfDHhpqB/spxj1EK8a9f4PUQ09POh+3T6tAgw
YupnHDatFwG5R476k6Sq2cSS32r5B6IjlZapTCb9vbwwoXtj8pnPL6c6BSzrPa55UGar33iCLSAf
rgmCPewQbyLy77ZlEOmDBWFh7HcAWfCfUJCjFBwjhv5j2aLO+vNWfI0kOpSqzaY6LSHPqE8phuqb
qBZ1HhaljIGPjZ/WWrt9wMQgpG3h9MW6s/lUYSWVbzll/BM710Alb/rdmJiTWb+OELZ8LcJ+N5Fq
5DNCn3yKIIy2JyY1seyOTVikSAMcj5fKK9g/kPDR15A2Ow6di/DED5kUeut64E6W0qM42aeWByA7
DTWtJQOjfGco9loMsLmqfzardITRyNA4ZKVsgICLPH6g186quUx7e7g8mrwS+Pm6EUE2xfd9NJuE
yfLhap2zYBtBqs2pQGuMhvhzChSZ2g02LBFwJ9XMaZ8ZLE/lh/jbJE+NuVzfa7Aj+gl6XY/64e8Y
uvkLAlnvSxhyYERVrTouJ9F3ty0mTRPYM1vf4qApFHWjG656bcpceTk0zucoRNbmfhkuN0peJ4aA
eaksqRk+CmxsZPSowa0U76wIUKHfknk/OsBXrGeXYPMy53rECUrKaka9DbRsn0rZmvplCkkOe9xz
twRqs3KNKvoWEe7TGjIsYPT9dzpa7vRjkEgszFdhhRI0EdRVYGE7MmWmzH7Et3KoX+syFYSn6sJx
gHh5ryRANeHbXU19adLJ4eKuq/jGn9y/sRcK+7kp0HRKJfniUxPUYVbS2gGLlz6z3xHPSZj0A/n+
xGHs436vQpXBjI1o7KOrVnMXFxlj0y3EGszVNR3dsKkKcB/yYDBjL+wfRyGgHqHwAbCxzR8DqfQU
zsABr/gM7P/0p3cSzDv3tNqtyMjPc6RLi1NcB2STLCxMqAti1/sjr8mJO2rB98Ex5XtYgN+aEmJ1
LFfmtEf2SMU8BJMpXq+GeBPeEsqxupwhz+F7QjFNhnwkvakDU2wkBVxgK1vPuXfTvTv0G3PmLRnl
2150NPgb9ajvZhP+GFn8dEU4+BNLQ2Xll2f2HoSb5PztA8B3JJmSJgITkg/ILBTi38NqC51XW9NE
UVt9eVpxkgm105MiAqL9NEExCKIPKkV0SQbBX0zkQG8gGsbEMNUkMCc/CGF9nnPFFCvc5Wqsi6Ll
QBKlfZ7AhaRXGgLbqBvrccFp8BxP/5eH2GJ0ZrDWBx1hVAie/763HggMphGWCRmAYio0CES5qpsN
VNoajJHgTogB45hKvyYxH1BxhzAkrl9FYkiCWrDUA8Soqf2yTczsQGtPzY88fTyQbN6VLTVm0ngX
pxC190uJpQa5AAp1PXDsMyRUbVSd6KXkp/in3TF28FY4QqyaMLW1N40bc0af9J+00VE+Z8DdJaz+
rNwcyKnnol6BiTYqijyKkFguTAAnQjE2YwXHcTHqH6RZ+DTbp1yph/dr6FbygSWG5UzkO0Qxavnl
VtX76Bk2XxE5DN6slGATD7nhiniQ4+pmJpHB8j9oZY82GjqY6X0hcoLpbl49sHBnLYdRcYiBDXMO
W9hixBO+lzzEH1Jb0ngpeMVbMAuHL4CExfUgwV4Q2+9K5Lp3cAeP9iBITLiTwi5sdENkdd2CXOh1
YzO3qgkEcqjNW/L4bkPxyh+bA5hINtAcUwWSDxZdzJTgY4m0+I2k4XORxvWLsNeilj1oKyLLp7pW
WliEuVcBZU5oLRh+U2ibIJoz56//Z3iPO2y6oLPudzi6hjWUCM4+3+53ZNW7HzPY475uRbfUgCU+
9q+k6NuENLgZyN7A4kKO8gekg9X9+I6vR/PUE+UQhNpkHHXKVrClHk8KwAmGXDpZhzWVZyAQ8KeJ
uUbIVgEA3ZHWtDwHp1CJUe9yIbdyPXoCGw2aI5dt5+KzcFFGOh+mes3DXRE2iFFAl/uRovK20tn4
3SKpbF+K9jYfz0xFHO9o4C4hajc+Wi6vWXXnBVUkNr2Hptqu4tI7iUql1jNfFQTPK8Awf+ltY5sf
drhYwU6OQm1U1r/CmffRSrfvbRltlaAMZqcxR0SevD/R3TEUyK1N2G61btPNnlXE+bzrKQJ2bP04
Xxf/fhL93DTEkVinuo116eoXXRmkrhdv6uz40awoZ9liNcHwdX9/AWvrkshMiOFGrlv2iLBlp8S0
no6Cxtxz9fGfZ1AzDFzDdwSzS4neMD7D3DE+FoWJwxCKwKC/8slbjHF1zHIwXG6mKUqkR+YbzXdi
XUNQknwPgDNbdCuG90laK2DoOBpw5gHQ8WWChgpMRzQWdT4lnGl3+DrLWh9kg//2QTWPyENo0NAw
hY7Vb6Vuxnn5PEqlNdgOr3mJS0a+igZOETtnijeRwh6jTD57N0Ahkk867jAoGy84IeP2A0/nP3Js
cYoems9F1YRal0ZqgoXNGNFnwRWinkOgVb9il7ye24VPXL3L9rHMT8AvS57bHsWmuGlWZmcSE0DM
jZ32Y/0BkczbsAo3LQFjgrGeVBIZ/VR6SFY58307KRqps+4dB+cDXPLAJhKSUh7d49ZhfJpT1aMk
V2l6BQmQp8q25FEKDLZwZ29DILzpB/w6aFFEhRfYn9H4H2/edfnrxVDHRly18Od0qaodIvaMvXzw
VeBYCp2iNCYCrVoRpIspDPNlVi76XkWow9EbJxrIaQPk1/J2SosiTGuGAv6BOaeCgawzNyW1yVLF
jAokFoSqMNnFG3nS5APAJI1skDaZLb/eBQPO28mgNIlZycMaaAn/21TC9UjD1FP2FtaGR1/QTYH9
MqRI4ymMg/V2o1IDCkJs7iBzvB3JBnfjBYTLbadW2PApqvL+iemqA+TFaGda41UxRsM88TJ8e4sa
p880KmXfKAtPi78YDv6mN4RGpsdiNISJFOvV3SpyRlK5ZA8lYbtD2scA96n/AJKacTSMplMEU0PZ
1Ds0pHQQR9N/0UqF33MOzMEoTmL/V+7Xixq/WbeOSJ9O3O/guR9/KcqzAD1cYTEuAmxspGe60Vry
sem6RgjO7wDK9BUZ3OX/KHc6DLwp5u6t8wJzlbRD1PvjhrJOxNDEyERfu/Wjd1YEh3DNzzsmqIT2
AcquQK6owILBkkc4NLagTbYS8OmB2xUvLVDgUAB0q8o6N/b43np5013OLsmDzOQPgFUsJHqqTGoq
fnOzI+5KSk8kLKlz/3t0H3DDwwQ8CpmIU8Wy+d0WJCkf4KbYHhQ363CsJwQKZpk9x2MGRlM/EWUZ
2Skd8znRvt2LuvyUHp/cn5jk+kbmH2WjFyvM4Hj6ifhuU+bP89DdoKrDZhBn7+mNKBDd1OqEsmo2
neyGssJjqH0ua8AO7rBSFM4PJmdlqSS5GUqnAz4+bC66uzpDToWs7PkseNnOHlmu9WrdB52jEu38
jivT+5+CSDhWokSc2kYYKCMnH/bFkZnf1Kqq3UO2RJa5l3cb+3BdLQsNFW4W5m3svuxnYCGvknnS
0XH6hiKAr9QCnzJzibni+G7UdFKAmc82F74kHlUknboFec8Zcl6usEckQ+cAi8cD2abH2QeCSTJx
JCde+s87BuYuq2KbmqkwMpEQ7WLLXMD/hJqB+NMjMHDct5NflUbtU5NgoQHuBYXBqqaRFEgUZ6lS
dFqoWEcouPaZa4rva6n5h08mCsKMvRyP58COu8lqFCwQL+AjXYsqt44IQVDbUxoVjRBkWIXP6h+W
MypU/6YYRYTDoyi+SGn+wocEYWiDzTvnbL3iGr3uVC8aEf87Mlpx95w8rOiWoGXeDoylX85XWWJp
P4mX9uZH54svVtc1vcmXs9+mCplsB29egVvcsiRBOKkLUKeprzdyo5r3Ni7MMXAK0RMjwph34Sym
p+w4l6IJtvhZ+sMg7IVRF26X3RhGWaswI4t+eDu1u9uAc27pr1qOD3D8gyCedjXkL77J7GwHx1E4
7At5BIjOB2g87yZgwKiqmShp8L+PEuDbZm9qVzPxQP/0EY3ej/I2SQOdIqQD1EaVecAHrj1jy8JI
dgC1XNuKStcDf+PwjEFPOxyR/kjCSPbJeF50OOfSfkGEk82Q8unDCNrGlZqJ2YmF70rDsgMCJcRg
m/QTJJL9PmGxZZFvvioTkNO8fzsM8y4YhDMbj9AyzwG0n04pWWXU8dLA8+kW7456XmljUAwPbSH6
2f3V2AqnCSMCByd7ZR49FnM7tijzJZIyo3kr4UsX2f4vGfKBkw1nxBFzR5aTNlCl6dlcnX1zaU4K
dIKY4pWlPFZmdUinnBOSw6dUHkUlfbjVpMaG9Daf8n36pKti9+0glmxfxxFsJiTrC6ukDYixVHm9
gmkUwW69inOdfNG/iRYqddu285cFpwC7zwZkNM8hnSgG3SDnhz1CM6+Vxe6nyhd94c+85I6cD18K
hS3iw5G1WiUy6KQH5uZFWx+LX/4FenuuLjClUBKrTY2DHakQA9OAsymHfD3P0ZZveW2T7iv3KVDP
vcOYOiELvynAHtX1Yl+tjptRxiSVyMZZ/QXuBO78z9a4Hfk2N8/VRHAOikC6ksqutAQ2B5XzSplT
rs7R42Pk+ZVMQJ1LN/1y1tfqKtJjjVs3CsvcctHRbWHQ1VlNeahAV3Hs/f4BcvRq3v4rPcBYHiZh
ZR/aTkww632rzJmj3YP183fw2VJZabajJ400a/jTkIKLw2F//PioDCleQCuzyGmQYBnUSfjxFZ6o
/IzI9fgY9lyjoeIB7fTcgy0ARf2Lbd4Hs2BLa9XkA1SS8e/lgV2qt3Clum2tkARsvaB+AMHmvx+t
QmwpGid+24Be4M1/O2IMq+5qVFFJc06tcxWwMS1Nw26ZftSUZNSnjOGZe6IsthQBBl0Ssd2biYu6
6Fv0ep74Bg19bgMqOE1czeJbzr/sTHKPrMPE5KZfwiDgxPnzqIJZuB0t4pL/e80GJF2yR2hK7Ndp
iSZSTv/3bfhMdPphoZc6zaAD0S3wdIOxCT2sNChJLdhPGgY2U7Hkxs1wExZ0B5FvGYJpsP0PoX6l
zPwrLThIs959SwZ45pjfsyKM6xZCCKZ5K9ZSe9WMaV9lYGFQWGbA8f5DhiCYvazlMsEHZ3SrB5kR
YkOZOpi/0C4VH1ya8kCLLoUXvo85/ahd35wSAsca6PbvOadh6jRD5f5YPkkXsj2CSyRJMNBIpLtX
UuP+rT4gr1+9JGE/N47gGVvXdmfHyVs4hSegjm2MjTjhG0BmMMVAo09bdU211poRu6TaOZGgro3y
unlIe+uiAHY9tAbbrZiIHMzzv26o5FD9ZIK/uKqmmC3Khyh53iX70Ynb+hKmZoqkneN2lMhb3TQc
JKxeymzK8lL2vT+3NJ3/XFqEoTsi/rGnp/ZI8hHjzMfIWiDTSyULsH3rG3cIyjEMX4u70HF04pKx
gzNdJZcCna3cr9QE0JjvvrToOYKLMKshsR4oNoGGDY48hpAIINCqhWWZiBGSiK6REkCAvAiNQpzS
UgeKB964JticZeDG0RjLoAI164TVOtkmf1FFKlyHeSFF2oOOVzfCqVYRdEehNADUYqM4QjpoZDje
wO5nq7chNQqAbPHfzBZkjAZ/7MTvjJG+qEbAVv4qLnHCSZ8jv1qhAzXi8rrpnfUwZ/TdAzPU3PnD
vsqqICWlEAp73+ap222NqNaA7R2EzlcTTG5HQDtx9K0klhdym1hBym1Ziqskzx1Hz+ablZBRujYa
7RoDWGNrJxSE6Kh8qd9wwYWO9pfiS/UBj0IQ9kb4f2KJyKxWSe2oOJk5L9HgbVNwztfLvK04UK9V
E61OrakNUOhU4YZjyvkEC3Lpa1dDEv7pReee4xiSZfTzJtvsFpT6MReoHVBTJWz/2hY45J7gF8C3
+FfVN5zYvNDBZchmbT6spxcjBNfkbWbkrz0+OYJs+2gffr6QQutJwplOLuPhQIrIinBO5HfSUbWA
ZSIZujdEu7s/YhCLx+SgUjgi/kc26jcqqY/ShKrcuxP9itEj4OkzztqOuEBeJhHDrmOmKJJwUHZU
1NUSFxIWytXztm9WLPUWlQccoxOdQaixju7NwoF6MoEfSBWV5KCStc8mz7vIMJY2tOipClCW9+gh
2dNssPTMqR+87P0K6uStCjPU0MZxCJJzfohVjuAC+ROYZ34zeXCZFb0+Jf7QPs1qHj1XKJe2X9xA
OiwQ4elV1cA6UrdpgtRn+92JGHlnyCKMTG3nJ7XXPG8XkZJLO57uj5w7e4hYdda/OAKbd1Ln8ip2
VJSLZo/QYGLH8xoV00W3cOKUFimoEmcjiQBdPCy5Pm78q+zRKlCztct8mjrmFYZRdQc2e6d2+vLS
U2IEFn188E+JBrjICmv/r3fjgAc7iFjHqmVtGJa2u6yHK/oNi/1a5oiYE7KW3jdiRkTV0erpzeZe
qxbiWPvQ05osSUPUsHHfxmOOGT0r6d/i+TsgISWXjHHF6uu7PpC4nH18HLftprTcvh9ff5480APS
aTGyNcyIbhQVjoBfrLN4WPhXzhBc4xHiDSeuk7maNrrl1hp7D0VssgLsSd+qNuTRU8TYmYnFGt9S
FijstXyWQYVblvu1lWkIqhbaX0SBESLTCopSQnzxACW3fYDrKVHXHDrnNpJnaP071ivuHfYj19WG
x4F/bGprzoq09gSQm8/KyRpvU4o5KdmA37g/vMDJmYP91tp8Mdgx3oRdPRu6BO1c4jyKhC8J8QkB
74m3FfXNNmJRq+OXCFO5Rf5qvOC9H2exQVKwX1OGCXnX0lHkBoXNmFYsgSUEBoytrJM9iL+e0OdT
Xb49wAbpG+U7ntycf2FapGEe8AAOtpV9T9pZOVysxm4NsJM56tQIB+QQZV8PKJLEZj9O02W03FER
V7du6JqAABgLd1dKtQSvtraY3WNUt7w8MJ4KvDIl1CY9/4XaiZuQoaHXMZbeTY5WFbhcT+TeE1ul
q3Jv3IMJsECTcuLbCO9fhbfgFYPztolVdF7vxQ3+0Hg8au+zDLISsPsxifkFwRqRxGBYcnrfE4D5
BJWJ3amtNhtVWvzc7ies9i6putL52Jg41xBwHxdaIwjHJ2fJCtgG02H5Ox1cgatZRSMvrg8hy68m
EIXLl7u8UKfPHlIYjiwpkNDejgYHFXwgp79IVHZiH4bbc+7ZcGZl6HTr9nW3v+CsWmLnr1fQXCu3
IbGLEhvX4nzj478FJlTOXHH48m29XflmyVXHCyav+yO1ehiO5NSd/jH69JwJeE/WjS2Chyx1ozdP
t9YF9sCAVjfqiejwwDWqqnLtSe+lnPnU1TrvkBgVWpmJku55Ih2OrsVx0DhKd0i8wif0QrVoxzqZ
TWk+qhV5+dyjmvlweSMkNqYn9++epUuJ74AkMtiEbFiz5gjv2J01x1H6sdO5RCRttZ4L8kztTaAR
jFF5+hk1MdiQyy5Atpq22wSsN3WsOvZtgXaQJvZh6kFAzZHIppX+2ckwTS7DrrUujq76/dCwtIGR
Q5PCpaB066CZCO57lNhDR+N6MUkgsHdOkQNGi/1sqzsLfycogZY2Gjtgj0SL1fI7turxycS3rKeY
a+z9ctArmiP9/2A8puNkTrw0HCVSDJAXttCv/iIuNM+FW1mqbKzyz3eMI8WeSaKDBTHaUJQdZRmM
tkagW/TdwCZzG1xdKtlZ8moa8cE3wzGgPYCq7NBPCF6CdKDrCUioWLsYzWRDldAdOcsn/UvY5+KJ
ovBDlbkQ/qBeT4ociWhx8mSzM3mRGCdl+6zhfOD9BP+4BZBIVjTeYzVr8x/V9MtbXBJf9N0VGXBE
xbmBhfYyMahtXNeBsSQmNtdUluj4TmFWjKRCSu4XnXmlau9LThtlTOqJoz5VtymXmRBE8kzKCVrM
loBklE/zLFNVGKv71V30XrQaVJb8I4iVNlJii3jP1PemYWmk1/+a8N2Lfp1kYb3uedUgHYynleRk
+jjH3zFG84i0NS2ItwQL+yjrJUI4jtGiuafbi/JLwI2hxjNKfZ239I7599onj03xwA76tznjGWwZ
DyxwFAg+Z9SjwoynyekUckACRcjgb4j5UmwLwDvZmP5TBSAOFWv4SmpKwYfVlueWYWgLWexRJTH8
RsOlgZGTKsq8OT0N6GLPhlYw5kJCVEaGgWb1gZ9/73/PVYrndA/vo5rfO84feX601T2cn/xcarvw
fxw/uQ6fn34QFAVUWSqBTVO6ApEPvzKimcx9agl6WW1SWQTtJOCdz22XnEI8YZeI3RuCbXhoSqhp
S0V1AUUi7lz3JHXfWBrsHTBIBsNDX6NWWs7+Fig318JySOmmp1nMAPttD7s/8Qwxp2qf/1imBtBx
6BmtQQG8gqaAvoxI06CoimwAFH0aBghkz4x6KxfCbuqVzhVbmu8KdvUNAUv6ETbB0YK9mlrgBZJe
afjXpajeAA7xUQfNNX16w7ycV8Csp9BZ7LjiGAZlFLXFp8W8WBogJeeAhHW2IjpYcNXOm7K2E7p+
Njwe3sjEUAZBf1B5/N3icCNDTVyzUc7Y+wIQoiqz6SweyDPcusAT5vS1JxDHVmWtqwMf4EIwkpGG
MDyBc/00CWTm+PI2Jr6PKdr45Xno+HweJ7QeN4IJMCTh6k0xszUkYxMD5JNSCAkJaM3DMBKbY8Xi
ipIdqlBBb3N5PAgNGua8SGxZATa7vx9q7TCTqcBamiocY7bYY8mkieqUuYCOrEab5YbOxSey7Tp3
HY0e6wN++9ViKnsJxVB0RBHGvOhGzAxQlLVP9Cz5ZFUbsCwL5B9p75ztmXZOs4bCzbea3Ee3raxn
pRtA4FNLNI9YJPxprjEt6T/vwhFhMvb9rYP8BhlS3gOgqHXEmiNQiONPT0kyAggOhYYGhUBEY5I0
V2lqFd5wth06jCWR84unfCw2z5bw6rqv9NP1vuYsjsHqbpzsK1kdsUKwtYQtDkXnfLPqKKYA7hJg
2rasqQue+9DJNiEAcnmDxo7CUhrFD8SglUee8EegMmfXwdoMmuq9X6a5F8stXozxKbj4zX9mhXxi
1AJpGPzsgOViRw69NkUCrbpdPBz4MsRe0HY/LLzJ3dxjZQ2wWLuFERTw+XN0lFUDM8Eo5kmdmRzx
xnTcOrUvFQokzD/w1GdLI6UlafWsNdACyVfYjQMsm60VWf3Lgj/EspwffVvc3OLvXWXZ+etuYssX
qpkm2bASIjqXbQ5Ts+c2FLlsbbRPgm/oeVFdM70lPqrxHy80jVPiT4jwkICdNpGXRgLHG5JttJHH
XiM3jXxnWdBSl9uho5TxjloElnfUJsWHd4rg44A9/a4Qb6p1McLZM9lqzXtgz1AgoA21oboSZZNj
OM8qpRqiebgJgTuhyHBEx4tkY9HrDecGratjI2aTKAzAWAuYvJvOTh/AMEUKKXvgkDdH6Bq3UuY7
p1wpyG90khD+afcT8dgcT7KIoYbMiqkm8+kMC1DagdNr3lufrOJhCOhEa0y+iW4FxeSq8e898Epu
geWlNXlGzeztoX3/nkC19YfF60Qic5aucm8jfL/JeJtMWkn1oI//coTeex5R+feNdDeadsgohbeg
36zIIAU9LeD38aIMwdt44gxJuB5dCaPlL+nHhDgFRoTJgMe6V2061ezv+JjGanz1FJWTMVaxi9P0
H+D7rb6fxQFodeaHeD7CmqBRNM0bMo0rKRiqNH65db9ePYuTdgBpuWpoBiwlgUfCCX6L2iuhFv7w
dxV1jEVzPo9yxXuGS4Oe7POcLEZzjhn0VnMT1AxLbdNXDlIxkaqBv2Ka7upIZzpZoDTq3yxhqjO+
EDYlRW0payIT0Hg9FDL3NhA6TFvdeWgHZM7Sv3eI3W5N9Q+XbFFHb6n3Zl8RLu3qN5ZLyn4Et9uE
8rFFyoHcS1wxhF5/hv3pMHFRNiME05fvzQJ8RzctKa2nBYR/I5u3qWwnF3kkGpjHJyqB2BvVO9AV
c3mRz+3dgOxbfcvRSzQpa2jVfO+gsjTt07I4BFQaR4t0I7VY01H1+Mr1b48+kxl63mACqV/Z/HDE
bSbdBlrmH5BnIq8H0onv/xX2QXfZat6vFFaYajpVFXMN8wi5thpsZGRrPOF6ZkDvJPmI1eS28tHH
N9lCIQnnqT3EJAME1YW52dPwJmRWkPs+RA+sddKubETRkD3k9H7hXOus3zmsSkUU28zRevxAayJl
nD8OuaBOXCqkBKKsOqttprTh86oVkUA2SpMUDAoJ6KmEJIzDiccnTOFjZVhOfNCiNk4qQIPBWo/a
+TUI2d5mNEP/0FNKPvUYM66l4YstAYExccRcILoZkTypDui3bbQ9rMzy4PuQlJe/lr0saY94F6Cv
7lpzOuP8JzQYlnMv9prtEuBOKywWAy3IXQCjwHYpFrOrDpaWyCdFyM0NPmcExLvJV6JsuxjiwNAe
2UnemDeVgNvD2Qamiusv3F/w6Ua7wYEIOWBo6/54o+dX/7x3BU3YqNNg2wJzQaUrIcsEUCidFGC9
Z5D/bVnQ1kFyIgM80Mzy+GT5sQolr0Wa4BHH0lHnzFdzRovHQJyycNbqNA6Ay12AYsytMbi/ORNA
SzEZ3brOZ3FnUoZNY4k747woBDW4k4ZqLPziWH7CzxucOrQJ68gCh/BLkOaK7FSeNFxiD3WdZGYT
B2T93NayZXLCXnUXMeQa+9ZRpL8IcEs13d68/eLrEk019RPf1z9gYhjexOJ7KZkMkG97pDvfCs34
AEiK7Q/RMD6r03PeALV0hm0Op6iKBkdzJyk1Z6D37UfYlrMz7ge+ihNFOeWCmIQ/WkSLJO/Fe1hM
z4+4CeXy0tUT9odRob05NU3F/1s0PGcefQOQ2exqOSWocSAsDOBXtGMQTr9c/MFUaB3Zy8ThxMxr
MWiFs+Ab3IWbf9LiIVc3+9E7nFWNW1R/ktMyDGFkkKHiZGRE8aLG5TMEuri20jx+SrGLOE6F7oco
uV+G8QVVrElF7alVMtHIwqKcWMqi2bTdKQ690uLiIhSSFszPkshkWe+CCVpBZNBcPKUzvHY8AZj8
VN9GF5c1Pn9ukUwafwEorXhrUmYVfo5hvOuDMsNGnz2DrGx+SMeDxanAxyoTtlD8Fj14m/cB4Q/D
o3RhY0QXLaQsir2mYnb00/D+1AIlZscwS3tBqc6Hv+KR6Ck4qCe/0/kJOOYvbkTdOXGrJcsNEZri
RCPXvixg6PgfKy1U8O5MZh56cv0z010BOXgGmwlyv4ZhFT6uJtcbb8lpzUh6ztt5PtKZ3H4Xlvba
jbGvSc8FARNvJyk4sYGK92pKijy0jJvTKd+1KzeqcrtXP06X8lg7iA12CpDzhFn1XxvYumlxuC62
90YW4egLnnaVbVBc7QYtelCyv8hjiHXptcKeAPeO4gHy6ORLeVMcz1biTfjOtE0Jx4hJJYZ0jVrT
W+nxPGNMzvRYrf+8KRpUqo4Tp7ys1qTM10RZfRUBmLUE4VUKPhdd+NKsOQ1j69rPc0kFMFNPj867
EFS5DvspzxGNvArSeKsFannm3J4ZJiN5mNykJzYFt8g4uilK6xgSPn8bnePCvUvxzgXYR6RtB/Sv
Pbr3/kboJWA3guwR0Cp2UL7mQ29SXChgu0/eyXHnp2F0jAmf0xVJK8smLcWGTP4SHc+ftzVZXj6r
ZmmEpzuTBk/+y6L83as70usgN56/1NIs7PtFA4GiR1GH6J3S3jXX8RiyRlwjQUHXO/W6kVuPOJIL
etgQxCOyoTfei+koRp09QAibpVf4tkPsxm4KBy+/O10efPmdaOJi7MUd9HxA4Pvmc8128IXrvWTM
UTntB0yl8Y0m7g0ZgdO94C35sFeubSxLUCQvtcD+s+9K5dK3rjuGzmzyrOoIfY7UXe4VP7ZSrAtK
ErdarJq/yXFAYNd85SGhK0b1RdYTo9uuNAC/OCPUzgX0zreWBtbmEsv0VwVR5DWDLbw7Rh2FumVA
bHeEjMT2rGtcO8MpX+/2yhwurLZrNGbYIxNdG1NtmC8nsyARPv19KsCfnx6BqTa+f0Yq6ptD/sQm
EAvz/8fAbsRGGLwlRK/KS2GIuKgXgm62zXHNae2DPsGLf5ZJm5RoLLdQAmI6ttydt+6+gSQGHnx0
WkYhEKoJlwWba+ap7ya5eKCML4xcEK+msU/GfYFxUrIVlhVCVwbzdeUfn4SKZcG7MDgzDkkZ7Oqm
SZnf8hEARDPXLsWKT3+dru0oHFSGmi28f3TbjkJyFxvpCurzfbFdU2RruAKAXiO3cxo/bEaHcNTy
xZ0I1iE/Sxsis8l329wGIdxMLYUydNV3gX3NwZZSAa4tO2yaGmN0orS7yIZY4A9Q35IXslfNVNfz
mghDCxB8J2fX7/K1e0mNlpdI8NURg+8Woaqk9MB1pZYJ4Cmy97VU53iInOZ03MD9KhTmqGIFKCWs
QVX0SCyUYLuERaRiJjqC6U3LO2Yq0VMGawLuwYWakrS0Jc67spOvdfZaVctKkibrmLuAJpJ+Oavc
KsZl9bkak33dNWB90jQy+eVS1wGd077yjYIrPpvaOCD9R9pP5OK5nJjfTtBBZ9jkk4p5KA3i0sA6
oQ5sMUCA8ccztmNH8/vHAyJypsxZPxWb0qsgwGPFV1SuvwKe2lpqdeJu2iR8Hb5zsykROtlSXatE
6WZ8WVXK45C4l2cm10mpODV73/k95rFex50iazDzyCwokoZoUCXbucJVnCt+HdcK/cnUH45D/QTw
XkpzqHZgbuYXZGXoB/FpTxMYUCm724LFyoTnCA0n0D83KMVchEWQ0XaEgtGgLy8TD1Zirm4cpYQh
XTMsXQeEvFbjXr05cGya1IVL9f0K2ZU8GTWz/NfqEEX68qWHEYcxkEQScReAwFfE530M4hNBdd5T
w02aC2T78fatg95EK2I/jIrvNsxPNT2rELC4chViodr7DsJENi68YXO6X9GbHbC628XztbyU1u3g
0bhP0DxfCNdt2ZbhAAZ+vSw2fwQKs9ojqYy1jWm74YW8DBBDQr6SuDZADi7cv+1CDswLZftPtmW0
6JGuKfztNkinX2BTFmjUCDhENtt5i8EZK9TclQU+91PqYPe/xN6sL1Hkg/WWGgctwKZdAxzMEG8P
PlTLAN+beUO2kf07iBKYkjOl9LY8eGxxtbpEIh9LLgSy2BhgreJ4os9RlSZr7MRL/KzcY/9kExJM
nBcQ75nDbX0TA8lmcsC/aX8+6afegoxGSNjGHZYZQKNCgJe/EEaenEYxZMT8GhiYWYP6lbil+TLY
Ldzd3ccKlGEjzHgOCT2rOkn8LUi2faSMCJSo5g45C1vCwdkKCrgKMxl6qcyBCGxqUTjpfUQK1xYt
B8Sg5C5alRlKyj4/Jp2HdD+8hC876SiKlKGxDBm9/mJL6h/6rmu0cWD9YdLKCTKNbV19Dfj33Asw
rRGcQsPrV5ebiRjaSeNPE+ImuKc7fOe7a4jGiIQdR8hc6dhH+Iu1qedVgRAsq3L6w4RONF15S9xf
orhhqYLV8GzsQJ+7hBpPzWn6giypMOIGrkul0ZwEgXYjY7G8PvBJijhV8xN6d/dcW86Tfw6hBweT
AMXHJLSOmhHZtrFAKVhePcqduo8ESuNfhPdv77uB5xxPVZd2eBr1ULMdUHzbfATNGJUmoFN6J7AQ
giMLvYO0EcxT6gdE2tjz/3nznSZNXlTt3qSCh0sTNhwHFWGeSY49jLBcT5QtCBG0BX65qROq0dkK
yDV/9UAzt17cAeDd97JXUWxKTLQU+n7252MDMCbohkSH8zCRS1WkSlQRif/QRdUWN1cnBYCfzHXN
6+4CFhXopkwJhJYLxg287zqXYYTQAyIMq9h3ptzY/1Wq5T1QuEpjf5+LnHx1MQtak/RY3tV9D0s2
OCWfI3HegNavGXT90+bW5n6ze0DnpAoYvfuW7ARsNeYA7x0e6fKSpDDrWlw87+ihp22NEzXcS3RQ
uMmfVnX6Z+gQQ1ADWLNdJ8xW48xvt8fdXbBNXK0pyqeXP/uxHkvijRHzfmMb7kIyuCELd64YbBr2
GV3dfuiHAZhaQRgEmkBdzO94s8kt0n3256P2uM3MH4OnDIMplk/rIkXH/7NVa5yvScRoEB8OOE9S
/2yjSLYlffcNPR9rwYLeYKGiQ/ii7invPwJ5MYZ/+pOiyYRjoZLkdAt0gAnMcT9kIfXKrbPyw43V
NA2e3JP9AU9F/IJ++HXsoVqEg24aDzXqkezidnSb41BY88Q2F0omN1Ih8206hOuOawetgnRUkoAv
iP8cuAQsZIIAsJHpieZhVww/21O6fjGUBp/1Xxzbjd3UVmOwXHBwYLzSgWGt9vMkmyEYOzGyYDK1
7J10XHiAWX57/0LCEHZsPPGQGczYw5kOlx7oPhtxWIGV++IsP24xZR5r5IVXEggljv3h8duBd/Dq
GE0MswODguVEs/srxAlYKXUTcEoeZvwwN3wj0tXhmq59Zcj1CDOEX8JMXCL/3aQNHYjMpkMkkKWz
8hNLyDIo4p+0JGxlJK4ELnSK4K8D8OZVka7ZXwGC8lxBbQQ+fv5yqx8sVGS4PF45nmwmMeYuAToK
r3mFERQr+ZYsaqbwsQp1E33FCYf05ij9/3Pim8suU5JkAcHvFgjvH9wuthbus6/CxE5yXKAMhQD4
q2wMqTRQlPfoVWNiRyoa3qkSctiyde7K1LO/dztldnFWMwhcgNwChoMHUvQjSHOrfPRK0vWnhhVy
Z9TzYCOAyksELWPhbKUpabFWzEdflix2lMbPDF48AqQCiqq6NsvNwaBy/TYrMd8IIpCYltiX1IcY
//MQ3KCRYELogj1aFOgvd0GNKUe71d2Bujqgc3qfgzNaR8mS7o/Yexwk/g+Pnb2aFLEFez6/okJV
5wvoriRhFdd3Be32QBdruG1qQsrxMn+hNdPEBTKJCuLxRjR5IQNZq0IQNzoFE9RqHbpdqbgu8luk
YN7Cq33GZYPcj06bnPh8DYv2kBnafPBDbl/T0505VB9co0kbP6d8V0u87AMNKpUl5JV+E1g0LzGl
npN4hHyspk9QEMR8Hu1cRu3PEULg1Qv069LJ/v9Wuz5qoeINK3/kp8HW4q2ojLzA9/Aisb4Rn+Oy
8mqeM69w7hAvVbU53ImenqOCyskWGTbvgA8cd9ikVWqWzr/Bj0XD+v+4E9dzjahNOGwsgcFmKrn/
aK5lzGwtAX0PBd3bpnNYPC0blBmtq+FVkvydrNnK32FVvxuIqbycpy+WoaWpfOmWCb8+njdOvqQc
vW4UbtlZeZ4yb5zTlCkaRy/v1bjq8AK5Ih+1i0mkwKkEhWbHE+D7k8KT7a64703iIqxQmDaE97Rx
hu9xNfPt6SxO+U9yhqBC8zcdq9xNyg67Hjs3KBQkcSmWkGot3+FXU8pChyWlA/x/M3YiprN+DVr4
oHYMb0YJwkNqO2F7kX0HTJ5+s6/cXbFPjI04k30Rt3LRWwS9rwzrDs2Zlgm5+oRVNR9CIlK2cg/K
iEsbrmOT5zvMZwx2IbBChjgTytuOV6dh0DHi17+xXsz23Z9lzdQoHWIK1G0kfX+WNq8iJAsGgP/H
1I3+uBXud0mqkSvk/jz6qnfU9Xwhs+VmzMqDvVInS+pH4lJjhj6Shfs79+anI8/0qGP8rYczI6Iu
wBSfc0rFbrQhsBP1usbCZAYZTIOV1kL4XJArJhmaYpNpSJrxnDvpigDvAtf6+EE51sH36n2D4Isu
P06o1mFZx+ndoiESbKv7kDiFNIa37W2bfq8TgdCSS2tG0SGty9zGHJ0NA2UM3qa63qJI6HV9DHop
YodP8G7+c8jc9z5uHiF2fzet0IFvlUmQDcioroC8KvZPSW1ied2l47ccqfrtPPToFK/5kR0qpSTP
op/B2CtesYUrK8r6Y9lLR2H9J8t0ERMHKnmeU6oidC5iaZZKLZF3onhrG6n96OXBB3WLjsXPG8W1
XkrQkep9N/4Jxz9WtsUJYTKj4MZSpDP66nEs/1oFNcH5kOhCOLnA+ZsHfDxKGQa3/29AYMADxOaL
64NTarN6B2xYbRYWlo2wRAKVxbdEIYjgX+yN4id8r9T6Y9aB6wVVuHG4gscQ8bzbVGsluUwDGic/
39OeqKNyfeFngL998G0fHnMlIW8ihogvnWIzWn9R3IGXxjxAndlDkHsurSiNgLJ6VJ31Rdv5Ngbp
eIupJWrOIhYdfx7W9XcnpG+5mwHBAegs44nS//Jx6mh1XgRLg60dPu5EG3S8sPoOMyVi9g4J21KH
6KszE3BAZ3lbWn/zeGlEZO4MhLcgLITtRAXK747dCmge7ulE5hTGnKpD7uHu+UMkfs7E1gyGeA6P
6hZV1O2RcwBOhzfEafnxRJBQ+O6Ybkdwq96iqr8D/KRipQ8ANyBnHyJZiBk73VqFNt0zZkCcGoTS
15n4tA+llUbDTY1FWUflPXd1XLn1iNyVxGkBFiMRE8WU8j/ua8ko/tOzI7qBDfLFHRO2xhMZfwjB
kLaxq+uYAUQT8p9LjijvyK1OUJO6byCQijCrvVv84DFVQ9s7ZiUokjWBWDZtmEjtiD3nW3KrbpWB
Mij2MQt31hLaUEj1kVxJwF7ZS7wxzEbxNDw7RlwD43WhUmisrpRdjb+h/y7elxNSfRI2WZ4dU9Oy
G1jhkqu1YxX7eRuMZRBzcIWanYxOmapkrROgyb7wNIeyAgKvDyuVbB+La6t0hw7yJEdDCesuSrOJ
B7tgYtpEKdwYmd7przVP04ghwvPqAy0ggEL5nHofAUgPlPg+kxvJX45C5tO/ULiHi9vviABe6XYs
5CWRjBrFzRl9wL53xKXXtQ04UH7WwvJYf5M7hwOtJav7lPPVV9EHVR8X33syYWX9NKE/QU3TlNzU
DaPXSkhB4/riWwKhMeQqJcSqOhIaoVACAF99DKrqNEqo6rb2gd0b1LL7hoFIhO8OeUy1R1xACdrW
BiQJoRe6ug2mtmME2serrkYxtjeLZlp7VfB9RS7UcLUhXJKeaqPaa52oRIB/FBXcjFZzifa7yie8
mPSFJxDsHclYuNbhAyp8bN/JaVwLfbNqmasqS15Z/B72yQ4gY6SvrTbVZykle9fv0jJJHHp/S6k6
D+3sUHnlT8F9UsJPWxipBUKdcVy2/l2bINHinK1eWXv4EPmT4HZYHFIZCuBfRC2t3jxRzZSyUJoQ
ToLHiLk1oTixJiNx/kzpQRg04SvhmgB8PEqgwkopKMJlOS/q8ugJLh4WFy/2dZP9ep4bMXTCOHOE
Gy9HS+TytE2pOhvbAeShwUFMi0qG8PVr3vqMLqFTTt3lNkl6gAhCuYdT+diWF0NSFM/xA1tFsj2U
yMyV8xKk0KyE3rqskd6NKMVVyEhCROnq/Fa+sQhrR1bnNIuF109v5R4IKupiCaoNbpth3JLZ0I4g
pEKkCq+XFoS1uBtS3FxCwXhHWK8LJzXX3fu9+aFrPxeWOQ9AzVgha0HFhXuM2fRJR8uPHHxth5sl
w2+KWZSKkw31lKewo1HZFXaj946vxyR4+1sKSZeo6RFykfFbIRgNwaFsqEnEHsEJFNvBIpatiCiF
48Izu3HcxRKiD2Vx/Y2mnXgjEzDjEBUr5cq1hR5iTf6nZTZKbu5EIqq5OXmIi1rG4MPuN4vmIyMX
dMzl8ii3GWFkhnF4WW3RvbzEGOr6RXceUSVuJ2ES8pq3mCR6sE4vYG7ZWqciKmK37FDwB5qYi/cO
8OvvCE9/ozrlu4MU9LyNNpSM8vabth0hhrBV9tB8D9gCHPBryByHLR7Szz3zrinKqoY2wRgpDlWU
DgJUyhPyIOR7ce9hARXbIYMANxOCPzsDAA7FGgwDXW+ecLksxxMpznH8bG57oyHQErTf4kK2/60u
W0QglqAOSSgYG8Ub6nbNJ6nEdQO+op/6V9uZB6HuMhmCVvZ1Kfo+rLwN3pdThAC1vKvmXaHgR6nX
3sL1tBwfUxsYNCCzuVTjwMS0NHf1z/H9X6rp25YPXo8bnQtBV2ato5SpWuVooXNBWf4M54PfOMiT
/PjhY8qPssHi71emL/X91gAtSQKKmrvYyXG9LXtAM/0+t8phDtVB98YI6bIhHu3dmwxueivaiyEq
lPhurXmkw1fi8jci6F+QSfK5GrZ/hNBq5HqbvEQOXAtbmXT7B7yJftGw3n26SG6r2yLBpTdS+TRa
Tl/pZz6tKTx8Rg9YhXiby86VeynNhzLW9kQfoGg/8BXYyGWwWLC/v/8pSrt2/Q7SCn3PExrNraeQ
hI9ck/KikFz5HJCx8zo6F9tMiISogUxWIGNdle8DFW+wrhqg9Jrgxzn7EDT0env3/gALKEwSZhY1
8tZI9Owetfq3CbdXYFUdZ7XXUSptvrE+qjyd6HawqnMyrtqHud1Wewq5kTzse0q0+mc9sdI761DO
/LePqwpHD6FkWc4LjdAioED2Pj9u8KAqCJvKWDritA8rlJsxmYbaLDpDOGWHdQGZ1HQa4+tvjNUc
bLCA7S9YwmvNjHlaGSTyiveXemNOuUMycAW43Io/4lUuVKCAFE3gS1r7IKyuF2U/vNBR77N5HOhB
dm9LUpW4tZvHJXZh7J5jYucz8BRXfiDT9okY326QFfhZ3z74Hv2xIkBHPnsw4w2IxRQ1M8y+ZjMu
rI/l9MHxhfffj55Dt/zTR3v5DYTdpKjWRJ4KvLD4oJCYlbitvEWRbvh1xClx5BdiBdn/tb/bMYST
r0Wnn0Gpy4pdpvNJGZvTYoZD+kJ9ilqCiXWygzNNLhBcIoIMiAZcnL9WhU+0dIe2BHCGpunGzjGT
8g77JzcnPy+/H2xLnoYreqVX9Aws6fsC1UV42e/k25MIvVL3E/YuQf9uArBk9NAZNmanJeONrycx
A5EzvJ/h5yryzUbR3Wm51SWNZ8vPzohhsZZ86AxtV85z426TRVHQsK0Zi7+4vSp4ZN9WkpIUIgje
1pnNPUcaFjBJE+SFK49TCvBhG110XQcqYyOGDCDe2Vx5O+Wh2zuUHp/ui8jtf6IMN/o0Be2vqVA+
AC4m3vnyDZHdYmbi6k1gDOSsO7WavvsKSbptjGenI53ukveJSybqMaZRupBq3lEcJfwCXntJLYML
LXejO/ZNN8omCmql0Ob3Q1w97f/wWx9opCsvAAzpSJoo13qTtEx+jwjncbClQViWd+7WnZtYFGRY
52PhM74Bbvs6spjrxufbmkoYlxRkFLihvvrizsnF0dJqcY61nhOnkcHClYpd0Tm5TrzqdBnUuSGI
Sz7M9hPqS4AoOoEmpnwlNSj4PUUT61LfQCjJWfPdXbT2tzo0BYPG6ka9umocBmXUwEasdn3pVfDL
1Frq0SixMBPdZa4BOXszs3vlu1XmyeoHM0C9NpX4B8txP293kM3blvjD6MSroOYp/odeUUrkEHbh
kMPc4pFAHRG9rIdDixtJtMBOxHMab2gi9mbfmqzcMMP/y5zxcFkvpruIWYuWesdi6tEvSXPqQyxt
TfnfYD27mrvQ0SsEuV6rAQE9tNF8H6ZzqXtWoFdRYgkIyyb5lvNBLLX5LFV4RCDwHUH2J97ugEnk
oSwg/uYnQGcqZBmiTFWlpu1M93yDqeoIoF/zmAx603SceGX4zP+4QpM1R9lWqor0HxtkRoWZ6bQ8
i6m6X0MJIUXyFJSaOfD6bBfPcyqOCoVIoGEogvg67WBVqBQvR35moVnGXe8BAAZq1WZpkqbINApe
cqQ1zFBOL7Btz/DTPRyZTO1KADmATZe3q8B7l/Vo1h+C6Ij+0rHYUrOjAZzAt0dFGw0Z2XpW5l5q
/5UJL7T6ms4tUm6KiaT1/kp3XncNAO7xIlDsEZRMqTgw4JG1WDeJo/sYnZ8RckWXyy6thpA8mH5N
O3EvSltaUITvSnjT72R0TS1CrelIvS+bof+AcRGMpf9OhBYwpZPUdrVzqZw1UubBu16yPrQ0Y6ZH
P9DCHz7g8ZFV1Xw/hOrVEzmRpq4oU7NZArPXswlJSHM4jz0GQRMKYJO7LaFWbJ0ghlW2r4Ffez9C
M+l2M96b4bbbFPBDbpochEDYfhWrqMt3E5qC0ijZaPkUbJfe6x7ySBXozMKwIAEWNhQNuemB2cKH
xBZRe4LzmKxsVOMoF2SYArDyrNJSXXKS16Mvi7ytdctm8PH0/v12Vcr9Bxr5oulPxEr45BXhkLwo
p2VHa8IPC8w9bvD9oyXtskmGafJZjHr93uDV6+GqLyPOQZUUNa/wJm2kVUebLOzB2K2ukLdEUq4N
O9WV/t1SS6VqRHmtG2Bv/Uzbh3Gx9EzZHYuoi0VJJ6egdVe+e2mfajb7zyJtWxpHi1piwy9bLvca
ob62RKtNt8kZRx85MLXJtA8/+Hm56MV3Bv8lPr75xuNJbi7BS7Xm4UHr1kMNq3tLiXWlGh+tBYg3
bqplYYtLZTc3FWdqAT8Tjnnig/Xl//8BZpkF62643ASiKn1ZWubnd2bhi/Y11IIbcXFX4AiLoR1u
Uyiwoi4kEBHU9Vm2y7fOI86hbqQqao+BZIRh9Esbj3L0kZ5v0zPV/FmBm6BWC8wax1BvYrqfYnql
/M/Qyg/PRPANk3aPBxQItVyVVoohF1f/94TLoLKaMlUdYM6/SIuco3jAAY0HbzLQVWfdXYXDFQn5
ed69Zq9vQzth65F6v8xvygJbdDzeXWt1V0uteoxzWd78dE83eTIPPZ3gOiG1YDYNMlneamEtrTEf
QkI9EF68C5NhQ69l3d+OFGyfLJZrivmIgwLkMBRWpVk8s/GwZMgCkQ/241X6bR0B3VE29xKgntX8
YapUSmag8Z2BG41QrrqDBW2MupGOol646JH/Fg+G53dpvzPbw+NSmUwJbC7GeUOPZksq28ba3CaU
4zhj/9EQLOnOy4jHHkRZlQYGTHBJdFuLm4G0uL40MQEcolA9GvSGpz+0BLpjpuhJ5wigOX2l+rCv
GYB6fMRM+flVrALV3wAL1Fq8I3hckfddp179qBKF3UzP0pSlHUBH6f7jJ+F8/oSSbehc9i5kFvFU
xv0BYrL2Ua5QsuLJDsFOtJDbB00Gq4ZHbKPQ1jZqK/uW8pU3wXUYuHnppOCRnYebYrlsPtIT0lIT
iJ6qvx4P2UgCX4nYhfZDz1puF8oJAfK4HmhsI+UrUKHpJk/jcyFp5Fo+TNUqKUyXgAQJsDYPMvpV
WCQGwCZ0pMxdmwi0lXyLaEsWhB1NlOZHWEHIVND5fZ5E5eohVkae55PH7JLtQzaUlBecN+HbRUAU
BeSgYO+oX4RJFFjJOWpCRnPgr1CYkt3tmBlQZxeHpUvhmHu5Fr5oi0LqPLBTJZu8XmxztPc7Nrif
4bUOrlWqzGNgywuURLn/yzocFkO858WAXbHCREn2Y4hfxBGcr/+c76kuko845Sc3zrPPfzjSCi0N
VQjtoX6GiHId+qyJYkoqzVKR2XhBidOQvlSRatki2Qn1qpGqkwIekp0Em0GVef2hPLPoV186dhlD
LCcczF5tyXQGyOiivBwqYyyJ8mH5c7CW4m96KhzRH+Bhzbgnj0txI2uCCY3WpC/c7TmMT1P3tYHw
v9IfhUooGMXUjtxHDvHjwFyGpNCjTHhU3eC0GpEd2A8MghRGc3doumqvtguB3xXqYVgeejBvhjxO
mDVifGo3ZduL+J6LciO/awlFnEwsDUMfs4l8wv+2ja32zf6uVBgUGQgifmpZgyHJgdGG8X4y1FwF
VSc8FPlO6u71BfIkATBIe3MwOgMfHnqIH2/jj7IoLPAhBtjvP09Bc9IKckzLcKcBUwCZLfrkPG4O
uEAXza/AJOUJs52KEzfT8vUzJsLDXJuJanz/OJXrqo1Lj5lv+PqvBCoiG/BD0LGxI9CH8eYqrUG8
SVRSRU2vgziSTTt+OSZlfWU++V0aIXMggrp9cEkmzcE6RTkAiFQvIWeE4WEy22j5KemtwfiP1/Os
2b6KgGJvAxNFyDgqt7Xm8nx5iejx9qqaccdY0m/LHIi+EeHEFLYk1G1DZILGuXObdUDdPQkIR/az
OXQMvBHWZlqYvFnHsvGRGwUAMr/J5MBzOMdwiLqde5P3OxsLygUVkkZm1TD7x3Zw/q65Yzz4P/7Z
Qn7b6TkpyQuu2t2/4uWF4x07H0EZzw1yfjKFQxD+gQdTszBZuqhqU4C6VZYEFrCj/lkNRhMCCcSv
cwA94FIrJ+6jHIdTpSgM2lIBlgWLQ85BTHFkAjxVyKK8FH56ON8gV0mv4qZ7ZtCvqc93GEznt+l0
kssfgSLgLjXCVHIDKAgk+FqVdfirTVNVTSfgpSHS9LgOansciWL8lso4pTYAKkk52tbm8TayVFcl
nBIVEPee6LxXM/TgYeyEpqCi6Yn3I+V5fdHoAKjQf1BfDsUNlf1LzkqjtzV+fjZxMqH2xkQ3owD4
b2GcxO6JXW9IiyVpnCaxgM4PWTWpJIL3NOl6DPZ5+BQlLC2eIL/LKuDRXJi18YNd/dACJBbIVbf4
B/etQtKvyd2PuEmlupV+/lfcHxF2GWjZ4BojOyiK1+tHx0ES10sEJl0SXLCYme9hBpJebNa4yhFG
Tpmm5MmlCoc0y0w51+b7f0tdJ/MFkoQUEI9o4s/DA1xQBqNVbOJ+XfhJWELlgLMOcdtI8CAVAypO
+vK3XNbpL3TSjC69pWC2EHGKyIkcke22+ExCSTYS5D8cabwT9HNqvjuNogMxLYBQxqf0ondxvfce
Z4G7Wt17+Xe8wBg7YAMmhcl4vIhBQXkvy15gSqVhFN4GwIdPRZ0ySPdMdTN1yWOzjt964pde4Sh9
Cc9+sAxat2dCzVEMKqEEniTHgA+ZPSidacVbg5N/oyaxguB8tfDmTkkMn08CSTTQ5WjXQf91rI92
zer9HTnyXRAby0zgiM95Rue828BQ5RWO51vNseEDb1DHiZX8f4xV5aGEzi3LoZyTklDURP6nCI5q
Oo7l0Xz3E+8EOxFUKwHQta+76yp9uS400fI2/yVGv80hgZyZOhc6VamLJw5JfaDrfKuBLvDxKzgh
tbryMy09OI+qskjBqcwgsXSKP8rE5sJWFWv7ciWZ6P2/I7OlO5jG9oSPkdlcQwxZLJKK90LgMFs9
ztUD83znLDqDd/eRG5jf0Ne8B20mOB2SsvmhaEV8gmlEGafIvkPu4Hv9MHWlQ0mCaziESTECuHS1
zQroblVLHuh+PjNRidtp/6CqJUOu1+MiwtDJ5nVU2F+XvLRI9D4NKRePC3b8rQL8PQK91Ar+09T0
LFhtf8IWyZ+YJ0XNo/2m9VE35napj4to0H1Fryf4ez8KSRUoP53afGt6cv+d6IaXKWMKCZhhW/of
ConLmr/VrdWo0eKKMhEkDWEScytYQBEZ7OBdsgGqnW2GqxQjVn3K5oJ3yxhOHLH8HVtA/vIIwaj1
PKIYVXr0sYlXX5yICNvSlHB0mhucUizERxfsv3ciH2nWhiMVbNJQhJoHsMErodKLIdLb7KqrJl7c
Rls4I5WeWfJWV6WD4bm70966NuWJpO7Y/+ow6ERpODqk+e2W0GzlNwnY0T183NztaTj56JwPW/7z
KNmWB1LY4d5JqnJZR9Yk+ypxYRUm6Le1YNiDwyjPdL4WU1Lva1Bo0TvNveUwAS1QrwE+6qSPnvS3
qPO9lf8p+U/X065evHRWLI18ICOEUs57Di0Aw9wH4VYtI4frw1p6dtxu+emWaq4vhVj5kR6Kju/s
hITPwy975V8RMngPohGWqIURLhEfjD7a3PgE3CwjddY0v3BRrRD6fD+WQsEpj77PIF1+7EU/+L72
lxA2QNw++++jMIVTSnwJf3FUu9kwVN+3uhLuLcFb7RLIr7/EY/HEZktWitYw6oSR1HSg2Rx/H30L
BPVI6s5WMpqydt0gvqmlieDTcTzGrn6JY4wEKt23b6Dzyq3eCs9vstV77IC1Iq9zeUEGQeX2goRZ
szwyYJZRQYMctbhFlMKTWWbU8XOmXu3CtHxBVZxPN/TK5dIaqcaUWSuIpd2/ny5EPfqgJOhO9Mps
kjD9TbNFy03ni6W9om4E/sEUuainbhQWrORy4RSIVdWi6FqtpPkP7HDpTm2MtiyVrH9JkdiMNtCd
XayfBvJ2yJwYBpIy22yMIOmDrB+UnrkwO2/OTeX+ZDJnALB961qmKyP68TJsr6bCd+F+UDA7rO4k
kGJIVIXxFctH4CnQnQ8kyhvzHOaDJbYvZxg5gF3DyPnZ0WhFhzTaOGkMQ2zPRMoR3RhTF6NPkIj4
CGs2kKgodHZ+yocr+ufJRAWnQ+g4dK/DDkQwo5eXnSWRzUWs2xNpmUNJ5gm6UxokpmdWEcwM8h7K
HSe9r78z1ri8YxYeJy8Qvpa8f69qAaNroi9FjE6ODTJWn8XLvgEOa7wjx103rpHThwsbgtG5vmgf
K8Ryarv+dJZnNZ+BNBA3VpjDleMsWkJ/29TcyM+nHV4/gsotcHRfBCtlDesT7a//sJ6RNsEilAy/
Ozoi2F/aVn2WTHSCcAiFPXas1p/c68ZXYrlgZedIkVl+OCL2vAZBmFLkE9EKeVQTz90OX0JrewHJ
65hA6zg0RvfATBB6/kUm/Mz5as8xXO88QTIABbHZYle0cm/9M8pcLC3XkkS/y/Y5+8b4A+Esp6L2
UnAltKkB6obYci/Nq/e5Bz1H1U+jFCQ40K+yTpbjsqEZqPIPW02RQQWYSK60bchmlEWdHrSMiP3N
E5KZlmaVCDWiohv96+c8eeZvQKLUK2Ks6bXdk1fJnSYp5RZoSabCmvnDuGQ1t8Nb6daFljFonX6n
R1/X3XAK/IePa1jFW6AfUFJe1zFAe1Kj+Lo/tHxfwrlvgj2gk3CDM55oswltjeRixmNyVaE58hEs
qQs00d8r1ea4EpjlsCOvTfHMDi9/DzeMCcqbtZGRSdjQ7TLFb5uKeWJ9CyPcSCmDy8SiVw5+hcqB
3TgxWFbRRRV7R04X8faaWIPCdsolAVwG0ZJPILcaY0Ou1RbhxXS6jBnpdNEmzfWr82buIpEpDq8Q
kVz5xE3/dLV44l2hNc18q8WvsiEk7SusLDCFaD2oqOBLNomA6gxZfUtXwQjhdYQjmQ4qnMLQW9Pv
WrpayEonuzRU5zLkOCt7lCbu5R9ZPvbaiLdQSSeMQ8x7k7+yIsQVkCPZgyjxNdnMSPKx0w7X7Pvf
NEziAhaGD/U/BY264bEC37LfexQqqYRHhhJTOZVvERWaS0lvKn1lNtPCWZET7t/SVJQINJ1SdY39
4lW9UZ8ZpHAE0QaRyZ3roKwC6d+o1RkYSdQOQ95h/6R6T+Q52v7gkjkl6cIxdprs25MyygzrU9lk
P2i0WfO1sucr0iv5AC0t8uzPD03MuadjHDe9M1MFtAAkVdXEvmEKWReHeTxJsHfw9cQ6ILj8PnZe
IzFsP/PfpKa5FQkFa/53MYV4zlx0fyCXZvg0+YAwR5nMQKoxQ29JKt+Y7HsA463pCLIUcsp1Wmyk
w+dpC3TZmy8NT34jGH1q5CKFJZbj/G14iFnKg5rAMlLdQo0L4sdDg/k74KLavqMX1WIvpKXV5LXI
sQDQ5kgviPqIbpubxCdVgxptJVhDfY2AhAFMuooMgFvtswEjLie3xVMIdjLzcFnFu3HftnvYmhxI
zYNatUr+dO8Pmf34ezXFBwCFY0kLC6oA1iZvsBczhCdAvrc3GTZQQK5rwLpPXLCx42llvhYS20QB
QFXOHhGOS/Zr9ontfeAyJ4D84xwhtNIt0+eHBYlM7eIz2LfXNsAo7S7SDW2bTCyrn3PX4fIIXPLX
40yzeGtSINerFllDnI00qQh9jXFO81fvqtSzJQB+KTrr2d81+HuhjSF9VYL7quYwqVJNhzkMpbA3
9ndaSmQzgNtO5wPGBBi7RcPjpTR85kEXmjT4EmqKwe0pRilc8cYRN8KZZ1NHGdrRXvgZ8kwGQPM8
aMQvA29LodCqoXl3Q04VXiGgnn2zbsEJt1XQ/KqY45meybQwms92T6O9eAJv+bJLtkOR8GEILW/v
gmNPqVbTd9zGbyFzh0TMsHjGuLSLgwm+gzLf+SvtZWjUDlt/TXu7gf+olXCWqrGIqopFwcqyXItB
zbSdh/vdrNHaJifQR0ElaWZdTKM0cs4BWJ/xLNVjo8rvtHjppBEHyI8gUZwN4UG3BBGOW1e7XmD2
iAezSFR8cLW5bA9DKl6MsmJgcps0bJfA4rjN21cBmX4lOaQI4BLuZTpFHd0GD2HBmHGmUI+ZL6I3
bm8H6ASWEC7r4pWNaSPd8DfJv1Yjn3raAXpxpSDnurlGYls0uxFb9+Op+zlWa6ErslWM5mPeeUpA
nfh0TgwHFNo222elh+F3R2lYEP0GkI2HC7gxPxrJDmFxi4vKFcze7AuS7qIY5sWMKaYD2b2B0ug3
tgTqslfaCCRd1njO8iNhOubncKML0P56uyAMemVaRfMjP/LX+yR1RRNCGJ6gnz9ysr+A6CXZak2Y
ltYuu5LWsNlGJxQEnbCqU7GztrHNkkv2XcXGbSegAnDiIoREzxTPbtPx5nUnX0lUzy0XtxJnzcJ8
FQuPv31bhqu352QAf05RkvkmLfzxvf9jypcs1ydqr27EMiNX5M7cVSNK/vzpoAewawPPOX1JYb5W
RuRYYmp29r734ShGTUmyIQCPFery1B1T2JaSxAV7UB7l/0mOk4XwbW13p17qlvjlNktJuKfRUE7j
yXb3UnIcoh/9Zr3gU4O0FN7WXgNnOaBgXpougtMnT5viV/h8KFcyr4JJLuVGBt92MWX7rfIL4VsY
uHUChTrsF2JHsi/snfbZCkLNgrxPOWRaSg/WLXSXl/mWc70ExpXDqVAM//k/rGJkrT+ClbV0L11G
Q/CvErtHMuUe751xS0sby1mSctJnP5LbEwqHSJUd4W3cd6mIhiFGKEVsKqmEPTnog6tM200AZQZG
EIXxaGLOUczoL7GMo4FqiVV0nvjU7wfuFYEbNqAjzTVJ+UhZv1EPtrePV3E5icBNPFze9o4y7AMz
gIj0K0JpG2kWb6HmK9T4Slo4ywgu/ORgQpO2y3TFhQpsuBpvCj0sL+9VrCR6M3qjaOPJxT9MYK73
7qdAayunKscUk7GNL9J9iFlyYM0WhWo5awheIeGUruGs89VTxubHwrYltfNgOB/ilsOKctChJJ0C
DguELhrr9XOGI8aGgQ8ed+wqETKcwrxfIR1GY1idtdrqrtIPlJ9kLtls9ufx6kZ1KnlbPLbTVvf1
IqRxqwORutvZCB6VY/NfmEz+xB1o1x/SiSLfdveXCuU8FK9Tf8PQYNaLCXnB9ArL0dlOIsZpqn5X
oOLk3T5zUOE9NAT+o9A8g4+oO6oHPwC2u7cBcxekXTqKR1aPcqWoWsSz/H/Nso/2qOgvsYXlZyyT
BKB1CIFSfT8RtDjzemw7/iFYj49jFUHPDOOXUMPksiPwcZ7W1//0SrExn9u22lxiwapzDgdpMjEq
3c8P9SBFP05+ktRFLsDNjBEfG/foVsOQp9XOk+036+xIZtaVrWLn+Rj59EnDKrKqRyZ7kwaJ4r6z
CSvFc4s9rKJSn2QIEdkJrPHs5q69ZEvXEv4+AUursuR3WYNV/wuPY0aJ5m2yc7NQ7mrvLEBLqMPe
TmEcJjvkvd3mkkrysHtdGAw3oTXWAa92w8DdwAqXlyaam28Km/uTb/w0+qwiLoWYkYNQqZo9qjPt
4XmzWdATCy1NEwJjT3Wz40w06rrLLiIObl1AaX8fbJTFaatvF51y5FUPadyjMK3LN6FtN8U4kqVN
oJZtEj4dmXUDfMQ5cL/FuySmn4BeOJirzMNZkXys0WloLVsU7M3a93OAsn/AgnardSNrmKqVagtC
rGFuwOTFMUpHpy/EMFhqTUSF4end/9KyC3bu1ipTDj5l/Sdhv/nfIFQVuh0sPQHTMRwmucHa9PQd
zOjbWowtbRtp4GzZjU3L6Aq2royG+RQjMAHvwFlX3UkALV65zl6XmVqf05A4htO/0yIxu3OZ71ej
u9ZeeBfwefzNU6hE1XxBkkAxzOCM6a0jUadOpqd8mda040jLPTOEKmYJ2ODbGyKjRpPjILe4FIAP
CLwI/piDxetvKC4iToIm4toJ4RLe9OLrKKOhYFYa057H6SSqBNd3Y9xCY265yHsHk+7KLBBqhb3C
2d5l3gVGbvLmGL+pUasgXxiiJG45T+SfggHyy0ELTy6ysWYYVkBuJSRbz17m+I5UU1Yttg9YX6ob
DpM2dEWlrnzNFwq04VVmSdnC7E47jGUj4vGGfSORV28x/TEhc21zgpEXcoNwNYLuJt5RH3FvDL6m
LTDGdCU+Tz0XjGqpV1SW26CM9/sav7GjIluf0Nct4lQPfQ1x5bQXFlF6PlBjQYI4vJppUzyNd+U1
ReYF6C+oUyQ2LYHIeAs/sqr+7f/gYN9FCKkyCkrwbC5VWYwELE9VDFcv6UX4AvxxgPHAkmbvnuqX
2QO6yZEFmGKWflQ1S8Vky0B/VTXRrrf/CFugxpr9al01SSyblFXgayn5lNt36+KVu8b5r4XCS6Ov
wf8aXKRYpNjaIyS3X4lYeh9lPKlXUjhauXQyt2v16ty/0DZtgiwGMwwif6PlE5Z8JzOqIRGrtN4+
cjA25sm7M9ycLc4CJ88bNrjX7yA8GOtvkMooPPseepHboY1818HbsX4eChmQ6+/KCT9mwswNWjsd
cj1h5Y7IPd6SzklT6YWSLDJWW7pmmQIW37rQ+paEztMIbIQI6UDyIuRfZkvRl2Tq/RW5ziUSA+Zv
YF5FV0h0dkQwCEcHWMWOWB3kcxv/WlgBp4lwqFo9teeSwxZniAHiTp6Fi0BCYAHDprQ3iBBdmWTV
ENPFdcDI/fgGD7QxixrqJc2EakZu1Xm4Cu3v6wYBcTIViDYgacVHCn7cR5KTOqeaWUXfCVEPCFQ8
csRh/6yIAnKx0Dyj0verCcSzIwQBoOlBOXQ7yK1M1UnTG6RwRwiP7+6l0ta1SVj6PLm8Va9oxrOl
dK8a6dyrJ82hycx21OYz+dWIeuNF0HlnTfaIARp5gY7x61Zy60vp8p2Qjz1rPXnN2Nu2SWBwhqRW
qeneQW+64pqniExtOgr6EV+/ig0Pk9vmZGrCVY/V0Mws6V0woi+Tkf0xNhl0X7Eb0IT8c9eIBf6F
HzHeyhmRIWN+wezILdvqvwyILsPsH/r/vvTN2rJ0b8DnEZzeftOHXp1uSDYIQtsFsC3/s6I0isG3
FyjWXbWz3bn8rdo+ZhhZJC3cgEhYAiH5FdAstHn+XruJpscb5Hz/OkXvtL+hLbiBKk0wY+mgI41+
Fsq1VPTKJEUQN+raSfS9yv56DTmVldzxrfL9PkC9nAP+nMgvOZyQDLHd8ano7rug2EZdwmklO/8h
fo04lOS+t9j6flTa8BbkJubxww1j6XBiUTq2tXEpLpC47a73llxXfCytBNh+r9gMq1JqM2z/zo7m
HvaL+fFLFezvliuOPom6wCp1oCSgIxQOfVM3O20y/t3XUk24rStD2aTmODjq83cOw1JZdqwDvLHE
t3Eq89fyZafM35yPE8Bjgj08XDcYsRjYT1sy+dTd4kDDNRNW4zLhRgXci/vAb765SozLE1g24QZp
dR+ziP6Q9LWyp5NmwoFlNAfg8xi04gOo4dqnCpP95K5D1LMzYbjYLw5jDSFd8+khgIGLNDRdelrM
sXOf4YmW8Zn1+OeZQzw6qd7StX6MkGo3KrwyzljCiQvr+dr9LxZ5BOdGn/eHJX6wf9gSxPPGj8Uw
Rv2HhTQGMX+Gmm5zAE/WfKZuR92muVo8bdFj8UBVOTibN5OxSZ3jNsNLwL7pMmCEPkQslW7UUXSO
h6v9yIMBbK5IFQiNikJPKuYA2pTnSH6lTlxRuv74eLoKwmzLpAeKyKl9tgo/1KSSHrx4KJgz2ZMF
RyqQfAjhZg5Ye8FZFYC3TJaTDW3NVd0xaVt3TJaaZ5icAVLbZCFQC/2hUOX2+l0OaGoiLNjX9fGj
TaERWWpGOc9LKIYsE5RFTP9R7O28KLMfbbuDdNBU9zFVHq2ticYlney5w1mbn0YTB06KJNLO6zg9
VbRyuOWXe213obgdOCPPtKbM4PdUTv0u+sDSyCxvNCOejaVYBPM232Q62c6oGEMUeanWWSeD5yjR
1+Y3XFQ+Zh3z/xj8u9jfNMFESP6rqi4THyVyCFSGAC84YeMN0BpUlwKFJsCAaOQcavPoTBDPVyh9
SO5t8HcpydHXr3IegH1SJ1Ilw1dIu+CtDgIkg46Xvohvo3S5m4+jEu6HeRX7aAVXDLZ4HilRM+ke
3sbGQ1/eiKgeHIYqlgtBaMXhzeRYSR1XeJ8haLSlqBwzTgVTvjtl2wRV2lBpv7p0NFMQa8e1ELdT
IGsPNeMaCvwnKeQRmrXW0iF54dBmEcuQdxZu9YtMAXi2tzrZXnSi8U007dVHAuv+m2utpj4OmCti
7hjV2eyUZKOKlqEc7zmxYZycGgNkEaIzCC+bdISs8qiCUgBy1Q9i+nb2f2jY5dNcIH34ehfeJbJn
GlYs4LdLmpSp9rVCBeBtJg89bCEQXViYUi/nPmb6NUe7917ux9LFaELN6j6ch9291wWanCNk59Cn
OEGLhX5cRQMmsP7v0nk41s8BK/SyGrgQfVzIlz6O4Un1Vv6RCywSz1uyA88gr4s1ixEAB4Nauenx
gGPhdf/DApvvVEhr0DS5WsEfcOSJ5SiQWXcJ6T6iK0KJxqKEfkW2VCGyP3RSxkihy6HQTUzuih4N
0NdvDfK9GYzMk1MH1OoJJwD2OZXUjSIXCfuXr2+37SezeOYgsEgOXi1yJYEMxfw7OMvraFMT9n8s
o62Q5Y9Zvv9fXl+trOtbxRKZaiRNOJgnnjsX33k+2qd5keaAH30PHHlZfPdFpbm2yt55b3WnfcJK
ZsGcur+MQJHxUf6582OdE5Y9pu5aLeoWANObzTTa2w+zlM1Yu1gwjjeOulVffh9edjV92u7Mo+ry
rRgEB0zrXTLzf7ceTcwRUBb+VS1/9fZhEmliObK5rTpBO79yMFy+zWwPzbjLcqyKX1LaGdGlQ+NH
qW6ZMUDj//6BDFxgYCOm2TrMTtMDinnVOtLdopcV8x17SeRWq+YaaNtOv0MfPnFcDN9JpGrJS5Av
tOO9FQW+AAQ/VgMiMga1JkK42Tjv6NRco1Su57SH6QqNX6ayrswW0yD/Du92ZPlRfZTl4157wMgh
nAUVrF8UjY90he5NnAJFNWKfy1QxwWrIh2tiSIuYFj4ZNOCs7u9FCp1rldF/3QabcLoCg0EHKx2k
015jkqQ4m9N9x2Ygv3yGBfOIwpMJYbA9Gq7g8pMoH6HCiJ+eG2N4PsxyNv1WhtTZV2xjmwWhwi9C
B4caoMsllpWJYMO/E5rRFLsyNTuIxnTD1yxARsuUw5X0kaS7RlB9X4nYrov2GEOKGahtdY22EWUE
uQqM10jc4WFmiucF6v2slLM/s9FRWRlF3m0nl0EEWvJpe7nrPX8kune2OvA4u66uXD/sl9Cylcpt
5bvem+58u3H9hvwpVNyy0uf4t6sXsZuViuh5lTS6cv3pk+G9jZ4tdxvS5ZnF91SRlLlVBHJEZEH4
5h9OLfciGgozLo/HsO1B4BACjFS/6uK2xIK/igO1rwnGncU6h4qIRe15cT6DEBAFvGqKZ57nMklO
rDH6Oj2UVKDw/TKbiJcT8HrnR2CpkidNfw+LWnEr/unyF6UyuT9b6u/9VKaIgmdbcbPTMhFjm8nj
BlLGDpp00Qx2qY/3XZ7j+0/bS+HrX/MtGnqQo7UTGAq6mtGl+DEp4QQMzunlFfUSyRo5Q+nvmHLY
iOyNQyYYD0yxVgZtFak988HLtdgPmf7G1eBDj8cPTxiUZpAqbqt1gVMr3DrU1lHLiUZmoHL2Y9P8
jinUbJTBgkpNP3yJunf4QHYWlMh77CRhayLHZWR+7rccj4AoTw1/fmtGoUgdRQSWYPhweWYRISOb
OyxsVcsGkanbaA3IzOeALAE2J7wNjIZ3l9C9PXv4L5mt6k90/poeJbN3+1BHsxHB1KCgEpx7RAOo
ADITDpM5Yr2SteReWx+nSvchb8DQMcm01idCF86Ekk43pv5U7bGJEZsY+XVAvPYm4mcUOCYPhZBz
crKRpoN2rj8YKJqoVDPRX3tuEa5cnqocFxbXHrZLDnMJe/d+ipSxQrSlIUdYNcCH2zHt6q4Tc3Ki
EjJ9xDpdai+ZAnNsq/5nHVZzLx35bgtQeOfDcqoqD10Yrmh1TGYlFzY0Gf/ikyp4aNXW0fh3zHKx
rkUgOwCp5KvkRIm3wlzRKjA458qYZ9J9l4cWVo0Uoa5EVy3yboQC+23C+w5l3yppiULjfs0RM6w4
pQrHtDu6HjXLTgCKRrGCAsXDaqcDiegCJwK+BZuZmcsAxbHYgVbQavSBPycctkNfDoRnq21I9oul
zsB8FxrDrxn7P92+r/B8BBzq3EYCZ3XsfAspocE7lrrzlRS04slibVZZSjLgUjRSZXQq+NpnkiIp
uJV7cpuT3PxmxsdYuZLl0aB4Hc4HNLWF271QlOFYwBgr0wSXrLlU3elnwvZTusmM18jKMZBjnruM
SASCRSOZbHjBkoxEqmR5HcWhv+SMjXDTzVpo7kxw0hSd2DvkbFBMAMaZpBJhA3d9NGEi4YCCQc2p
x/VULNEs7ZhyG6zrr9XkImCIxwXBBkAKRs4zm9s7cFsaA9rhb8F8pCmbRE2qMr/T7AX27sXJI/L8
wTis17a5FQh12c9aOUGLnfM2KiAaTMAk+zE0m3UXOwQNs/JyHB5Bwy/SUW/yAuBHIcVSX+TEQtKn
IpKeFcwErsQo+vWOO+ogAek2Psv01pUPybFqkIpjmPJ/FydZs1n5x7gnjc4V7IHybU//C56BF/k5
Si/pVBYytO6Y3I0P5uURw5EJDyQmA9fOJfKHJvvvFRk9NxHK8OiIVmNZrn/FCtrGmxmC07E7Eckj
G3C5w7YgLDxxLzayqYEe+IbHnvjBHdEA9T6Q8nIhM35VJsTs1/kg2JEggTKIVkfUZ68q6A1om8IR
yGgHSEEENAyaFGO86NKJfoDuob8npPNCFO//umrG82u3ugOAKmb4Y2zk57QaDl9CVaOjjFmPHOMs
yZRmeIE3cuz2l7w8WGryby7CWmJnMaRTHaS0YwE3MQuk1E6Gy2By5UD/tLc01DQXspGHkEz5XfMp
7FDLgFUOXJ+2xjAnLfGRnvNOnra4BphSrrmhl3EcytRLRStXfhkXHiDKLz4UcsvG4wEcafkIvBqX
dxXA7E7D93iqBhc94etThycOhB5MevZJSotX5d/tw5OxQOhDpCdjbzub7dmswayzKht7MLRvAm/I
Uz32plSDZk+HTvqwzrKquAO94JLynFxSqh2DoySfdYu+RqZ0/rUSUIcFJeb29B0UcYbBzjA9RyN1
jVmqw6LOij0ExSQLRsyMgSTS54g308xaS3XuLuonFmvnFDIUtWg5YiETnMnILDyH7P1UWHrtEbc2
AsqvEiTeAgriAznyzj+IrCCmX1UbAPvVE226uqsJASe/Kvf6Svgw2UJfXXXDyWqFTtN8M01AJA07
9BFnKn/TM9V6Lk92HWpFuuG0kbiZsgLGG1b+n4aClg4NLZBDOX8P8aQydTbD69geR03nDyYeCy61
WeofGEpQPv4WmC2Ud0xRm8Ny+9QMCgmS8ypyefbbCCp0ros2dwz4Ibci8ddun2jf1tKOCyNiQcMn
AStg6Ptzsa1cNlTKf0rOhXd+QbgpJfC4tbZcADtW98A6McWJ+FeksgFwT7mVe9WsExtzuLKvaYZe
Z9rL0CO+BVVUEndH46ufSkY/b3ZqJn3appwfPlGrAZUymwnCSgo65af6LosDA3ZivTz/7RCO30kw
fc7V/aZBpZTHBPGW635/hETLLwApJNt4Vypf+LpRigUPLabGIuKQU96SlgITSAHS5olpUbeu//wh
jqCofR5auWPjANYRwadUP1v3hRaOlklfRmhveQZCUqZtHZBK1kOSiI9zc7oR70BIsBdzR5O8Qq/c
ijgf3MXcS9zzNtksb3mDbJ5jVNcYhPxxPu7et0xob/hky5Tjfu2xJ01G0UVQAlH6KZ8ZLcgK3IVz
HvVfTJ8e9oRntev4FIzpWU8ztrPaAuKNwUmXjBow62VbhsgvomUEyKYacpIKzmeMZ84eW+1TlCWc
roP+Z0AEI7tC+kKhDZYT42o0k/vGFpUv3z0nf6R9MEnL2+1o0pXXvDgYMy7S+CIZClQOHOpiDc+q
QEwrjkzVu7+xy1v5NGQ299sp2DMpF0+ln6jx4ozQbttdtzOhA8Yuj9Gj5sIqvy9PtuaRhQzxJfqk
3KsHHQaHvFUuvMbJBd9NwX8kheOAUFZWW4isbcvQchuibW098br6Qx5ac3kQ6rxgWKx+AVbVFIZD
YHW1Kew+kHANJWwGBEwUGWmVJQcVNAkeHly/4sxuhXnQgpQkfh/oM2tnB9ehUSe1xMB5Jx9+Yw8J
kwmrBUoIL/XsUu6vEyCuVN/1/XZoo0653PFZ85FuKfqImXPuVnzTLspsSaLJrADH+pSFRz/sbqu+
/XSctApg19WU2+g4QB1DgcBXRhMhFDkgJLxFZ7JlllQi9GK5FWqQtBcVHPpYeoPFpIF56xKxWsTq
P/Vqb2Qtsbph30WY1prYTE4DEQ58lMzNUV6b+jKOM/u1h9tB5HLoCJxGmBa4e2cHgA5T0bjv0L/T
tPB2U1eOZiZqUgQAsepKNHvGTOjqI8hEmZ7FrToBTOL181KaqkX6+9B9eIYqX7cjICzPq6lrrPL/
4U0JH2zhO1wJssWRWWPf7CECAwp8GXj44EWfdKgmmuIHeHiZTGYutt7BuyVObMSFg7PAkWDFZ32u
NxFkDIM020KgExFkCOSpyI6IL/CTjOblkQLlCUP4lSye5MPA00RyXp9y4XaAfsttHm4zYxY+rq7l
xfApeN8xxo9EhPXu4snHsJxEZryRRLs4otAEHcbmdpk7W2vBJwboR4vMp0cBSmRN3qZPzOEltrid
otp4eGcvLbNXisknNBAyj+rEgu9U8/a+LiWnSqvgdRYZM9iIoqOltuaT0Bzry4IdMoZc6eWtqeZC
IFaOTbzrs8ESSAGQ1pbJYA/QRVAcd2CTpU07A629Tqd/+scZ0GKBJ3WLmcy3wu1rljFxnthmd8Sv
6AEAL55eKleJPJqI3OpHSpuTgt2fGNy5bWKcDN96LLH9eXC0IghJHHst6zWrM+MVX3gKYaaAclue
dpyWtSXTlAwbNGiaTM7853McqsxU54SLq+39dtxT0YZk7jDoiFV37VHrkH5g6v8ggXA669DvKLLa
o7TZHE2lzml27V6svU/XYiDZTRrenKs91/O/Vp9Wy+QxNLYgvvcffpKGaSuTKL/T32isxzHQQ/oL
KF0a+wVxn86HZULyaK0oNl3hds9euO01WM6+T21ZPLo42DCQkNh6K1MRrYcZka6CF+N6hI35sz2u
KhSQRLdulEGcQXtQiEG64xb1fAO4MI0UxKyHFKAkCwn4fh7io4RoqwkLGMjDmTgppCO4SEHRmEsJ
KAtw4mFfHzOekmjcC9tlb1uRLIOnXyDgzvyOh5OJ3mKSSTmQewRVKC7kIzZzSkFjIzXzjb7tj3zb
vnyZNdZRO3lrHY6JWT+XuUlU2J3VPgjoXLqK3mgPnfivPnU7w0CU0hY2iByg3apEsCVWmV2bD3gO
RrzWtO/dRc9R1Rg/i5UqT1SJMRx0/khQEtz4UQslrO0KlHRhl8J0QV2oYTn0otlXHox7lj8lSp8p
vR7pKdV7eFgxPz/gMGaUQI2NUtOT7NKYuby2rioofHgq1kAvjDMScpvs4ccn98p/cN+XPpwXzdiX
l4KA2zVyz3h/xCIYcnst/YNF4AqDDh3IhrWssFBRN8rR09zJtlTp/LUvdzTaa6aLXRgKdf4GvSny
trwdGIhiRaY/HHABfnaC7kKvOZ/+2pEMjB5JJesBQYlDmt1yz5y89OJGCsxlBYdaI3PFxO8TGHOD
FSzWCIW23rr9Ia4hGD5pgVniV6reRDgDIEJmhAuZ9HWgz73ICFVFxr1IYURAmTdg1Yi66kk9OhsG
WI5d8WtjAXqv52QJvfaA0B0PrTDkdwrTDJWrInjATvSpYMVpdcS4OBFDtP3Zs45POfrHE7tFzqcG
Cz/bcBzqpePIKvkz27uHdqCrK+iH1Sg2RZTWGs89is7Sxt+ffpi6KdYrFOjRza7roh64eVRO2yoJ
3y6npq7fdoTbVpQe2wK3X5yEcGPXPhCvykoPm+/XtiPu3XS+FXnbSEMnXRZ4bi+TZh1WDp7gN/0B
ndAvMoN5qfTaoI5LllzzOnLkZIJmRcFvotWHLNpHBqZ16dEBWawCqNNr51Agi56hxRYLdrt3tht1
X5UHNXSZ9WLd5CvRmcHtZfhtc9/8zR9U3QQPtIxEBpFC+55GBumgfoeJxfgLGQR1tfUcg0KCuFxs
0u+FYvAgQGi1HQKD/PH46i+9wsr2mRr2BBRwdjFmwvAEwiyYLGYq7bh+zqubJ32G9qqVriD3Hzse
yIpEDPnms+97JJUa6xwoiUq+1VyQ+Ez2dUaOi5PujCqs08BFs+gI9ylcw5W7DqyET1Y6pk71Unbz
i3f2czgCB+WAJr/cLtd3l/Co3VZBKVJm7WFF7p9m/DCiYCebR33qRJi/gI3cj1PwkquyQ6dYw6jc
J8q+T2PCXgFoIZpLyscz+eJvJvJpIvQH/mKrN0WFTzeei8UCzax7fpzsVud0WGzwET25Hb2zY2BR
6sRqUBrDfHzlM77iyAGU2Coj86iFeOthFpxOZ4xHe8JxiHFBmckWTzLHA38izHn5tYz60KHt8gp7
DOmo0W77HdBfythsteAl0VRWN3ddAu+qxZeaf+HJAuuOf3cRbz2gQhe7mcLkYy8HSoJt7oaqEIxj
IZV5AvRHQ3YYVMpImziX7zUxQJhHTHKmi/sP/wTtxZy3weG4ODI2xpFySBfWEd3F145sgsMXVkne
h4Rp5t99cizU9wGoBPycDjW32Smtel/yWToYt2pILl6/QXqMQNJGDQbL179LtmP6QTAbI3ba+9R4
AAggJbCeWiLP3bXPqqLv4sSnMhLwk71nSdkiSWY/Kq245mE+QpEADGOmkqAW6CJiufoO7jqz7mlj
zYgd6N6kqzWN200Dj4duu2IreusNk5F3Zkgd7ALIQUpwshTsROaAQY4Lyf3nVg9RNuRoXgaj8NGr
SMkNmy4PzyTd2xOwwUbczQtCgftFIECWc0Pe8fnyt44hViFhRrhLrhWM91CCNaWbEMLgtUNAr8q1
TcwfgSIIgbHS2LGKK930AAg8glRlKm2hwRMQK5A6TGuo13r+f8LI0hU/zAqEAHZgdCJWLGecKlwc
HBXhxQuiz2E3e4ox2GcrbPrU4AsodprrQE+Fml97IDIldhoQaMFDU+sd1o3wdf/XxpXVl8rp3MN1
Y9NlNCeeaw8EBwjzxhPgRloc1YX/VwO//A5/LtF0EOJD6zkA6l7jr0+p6IVw5dRdwk1rYrnXAP9P
QkJYhPnbOYkKYGYuh7D5wWKnS6LTHdNLIySDWM4x5vplCmxzqOyXY1JlL+dJGy0mlBrgnwYscMat
Yz0oqmU/rfL7LpCWDETTLrhOEu/L8Sk1cas9JGqEJHxWMIdtCEpbehq/4im/JeapfB1+AS32g2yM
tdv5Rf3KFOtjpBOBAelZCwJFqOAauU2F8cGwdAbEwtHYjJ8ZYY4QqhzvE6i9SnQoIsPm5v2KoHua
+Pd0rC7Pjw1HWeawWl6iphqOfa7G07/8Bx1leYww6rFOQegx4yzVA1NOyixo/4kIIZiPHCplkbGo
68CF9cCpHpZsFGRgC/ZGs6nygiFmpb1uAlIh9B8VN/jTzsvoF4OzH7If/3BvQnVGW0psThAJp9a+
vPmZQrdtAG8sMDlgrGYZe6mxqv3Snk+RXBWjf77cCo0ZeaAQQff4ksAspVII9PfD+NZy69DLcaFw
JTKqE5Ka5hVzmkQWxSGT9pZIWANJmvPNyzBg1hHS/vjQa2v0rrSJ1xeGp5Ni0oSCe7HpOKncpAQU
3u0NR9It+d13FclrvkC81VYN8AIKVcMLl8czqGPye62nz9K8qULjTaszvO5LG4Dg7dSxgpFYo7Fv
1GuKaX7YmKlv2+HGna2Z2xxSobwxHFdI5GTmE3dmGMYZLIVn0roqqU6dvhaMAR7Zzc9AQsD168NE
PWUh37sIkE+dIXVnvcSQ1I3bRDx1TbA0va/gxMBHo/zgyRwQdwaghZyhR/ukEFNWx7J3rjWhVERA
4EM0Vd7NjNsFfOCHMjkzrB8z9ciU7MGfwL486u0+VS8uQzvEASYpP2J1uhpTQm1rzNt1Pc1Yt00F
ILwA1J8E+Wk4lKgVP5V+xPSiBul7rtWraFnEc+NyVtbqPRYjXJikHuY7YgVVNQGtw+tnVb3BbIEu
Auu1Z2QN89VgzlZImmEVNW0VUwoaaR1r6rot4/q9yHUZjq5bHZFLBdMEjdIIgCm9uQ+5dxWARDOU
QDI6pgikEL6YuqtZ454vNODO2wq6bdS9c2QlMl0O68VpbEOZTIRx2JLrYpZvIAj8JRVpDrxe9qK7
fFWcOIaowrYKREcExfi/l+BSnsY3U1ZHen8vaym+ZWMhq0IJWO8K4c5Nt5Ogzl6hXXwG4u7pwgWb
WoYywdC9ssfaP3ItsA9Gdoe/jrYz+ojAmkcUsedpZrM8wPlHFCwPJLaNCSrPnDKNE6sgMqK0RGDG
zXegxRhCXWQkEYrefNiMWB9JyGDlX+0/LqzorarTsrbjRIOQzRdQWFK1a620Y5HJ3IXyDnAAfRFV
hfHV5dJ9nEs+TcjsaAI4Xp+DsTVs3FBT5m2JagoSU2TsO4MN8jQlLHmHiNsCckAp9GziHLLsWmA1
R7cTf4m0Py4lT0arsA8+ytHY9h3iyuLiG1dx9UZRW9c0grdIentlBjVUVaGxY231rblQ52S8KzsB
yQUcvBb6G7Y+KE39rVqttAWUPccyWMN08h3GfTFDoOvKx9y6xJUIUcH2PCXnkLcQca8Oqch9QT5s
lNzVgZjzjm+zbau+kvh767jig9akCc4q5hlm8j565RDnwtkE+TTgCaidcpo0YNLI3RfppPMb+uf3
7Mehlv2eYN507qT7e+T/DSnR0BjJ6n4BUud9kDnvOX+9NbgIGJSWiYuFhPRyU49exrbi+zYcJXxI
o9dnA8SSoNdARhtdyxyvyyVy+VFtELH+vEJuc5++H0yJGfXBb/XeVACaSp6AF3LtkGavRD+UUonK
f3ntUzWJdgu4bJo2rkJk0TlAyb0QK5YKa+wExWzdoKDKZjdK1m2PIv+fo6dxlWQ3LfozFZZrfT6v
6FD3QzJXxVn2kCf0eP/+KO5yHTURZNo14ZrO1B8j8qCLGKOLu/ztEJCRUXo3AzlcIDnS4h5umvzr
PX0oXMbFfmU3elqqQn0rFPu780PjovRD44pOnSxeGtBqu8L9tD6Z9bKdaDJvtRfD5NSvEnA0otS2
NMYn0S87DiYG+wXYAWXq50KGj72fC6fu6OhQPoZCfaWkvodK0stOD6zgyEAG0msJeVIqQ0kKtvYe
R6Idn1iN2ztuGmmF2LwjVjKa/C21RzQKpe6JEf/afMLdcSsPEt9uo4GqKh/4fCVF95L2+zjtNYYg
SPXP6hkTCq22A6Qnp8t00BghY53XFAk+TU/U5KBSoIRpGKfsCppl/7glIQLVlaMs4ISiQc21z0Bc
5NfA+/V8xIAunS5Yj24+KBYAlP1u6ZlAmufM6i1THnnLCG+BRrsQuOmrXky7Cpl71fQ0xAnwqa5n
dlzNKW3QbFIZ6MrrBlEwsoLRg4AOKbQECKtG7zbSkDz67bZmvScokjjqM93RlFw5G9S9nkMxKnOv
cDEI+yqTQMx3WWtap7x5n3a7cc+TQ0VXtb8ii2/1C+kYWft3bVRos9B4h52mggEVkXprGQ1w9767
+cSfbmjcmCi1Fnj2MQ49WtXJ1ntWURm3ktVfgqRHz9BUubfgpkcWRcG70QFMottbWcWb9a/wBhCa
mwiJFbYe52h9F1vuAo8GyajTFujTQeCyWWOQCWrsAS/nucRQNryuNTyaJBjl+hxPhK3jEXjKmQv9
MiLwH1SMgXC83LyO1+lY/xaAx1miSjIkZ2SH9e1ECeM8epSc9wvC8eO4v7jgerjGAg0S5rxVlo3i
mt6RSSm/bCNP38uHSOLU4+h85zNxQly6CrMIQ/8aPABhBBFM3s5crRpd2JGx00IyeUzg4EA22Klk
VnKiek+lvY4MzheRxRCpuPR3Ma0fVAMsGOOCvb/j9NQ7KBz8azvcMj3Aa80CzA4P0n8047aQPiBZ
lfsxpthFN0qpk83kvxudRA096w9c+judHKVE5vqCc8lp84jfArn1NqyAzxNuTzgNbspR6Fp6ewwg
5GBzdgBNi96A1gxfN8aLUrgpZWcWXp/6QS+yHck+vnyonBTl5dSzq8ccTbz1UOA0yhQLUY1+p6QG
mFYRJkO4lCnY+WyxsXzGMTkGI0PRAwQtuQkSkMTNdCuynjLmVWSJlJYJfK8tLCuC0MCKQUiUJset
grdVbal4M2CrkKp4Ianx+uy5CPTbxUq19hbvdbQP7ToUvBnZB49bvTE7NMtrlwcwxH7nHgVJFGD+
ow1J0MhmDhmlERghypCa6cMAqj2nr4AmwWZG1g7+guhSXwDPFBeEDPt5dTr04R7hiPEBP/C9C9S4
ukh/X/fz6aaC6RygW/2NU5nSuK9IP/TULQn14dJDkr4KQKSmPsBmNKf8waseSPnnI1qVTUHnAt3I
WdzBBgt7CGqNzOscLMeF4wY4imGQCPq3EDwuj58z7okOIHcLKISU4fPquSOmnBZYrejoVcMyb26d
YwsQ7mmDagHbwTymjOsUTjpbDehvQHaH/drNr5yHtOZvp0ekWPtmGbdsNm9/Ce780ciMSBN/TuYR
BWUer6ebmQKyRevCB8d2mebfJPorbrV2sGu9BENrX9o3PFxqs5L62Ur1yb0VlXJ3dSquWeGegV/r
+qAiKqJ4jNATZfKY5CxgnrPlEMefDvS71kBDWfkrBoWyoWkG33CEzme6CsaW2Gsi+GNVGHcbsZ8X
zApnAEbQbBwEe4tK18F7l4pWF23L5uplyr3y0ySsk84cnsSAT0x2+GaifuidTHVYpijiLoB58nRX
9qOSGYdHYrSZgllHvyXtUOJgtbjjD3PqR7OPxqloePAy/q+lBSC3y4x0BW1ib6tXmV6b9yxzdqRS
vA+RlZaD2ThJTrmTRAtUDKATV8dnaq12956yp75PABQcZrqnTtDAkryLlb1fvSiBBr2IHsypCIA2
L+O8QZOIuC6tAiVWZBztGLrH4bspMSPCNJ8giF561XhY7oO73W13EWfkLPlR96bdxwc+BksIKvbw
VuKLkHW4lmTlqUvxiUyW5aEq9lY6Dsgp8aDd2r1gqQK1V42CvoAvqD7FBYbYYqtwM2s42iwXSN3Y
Fq0EednMdi3TEGKNtM2hnvI5HkK1HIqvZV3wj+QXyMO+m3XnqmbSRNMTnu0SNAkpKqX9lGIdB+tI
2Ta+PX4pfGz06u+yw18GQ9d99bTCfaIFXbR56tmAisheZ5KPTlOb0/AWmtoY7yjeNUIozMiuWBl2
2lgEg8EMbsPIcmSwSRE1IVTP+6UO/KPWMOofdfGswgG2rb3IWK8e7jSiATuPKSE2OIN++WAbSoUW
3sQ6swYIuuhtjn11UZPmLQtPoQVvSg0ERj3958XqawBm1HXGtgwc0DiovOoCE3yZVfS6jeanHMud
4kVlT63H34TrE1o8Tnly03+8izClOP1w78dx5thJSbsx1KQ2oDxADhbWLCbWXqVtbCU62DSBxkvE
PEs4eNmxCv1P3pH5Swvq6dzFcBX4InEb+HaBCztgsRHlDxmCwkcjr+D4gQ0turtpH9xq6GbhZq4Z
jU7Vls3xZZGmPu9PDNJ5XOCI3h4599lqF1bGmrIr6eFzCwq7zs9p2CvI7Uez+9vrGyfBptXkEcFZ
OcDrCuCYTTruR3JhkUhXPPP6AfUHEuXxsaDDFyIFEZDnAiyaRRQcPq7H+0BYVUOlwKNcallZpIG4
rIT+83u0zBoDHQlEZufdIgJ60YBvSN07ObEs4d9Psxp0hUK+iqNH9Q6hpEPEr+kmC1S2LJtL77wq
ZsckiPDpH72CfkupFTzNXTF78EOPsTJqyvM4OfUAmn39MDnttv44HLX6UKUybqbCoyndi5T26Vbh
3g2WEn07+sI65FVTE3TonIadV4RqUJm0CfrYEZdKZDpHgnILs5FOlXDXU9vl6YVRXrbAmhtFUI3n
SLxw1/etZ3M6r+tqxkx1q0wzBezvplDFXyvWhvxTuhMVJBxl6b6TkNh/H36jtrfFcF7OF2wkdH0z
DMAN7HiYsZ6gsiXzY98jGbF++w5jM9Xxo6kHw+ucnOyJL0Tw+xYn4M1nF0sWdnf+OK/7Knjg7ml2
NXbcuJMwew6WptfCngoCBYkqA3DhBUyCEdgNbie4RnvaiOot4kFIb8K9YzuWNM5Wni7+f0aWxWOR
frzx0QjFx6XyOcnTuaXAYeiSP+xhYgoEikqWBsx+D2OQEByA33nK6Js113mUfhf3NDGufeUy4tNO
9gSOUGWbXiib6FyfMRQu3wWNziU5S4g/QfmjB3+YVCX5yZOzv1/jAQXmsrw96u38k7xxE9+N22mk
kzpA9OwFkTFix8iLW9PuXcY7JQmj+W7JfJ8AzUivCRDQYlLeKAR6DE6fOIu39RnVCZCtQAcMJTac
W7HjvOWmDKdOzvsseSccR5+rIL0Z9GXp182A/7oK/jSo1SWmdT/8l3uQ98Pxn5Mqb9ZKMDdWvV3a
1lKxUpVYppMDx0KVw//RCQHV3EPbxY/Ie1hTzAQHly67ujg+aleejFY63VrNiI70q6AdNKZ4J3sG
V6EzFY2S5QimEMDB0jjr66cFwnl9gsKEs1xbA2CXIv7LOhyokyP+OVWvjEpb6F9EggFZnZ3pg79p
Ekz3nDHMO5KDCiKcKtQkqVf7LYkOugyS4fs7y95oPWyyy5ZEHrL9/t0VdAKRDmVlNxj9uH4AZvZu
/sIdI4ZFE51lXV2raL/vw1D7wBY77m8ovFRgL8msEOWHdX9Ym1STKvTEesKKilncW/zLVEsW2B0G
WkjZNR5M4NgrjlLg7Kh0XWv3p2cM6E4lR+eCrTIFPgEjgUCo8+9Bhm1GTEwtJRFuToZ/lbI3Ty0H
uwl7zrqIP4lLdasvmIep+HR1MRvwsSURvc9oDsYiyJBqFVRK4xsHdeixgN9Gm8OQFeggw817uta4
rNVRt+JsPIDepHus1oPTGma2kiN1U6sz3XPaItQhIjreSY7JLsMVt8OJKq26CHB6HnBhDgaQiwSz
WefTq0YUaQPNgC3Kiq/Wvgg+B3C5+mRHC17m2wx7PSwHv/xiglal87YDbV/YGOnIXc+3/H1qJb9X
8Pm8f9g0MMD0AuIS1Fox/1dmb2buSD935RrLE46MpKc/facQDgDGg+O9Sfjaag9n7pH33CWp23wb
u5Fmv+qTJaI1bvCnpBSDYw1ztxE5VIWzBftWqXNAd3eqRYB36xop1M7+asbX9eNFYrrg26im4XX/
G0hRCcNDEmzJ8SRZ6jtNVc+i7EEe2li6SAgdjT7fJhwoYunbqIW7o/Ev/mx9WUZCjPUBiJx6UEZj
uL5ZpkKzeiCJRFvAhVUT19tVnf0hcQxxnJIXS7KMKftkFOWmwJ4c4PxNB0lCWH7tBCzcNf0N0ZQ5
vEsW25pH4lEPqLkIL3C+ZhEs/hnWVIv568I2rocMTw3ICfPJ5FupH0n7Ig9JpuknRMqzEYL6j8+Y
heKxcstlRvIz43N4Ji9tDmaZQOMnIjW4vsVFfZmMZfoiJBK1lAiNjMjd1ybNIDV4kjewLxCti5GL
bI6EqVjmv5hTlbF4wk58mtcVnebLJkqYSwsAFlP9Gs5SkNBcFgA7uCKiguumhQlSkvgtvTsZjFSv
eTj4p5GZEMx37uC0toMqQeLMU8HPyOS7MZp1hm464k0lVjdvsvArZ7OYkDwVk3avMTtl1LJ2nhda
ldVdOhiMEJTlLMYZxNp3A54M8tDwhqK2izoi5m4TMt0eqUR8CRUgFyqgul/AjFJ33bqp4sMzNYHt
4NRHk/eic/nsDxhJtTTehtEhJk+i6teLjIyMo9jzUr0OSd0ff4lQzOO7v9T3lB2xE850FEiXCIgr
brjJfJfUW6lCb3PVKQig91HIIm0XryzdtcK0O4jPOPl78Xb+zalldkhW7PEgyq6KhfUEaFeJCQdP
2SCl0zEK25Fsm/i3knaENTSFQt5bvkXJNkW0uPpAYJnBJ5WE8cwcBWWLiOG10IfuXyGc6Bto2JQl
tCkYNHMSD6x8azCwymnxWCdLkkQWtD+uLn0jIEia5nYDFeg5ja6RX6rL6aZYkQah6xczOVygfb7W
wLjQDccg+7uq9m/Lcjj7ue+bXa9D/0XAqXymy0xsxSsTM9ZLbakMlKj6U36BWLsUvhIi+RpQfw0S
Uu3rA30Khm0TQ5664JgrQmr/6dMRB6kJd9X7khtEsVCrvi287NAuNNfWwBuSydi9XAh7GGUll4hB
W6lV1hMZOrNoK5CL6sK4/QyBl8y8+Ud6BgSaww5qEOPynFiQIUz3KS+Q1xwUlVZzu67bp1pbYUfs
ePtgs2RpvkFpZQbeX+eWXR8txnWYc/Avdx7MTxi237lHjg/OXKOEy6XTtjlSlApj+6+42k/oB/Yl
dEqrCh1LXFCCjdKjHSRjNqVrqENjokW7KLUjVEySNSs0RK6Xyf/ldvq2RXTv7wTeyimFwjWQfw39
boJ9L/9FUfX8oR/k6zCzA3B0PW9z7Dtr6izoHInUHWuAyrFsta2VyXksvWfNkNyGQFYBsR51C3dz
2nvnWRbQ2lVbcTLSS8Dmt+v7f50tefb/N00onU1iY4pS+1Uv6H+X6bzD/m3ddr/B0vd0e8IZ/ET/
hJGUEUkJBmahcmTrFgTbKCMdlTiXDMagw9mQFH5mBxAzy0nn9MwgObyjx/7D9kdgpL/1dFo4tMST
eIOFT34DU9k1eGgE1/6UbFzTUVzQsbjEg1UdJCfJm04duSwW6xkf3lZmLgEjy9i3mSeJJvtgXjaV
gR5iKT5P3HsVyavEMzoZvvhjj7Q61egdCwbbe+GujaYoM17DlMYSFcJ4912jlFFbeNhWUefakT8E
4nS6lPF+YxEw5M8OVK52ofgUEJ0uElwMFpTDJsz8hsX8KfcOIX7Dani5te25QFasaZ5wBiu8sr67
Bxl4sA/vZZjvPfYdpUVp8rlNsrtaaAdtFrSLDmuEBFqooONuqa1l60BTC7tuaV8xohqGEZgLECpx
kGrGFe6u16LACeFhzD1Pe2cRpus9yijTdms3t8Hdyibavpf+iAVigylAgylzaewoqMurTF0AZQ/4
CZEpgSBriVLT3ahHU0Ct2rxpbjguIsCB1D5gEn7yIwlllcUnY9cqF59ECeYbyWTaYYXzmkGbNTmv
BHL8hliLUkz9n9/BiSdesl2Z8aHpxXzTv+/dNCc4a/7yWSrThXj5DWJOpfMNWGSuAjslfTjVf9y/
xiEoe2aQDAP4A67cGOpt2vFlJ8iqcWkfcihsr6ZlLz8CnWvT95EbXEMLlmAGVbxRJVhGs5sJXIMy
c31q4u3bHxwU56ZCp5e5ybLewYI4kTrS93HFeFnpCNI5WiS+0FGgTOWwMZyRe1UE+ysvHRb/pm7Q
oHX7PgkngMyI/zX7zzpxYXEJoXAAdJ/QUbsP4AKs2Sr54QldqrXIh3BlQUTrBntNytG5DyrMjD8t
Mqnx6F7m+kKL6eV9q+GhMn9SkmKjZ+druYrmsBIFRpm39In2uCP+aoRH9RFmWfmjSdmB0ALaJuft
5rPUiwegbwANdLpxCVv/QjITj+V7x1TWGIi2Fru1+RDY0PJ2RoPeOl+HFFq1Qxwe8ICoP/ZBnVu9
uMLsu+4zj881uw5IqYgXDjOZcHAv/zK3yBHMenh/jBH77xHMCe+uOzKY0QmmoTIcMLS3MWZ40tE6
TmFHKfhslWcynpAR6pXjz7wOZYOvX+TevJMoEFjqsw0KP8kucWVE75vvl+OK7g5hoEnNW8TijsHi
rMDPN2l/O70hWqhcBzqHdTE0BzcnQMNyNyh9MxDGMN3830UibxEu1an/HIDHSf//t28flWpqAnkE
/KYWErjlhlIwy1sB3Uaw60CRsGu+y2FnI0d3sHxfJnXm01Uah5oYK3oJxvRp+olMW7gQQUp4vt43
lCU6ptIHys/uIEyaGKWJKskSQTv07JQW4H5uhy9S7Hdon1593mhBAp7CGQpYs7ctv4lKIokqIlfd
snmxmeirMtV6V94QdfudilNv7RcErfteQ31ZqJYUpHAnp55bCPVHxaLRtAp65KCuTKUO40og3hJk
yy+HPYfEV/k3P9o4NaBNxQs4jSpw6Om8Mj+YEfTm0B2bL2az78j4kyJKYC4gBnbjpXz9q9dt4TNV
wuGhN3HJU2w6w/9/ewAHmwj4g+edp1eNmRT7uq+VVJ41AwwYTdK1sQjdwcWj4uMRqWk8LMDOYdiJ
oRnfhqMC3A5cabv8YPYIWMArnRi0KdmRdNHs6wgbUvee9IBsIMZaLmdB+1JA8y/dqZaH9gCbdT3j
aeG6MOsG791hB1rHIQIaj422b5+GyjVtzFzSZDpNyFZ545MD+WwPFpqxDKi4JpbilFf2MOfId6NH
9PSFqRbsB8Lw7QjUPMaNaqxgpiBtEImPD4GF0sxgDW6phv2s9JbwKHHC8h7oq+2dqGa/Ou3JVZ5Z
u4P/NTSQ+Yr9UgojoiYQbaJGJgeasQTjb2r9zDxU0RMDUsWUXeF7SV2WMUhkkdACWXlkNH4KRSru
ppqoN1h1KrqudZvSF+dKtQSMlbvgGVmTnlfngWBUKVD9Fl7k1K8L1u1800H6FS8uTP1ycFhi6cav
ZpG4FWchTQEP1umEiQLi75AKwIawapF3OaGz2eF0cEwHyI4URmsuBhaoqUcPfJIW6YIuk3cBuTn1
moMQ4ZlBWK6acVuReRMH+V7nPeiwkVbZoNcbAJQQY9TjqQ5k1AX2WhSY2fuPYucEpHsfkgKAuYIK
5HMKKJX/xkWmnc4xNaoty93nMbVZZ+wnHajjqMp5mt/sEzQsrCo+cGIwDi2P6JwNWdNHLe0CxJfA
gj0yzu30JgG6yPpd0PIPu8CUespo+WFMqSFDf/shazQ2wE2cnB3HvpR6N/2erjRyiDD2fYGYTnPA
jlWy7u4Cjj48WVq2cCM6ie2Dm1LEQyZbJcJG4wG4ZoUfAWUxQxTde+5NBWNjp6ZvHiXnWjUeyjSv
642DIRO/gq2bgQAuabP7cMvt/W0Nqi4S/dboAO5hRf7YuoZiOtxuQjgBZufhSZoj2kUiiQD6/vmR
MmBYwp1QTL+4Zz+bWlGqjKzez4Wi6IqMaZGhAjUDrXj1+HZlE027Rk28C7nFjyJ66e1a4V1PwE5w
MErXKeKXie53RHR7spcRkgMGRZkC55DuKy8HeB8UkzsCdvggBbbqA0hEVSuGx9YgP9LOOY79Jevh
T8UPR5T2I7Rw9zamuDeLgNBt7QK/uzh5exYnSnbG5CocGcerdlfQ2XLx2ubapg7fFvMwHHT2J/4c
Q4HV8W5FsQdzEH4FH3H3rQQDB+WnYSZSesNmD9GeY+90eCyV3dFmzOb7aS7A5ES94EDh6fZS4AEH
hN6dwsCT+tZjqZCwp0LiwGbWWaBRdKODbZsZAv75JxDms7z7hr4B/Yp1srofoAmKzKp3tkTaIS+C
aCgTs9IPy8qK+KCKUNNIhbWeXLC8KB7k5E+UkkTAHJxI00oWz7gk8WofOq4ESorMTiBNntpXzY2o
elNRR3nfn/oyiLSUjj7lW7x7cXwYMWpf/y5i9X68zaf9jYDKF3S00UoFFxCNFmglgFIMImPjeOkw
XulGewT5ADMNZhKokDNvgB8kdWKdqbZJrZ2ikapd/dxWxb3ZpPFelNMpmsITa2dukLq3WQ0/X4bV
aiIQqWhD2y+F2UDb8uerAu50IAwWWVH03bR5FDJztZYZCoQHux2+LV/4LzrizdalRnTvF8cwZ8aZ
IV8U8fKj9ta4uZ/HCkCbJ+rlvd9IltWDA2i+kibtMQ+5DVZ4E5tLixpMLfZZlBrxSDMIu4B3x0o6
tmk3HDUHa2c77rdyPY4kVEyhb1narEPxO6JS7gEJeLWzGcSfGDZKFYn+a4RlyFMlcWaQTrmD/uhF
xi5jy/DmXPE/WOwPahhDW1lYtQI2yIASbqBr4HKTeiu7DupDON4UttUIFHazPoc3ZpnXhMJgLsGG
707nCcbr9OesMIls2AQTIhYd9yxLxCRyRxj8s3rDviPTFXraJn52ORhs08E9HrBa6kwc4Bulpb4o
u61Ed5tQUv9m9tgZ+m20rsZY2S+UdTaH3NdqcrTB/wvJdhbZF7S3Tkowlvt6xJWyg7MF7/nez4CK
u7oA02xpvK3ffw7oztC6oLNH4K6iKVNgangN59BwJ9bjtScS5ffoPUze5w3E4toE8Wtitvr4wmZx
BxfQwf+kS097gqFKvvoGEBwKdflYUKg3V8jm7KOoslVYs6qZn+afhUbx2kkKuC5PX7iJxIvcOo6n
PEg55dzZYNT1+jNadekRidcX0hHSqCT4Q4RvQlmXAhYRZe4ePE6oza/c1/uvWh7Aw8fAeqN+7wv4
L1OFvQYa3wr3gt75ufvcSIgIW+1587m/VsOk7maHkNeeTvuY5UL2TS5/AdcLPB8P792Y5XdSzvjA
37XW03Z3rq8bxBwaqCz58QBdTG8SZmfGjS+gZ3w5WiJn6NLlcMGotSw5KubWpjh+WYmX0ubi9Pih
vPY0fgbucP9IFkU9LQsXd0BpqAHvokWywzs7DLxdlPfJSjggz1oOF6nheHnsKPgZosYptbP5ehJD
ITSFpQZVL0Gny1htSdBH3en9MTUgKTUopP8rEWTe75WQXbjDhV1yUASzczZmOfV122UHGvCwb7GE
7D/ywXDiM4FwhPvegGS0Plz8N987+fNFCHZHusgp1lPuontBZqyT/DRrJYxQb8DyPE1OY4kILudR
LynR21V32nd2MnIDj/lu578hSPrLaVYZ6AMdgvk1JC3bDeUDEbMWxaBRbBqrifjKKLUv5ofe0Qju
oFl7PlZJNc4rcybjdrMjR7xhLDzwvukd0/PFdwRmURyAklFi7oWO0P/2CS1z8K9i9C39UzBvDHhS
YD2FkQcShCGHrI3MFUB6W4A5PDq2lHSl5Wu5pACdc9GBtustGzHKFI/J9+2kWid4vKnug7kRjhDP
xBIY4ueaO9pACBjfs2diP5KetbOJs9p9XP8R654tSx6NbWNtGKf/eqh3W/gbQY35g2FdxzmlfCJh
DfXB56mqoyJtUqk1TZ30PBfUhYEjyUA9Z7pEzOKNQCbs8qBxX2DVsq1G90ZenGK1UTckWZbmD5Mv
1Bqc4jc1BWEIPBIHkzLNMUz1uVP4o7Gh4JtRsROUmJACCt/YGyP22Kq1bR3brWdfOIlqDfeuMiiR
z1pNbqiiULsMpRUxQDruXpieUs17ndUDZGzp9axTgwUaueVc9QtXKKYmL9qxo5V0CuqqFcU/iU3e
I+Ayf3CBmmt6Wxg8D8I02HhjlgsYvLuCY4XRGyLFMxF0a0fS90zvfpYFwnKgww/DNapiDLSLFD/O
A1uWZHJkOu9pDcJhHm+5xSfqo3o5L0G/FfJh9XuL4ccauT9GFH18sflMk04XSf9JNfB9OC3ukABe
RG2oOdrQRE5zw2c/116R4QiCl7DCZuvuVoaKMu1qgScD2tO0R2xT2uGhoKXhxlDStXWPWflq4Ozg
Ust0ZBltlvzzfI7pJNqfhijWT5L7ApoQt8SYSsQmpFNPqY2JeWM0PQ8POKbak11VNHlzZqBnn2RW
BNlujPpKagvf0FhoGxiPFsQFbgCOFF6ogyHDcO4OqbTwsMNgCtnbZkjtGrvsekPN43zFMsBvKS9X
bls7IYJXC2iWLTOwYggqCSCwDiFG40ouay3xdZSlgMbbkG+1eTBtGV0NRoffyUlf4w/AGKR0Zn+F
5Ei4jHek5CXB1eAG9jlnbgNVvXQlkfX/h2KkkeOZZH/h836MpxXpuVxvVoHC0gjmG+POCupXZaQz
BIhBR0Dsgor9VdfT+mMKrnwwEmN94FFEvBeg7m8jlGHhyDCzdX8r4dTluQahBV6KCMuFmKWIwemC
SB34dFKH00nV1gfZkllf+K3e3J7sXIA9b1W1YgXdTnWNtFa0K4ZkbOzpARCbpPulZErZWRY6QXDm
xNiVDBQx6Z5Ksu2DHQJP/fPeKQFXT4dJbVZ0e2MJFOMV34UyXlxKqHK6XQrXRwI3GDLxyKMQ82Bd
u66A+xlHEmndD+x8hqqAw2y82Ag6DnfmLDZL5cNsubt/QfQGyryLb4Bn3Qz/45ZQ6ea4ODEn+O/8
qmqYuIudmbgx8RhT2AT3CTNjTGkQ2GfGY41BDaGwA63rryXWy/ehwMtUVl62RXdqLh4Rvel6bGXY
9lzSDsQKanjJS1qCEtYl0048UTHy3pNZav0oopjbQLJOlbXsQ2Pohl9SIKJ7FU1PgtCMFveSHvqu
QzrQ2jpOPzJCuBQzCg+zAAqccl0lVdcR2ys0f0wcfLGeWaRxksQdA+NHgQLmusdfJ2uKrYVtCzdw
/mAeJwUQvq1wiq8f4lortc09tkpelJvMjtgVPe6gBYaOMMQhfuTlRCsJDInj3rLoWMIsC2f/7V+V
csOiZv4KYOZ8/YMydju7YSdR8e0ti4fSyLoD2c+UeFvIDYshgJ/zNSTNABL3OYZ37GUpnqZXuxVJ
WAE6cS3w4JZiwIHXlzURTEQ/sGKgCFRrCh9f8ctFmY7aepoIeNjB5bdMrZJZLCibPRl8KbRjPihg
MkjJcxsSUc8U4lsPOYQj36IaOQIvNO6EzCSedrbQeJOvRonc14VwYb92ra51QW8hJZBNRzenvZBx
/mB3EYLO32y+34w+Rf48SwLy9bJCbZjcsHPTtvtecYnmkI8nJHFN9s+O9ODeTp0WUk7N25mBz27D
ogxCLiq3wnIa0nZGRsKiFOARTbAG8+BPONcOMz4d5IqWprH5t6bf/pFpKdi2c2DuU8GKJkmXmcy9
4YbNHsx1aWqBsXnATa1C1elZwY+sOc4jqEIuy7YldsIveiGVn9izUEsjnYcQbcUa0Fa5t9t0RDDk
3xUdlkoCqSXgeMzz3fREvr7wkjDEQnXonpfD6labBjNvikfJV/Ou2Gfqrqe4xRuJk23+e8CjNxQp
gQwiQH3rGIinaMvPnvjlYWj16JidMYijfld5wTLsA5N2ZfZxPyk8+A8k8LnmEv/dxOHnOZ50MMSm
nyi4VAMKr/DtftLwv27Hwsq9ZR2SildzlIdde0wfAhAk2liselvEnmVj1M7waRy5LJETQb4AYl53
2BwFDBn0irF0iAdfSkdd5Vw+lWhlY/bKBq85cDpOYP/xwb7Zv0nM8u4D1t3qshR1q90UXVbKAHxx
M04+15G4eoI5Z3TPMHgfot85kvpjU7LOBF85CueoGsXQHNd1LBeRa7RSs6FfTwY29PAruShiqmiA
CrVkSvasFEjfRrBd0iCiLQ2eF9Ug/1vCt9LYM1xaAf7+HlJHRqA/iKj5mYvZLfxLjv/3kLHY64MP
je5n4fPtv3sHIvkXLKH9bzXurTirom3XqTKNafa0PRaLlT7ie6KjZzowFI+cZcOCa/sVhyOGIegP
UsWqnXOGcFpQWSimZJqLIKqkES6g58miZQRxkcUd1AjrknVHDbvog9BmjIkSvmcXkuPzQ2o2XYsP
3UqSwsliUl77IJEwDGiGrvOkZUX9zxlVpiTOK0wNogVjHbm9iIKRtNx8JVcTrP+EZvZ6DTYyNvzh
56CQOD6324JGDl0eEjFTOOmkNWR6XlQnnRj1Z18s+OuBegi1ct15bE+Cg23ot93PgTeyMSAQbVHg
+kbEKe4j8mJWf3rL160WxLr3sLG5Qzlw3PB9mofcSx2ogr/6mVdEFaaTnZmobYJIX1PML4vjhnRr
GIndjFhmU4iDwodvr1ubvdvcdBUf46XHuD2vIv33JCixqRocANxLFhAuag/QcVA3DxCD5+akL/Be
cDKyasqb5ZbrqnlXfN50VePYO1QKR9PXyZbHI22y3hEdlUdcNeFlWM0uBgozS6035tab5VIundr/
XpHck4QvRHD6HDi3cw2xd8xmrfAiTZaG00rRcL8urdIUJNKacYtIbhZZ4eD3BfgHN6QrkCe0elBv
zYXtQMGEkslWCbqBQuW0iqPmopycDwNiuAZ7jitG09wRxlMyHVPGdv1hu7w3gITWj/ZmnqrREJPT
X0j+QalDY702t0eOj7eeLOoxQzm6Mp3zKVRxB3LZzFjxgh66mcZbTG+eF/B49J6PxaUxW+9rQffG
H167KVcdNLMe7guBHjkjZ8ti9bDPBY5fOFL1lg9ZnpRqGvv9G+HZGEhYQ9PWIk1CJv/AiIvvuSeP
YyzWZ4JdwhWcPzr3IAgq09E+qWFHxWEMou4EgTPJhDD1rQq68I7vXT05v1+wFpromW4tnK97AvcB
t7GRuZHATEnSt+ucB3rIZJTKjYmedmkmkKM/EjkOh9Vqd0TsUKOPt5eOzFoInMo7zkndbNQ93z4q
8URf6mPjFuoM2/2iBYNGes9Aq0VB2H+rzuWHKodU7+eys0KQsw8EmJQniIBBaJDOP32mjLZTpp8e
+h6qFdO3gGvJZMt/O9wK2YgLmEgt6TjbxeAWESYLRyyLWI+2xqFlH2BpdnjZ1C4qFJmzX6nmnaQ5
tAspGIF3vd8pT3OBLjpEgGX+rN922AQ9ogM2UKy2UsnPKiU33mJqEps8mcU3nKGtDCYWS0ZjPvWR
fYbhzsBmTcz/ZqmmrkeQmD8W+7h3iM2qwvfbtt38E5PotNnBSmjUU3TtFPF4TZ8ZMH1YTn/TKBEk
uu1brYYpc9MEf66/ezaONPplBVOZdOpbdtQWQaIdh+RS9ki+Z+KbrhhUlQquhiW9orFsOxbW56vn
lbIKv+nuyce0XhEEF51NYBZofBSGaMZCXOjB9KE4Fa8j/j1+AvZwPHKyTZ9gY4+M9Z/obuIX86QY
Z8f6bCLvhsh4Sq2ZS+eYXv4qKnVIy+xZ8VS3GOuU/suwts4h2yrtj0aaTpha1uSwgbNj4DkASkO4
6xSXdBm0ZagkjEuDpmH9T3IpwxDG0FI2K9QH/PPrpczI/D58gFvNavyAdalUlTNn6WRgAMTNhiUH
Ers8Ih4SWMP7ALWdfnoTfBJpuhPPOZI88EA0G2FuO+Ltk5XG2y/BcRsXmMInlBHAI5HGhzFRPiyY
FarA8z04J02EyFejYbjnLgZ9S7pL2+q5RA3T4m+RhPPTrrVtG/USYM+Gw1sXwVjZVGZDA8HGG43q
D0hwsX7WbD0po/A4VtPYk8ALw3lrMg9hPRxRTFd25l4RjmNXGiqZIKEkOZ0uqmRhSlZk99naM4UC
GAjd2NhXFnzdkTInUdkiO2f1+ryVA5IaV1YnJOxvjtj4NJuLN9xSZWbIwGW8SHp23HBJy9u811yX
3U9rTZLJx2U86s0ulqIlbJn95gch6F6MNsFx49Spvhs6C/fCMJ0Hr/D33+TG5lUbJgQeTW26NXf/
48RKPr8atp2AGBa5a1bHCASYwmWYSJMAfou8heYFgjznoiY+ElrBRY7COJcbT4BuKI1wloay+A0E
uLDoIe5Cu0fqUIFJAOXJXBNpKjiCUgBgisuIqylTFq7XraZjlSFkVWspORkPIS4cdnoNGOHR7AqD
wH9v4AQQ8vouMgDFKbPVgfYo9Jn1UCMbRcxK2wfV4Xxig6nUUqDmDSf/13PvpA9j41a+bkluCwAQ
y+y/QJKYjaVZgQ54wzblIMKtafHqbAP6/tw45yCDL4DK7DwNGnoPiV1LRu+Ukjm8KtUQI250sHxG
vtYw36d6fA71DXINRCiGEiwu2LwLQlED8jhGTdcCdEu4rDgQiWZvViLL89ZaZjBuQyR9XT5PU8hD
uyb8Rm9IeC9r7i+oPc6G9RwPyv9TBTch3Q04owp9p17yx3NMKB5XkdJV8xWcrg1tjhfo0hTQux1U
e++Jc0yYRbnLyLhGPP6bPlmBxmtDbzYFAeDF6hOumdrafkWkYvO7ooVcSeCAW5D7Pn+1URPcAVDP
jDPZOq30dGu9jamdteEPe2H0uvVxmSnoRM6jyNMv15tg6yROyZnW3W7CxybzepzFpvxk4uowPAqO
0QKzYBuCcZyllgZenZ2UzWj2aMs8OCRaYGr+GFpqGCWLOagWQgZdkKSBuoaX/GTUp+24AeTtOjK8
bEOdrENV9a6pe91ZLCSbkNn1lVwDmh2rw98xqbJuU5b7ZtuG03f4a2VrGb1V85nTy6lg3A2z+H33
44JFxICb/nPow7ccg39zo4l6PvlD2yxKWcT1Y2NNyFOFcG+G4ZkC/TFK8hcDLIize0J3YttXes/U
ixafCMTELTuWEj7jZ3LopfNy+8UqlI9hVCrpbDTyvk7bXlaVv+xgU5SPRyaLymJQ1P7zDQ+4gQxU
ADhCQxOCYty1U4K80WAACYCJAHYYbgjk2pxdfXVyslXerwthEmlg821BX0ndfoCIfcFgV08sdsTF
7zlSn2S5Y/b83SFlzIiidXu+9XFt0vlteqSXjIKzVBeGo6NMLhuF9kbx7vxOp0+S/i7xkLC7Dyme
cF417oqAZsOX51bAeVkLDILDmXSeyQ73W7cnNoXyMCJgQGWKQp9EZxpMeUgQrn3Fbq+DnixRt2k7
icvf3S2P26D/h/aPhzWviDV375SNzRI1OKQdbHWcZCcbvjQTLNdKmFjMkz+EvmRg9IksvsxXtLjw
AU1U2/SINa4Y/MEfUPElP12g28+txgQZbMT1dJrgiRYdgNYqCvM9OjS6AnrfdItyuiS+VTVhkBm1
1xyXT12B3C7y0+2P6tyJo6QRyGDA3i/GrwkgwC4bwRREUN+ckGYkrksHyMrXDIYk38JZn8Zxn3Sq
ZYZf5b7E0MbpY1476AXqtuSWD/HDozgs5J+DvqgfE7n+M2sXeq7Vu1eEaqEDkHUqKGP3YwzboqAA
iRFPPt4eJsf5GPonak0ZWRKyU3flZ2lSndsvGjTTMDppitqdpQb2t/IKFH5tgXVRqc38Qv76mQTa
kOZ2NXIYUTU9cUN0JapGB/UlylYE45DHNxqpNzRhaOZBrrPc8TAAodtKGN0JrO5InUFjBWgvzbjR
8RQTEP3+lPJmSxncF/BJQGQhc7uTnAGQp72ZfcbxrbJfPZ3dGqegHqifAj4E+2z7onTlb3Sp5TPH
QDYQPv8OFSBOfeoHkUUawpnMKcjnBu5aT5R8CqPKNWyy9yGUVHxxInmNSMrUq32hdXAUR/RXg8J2
vkVIcrdbI1xiXKwgR7Ap046Wqol3zdWc6fn621oyvoA1TvP2BOSyz4FqchNDULlqxDKUIE1VSIgO
8R6uTjpc5svm6kHdd6MnnLRoeZ3GXF0S6BCqf7RtNk4gywvMm0Mz1Z4tmsYZKhPN1XOibIFYl/P0
Me3qGpFiXVJ4trcUNoeo9IWQIEooObW5O52dRnZX0QXqeNo+XirCOt9FT6Z8fhQ2ONKopFO2PTMs
2dnESFh3bV+p+e8oBzTsHo7PY0yvecoYhdjYl6YgwcIBKV4lkL5+JUwPgSAB1d23Ed1U7Wun1pCh
OSuFMSGlN4lqNh4i+pJA3wQgUGym4LSSwP58ywtfkNwLgWO6afdPD1qxQD6ChjIi9s7dFV9ZWk2N
PAt0wa6pwllL0Kf65qe2yZjoei/X+SGdp0GIR0XqYNhwyn066T7z3HYLdeEFUBayg9Il1tHY7rVP
G+nqLfkV/Lc8OmrMKV7GlFuJn4Cpmd8fmONd+P9D0Lr3yrekaih3opL2VFxyODmv/qmkR0+ZLwDO
3pt54q2sWebVezcAwEz8uem+z0/o+tKDssOo1kr+78UDdaparG5Tzruqiu9H1ZoQi9MCs8SDlCui
9yoBZ0RDuUdyIR7G3RTP10iOAt06X8nTPx5auUakusI53t43OFQveMMtfqVw/JE6rMvsWxkPs6Pt
684svt8tD07KsPQJIaUi+Hz4yU6S0L/Q81rfBBlesN2JFa4R9z0YL2KvB9iIIQKezNbMpwrh6XFS
h4+fLnnwAaxOYaKs14L81baoaonmPl/aBlRDSgMj4vGlzc0G7iBdg/JWVgsUtKGU8StXRYNNJ5Eg
G5Xk34+ZUEJuuwlYoo2rdmrb4g2Gz2w8j0wu3025hPnTBhHq/b/iGHTLiqohDsyCzgzsHdvRix2C
YGsYATDgvaI7j17o0JKDjiFfAXAUckXemwD7ithKlTnkCyv5gmcR9kFf16AVC3gyY0t0oxbTkErS
zZ1KkUUtSgPRaaEIuS1NUZg28dDkhxaudabbHp4b/Wzc66Eiq7ZPuyl9jtmG1L0NaJi4pGJGvjkY
nCLahUx9wvEYVStJOJbAIZvsnhmndnWxAzDQu+calOMg84R5zANcr7bE+ytGAK0pmLq3YWJbhemy
VxNDFLKK9fdiHh97V+uToBx57JASiqMxg2joR3Auc7cygfCfn3WBwjqoNPdWerV5v/fSlmLY31hA
FJ0R9Ej62YLCZecEn2z/Eckq7AhSvpQdVOVmYKKG+1A2db7/R8KRd6pSlfuc3nXHhuG718naMC6D
bF79BNXS7Dqd7XdpalW6Lyk/ZDtc3eck+Tj7fFvBxHDsOfps39E3gQxugQLpWHqJtjvx5YviAHTK
opoo8Z04Y7OZySaHFGLXUHNtd+zlwQg6gaLZizJODbzBAahN5X0fcF9wCM/aAN/+ckIT39Mc6vOz
0oajFQcyoYynL9YuTVQ+3OB2dWpAGPywIM/nEAKk8UT3fj8nO9OkILMAMz32r7j08spUSVnmhzSE
iQMopyK02nRBQ5e1KHv249slUIbqcpkemvwP0uRKWw2PBV+AhKPJ9ctK/I02Cb0LYzqTw8qvmphD
D8oZEaxIYZ2XETwrOdXZg5r+GvAC1cQ1uDWld++W/SgvQ6lHeQNLoEeWgUSJ0dXtcnulfZCEYNtV
GHe18J/9eYqlDvdzdpWPRiC4i2cRRIz3jfx7pFDRzk6XjDtQYVuApBCKLOAN6zMEKHA14P+HgKNl
fZk058BmzdyYhIIbdQAw/8tg5gTcp1sLOS5/grXJ+/lYTiuOOJngjf+QDrM70f09pEhBHqsTTIls
IUUmAAAuZ1vykj3ZHJalyqkn5LUGpRbA4MTOLRDAcvahO/ZQKjADuELsi4NomfLWhy0bkG45P/pF
8943lP7abdCFm5tMPf8vMxG102wb7y9vbVt1qaqByQpVOgsc8ejbFtx1y+uj6aWKaruOGed4w90j
Tg0iHwDxSh36YaY4Xnt2W145t+TTwO5JPW0ijdA3Hg2EowKehRodAcdDJ4CDHHKOzXGTWeslS91P
k3E7gJFuv2blFyiDP4fTwHqvftY2WcpYUUvi+omqrugnoCwGHg52iHueYaJzyZt7lpErpqBMrWc/
9CY4Bqh8GWaP+DB5R8mYYoL0UpNkKEqhB8MWG2Vmg1QtqBvq0psdRYc2ijArtOefZegTD0yOsfmK
ko4xGtVmHJ4ic+ajbj/HAt7kKRdE2EEWny9ZHz4Tf119bU3SjtkolQXyv7U2CtBCextPy1FfJYaB
wtHWZ734zgWWCJEPX3wRv9ot88jiAYUpTMZ2IQZqDy1Af9f1ct5PDs/tELsckkBWWwynL7liUY1X
QLLvlLt+MCbhzbUB+oPuLYXJ5C4OBAqglflihkUKJU+HyNoOeGPAOginT35p235aXB2XUM4oKJDR
wgOOGrL071WnFR8Bit3U/WiTdj3AhGRyPXSp3wFNBcJV5aIsVonjZ7c/dBZvdaPxhHov2euVb21I
XAYE9zAgGfHHrYw469DyfQtsCQPQIGqqdtRkoDv8uI55YOrR5UhdFVA0CwNFCkv7ZkABj5AvJuHE
YRzk6qUHiQF1vysIdEBiXbakDXymONn/OIjNIpujPmY9iTyntjidQ37+1De+x4OFD9aJWIl0VrVO
OWi8AmMrifJWBK2j/Lq7njm5VwyA9+L6HLblC0hh1IIGOfkrKZlqY3w8/marEyJVoZ/PFiUzZ6g3
NIk8YngWtFeBUBMOJ9nrfW7HvUa1yDpbx1C0XZYDSQ3kirkod5wUc0N20++w+VeM2SjoEDOb3+Dd
fthgpNlb/9tYi1fC/pUGKdLOxyTpmOoxnGyTNnQqPePYEvwK++GiN8oeGyiiXfXclKrN1xZiWM5y
nivieTSVD2PF9UStf9O1Qm+w3VQyLIbGz9K+ONkQzLabIf9WvwcgTGLvuhs/Lxa/Ecf4+Xb6CemR
D3s4jAj5mLZmurzBCc83AQVuvOocHt3t/1TtxQKOs/OU+l597Sucp65WHqtrGDQcAKIqCHILu0tV
w9Ht8OUu3QeNkzdXPF3MZWb6RYiN+kuw8zd3YbDwLM4eS3vq0gh4qlvqHQuzoOCIyqT7+f167Spo
NrJZH0eIGPfwBjxDzivgu2GJ/P7BDj7gXrINP8tpEZokDM63rtEDNFCtPDwOYQUUzpiPOnbZ7Osg
8jGubrRSvIQaqK9eIQW9w4Iz6Swfg8hqWURT+ExzSES0H+YkGfKjk/ewBQFrVRD+WA2/1s4GFz7e
XSeGSQH1XG5U144UM/x4bOf3vYAMDFGNCZ07t5RlcuKeL94pDajjpj0D5IdAktxJKObFLhzYQQEq
IbDxp65Z7X9tAA08UlQPOQxm3i2Dtdg3zC1G1lMtL1MmypB/wZvQZLtVfPH+s/qYHqxbSNE+WyKV
XV70ICNaghr9axRBThxliKL4OnTUW20GlMPB+CNHTGBtUyDE7wku7vLvJqX/yAUHbQdVEVebfa6E
spPFVM7MVN+qDuDkCy6DrMtDsGMhFJp6+RZGg+fsRPEdo4zED/zfaQ3wZG1Zww4cLxQNmb66E97b
eQlnqLbawFjjsbOYsCIa6Lp7rDInYGKhmlIHILZLbprpUmKT59GXtdWNuHQNFFXiKGmr3CdfEcKa
WtuEnlLAcYG6tA5NXu2dlNqKHGiDJagVOgJ2Lj2BcXZBWGhUtUB4BRAm6TQDbTqPzOKCDp4JuyZx
LxYpT5woqkP04wVkrzGmlifex2hj9EPsTL8AKsElXsOAxIzEozox0D7Qhk16mIpr85mwu7W8F2JL
8SI+zO3vMigyFgjQwwWogfILihSZxOa6gQjKYWwD8llh3vKkAbEpyLgQayYgIdNC6lpNHNVr74jr
/bY6dJxDFuhzFhwlyjU6oYH9b90jstYH1fqvC5wfLQFYFaxpX3WHA/CgiSIMGFRA1b2lKxwXnG+w
CJKx6sHAeJL2oTkCmb3MD151fLnj1wWG9RafjN87xWmh7+jfSph0prUznk9hRzu1GWKWvLNPmc1H
clJX2VqPcoN6Kd/keRSVweextacD+EN786frCA/KoclNehEdRzeE7CEwx7sTwiA2haU1BbZ/bgU/
2wQdUA+DPNC8fVNpnnzwDgcTLAfuU5wCED3qERV6oaoBcFGtnDaU36G3tgnVkPoPRNS5pbK21cp0
m108BrMsN1FChoFc7AHf54RH4fqEaR6tNQRc0XFg7rjbCWgzZiPVEtIwYrN8vvQjiKhFsk82zjuH
WEWSyuV6vVKjUSPNxmNZ1aK97SeBJubLzczkh5CgxAWcb1Vw//vv0FPVa3GJH1TZSDszdk1b3xFb
CawdcVG9Ox8Yb0sjNdwg1ASX5PR3HtSSDy6vseCQU4YP9LXcqfewbaeqAw0sgjsbuRx7pCWtBVT2
g50RoBzZAyg5huTmXvJRQioqTs8OYZMxs0pq1ND+QLYGVtJi2m8HqU05GzcdbYyHUMYTagDlj32S
oOCH+KfVlgFDjZrhxTwq1sUzI9AgTCP3lfaxG8wl3DcA1hAWxZdQBA5vDSX2YGGeFRRxHBVL/jRn
QQrdKcrDAdcx7uu05uoiv6rq5Yxhdv0J0IsebcI069kcLqMVI0vWQQnpjmmb25qa/h0D88d7gtir
kedZL1daa3Vs4VLWOBPkyVxIOosBnwnxBncXTjHIqoVp3/c2dimM5S1cMfbLzwUmypyb5bn+XTTY
PoPdDznTwPOjWfiJ4OrrKveiBbVl35+XTvH4b7mCpNEOlSTzITfdMjFsRSUbiog8ZGrUCDRzfAP8
HEo48wv598t2+t4pqMIBHoMrmHjhX8AHkW0ttrNjTAHAac5Vz6jHtNV7fcLpaU3xKnsxZopi7TTS
7R/PbEkMPuUqKq7ZEpycqmHanU3jZBaRQxQDt55VN326CTFVtpf5bRj29FBhOHnsT5GEhqSw1sPx
Lr4XjgxNy5xXoyVPeLTfZs8pZ4ZmBW4xInF14cU4wtzoXV7bwdvp1TTMbCRNetfia4gXE0c8dxik
nsRbEEqoy5HNn9aegS4TN6V26HiWzL1MEseBax8UOW9V/nRaE1f9DrWJoSUGFw4CjdGXqFmVTEGK
b6683gn9kmXPevZfQbyIx/lruE+jFKF1aV1vqYI3QZExS19Bk13OBBY6OTvNZhDPgJMqfPTfuhO3
hdqmjkwJ6neQtAIev2D1FmWmebkV61Dp/cgAYqgemDvWol5hONSzqC7gi2bT6s2epdI2LQKoWz7b
8/rSyAyzUA8DL6CwylqXwP8ahi9oa6jXmef5MIXq8VIdnSGRMxvraXaM4O56tY+156He7dAG+EAm
SdVHkQBg2NOdptlUUryKhZRGwCTfMrESs2rimui0aGFc7ztIab/q0U0GGnx+9gml18LoLtKy0R1k
f+gtbvJMOLCyN+49HbFzKGHRyPeo02Vlmug5fn+UJBQrHeMWilsp/dpTHNrm+o5suETFntT6Hukl
HzvdaoLrF1qehjFW5GALG+k00A4BvGyBwDlf6UNZY7pxus6QnROYk/LmS7WMWi1eaXW06slxAFYT
BSd46qZwyVb1TD6Yw/NQL6n3DURDKKUQj3iCa5VR4MEhsaBsgrjdsmLBZrhadkmMXpBJpzvhKFad
Y393TrJfDfHIEZ5kHirM07LgPU+Bw7kfQ7ht0BtcPYmDuC5bqopwbyb8I0bHqVephGxPXBohFser
Lotpwfjz3XjkP+3JTWkzwjN+gK60HGh27iFOuzuRatU1VuUhb9hywqTQ789Rib+vhG8ZxaFRqSiM
KBNjlwxRv39/vxqUmP6Fa4F12mpXJCRlgd5uVgdkWqyD+rncDuoqB2EAcIjhZnkcWcMZYgYMhM+S
tZhyKjf3+E9OpsyAksy7DJ8Y8QERJcjYpPc3fS6hxZXgzKiZWC6o1xzEQcQ/q5WlwW4f7VeiRqTE
NUZJUbAX3YsNZmOYwxXN2H/bpBJYHgWGJKghHCOLoZNjpQ3tVSexFGiRvytmPfW0p7MHY0qbc86l
dwmtNO6nwyP1g2Q9+/Z271U1OTasUEslQ10IRttJBs+Hab/e5l0M817sbnFx9D9WcqowsoLWH3ye
mb0aIfgc+R2gTKRMRdd8xRgAuVQ/7oXc5GU5jL+4Z2kX5fEco+RhvY2IRJ4T26bF0/SskOiN+UVi
BgpQoxfBzeV9e3hVM25VjPbddQK5J2j96iI3Lb3WjGna6Ae8QGL47NyFvjOy2Ur+LSiSqdtDpqHq
ebsR9mt9+tMZ3V7pNi1bXvfCDpLg0rVp1GiAo2tTlm34vr/H+SixmidCCCfPRngFf1fkC2LIZKp6
NuP1aVNDuzhJcPgYOKqUGwE7Gpme00jjZpGfM3aNhOK2h/vcihcRP0CWYyG0YnRHqm8LH3g7JZee
W6aoo//tUXln5CRU7eSk98uo6JnCiUTKov25SDHivjoqvvNmqEVzlmQaaYvyW8uDCIZ8H252Md0f
FXMFFrUkYrPeD3sJO4ZpFQEusMEA5Avqw2o3DwphO79qLPnyHt6k+WXNvksbadjF6+tFxWVpWW1K
jguyFOe+4xF3EmrBMI6V6E8KCJ9z36JGagmGip0F8QP/NLZ20VfoahE1m/q/4MBl7DHF1DjUB47G
PvEcz6EmqP2w1JNToBwaegooXa8P8V5GuW+X3BrZQnQ9W22Hd7pz0IBIJSuPjvHBz+nsstOobDN6
tmBEectVq3/y3Br61YmjZYofsgjOGxbW+UN7bmlGQLM5NU/BNaduqKWVKldxPSeBwZw3d1TKD4Fj
liQENArV4HFMC1YxE++a4N9P3brrqm00Vrz6Az8yukBY2A/jW3YtSbOVpkAjubCsO1mKax0ior/Q
b+M8QqlOCrb/LQmjgvZvCmsRCNn16jMPf0RHBkOD/8Sj9FB0qI7HMaX0Fw5mj96IATOnlFehNg9i
H+KKhVYqS/HRcYV0RY5wYxTivA/eMRFv6k9BF+o+nmAZw5kDXLnboQieR6UjAshKpLBpX4YPa5y/
nF8Pbj+QHvXSY4p4VJ8ZV8A3Bg5+bZJljHtsT6hAvGFLWUUv0wYkVfXvoHjQByfK68yS+VC5V9aV
rFD3C4VJgbg9Ji6bKIxQ1gxlrzBUMitL/FnPJheGZrv/A04QKYWO3xf3ibwtHZyEIp3JR/WprO8T
Cq3DUbeZ04ihZH9/YajixsZGoVSCr1tVnXCcu0PbWXt1KzT/hYb12JWIKiQV2m++eqSYZzHUutZE
NlZvTQjyhcJkeRA3vJUNYiHtTcEAYFRwB/ZRc1N6RQ3mC0562i/XF4ZpUeI126spSy5QovxGyOSN
3X2aP9zPcwFDm4NIob4OnSgo0tG/QjC2OveWS+laJu1Vr37CXADSz9ggoduJIwMM0UgLQr77fgX5
2F60+3KveiSlGO4ncRemggRMc/yosy7GvKsAfhqwvbRzqzDpy3xQzFa38Th+30jxjUI5jtpp55xE
9s7Ut5QEVOKufjB6YVPmxzsspPBE0YSxSULqqMIThG4mMPvMdBap0iz/81CWqCzvQyE7VcION6Xj
QbJPB44l4qqgw3So8HnFBJZHRzmyreteCQkVBGWUfXfzCH2OjYBxZUKKWi0pGTPyBgHn//fAIS9i
Kc1K70yyONCftHvv7EtwbX2XR1LpmEDIAO8NwlYKnTcWtZqFAomD0RZng3ZRfkbsTnHT268o5YD6
XP8QqhTNAfAnPEe9yjgy23AVZxj5xgBEeO4X0mQ7smKFqTkVC/+vsEDpY8krmMWqbbGSzry+axbv
iFfLXsHjRcdaN2zle1dmxCJwDDoHXFIZzaU8B+lyJ+U4Dgb3jIS92TePtHMpGG9wrbhHebf0j2Li
JKTDOoWmMvWDnRBmKOPX6l8QAQC8DucfpjKT90CzxcoPtfIj9vU+j+hwbtvCH9KAp+ni5mWrR6BQ
KKSACJPr3/jm4J8gvVN4d/riXd3l8Qz7jqZUqeSBlxvM8LDhQRYcI4+LodBsPBNqDdW1XK9wqH2X
fK26jbfgprTumlXtFWQHhbvyY9ZRa2Y1lEwywp/4QcZYsk3BTZgt5FPN/XkOjqJKzISd3WYK6KLS
zJRcYBPcgpSKUupHHLkXdhgnC5vxB9DZ+u/QSbofPXS99RIFYFW59WEyQNpQrHjo4WBRMUVD13xj
w4wWj8+eF014e2AVbqvYT8Q7SIZhjxuLcRHqgCgPn4vmy7c3p22F2WbbEyEwjVbYXPbzXjhphxXP
Ddv222yreK6bCQU3JBeFuI/9NHFzdLK8UCBKPJqt1u8akZWw3NPG1qFFKAjBT21fFODKF/aykjg0
fKeVA9IbjatC+5Jv/biXROrjMbzak1ar1m971lypY+KbQAdmyNl3xKOM+JUd+8XdiS8kT4+q537w
nR77JAivFasCXidBC/HQRDbo3e9gFUtD1vzHGGzU69+4/j8Q/GwBT/TI+WBShN0YP0kS48j+Him3
sYY9o3zHjlfByt7SzfyPWkuaE0obLT0pjaC7lJj3NyUh2/m4njuobxORyZotKBQWt4MtyUhAtDz9
W0AR1zWQ+JVeuiTKY5FJ87BZcPoer1ETzE0xXeToHLRdrkM4QkoOSySOYIHxgD7hZvBmoXgq/MJF
M8shUqy/TSqMmye10qghOoF+/999FHBihzqb3afXAu5+WRkykqvB4ToLMYRw9fJvUkRUdLSX9sac
tECJW8tTejxX07NB0YF61a3KvwDvafLC0UkLkZlX4S+1pUakt2PHcM/hZOUOJ/BvlyYnr6HBgRsH
n4eEFvVYHBwW7II9nRgDocsALteSiVoALGVfcxUZ1hyGPyBuwyMVMbIR5uiG8+gQfYKGBKIw70ns
1gATAnacj2+gRH5DlP24X1GIxqwKG61n3n5p7WgFNDDW7/4+udFpgUeJdVx5lHMNpiiaWYOYMevl
TJqgNa2qJcS5wihc0eLDx4QRXqIBFH8EOfdeA/1fxP0qXF7FrEpFU/BrEmbaxijXGPni0IwIGauo
H0vAVpS4pBC+gO8z8N8krrPfx5OvMk6oCA8cdcNn61z9DKSZpFehqQJAeOYI36ScyaNx9Y76KFz+
y9XpjYJHADadYVco9Sssi9LScrB7ymt7zrE3ZMtnvRbqYKUGi09eKj3BY1PxPBHijPBovh1P6meF
NjTmhspm3ZiFxaoC51CkKFgnI7E3p1ZA+3KfKuVBjKdBRoqem+F+ybDQAkOAzlvsQmRbHwDc0RfB
NG0ISmF7IN8xzMfHbIPWQr4ptBk4FHQ0FJuaKFoe9nHgNpKlrt/9zDZa8vaN2M8ZCHl0XrAS05rq
5sRGMiAtqq6aPybFi+FtkXY0V6ZPVAzo7rXnkRPPDqH0lG+pzAxLR7dQfOXvylu4hm0LPOQLRo+1
Nwhwn6+C+YCBV4SEdXSmR+glHmBobGEYFcgWm+kBsF5Q/nJhaQtxJdn7eRN7kz4ZHPUVYwWQsTvQ
VPG28VD6rfp1jFuqZu2V8RPkYc3JFRmVJImbaxaLD2ItDWNUW4oRl3x/doesYQy0LhiNdwXUKgf5
eZlblSw9cfxPO/mfKUy1wUUXe3Gk1q9Du8F50KhlM10D+f7VQWpmFJVdvmCDufk9ssTLhcXld3c+
BrR+UDLB2QQS7tjmR2xLkIuMtRndBrlIGXKJXXiVd1cJu55dM3YeJdk0sFHCButGfwY5QF9EQ5MW
sd1J/NQWPlYoqoxlTBMB4BkO+4I/etS/gIspdQvGj/Lklvct1Z0R79c5+B2kuxQcp5lNR8U7FBo5
DbkRksCj0DLsNhUCNz2BpKCB8KUswSGmsg/bAVySr6JN5Ktrg8U8k9yv+37crwd+3zKQaV5D+OT3
VAU6C6PrPSCdRcwo7YVQRsv+YRsFw2E7nBApUcBaIX7ML4lSjrtArwg0OdLCWm0Rdn0cyB+eCeN4
nE+fgB1idXf+3sFJEAGnbh7vQFM0f2wNtlNVljSOOsbRA5fxUvsmK2XAuZKxwIM+g8Los2P0A328
2zeIcO4yN5EXc1MZyeMw4KTtA08vob71MiJOCSQwzv5sNC9fJYqeJ/D61iikUaBa7Xkp8hqqOCau
0bMtdQFq1rGcUKgxnqrC/W2rqVoG5JRK3GYLWvf/CH9COk7eXfsK+sDo6aLM5JpLXFd8gS7yhFCe
4r2UEByC/6777VxkvMOc7NtnGhBPPObWQavPY51Qvk6gzvEruGCaHxC0v8mqGB6zHJD0VkVZnSer
1tFy7brYxoHE7hqQ+Uv6XcWGeLacCvjTBy6F1oyBVw3QoySDYCTPOFORDz0N/hwoPXbXVUV/qyry
zNUwqG2Pj8kq7nGN8KJjx9LjbKFM7Q9PVxkQAnT1AjQIYl2N5HWW8XnU1TgcZBXvx2BuswnAf/vX
zYRtqkIh4BvN2CiZB0hsB9WclsYqW8aveUrXy5QVs4gYDoBYTnw37cmSqKYgTl7ekIeiz41m3mGW
QeBsfCJbZooz75v6hgK7Phu8U2S0RHuPe5/Fxtc1HPFbnnF91vKNh3Lz2hQpj6w8RphSD37vl7Oa
JPvkMnQKm5Ousdc0vBbdAfFSSFCKFqqYSrPK/Nv/nrrrKi9kO6Yj8m+ukGJAObpifd1wQNOvy8hv
FvzOgzNeN/w1yGVvpmFo8nJ6U7Hi0mtlYBO9nE+i3TX80euI5HbPxGBqX00BNmyMT+5ofCYZ6twW
n8oHehZ8jxrIUfSArlDsgfnZf94WAIVaZ0CR84TbtjbuINSOMtntEi3WNLHIPOwFA04V7KSx+U6q
bSBxXOBqUs1VbqcbIG9SXuCk/fsVcdjhY5jDTmvptt8/XduqKBytXd5byLC5PisO/Ugld/e9+GIL
pH42BeuM4qH+bAW9wromUkjwQ+52S8YmTZK5o+oI/lDoyvE6A1a146lF9D/4moPg5tOakaI3HHga
45vEXuNfnPwSFLPYxa+bpfDV2El2Cprq56jtdksVPPQkmhF8Zh6BvBFKVr6ZDMzfZ+RX3wSL1dx6
y/wuDjYX26w+8JlqIaZRAG5P21P4UM3pzsopZFgtAEZTGkCfh+Fn9WyMseQdTRgxnvRdOUIZXMwH
EtugoxtiYiV5WjG5f7sUNFEIucBnjQB8TYcC2OE4iS4RiI/sBBBkgZpdNYHYGmgFR2wJjamiC190
7Tuz5iJBtqjjl9Bgv8aWL2wwAb3ijT7g7XcTYDuPKdyNA2vqMvQFYvDtB0IAGGAYu/CPS4gvahmA
DWFoXYlFZoSQooWFNNVIwe2kvxWjtsknq9BZ+EkwQZ0dpOYPXWJEzpOR0tQDuvYOzaYxrZ8os81T
kjf0lmpI7hGHVAj1txH8f/mOtcx7TlWC1gwpcqLAabVRktmq1cxyVFXzXJg+vwUYfW7yGsp19233
Ak14zPCTVXvoMVJdh44VdaV3o2CftqeSJdHwz8OCl642VG2xux/hp3xGr+3hG4kM2pLICmg9Nnl1
Vr7gYWVnorGVQBED+A6MN+6TPjtWYBh7nvWuvKXFMqz2rOCRH2C9dPCUdL5u4ISqVm/yt0uSdW0G
kb7BBhoMQzBdIuVk5zY6fTTOlGp9jWyKsxMl4pXfPBJOnw2dW+5lMrOPG36gH3Ei6Rz1AdAgf6WH
zRvBoP3ER3HDEd9aqkp2ehi7NQgMLMKZvN+5Slc0DOU2/IvYp69la0bNEJkT5a3VdE8d6fhLWGcO
MM5HUNmE2XHJi82ptL3Ypk1pfyxhQV0SDFJMx3i5MmQ+qh271Oyp9m1MtxcO3Wz6Jwg2SzoXjgUl
tU9XLmJtIKXro0prwR1tUMeI3EfBuG++PKyCuuZDKMB7iiDiGpNPD4DIMdHnbYP/+rOqHyYK2BG7
JOvNGs0WnqSMpD3qYR3LWytNRu++pxNinHJv2AAQhEGPJKrbgKCtUUC2XO2xwxmeNpG3wY4iaMia
kNy191p1crUVCRIKjWPWNw7Tm0DH4ITU4wOpXf4VaOkg/Dv9Gr4flillnYEi2r85SvRSKeDM9tvB
4VnxJB+Tei5C91qUt9HNXmQ2n8sxfRw0/thwxKgt/8/b/d64tadSDBScYzHoBxdpV0SpsaXNJb0f
hQSd+1kvvhi8QPxgGRXH9fPNdwFSd01aK830MaAsL1tWRf3ZM6lxRa+zJ+sm6zUB7m66WbMcinEi
+99mAEB7SYLSiUB+ZtXywmnrzUJ78wmbNFvGiSMQ7JEvak+kg6+WaWGErw7f399jgEguUP4n3ou5
ACkJ2U6EHTAAimJRXHEb32PI5MrLhQTQtO03skrVMfJsnX90tgsXgOc3kkuIwdzYUdtcDWjlp/L2
QH/JlkSjXdPvIQ0T6snvESJ4ndOJb3LqKUjGUCe6wtUpDz8apPCmrOpe3fl7tHZm1SLTZRXeRfZA
2P0WpKrZ4Vt3+DnGILZsswbsuovzYVjpEAB8VkpTTazf1iNyAA2yxFgPkuYJyrjukqpTNozpEHap
EbxKrJ8as7ccU57875JvY08biviY1Uay1Z/yPAzTI8INmJTEPKN9eS5LmuXIzRtCMmGRTNehdx0o
bswjawAjVAW73oM4R2BmgY17b0i6g0IvJkgJpM6oFkqh8DdZbnD0wFj2XMfhSLCteqLkxsIE9ejy
g7mDolO7Z3ePH/eczoqiOBUuMf1fLmFXGqvwsdZ11QP6YvC20msP2LiDdwOdIoNT5ANOsvPQPMdx
ffcvFCOfmfu+RzcYnOgaL3Qp9ZTwtEb0SI3WaVyYsAn8gZKJSr7LDNolfuVf/XskJa3vujvpezXv
D8yN40xlpz9uLUz1pDVLTjAGQyGfXy06RP8cM0IwUT6ebIZLS+/1RNeqlf/vVkohXq0aeAxpfGfS
ZBwFuymPWQqDQZLUa25tkhJtBPfkbnHudF/t59MBQpmmGlV7TBKbkgnk9uZUJcBhUPW2dYXSD/WS
hl2PQgLhNdf9cmTF03gN1p5fvKmGVQ8t/fkxnQW6ltnrDt4Z8Tm1HFJ0rVsxNU3Zr+fSN8puJ445
lN9GXddoHkpFAHupDGJDAqv93N9RGb/n53h7WQcwVMxB+qRpos66u/k9l56mDYDOYk0eY0iOT2GA
IwTkDFbTh30/a45i1SfT6V70O11bDue/4eiwLV8acdpxKlGRLa6xQwLH+rISHnd1Tab/xq9a8NVX
8DY/x0p/piM0+tXEwSTBw1M4Cbp5tII44HJ4Bp2MciVkeJFvSTxPfmA3EB4NkraCrmmTYeuky5/Y
WVUj/P3ZFZIY1r9EWmHzO8V0GGFEmTxzhlfOUPbiPo+YmIyifDFVjzmTclUNATQtRBXPQOu8UVqg
5Z0Iz9/JCw0IXK8qbVrPV23upr7n5Q27yxtDwE/GHm8llDr02OTQA5QERg+s1MNwqjIANyrI66VW
fouWIrLi2i11tHuFRe313MLYPzvIr1IrW1n46XHL6dyzrtXcM8lrk4J3aALxAsz/a0excsRqAa+q
TNY5PR22//7vsFgqvd3w60J/gov8RCSljCIaDQ/MpwEikdKFxYRuh2UVJTJfXgFRY6O8kPZGEQj4
uzUNVJeVht5VZOXd8/ez/JiAE02hwLu7AY+NHZKoPgaXw2GWHwlvIUYM+DYCbCR2TsZ5MeFotJNS
zHF+rU41PQYlinYQgK8SjzdX6j4i6mtpJZ1B85vgCSfjBdxVi3mFzEB0PYMUo6ecPBREJ7D+YE+p
z71zPhK07Cuq/1CnkYyr/fY+Qag8E+4eCQaNjSrS06zzyk9oXCdr0CTEUIiqmha8nxIjF4aUf+rQ
/szntk1Zg8Nj+Blofnd9W7QMhelWd2D+zRUrq/c1BylzI9bYW/GTJkMSa9GwuXTWN0bNC+V4ZFBu
D29lChGOGeg0yaLAg9MjiABe8VTaSUTRNhdAHrDS1Mlxki6Z4kJ9CdIPF0TH8gqqJViBbx6alWd9
k4F7u0CsgQhoKn5/TxuzGp4csXsgP8eSMEnIscmk3sgRhfn9hpCH5Ccl+5iiS1wUcrwzDOxoHItb
UJjfwg3scZ5xyzrJ0CQP1qzEcCNRiz+LNpFRLpWL2sp7pf4m4tUvb3SfhhKbLsLXaRTLLmFAqDC+
8TitB8Os+NB2lGqMXCGmC3hOz7A9p93UBcDwq+TV8V6KQXzv2TkSwiipkVLUnk+ap5zeUZEWSfjU
+uJwDaDbjWVZoEf8qyw3HkSbZ99eoSXR01vSM6nwueH9YRyrg6RX6GtTmyV8pLunEeMouxsFmojQ
2sQwU9z3wUYTqFmd7b0fGrnAtAkt9YhfZPRLQ6UYvVGCL7z2ie7efYYjMrlSMR9PkRUvRoAuI/Yq
vp6FzOr37ZfTQY0XZrdjaz2f5ATRdEbghLTfuqGJT6WF9zaPi5kXD055HQ8cOcEi0qioJ2E1aUxQ
K2d49eTGvr4FMPBWdK6lEi2SJTai1cKSQ2ubWXPCM8Ayo6qQvGg1MP0adI5vhmJMawj/Uak90lRZ
EE2RSg7bA/2kzwXLs3xqC3a1uj1pLuVOpYCocv8xtQZgH7OVHD4NsvrOH7Byb89mmnDgC5cV16Xi
+gomZKfU5ok0OjiOhK2w9j+aC6QZfkAvLI59+as8jM7eeVn+QVYUzTPQ5uusdXVaKfIW29YHOL0u
XA3lUpB+VQh0TjoqCp0En3EnCEg0qp04nyl7Yg26xiwEVmJFjCZjpKSvDQjoXfI9CH3pRQgnK1ns
acjRyeDDYhEo89Ke0th3T4zyNGQyP52F87nTTURD51YYyo75O/LLeKdMFneyGOyz4/cVvG+K8tEc
IGnIL27SxTkADVBuNpjze8QKBTuj6PoXUqfNgl+hilJmVclpkPTX148DQ7XkwmGpppbxso5zQjts
9o5cGGKUE47uqXm5NoBotcJUXLiBJzwQb/FWIaco5U+b0pr/czdE39DCxKTGTfnOlzoqrP8P2skV
JRL1aCAP9RJ5FUHcHY54YVzZJY91HLqxN1Pe8OYgAumOFEKx5CBixHvAPgqAZYvb7HpdiF6inCCl
e0jeEqo/6Bavtq7ePC3kD6kevkI0Vwq07THsFEouIFy5dbRCkT/RWm0tmgtT0FO5HE3HDT5hwaLM
FwykWeu0Az8tXD7eDpwn8J184CNdQGt1RXygL7wmNt7NgFtvsIbJ0j+xFWaWWG4jfxqwN8H1EJWW
0qbvXbpWdo9VX6egYZrZ+zJauI7lYAvayzV25e1aOQstAVMi8wfhLcE6KI3Zw1rVI1Osxt6Exy/F
bYWVOuVNdn7eSqeD4/YkJ+8EOctfZAPiwYh35HN722Bn7jTEn04dqZvwB0ZCu+QYGrYcIhU/QBCV
LYSZtnPUIZZleoBFfWjSQCuPWNn0hMj4NeMXfT5oDD4BUYumhSWeUVc4Fp8hVvdz3HIWZxUc/BuH
9NIK85oxiH81RfqAwQxGCCPN9ezJXwu1UBmF2+LAXrktuvCnc7DX21q3FduHNtqNBAMEaPVQ9IGP
0L4zcTi0RKdr3aH13SxBzRdqHkoi/P2FA/4mtTbvz8bFLoOno8pCWOs+zkD01x7ugOHZMZ0P/KI1
LgqTsnOPW7crp+0NxtNxaxuFFc6A0M9xj9ezwMTFHFs2OvrfUXLeDQHYQOl3eHhE0Qfh5/0cqN4r
azHrjHPhWWK4bMdLqKwSFcTKv4A3AQ4FaykTU/rMsKecY6369TfhYd4/ezfUxVsG5Ie8QKYWdS9+
KkFxsgLAqq43MFE3UjyH0CTjFuteF8rIiDmcJnX+m2wy1GcBOfQbFm/jWWjwG5kllcwupBYEt3Uy
yMhDQTiaAMCvLmN8y3YfPLw08d0eFxnvT48KMMPzyyqy4ZtKpiIlbUKFESCnglTh2lCm1KjVkYtn
kfnnFMEnGCHWe4fms3OQcYVFpe+8HeNh6zn6bBHvjlasetVjWhKjYVrWCVmpW0s0rxAfDOH7g9UC
wJNmx2aflrcxIjC39+LjLv0kQlravisID67i6bsdWkYVA2m6c+nvHuEVo7s9sVc56D7/J3/GMrli
5Vqdyo5ncRshsZuNCtokaH/pK1sUlrljUQlw4Ce34F+DHPoFttVG6WXO9Yj9SyEGEniupyvBBxvs
LOGPvvpYushIy4MRSdIu/zzDmdpo0qm5JogXsw6LPhzjY4deIdQ+2hvypGz2RPvQjVh3jQVtamUY
LbYo1OdpqvjmqILH3NtQIY/Kkz3Wa4WGIqQ++EXghWZxm+Ep49TYYBzy6rTJmZUq6p52WfqJ2Dkn
uc/CAbmcGASrF/z9x0PC5DYMPRGJ14+Yo0MPGsbt5k3HBsjHvCzjMFuzpejG9S+rztlwz26Kzp8G
75xN01mQgnruYFmZGfYhJp24l+2s6tYRsuMbtIEr+lb/E0F4uWnIgUuwmcqtOQ+JWfYzop//+9id
bLWMTEYoFnxA4evIQdte0C2evd+kRxf/EjyKB4zI5svd9G+bu/zb/yvtIhFTLRWg4ItRGM9moEd3
koeydv2afEPt+UfuQSaU2z0AJ+/exzjHFdkOvw7QYCVpX2rzxyc6YgeHOfbTrKzn98JMxh2xXQvW
V28Gxwy7ZaHfpwrxiv6SKqwi505p+vhq+74qqGXx1+cnXac55RR35d94tzPo+KzN9IrnuiBsOX/D
RjZOSidYyxH9IDyo7K1nZV3NL041BbQuDNJzLMeoFBram49j8eWjundvh7r3h+wzYOegcgIJxkZD
CuVQfM3cvx/IWnz95GsAUzuUDrkcTX+9xJjhHs4+1LhPMwMKhSUTJ1+7Ls3iHOQBmggwLAUJ2uj+
xykwvgKyOB61RI6j/hbNgXq71VpdGG9Ct1aSD5DM+D+z/LAOUCGNC1kZy2pG0cd3M7Q/SsarENqY
g1s8IlSxmM7hVipQuqSou6jSIb3N3MLUlp90AJix2JADCO16B+p8fCGM5K0vvP9lSdKED2ooSv0u
lOTrBpcKi3av0UshRYyQ8JLOrwD8TtNfdhjZyaxosEKOsGEtnAqzcFY433pZtu1jRyB02uhaeZRh
Oa07rDyB+6ajed1NBTbiEw6q17YIXI2NW77D/1PJbeee12OSV3d13B83zZsk2SCQHqk2lriZw9/v
k7vcfCXZ/pWoOLdxKFFPWBCBTKZCrGCZxgEH3TfsWmfQkfGaXQE+ELNr1m4brcO100+4CiOubz+v
60qeJxWcSV4ZJNfABFZ/fl7Cr0DFaT86Iq9hiVbG1/8tMxtz+VF9mLwUGveqA+2HP0MoXvHoQSGA
ABHPf+zi+ZCyPLyKfO1LgWppxGEPOksi9gybOGBwAAD9BeF+q/Fq5khWIKaDI1bAK1piyks0ivFP
tWI0Tx69G6F5fVg1b5lBEuVzwZbXswsrF23bynD/cH66RiGneA836coe9Fso+J+7C6I0KoQqSk08
fVi1AbxMtUGlhpbjl/N0U3xmFE+YG6cv8t20zXS6vf0/NA4kqup322MQb+Bg7GSB5xpoVRXg/Y34
lLRAHTq9y9lK+EnofxR4ruDjp6J+XJYHxoDetOVO/ia/JNq4gr0BfBFhI6kZvxUxe5gDDyL3Rp8C
cSXB90ebmtvdyugmOgbpoHIfKc8Zf8IjCfkOe9dpqkPuoQEGWVGv6Zqz1v/XOPv1M85hBcNvZRcK
tUISUoXONzyxm416U4JI3klxI+ZkPpckewag3MiqSfEUPxfcq6aHuny3TE1pFSQFev6cAbGGIcRb
NZEmzlJ46oy5RE2+1hLCu9fs+jAohOech9gGzdubfSYV4EVkMPWGUY/ZSuSPj3YCZdcNKQLKsTmD
D1soVX416czY9AsWZIQtaAaEtm3lZwQRY2Zub3z9fwDWcd7qazNZAA4xxsxMrmE8jOY9xkv1zyoG
O7rkFKYv7B17wffIsuqm9McUmJFReFsN4zBJh6JA9e2MuIonFl5fnS3oslw8/IUQsxdBLxhm5lh5
f+B+Qd4nAOUqcD+B2ZqGtDIWGDGPNUh5bu9+vU6wBf9Y13dAS6Ek2/8f/HOwrr0rm/UpGXkFH3PK
zgDyq8xeuEN1juiKjLLpq62XCYwt2+rVOaVhyd0u+pB79y4rWzNtjpBHmhsrT+Nv31qgZn5VtdwH
zUL987QqFzD3zttm6Vmg7W6QTUcLFgqBKA2jyJgdvBNCdUIdT7x0OcrV57bGgx5u8Xu9+gWJx8J/
MbUn5sbuBHYcg9aehZbqhuj2mACgNnHKt5WAhzO2PZ4Hq8VmNbVEpY5oLMwIxF077219cHpfOIjh
QMUC9iSgUkJDXMCJzIInHcZdSt9KnAJvHTAw7bJHLTlCvtccv0MugzALfNJI+qoTyf8gu5q0nbNV
DOE1kIGzNLb1fURPwxWL7ob4k3TnVMNWOrOLmXSzBW3PUtOmC0tXzrKjdNMtDjyvkR3bngByeH13
zC5Sp/qabqSEgH860QOpAZ9oeqDX4c8r+frCxLvSXIj8NhJl5uypOk5bt4llhsjwzazsLgEajuiP
Byr2ZsKmhSip6puYPgfwzB/9RbN5fZDi0BizJ+vdis30+7A2TN3wdEvel5wiZOmerPyhK+AapDtW
GeHLjsSplCgkOOPlNfJ7qdUno+/u/927xDbW+r29vwT1bKCJvid2zV3YwTIRrJrvKX1H/9kk1fI9
QEWQicwzLEM5wVC5zLGn9tSYqh8/s8xwzx/gkVqAFcgxrio3ZO6iSg/eepuIcAigFsROdC4bZsdN
MpGY5lKL7br2iGEJCUWkVgLB7urxjb3O9uEgoyLWjYbB/RbH6jOos2Ztw7wP2f9gD6o/KEhwhdKx
S2ZYK3jVlc0LYek+5wNyVQmlOzCia40KtudSAGtdVqo9WDipMELvzGb2HAJGe/1UehrBAe+6fxuk
zKc2hQcBJaeyBOiNtpYoM7crh74PJ1Ip6LzHRdiRKTZl/LH4zJrIVn2ExzeWkZjXHIhNVnBGCmhD
yzrd/lYCsGNvjg7JD220pfjJ7czbv29kazHx6yW0RuqoXIUSjixjyHP/xNs1puCvXlSF8arG4l1a
0DMBHRvca8FToymWMw4cIQkiDSo4sEoxeUGeEFC7lMMzvalVBYl7GryAvkqie+m09qBlngxSIHlN
wZ4SKy4ddqe73j6yg1Mmq8gWxNfiLir3PGBQe4+xx9jDsuYs0L6614AWEyhhf/WKN2VbH27G0K1y
NxD54gMlbwIhUYoVFUMmLtsnlIljPpg75+4ENDtFsWgAtbB9n2pfPalDquODTJ2XJ3mYfbv0javS
o0DnpV5sTaPiC1r7BO3G7fClVpZGz7/l4d1/4oA4IRNUWJVd3MvH8iSiSkbKCPjWSJediu3DXBKT
XK4X+sZbeHnwFnN9pkG4H3CGOUawn3id1QaWpNdw6kJKyzZigb86gys55ABr12PA2W89OpnsSquk
d4IxJiK0sVW7YhjbjmgJaADLLF0kMlIjqUxgVw8m51cIGCJZS/LZHU900M07MLofMLjPyd26xdp8
6cK+OGEZM4FK4D+yXbOyLnpqgaKobx4Kxb2IudUaC7MGYOrj90XYb19WNWdO28upZlXKyW7vG0Fj
1aEqb6E2HJ1ZUlJEy9DxolirNCLwWzxiAXgp9IrtXZoTK/QCBO8wFM7fjc471FVGBvmDl+psYeH+
ckl6yCi6c/a57ptz9w+BiJBFSHWmCkLkHVs1DuGRcBQqo9TnVbAn2G7qhlXz2OWb+Vdjqxv+BT2M
8CXHK9CiTr7+pDNJtws9zmatkdDZ6bbPEANtQat25wTRsdRcYOq/MR7AaeBNvaVc2oX5O2sba9V5
yfUwJYFh+SI+z4J+xzcSrtmWhCktbs9iLjWghya9hcebfmGI0nQJdIegZD0QHofJuAIlI7tddepK
1b1ddAlm41uhTtFDwlbHI3Q+9xYZs4ldyezWCe1SSeNDZm0hOzQW4me4lJhIgxoDePY25T0cw00v
xWx2Q1/n12E/CSCmzwMI7soFiCT06w2UO1WZzogUIH5nk3KBCIsEeRP92Yw5EwVUs0XyUkjTza2O
i5jIDNacq0ITbkfN/O1GV3nF9dPEzIzYA0Fg0nYAmgyUHV+dna30iT8PJ7PcSRFaSkFMRH8GKZTP
AHW8XKbg5Phe4NhpIjI6CBPLXoZSCMuwePPmdkLbXsalxYSyHOAwhdnSGA7vLQBRK9V6bp+/iRW0
85f9gR+k/5MoKP78hmsfURif8I9TEhi57Vyf6Hw/vlLM19PtvGpTvd5RTFu4B5C9dca3eb8/QU12
bH8HEbNCosPn/K8D4Gpop1wFkq990XHag+I/jDG9joL9vyrNcz2sBd9wxUZZ0UTTgaIxzhZ4AsP2
Rn04CSDtMEUu3tzP96ZYgo5nCKl5R2L6hvKHJ9E3FdgK9VFIvv+Ji0z5ds8+z6yZ5RjPH5KiWZcl
bpGRR6HsuODnsC17rRpRyXP8rvOHd4EuPMly1U1Tcv/AKhaVvsf6ectUXsCS/p5FEk0ORQxoOKqL
LaJOfRg8ib76dWDMZ91bH7+atpCm5Hzb34vPCL/qX04sRD3FQ6gyMTNMmy4Qsn7wqWLN2vBgXc0w
IK47QuCKCmPv8JqRN2dgK29eI/XAtT4Edsi89z5FMhD0Pw81FvU0j9mwCiEylTJHA+Lmhhovhc6i
nNntIa9tWypPzzstm/1XmZtaq8UVc66R7B28igJMSvORny43tZvbSTH/Txja4AkttWEjBAZ6FItt
9OwN8wqf/27pr2BmDfALH0f+MhC1UQOTkdbQmrus5/5xgh2qm0BlrAtoY0+4uaWP+yMlLhzbJZBe
xxxPp/T3acDMBMYxPIfywI49vxUgWpyQMuqP3KMtyXpX0Hf518a+wNDtwzXtofpAEM4OVriYyOa/
HbMNK7OMeLv7ndeKwvz+WygjGeJnopZVSSxy1YCvvLhQ0BWHujZD8NfGObSmm8fo6wKobQ0uREAZ
yT1szi8ICXr2fVxfUvzE5K12Y5axVVVypKKHxyUqpC/SAvDd1LWN7GdxMWZCy4woMDX0H/D7mpoG
1T2J+vSKC7ThscHy+yspGgHqlvkvFYqrlmj7zpYohKQR8JVoUsTy/dxdjl2j959kzXbi1TOc+v3W
6XcrxW8VO6dd6bA7LeTama1U0HIQSojDGNRVoUOq2Ki0QV3mjDiAv64IJROwRA9gTlZa4Wx789lK
n+7BI6bnooXYEgP+v35lRGmqdziKKVMyUbdgJBWZ4vEuED3K8GJ7PnzRSH1qGDbVcHrwREkd/tT/
Q0GmCLRcoTE/qmbYUrHKy40rqrfOc3jg4LA1y7ENQtntFFOfGpTJsCps77+wAz4DH3CENX6YnAgz
Rm6ZW9L5R64s8cgos+0la8BqMCnxf3PkOVKf7EXF3ZIPb8HxUAyG8Kw/3m8d4Gq1M+xriLGtrBju
btza8bS7Tlh9iF0f0mTFDryZzRGMKhhLRXAwgtjGh4lmrXXJCCSwBYUjSTIMAt2g+KNAdQMOnCf8
PzU3LRl4bKlsJJUIU6MysxP3QRO7OU60hNjT7YZ/9LgtA3sZoM1FvaNEiAy9YA1sft1CG83Mjo2t
BgNqHhnOCvBJcU9z7wlcYJpLk63KU3OSiwnr6TwTsgQOxpqotuUBthDQuL+Z1EwCXfNwhl8gIJW8
Ohi6PjxUhd/nvCRL56qD47xjIoclHx8gN3wcEM6zoZ2ten3VTh0VA04M+21oh96v2t4nxREV383h
jQqXs5y6QEMKBpFddCoDL4ePxjuKW0YlCDwomHymT5BT1FTEFzy7BnzOfrQ0X7vPtS7zN086FAAo
pYKtmOTdC/YYhb4GAV1VpA19ltltajbCZ3kjS/z4v/xFh8PNs011T8bQN35wWxrXKLZJg21YPkS1
nAWUxuSKk8BAQrTYxeFx4HUXYdfAOmxFKYOw6m2g+cWh6QWczNyZl2Drb85uWC37YI9D6xO7u2Pa
iSoAXwzswoA3FPQq7jwkc5dBJ1yK4EEdNozhPgIkjuF0ipoGj9v2TsJnmSXPbsGf7EaNRbJDp/Sd
/pskAVoO4tD33xOORuz2JtZzk/yt0AV6LlbGEK+kFv5Tx7YVo+tMgwkgEn+EVnsh+V9lHjF+Z8wL
aLmXuLYiEhhzVhym58Ozv0xxKLiVrhf/mSaxVSCyPeBXBuc9HK7K9wGg+tI0xuGMC5gcOebrLrR9
hCkCHMuwe1TvD1kyLlc7PHS9RaTWWN8TLBCrLZZZyIEuV1ZGc4yO3JOTokQzSkdf4y7mL/lfc1EO
1Reb0ZXSsDl5/KDPq67OZejXtxsi4lKp83TB25LOw55guFlL7RanPxdHlWGrblal9GdBISaKk8Am
ApP6Jl3CyqewxBXkobfcXu5RySxPUmiBzJ47DgNqPOGxYG197x5jWQ9rnTzycPvK4QOSdeK+Mqfr
JP0DwHET/iZvqDwkwLRT8RsocORZEs44YXq+c6enKj0Ui5MSpyzferBQxo0Yrdih+HJHoZ8TpU+m
rvyXzlxF0kI7057Jt7uU3k8Oe6nnQvxsFloHQYXvZHpaEucKqEJgOk4crREpYtSWj8zFp7xnyWeT
Y/F+SxSo1ZslnWv+42uPAepMyBOxB4GZOf85tqBsGXBH7tHQAVHFN1NjHgEhAKEYQX2geekCc9qo
3et44TLnGKaJ60kLjSNB3aNd4xmudNSKkeiVnbvfl4LJel1hinjIgMgg7Np4gRcJAWXA9TYbRxZY
UTANVtq0Qvr2GpbPk1uCZ8qDTYUDiRYO244/cCCR0ftbNwOkdxK19+bxuZJ1e+C9l8Cfum7GTLYj
NUHRSiPj2Ls/Zav7ZDo/gcqOBZ1W7qTyxmWTANLR5ftcCiPGh9/+91swhxVeckXPH4GjENQLh1ZX
L2t2ciWbFCF63tUJLgICJ0K8FJsZLWA3SdcNjH8x/BmWsHSrkLRg1NqwZngEsXJx1x6a5Lic86et
radtmGKiTQn2pj+Y9iUuIro9KRejKe0GzsIQNlt1xpsc2LoWpZxhSYSOJdzYyFG1/bG4OhUoe7sE
NfR5WghEvq8aThRK47/xIKj5/2Wf0xvr3vEiqhFk7wxMyZuF3UCXp5JA4TdgCZ7Jf7weLzhKxb3I
TSGf4ZHM8VU9lB0Lh5xF03XSQ/+1MobXYqyNdYill0ZN2BNysq0zm/dBdmhLgbD6giu5DfDQecYu
UEr9dcV24axBzXJVNwTvnWMgZ3p1rQkgulJlkCUzlaCIXC60eGInEMhRvYXDWHT85vW78K4tHmLq
kDl5XkyGT9KIuFBIfQV+94fWB3vcZb5+Ihfrb3QVb/5SS8+Q1Ffq8k5IfW85hxJfCVgBsis6n8pr
dWQo8GpvcMzSJ5jRG59auAi9UGDhBC99u+8ScmurbQuSQDoByyw2VmS9BxbWHPq3FAFsJoG7XYrK
3lWw7WEIUOIhjZtnhr0JiPzS6sI+Ss/lnTMVvxW8kS/O004jKgutNzpxVGUY/hhuZnF30sBBRuOT
JebWduGscvS3Dp+qpcgjF1tmbxuzDXwmVOmy3W2Yf49iQWpTxMwX1GveSobVM3LDstd8gVcNJ0g/
E+m5p9FGRGNCQOfTDJgCmjnABrySHC+udLFtkqhGOniLWJxpowKx94IIdUb/Pvtfgqwgflha8VLQ
80aaAsdPDzISU2WJZeckbHTvS6ssqcHW/zWjpZ3hSwQJ9TsQgHMDR7oX2E1akZ1qduCyaocfNTI5
9emWzNzmyPSrCXm6e8oltHj2DPusSPKDXVCPBZH8yOqjCAGKKTxZci1j5xpCf3siZEfkKkshz1kE
YI+/twc2oO7h5ojDqUaqiMuAaoAQnjTE/p7WOxtoQ4g37mHB2PiZxaURx+fZGDuGsJGSfRNlMQby
du+1ZllBi8+dSkPCvNx1cNWMfOh/Tu2/NtgYEZWzKp7EmlmAljoa0cMj24hks9gFXE0h0gIAYv26
fkhS1ah3xDmMD/dZJ/oDfttXkCzoayO3vSz8lwsBAR2eJZN706Zhy26jB9chUtqerxWA28043SDq
8rGrA2YgD6z6vwaqtONqqROC1scq5w6Cwm+gnom8UgMUZhf5pp+oZ0k+QWN426ahAgzc/e4KMSZj
cUVS6eQ3h4fEPIc1cWu21ynAiDP4ePNM2K4H51ulgFR7uwFv+oBhnCJJReT7Fk8FGfR8zr9Knoaj
6SZTzR1JaMow8fBF/Bg1CGZrXVG+6XuOiPRcfxkOxJztPBmjCZrJ92c7XMnehyTrDWPhyYCJSDqi
gdbegb7aNG19Wh0q2L1rhK870yTIGJcltDYmPG7ApuRLSdrUHuoVFz7XCZcIbg8KXWHigdutw7lW
HWsjNYvedMAlcXXD0bUpJF0SL65iY8cLKhXDB9tXG4spOgSqaLSj1XTRTFuucdGMaa3ia6rqaVHj
3lIq+YWZA/P9kHEQhYUipPDLEztf3XuAEkfWLq7Te4RT3YJub1NFeYVmV4Ygpiv9jJe32juDqde5
nrfDKLDNlNi/1KFjq0UpAR7mjU4UFwmjdIeO5uhkY4vd5nlh+K/FbhZY2QATZmP4j9RuVpt0UkOv
5+ZSai83bLlq28bkFU9Bag6qgWxJeGucf2a9J1/EjiPcjJxucOK4lzMa16h8C6wSpl5k9OVQDfIo
C0aT31k9M7Ihhv2hLr8vb/hXrS80ewNkG0mBXbz1KB5f3okJxUCXDHHl0eh0WJm28/pazme/DTrE
N9vJ5G858z2nVuqEPWjhuidMFZWlkKTMBVCJ53ZZ1mbWyY0xMb8b0HBpme9Pl2qU/Z4AFW+kSSQp
Ww/OtDPZ5SkdupFmttmZ+sHr/oxyA0p2DWMffZzvz0GowPJcMHg7CjBSbjae1k/XBow87z5OYHnz
K7auHUYGnkgm3pnpF7FDGf3JRxZHwYzW5Sln2737gbKWJv/O7EROTyg4/8c6GVj0kP01/BnSimAS
srYEYp1NXuoUjxJ+LKvvHq5vnoWwhVdFrMc8ZkDwXLszTUdxcnPiwfVItEyCB1d32ehzrDAVfgJZ
ukASNswthwAcJhGgqIbEuRAO4X3nkC6w9ftPD7Z4KIVW88jSM0Nu2JgNVDurECYfQRfwiIufF1Xz
KU5hIm8/4Z+tMGNSlrRspkyJeiNiaQ9RHFKVDN4i/bTzFjAZ5UctSPjDkVucIJ5PkZ8YVusDW6RQ
o9gJQA08I5bFWeZtFyXMfuUSwbQMHipGdckXmLQFhCDVdbJVNRjDBhIrk//Ew0l0c5bshaPOzUmJ
43JqUk3ixwJh9phLV1uovPp05Lf6CILWLgETLZid1oAqB7ShmsZCQfb2bB0DwoDvCwNTMwEHKrpB
Kgy+GKnUrqMU2TzdezRkuBIqFA9mHO5qGTqw9I7BLpf9fDZoVAkvon7AbS2j+SXAaE1fRaGpV97p
YxpwVxK6HLgfYlk49MRtxjDZ1qFg8jGMjxFJv7Z3WnwjQw0Tmbtdb/fAaZJzp65GSZ2F1DWkpvYI
mIAByFbwN9gr3RAHx7uvo7zYc+nT224h1slt2mgRc/T4c5hxSNjKfmF04n/x/GpRS3SI/gy6WTrN
JIgOlTdbWz6At9EoB52si0Ug/F53+CnylwuV4vt0dURBccdGy66Y0cAtlwLhlbw6Z6TGJRbUZAgZ
iqY/LHkly5pto9ciRxgQqvFOTQGPYNO+pbyJuxpijKXktS4WbjupnkPghdL1BgfXfQ3Rdg6y/9n2
Jhvrq6kVTUj7/S+aY4HBhJF58d8YPINxWfLRgyB/x14BUsIYClS/MJkrbe3nYyjuPDtrNiUfM7iN
RlXGV9NX2Bwx/FjbT7oNopTMLV2ivfoXkf8HzBxOjW+XsIyUGcIRpJ+R2WDo/wGou95yo1/T9uP4
NgTNE2YPSuViH+wUYgdJgAhCLAINOP2XOVQBD0tCr46JoUviKt+dvWkSKTIK8ibBE9zHkozD2rXY
viozwfGWKN6LeZmoTTD4vcsWXw004/K/FWQEH4fJ5envUfjZpeH34vFus+NNqOQElXy3kRNKG/re
o2nzwjVwfi4E61tGd859Y20IF1M6xcUchXni/nxyEFzHUjJXwk39FikD+eAQ+Se4JJ33AaKJPBzB
OppIP33YEfyBdrsUEIDDqzjZv4U6wbGiEsI4kI4QCgQ+fs6XKqwYF7hbfShr7Q1qwrk2R0FC/OCd
SSFpOAMCcH/DtlbMka0HfgYr67ng5yBlgGV8rolW8nDdzQFHgCG9cd7MIfIe5G3MWckoIQsQ3L4P
P1JUC/s3cGKLM73Wf/7lxGFeuS8jZmWdx2vniw3P7gigrY24IbobTXHMzSfNqpOodV5PwJ0aiegx
rLuGBXa9VBTGPb9vYEkZmSLmzMHwGPXVIPNf/GxehC4fYeelS0O1iU104Bz7e7fYxLxxnpf+HWHl
HHrCaSA8pCYIU/qDzXWaT9nD8U+6u+H+M2RSKUdyH7cc6nCKow1HVLEBYFDujEHybtKgq6wOJnDV
egIBeUQ/fYvkoEhvUo9uZ/oMtecRM1FsEgd7V0u+Cr06POnoxy7s/LBFQBcirHIFcEms+sskpeVQ
b9voBFcGdIeuMcT35V7Ilm6BFDMF77kL3n3GKGSl2z/hpoVDWeHs/M3q/TXh+shdE6eFd4N521n1
qKtwjyee2MitnbeI4ZwWI716caEezxUGR+Nond7h5UES5UOUFR7RRq/BDG3cKOHfr6Q+EELjLgxZ
Ugp1+na6csKAGk3u/92Scf5k+E6jJ0T5nMEux8HnWp4fsKCE5ZPF5I25INhFNYOaUuCmadczd5YM
h1qFnLuyxc2A/WlLvTiZga2JoAoeDfnXkjZvDggT8XpCykr+pZUV13haxOakOkKzWFOob7gRiAmX
Shl2DsMpQIGBeNwTqBOpGtf1QRDeHD/lgwSNpq9iKQ6zpsWLtAba0IpB4DNLHoLO9tIRmnPWRE6L
pQHrO9z1pf/KK0WbuwCFlLeUIpH/7JE2EO65b0sv+EtRLZRfinwAQ++ZbSaM45la/TE+HXYSF08k
tQ3bU46yVOAD8LzTCPguga0PrYmYTJF2KGxBDtYkXbVXTLrsMU94DpAnGEetgbzXJf0MlJpoaOY+
Ryf5fDjTSMD02Fb1aTum64NiWYFEi6SuVVm1mDG42ubuWGz5F1Ov44oLeN6Wxqd5BqpGgDpMTP1T
Mk7LEwjkdsCl1BHcMYT25IEW99bYHBngSewLDjLhjRtMKtU0R5rEIFjmTkNcdgM8u5Vo4fidA/7U
wjE25FLWLyqF47xg1vN+XTOppWRhNc16MbxaJW7d41Wk+MdPAK/1M+lMLOaRENRUOyvyg8SVFEMi
6TNL5yIwL3jbIQK1f21pox2Z9ZNRyT0Bc+36pt9gfmbkhcD4Z1pfq63Z57i6A6VgNyeUdLsOhtXg
54R4RLpX/EYbkic6Msmwl0giEe++dnFRfG32rCQM36YzhjSpHEdYbIYvOjo6z4MYhkjj66pU0uZ+
vIXC9TasX3L6uO49aycuVBzu87lDcjwTydsKD+i04DDAAJzUO5OC4vJExhi7BZKDlEXmSQKdLCVj
0OaSyeCp5PLsJYU7B3foufIPGQjr3NpHQs73uxSNiL16ozvaMBB2qf8rdkVj5bGg6YcXpl+5j8W5
UBMBp6XoEkHKqHP21Na6nkJyEqLhExqe6wBXeuS17t0QFcepL0NX466eqrJRFYD9le/iMQPgt+yN
BMWSrPBwH+iwekig0Ufh78KZuQdL3BqJIMlaTamfqgHlKuaVnxa+Fz/nmLdohcWZFmEYym/LdvSJ
2RazDhIyUqYaWEiIgP++WSWcHbjuMKtjTxG4GaEgnUWiaNV+xApJFkAcYD5z7uE66j/UfLFIewg+
AtCMuVAsJhoqR6Yz8vK0njmjjIH5PpaY2it5j4sw65kzUCsJzOcEuomjtzrI4YBFXOISlfm0wev/
z4vG8g9uQ0Mr/D0Qk9gIPrVmtrTiDBixVZ2shaMgiagYt2K8AMMDpTKs541MNZEffsYok3bjNC9z
HMOCEpUvzM6HyDIoTndBLeKZPUPtiPuXFthf64JoaJfH89pg9mruUavwnxNc3ayBUUIX+wgrOyrb
GUBSeKvVnVDbJEVzKWrKlRrjstxl6oi7Pwt702B+LNO/mvWNFwakZeC8AXikhk+iRlgMT1hwH6zh
+qNkxqG2R0KDy6EdeOEHjTV0zPxqop9NS7HuBhG5Ggwf8tZdpKssoDol2pUIZQyMiH/k1Ys8lLwp
ILIJR7f0kvx6+m06FFVNCvmCqj3uGnthxC9QtNXDZ52+9CKZFFVovZhFFi5Zgod1X/ABq29a0JhJ
18osHk+3AYDuQrNj9MOXAxp4sZmxdiid4x5vWJnYpsDhiHwPhqNA4ZNhcBOOyKEiupLLg/wDB6PV
C25dmG0OKhS/Acieb5eA9A2fXEJbDB7Ur2ElZzB/afwKOjZ2bCp932tIkdDdNpL1sts1qg8Qug0p
I2+HtBpMfsDGRJnFM3Tx9ZqNCf9IrBEga3PWHx8xCyfGFBwGoXsjmrxVsl2q9a7BYm7FBEG2u7sT
z6lIgTRRqpG5YLAwWpC3uOaWrkKowdClhHIDR4CuDB+CQvhiNkDd7yECHwW45EVnTH92y7vyNN94
rPcgicaFQYhs2F8h3vvAp1EH02qQ9h3WBNttE8CuxwmhT9WAihKysARsaLFuB3CJZelRtTEvHLu9
P2QK5OeqCegxxw9RENPjWmhgDG0Zq6kNYzURfwC6xC/e599K1yWpFRwrNAg+V+k/Q4ay4o4wY4Mr
tZW2AvuDaPxk7NIMrxLe7eJ7JfrR+mmjc51sl9YTekkMT9ateyQ6BBLOgxGzsizkr1u3hq+g2jnh
sZuRK1IwH7J2X3cqLPMQPfW60tB6/GqjXNY0acxA771FGUwy0vN++JIrA8WOF/6FOi+Jj0pfj+co
ZGYllLKGD1JJMCSaA7R5l4YGzMj4Z/EZZCH9+dVxeMf2gDtqoRegX1gNBpb1A/jHXupmrQosK1ht
3CWKfVPNowibc37zjFgcZc8p7IjejfP0AmSrR+E8y31z1blq8xdKYOxNZepZCdB0aodz+LibvrGs
lV+EvtpJTf9DXG8yzaHYir9agC22AnWf7044o5+xwz4ao9eeLT9+jL0kvJ3tGaWjY87syyFqsOky
/BfqYrKPTnQLE7Mjgmbg4soNCOinS2aygj6JGkKv9paafK6ueqPENvMr6ILxwaM+JjN6x49kESZg
Q5aLvHWr4rNrg7i8lpXOfugY2fUfrK6hh94h8OFdjfj88PZahcWhXiW2PyQZc4nnPn+THIoLogbU
VDxs/CWrE7w+zexX32BIjqlQoLbO+CgCBU2O6fvM+ivWG5KTTs9lA0k5PYjF0eE0flpIGvAw/zyN
mNewLgv5U8aKJ+uvauAOktrVDW6bcZtGyFxhViHWrPuGiYSRs8RcHRmCIBjt+s9rQprZv5pa76ac
ihdsoBZ20NvVFigBJfv0Ilt7wbRJMjYH9Gs1DXdTZ6MG5dKLmm36qx7S2ameU08mMlI/u46W9Cvj
84aN/e9PTeC87ZhpK2eEIOuo9r3E0604wuo2js5YJReJ2AGdhWo4fEouhsrxBD/lWW0aiNq6aMHO
Kt6X2sMTGhegDdpY7PBbDrwvF/lPhjTJpdXvO6MNJIYPUZ9O3pw/d/NMPttgqO4IaACdeemUlz9F
6/wMiiCA79LrL8/m3KADCIpjXK0Al+X2ok9JARs21wulUGU4qEFJvQV9aIPWUGxcvuR4Dj3PD5Bc
QHzEcxuImnnqvLeG7gvhCzqoD751hnZ3OwwgGgLpNv3Gk4BtX3iO/3TFsT+gfyhlyV8et/AH3j+k
zG9SI3bq4cYgU9Q+fVbaDLNscVz0oOyGnFKc2PX+bMostu4K+RSpA+yDiKisMVtutM1rHOQJjPK8
tSsqWeMoi0Z1isZSIYJkov1bl20Ti7QALS1xmTztiItJv7BTT0yJ5MpHp46+fMCtC6JvyrW+IDaz
IaTdFvTCfTwDFtDoOUN05XnzpGoSJtX5OWT0uCWNpq4x9FlAl3hR6OXHe5DomTzcYGvvcNuciujr
cucvjw0KAQsVFLI73K/75AkOzC73v2czdQnUNKk29CXCVFGN+VfgWXGxeg2nCGGG2WDeJzRQ20yu
Q9Y6uziVcNLs3pAZvelAadavt+gefc+FFJTTPDNAhL/3O2qnTcfokIMFlz9ba2ZGmcciYTWF1WBJ
EgL5WCqxsYakj0zv/yUeYrLkDHCs5OCxoMafFAXVfsnNcEZhOkS1XAkk+h2/9c1sdyosypkwiD5/
saFo0yD1YDrJfUX8UKhkvC6yFmGf5QhdT/l890G76SCeg3bC8qLBm1K2DyouMzturcmRLRJHVtA4
PAZTZqsq7GKWQJ2zK3m1lZY+Q6jPF0tlhlT/BJEFqR8MFIqPIqGfSPvIUbM84/+8GRVEsaajDo6C
/18Whu2TwymNX/mRvWorJeIXzUUqcvYbC9rTlYiWJWF60zyB4cmCnu4yrqRMEI+p6wjC4w+PkWOL
OYDWHkOtKOMp6o2YH/jAqH7gabGisEFdTFcY85tyLdDLv4ZdjnfcI/FkzXQaaSt7ynJntufWRIct
wdM5lRvz6cxpyEwLx+9pqtlHAUXGDmAz8XDOZUe44VdwlzdvH6MxvgWO/8/JSQ9KW/3juIrSz/0B
K4+Yolxh8q5L9V1zAz96qpMlNZYEo1nE0BDHPvypu/7wZMMftn3DTVlaGA5qhyFTsWdxQeD45XNC
vuBF1Bo3zA9Wdw4vArT2k6EiAy4DewnoMhYPilcxhmNZLbhNkaR/mA9p0eHfFsMq4+Le7GkcIjde
AaWePAnqX0jrmHWyhUSZl8Q+dZQeXsA2eL+mtPLvaqqmjuSaA4NykSH8KIYb5Yh8yXg1oN+gaQAP
YsKDptKfxHrCpmZCePLu5RvfLldJc0q20f0t/I88OgQgFHibA2IYzXlhBgOp4/JK7rLACWAf7rle
H87lNogt1VSx/aUab1PQLtePRGtGO/RNp3zeT2duQlp43xZnAHHrXrdG+tLQgx3WFaoGpLatLavS
z5y+ezTNPem6rPZF6pD4KpDQsogObSfpsEOiZCyOx+D11jUVtRRGfsmkVC89cmPtE36ChCu0jFjT
ofxCbjfb02JeInWVrK/Ligr3oZ0LPDZr4RenJHIxGeX/2DS49sgkJBLeZQYmlGeKIw73HU/Vk40z
0HZGoz1Ka//j0kR7aKkrESRottZ1NVd8HCB/Efo5/uhMLoIwUjhLibGyKsWwA3TlkmVVYUnwIh55
2fJJM1rdlk6vGTDw3zO9PfUgXWWYYbjGYz2TE0GEfQzb03JGLTexTh9VC8ReqDyVw69/boEt4WEw
pjICQ0XZTN9EKMw4zj97p1kkT52JTOa5HwrsHTMtiMNLnkqD19DomXa93lcQ6b4JDVsCGT7ZgpOF
mG5hOLe3H6wUarft9aNn8rxzdCVVcpBOg/aG7lP9LVfnKMQffkCuYr8GdsW39xNjOlwUu5p0Swx+
GIvtKOgd8cEO841OGIOdUo3VL/3gOBI06d5NxNQAzzznbPzoVyTj/t3nGrqI1TqrJb01YRt5Spt9
C0RCUTxEjHI+ywLVnqLQn5D+ICT0P/nUb0Lhj5F6WWN+GGTtI8rBgntpDRUSTF9JH6QYpEqCyGiB
BUCfogqZTKkM92GFn5H9/Wj1SxPNJMzggWXhs5p4/QBdXDzJJrNzgL1Ivwe572NeDX34VhPN0W8D
p4b3GmkzrDe3dZbKZPH1cXtFipT3gACsMUJUPPTWaoaKz0EhCaYtL8jwb/7vmfcdcg/d+f84tFfw
L9FtpOz4TLdWu9eWtnb0GQi4SkyVAeZVNuGaMuqv/AgClq5GvL3vo8tzhQnk9NTckOUi3U2kXM0q
zH5nQzdEEP7oPYr/HAzcsFw6+EhTsZ8FW5MBum18QnEjLzzHoMWmNOINi9Bv2WY2KjLALwdbyOdP
4TaXGsUOC9pwhZvEEsIcOyAI30eAy5fuEhT97eobIK+MnB+7ro0dYLK0ReAXEz9creRORT7AGY+a
rPqyU+OAjS1U1N9YGAqiP9OeX4bQL5UA501g3m+sgl/CNtZIG0GrLDwEikIsusfy11+vgB45mvUW
bTLHgyy9uMIIGjZ3RO/lqj8xlRDH5QeUrSRGZlz3jgvw7GjeEEy7q71ldJYy7mFA1KP7cngsp5DD
DXW8dei9Xh3XKy+WEXr7YUxdJrEE1d5b3FNZ1SvbofSHTTWbGpcXTb0dJDzxsbqYMOL4HxpTle6y
7AX4WuDAOuBUDG37gsujzopXMHU9gYVGDqAHjFocBewkhzpukHbIbdglEEPxu15frI+xfUYl7+MT
rqCBU2iindZ5gCoAxH//+Upo2sXdg/s7hu/JBGTRra7WE7l78scNZSG8yIuVXn1SupKzctOCaNCI
B6PB6TmQdu06g2o/A831aJPThe/kDW5n63z6yfV5TCeZ2uyBD4ZsPJ3+B0+PBQygH25Q88WZwvP8
5huf/CFAePFdRCNVdSpDchrRVmGywmWv29jy8swfqDpl5HQwLxBmIO4zwkuLxeQGmP7nhTavZLFm
/9tniCAOs/cl1olN52pjsgLML4d6ps27Hh0K3/l8T3TZuxCt5GdFc4TMerIfPZ2eQWaEdsIM1G/4
3ZNseSMD+Fhd4RKcS9dEVyIHsDisjrAqR4ZVXlvR/VpxtTR4KEuJD7sjHnYavfpIfQXmP0IMkZrG
pm9FLA7ZuDxJK8U0B+bE/8V926Uc/ZJSLMRYRJ5GX2LzrnN9CJz7hKLI6EmPktZXG7T1eEL2OLR5
MnAvgfVxFsaT9c1NyPSp5TUyHgV/QzgHpnjIY/gpyxBnzS1rtlcQfHDKTAM59NTEkDj2ytbQMlo1
vvEgtbVCbxgeuxpEre44Kek0gPfVB0behaRaKXfyqaNuD2vW7qz1oaMsv/tHpsQEkGwHcJ+Rih/x
t01kY+7ydAepEc8zs4doTAAzYCImOV5+GIh80/Ct+ycu7hYg1T50YHLe0s/McZlJ7n14SeeOY3sC
luXKZFqd9BMclVu5d1DLp10ym5IM0gCepM261AHA5sY4tFHr+auoua93MDJWq7GIKukmAtm0crmp
8xj0zrLEwsHti6zdgKQu16ux2lbGeuOAvGj8RXJxc9jtw0ibs8aV0JAwjDml16etq8lVTVaplzut
NAdk7rSw8oPhlsoHWuBqqC75MQxxz0YpvPJYkcM+0vhe9nFI64N2zoSPHlh1bBdbtgcMYpguOSEI
znzJrUT+tJ0CrcWb4dXOZvw0HKtOWYBZkf8aFc3NWEinDOSeKYnKOE6U+mgoBSCzHNH0cebZYWVY
+Pn2pYUNv+Pk/VaNx5vDGo0vxgVjOXbNSvAT3+gOnOaYNVpIwQhoidDfGJYmWPhpCQa+v0KEcc3q
m/pV6UDz7BlseJbyEmHNgXOci9rSE+teaHvwx+zkIawkMDT4295r9ZnBD12n4L4pOg1bBcYw4n3H
RXA5VKj4J38EvX+iwkvygp0BAEZYyXLiEMG2GKcp+INbVbQkW8bPRHh9Z4Vg/CtEOZhVCr7zmC0e
V3dNvGB/BUkQRr+OCZLuMUhqr9l4hNcbK5pjxJzEW5Tp4ft3JbWBxPlRy1vtiqyu9EwF6b9bscAS
1/DqunrTnw8dgv2Im3OiPxlSe9Xymi322Id4NLTC7joWpGBMVbdAEjyp6WRL5eE5i34mK58pZg2H
w0lEybHTL0yRCsFJk4HZixKXBT2c8FYcy4SeoQwWr0D3nQ6S9E0CrlEmIbRRRe8EyRQCF6zKieev
yln1Ffj1MFqISPVmlGrosqsmaIgBgYiqiEygoCYVrqHe5E0dCfP8HIbxbzVJ32+K8MKyQjLxTeA9
HYoUT//hra3n//xSP4mFGsGwS4xlfknabp30xRHhdvI6LwT2q5oXo9N7w32jDokjnp+K/Pnjd7RT
338hpFT2bCZ+NETdgj11PbXIoWZdKzdpJTrKW3xriZl8/dTi8zt0rDKEsl3X1iI6+uEOXkF5WHpF
6q3NVV9bjZlt6xRuJg26EDTzL6IRTFT8IjugHzPodOkfRMvhaTwn85baWbyZQxDDHE5OS32SW4s9
tFTCRHYre2hnmHCjNxTKZWTifVUsx7CnWyGGoFL4aYW2DKqVg5d3JWgIjh8ZiyWEtMIkeZhHbRo9
mNVxenTn6IbFEu41PgXzgfSVp/FGjHFRQUIycI/uFWHofapD4bIBCMf5/5SNqlHu5fqdpM0BapwY
zNHNvAH9r10uaYsywy5EpZyOS8twdM7GcR2KywreDD9nl136SP/s0oyW4ag6rw7IKb9D/0vvbltI
2r5LCJ1rNtEE2q4Q/AH7LfXoH7P/8s5KTVxWg23j6V27kFXWPN+aujss++jL2t1n4bhTKtFoUfAd
S3hzww4rhzyHUWU0ZHrJ4+UDJM6PN1da6/C5itcSb6Q6Hnuq9NpqKyb+w8eL9gLSQsjnBLXc7M1G
wjeg3iI0a6nhZnoI8skksscioYXFZU/2/RIcsv3Sn0XMk4sFMsWL9yic+0NnKYBs/ztSUobIZ1sg
XQjwmpC0QXKKv1do4D4q1jGaZ2dpqeEWtoUL0O9Tkx5YpIPsGaMNCiY/w6IYq7Yhl/E4XheYfaDQ
Qd1XqXyUoAgB9pUrhLbMAfhPOVIj42oHtdBxfTtdr831a65WzEHdR8Ec1HFmGL0oV9oUt42ht8Bu
vEspNKPKkXXNwCZ4++dPSHP74M1VgJy822nChrPE/e8T1dDMqesezxqPqGd2DTcqa+eEaoOdF7dz
q3jBt3igMUjhi2o9jjSS4EMahCdFdbu9wAJ2h8ErzjNKeOalngyc9IZvtyFzdp3+gM0vaCL7f9st
WvID0naKoZpWjU/UHGJw2enyk58rkoZVkVNuXXWl9SpO9t2NJ/yDLjTMy8LcnJsl6nwgocGXeeaq
IC2mqIcdwVo5Av+i5RZk1HaYt91ID0sUmzUSBGWDNn0uNzQVSqU2PsjvFQto2lZ4RwEsy5pYdX0C
3NYBQx3JGP8DfQN4ouaPVTMUosvFasBpwzpAeRHMW5pXWnhsFWoZ9tCtD+zHro5+XoOLw2PEzhMm
hiS7lVbE3PrwUMH96kobZKZ23Cy1WkBYcmYqbSVDbP6tfLEfC7Koog5wfosJbjJvduLiXVJFhYSS
dt5qRyQ01YS8O5LfDzCOTipjYMqr/pGjC6fS2mb1YAQGboBDE+076UqKouoIBHLESYcHCBoxTpUU
UbStmKq8LBO3YFdrDvGmtiKvVJ/hKPTEFT3sSLhUTDK7NyghRWIAyJcIgpAtQasrZqJuSItGFENq
mKlLTSpNWbbC2DXJgWJGa9F3ZUhKgjbstR1oZAEb7pWodPYiMUp2Ao1WfOEG8MffssuZFv8k+yxt
f0g8/9mDcohw/Rbn3NiOeOG0Vs/3xA72zP7Tn6NuC1qjl+DuFVCf6C/EZ6K5r/DOdrigu9b/Dlcj
hPb7u1n+TCWaUwjccyqRF3PnswH0bUOehuLkPCQjvpeT4/+6Sw/+Co8rzlQVg1I1AyQxu4UOldcl
2NHZUqIliY+OoajnA5KIBA/iXNJOTzeDA6L4opR0oRGExMVDJSRMNaXVeX17m+G6Lbp85TOZOs/E
OsOSCGLCNnqaHEqEsZ/I+nzk7hMk8agz22KqrXV0tiL/ge5GnUXOkBQ5W1K/rJmUqz3xFNAYt8Xi
eYVk00S3NJfYOeKuezA4EEnl5arBQIeYT9YsIbKAy6kNroTLUBi9nFj9YV2+SkGynfPFar2dZEui
iIBlXCjmqhSgDCRAI6WMjo9QmRi+rlfwCPoEq4hDmHZ3N2UB+Q3OCvRifo1CHnd6GsrBxA0HQ/2L
SyV8razRHHccjm1yXa3Aq2DhlSIl1PyZTsQbiDPGN0eDe1T5bXsbvm8OnFPk9BuVewmFA8YkhT5P
H/zRo1pipooiM1whrDVPsGdpkrh0L2GlWQtWuKJJTfrMIfmodp51oyYs5vsVxhjmdY4vdHKZichC
NkH8LI3tjiAlCga7PwAupo7phMOmukmWEoSFbGsHQOPkZfrm74ePsmQEPg/U6vbUbt1NwmbuKKob
Ga7g9Gh9C7gZPFZ/LPvPgEXZi/Ih02tyZ0hSP8YPUOmOGI/dEjkOAXDQ57YKdnaQxtvRNkdE4Vtx
zBWOKBmmtbh0r8jM0G5dnWgzAoXYtp/mYmCn2hayd71NfOi3F0hge5HaTq/gRve4ZUjQoLtQjUOq
AvA0jfC239sEz/Flw6EflA+HMPgX3M8hie9XCyCWgoP/BGwf1fPXFGvxBFxMBVyFvwG7tQ90DL64
0Yyr1/B3N6UbkoxYqa+ifxSAOIXsM9hocaCvz/4SrgZ+m+spu9TvdyNe0aqyEeMT3bgsik4s6QUI
XctMbIJnPsS8mZAXOXJoyap8PzGIsdoYNW1mp2CmrjAxxqFgU5m9uTO2DQaOfYswuckYer4YQXkU
pdmRcuQ93F8p+mR7Qamu/h60NYbusr7K14vUBwc8t7lcBEBX1j2I99XPVAB+gCIQmCf6+WCfIgqA
Bc6C7UNs1/57CmwYKKuhaZAaGL6piuik8EEFEDoAv48HbVs5XJxMsyc8V7iCoJkTu9JqOdDWIcZT
5KRayUWdx7fLdzfEQkioVo7KKwEYAA308RClaOgNMsV5qITEfRIC/o6MmvM9JYtGycsuLrosIEgn
ONC3LVPOfvLC1aJjewWG+M5hk0hbiPjnzkpBj12CS7CuLz6Asb5RxPPKCULyZwNhY1Ml5yYIDsG4
EHxnir457a3XiVoRu2iBZU+jGVIQNj4dBIvWzqCh6HU3Byufiba7DYCRAzpE9GYInZzcSDZs7iXe
dZ/quoQ7njHjgz3EpsX0MHJvGleE47IEYx/pWeAgBcl4Ula77dZgAv4HZJ/N0nIq2Km+kvm5suQH
6EiDehg7UamoC9S3KdvVFsGGYBBHapgtHX8MOZ+A9c44c8TNhZstDX7cthKOuaVvdxSdrfeFuBQ5
GZRKPwp0sM3zkHAU1QNyeuz3Mn8DRxurU5Ko9smoBukpsJDA7c5mEfr9oNHjt3useSiOHnsYqNAN
eZvf9/j2jPfIXtfGmSmI7MJXEvLjcUyfpYI8aIIOhcFT3ZzPOqYcZatdWLtc7PHi5wgSZRrL8ONP
Wnfq4Ec/5HxhVeTvXwSNw6yn4CH+K37hNvTgnEFz23mEXv7U61epcMFUUa+RbqQ4t5LbqWrYqAah
7/9ebg6ZJuTv+SlPnQKee8lISl/ozgd4+Lq+t08JjHPYYr+4Xy7FzhQToMFE+Cc+jvyIPSxPF6Me
CVHNCvWY/SFBEnMEkIsFD69iHj19ctkD/Kih6+CY+o5I+Tc5f4vkzoGlFLEHmZW2GmmuBMLqChmw
clJl7JtT3OuBDT1/PiM9JJZg06JP/O+ehD2DDHxN2cGu+4CduHHV6843ktoBETFvSCXkqHZktigv
T/QEqq7/CyCV8FSNiDBlnuFOIBtfeTzVzkIQM4JYGmCLvH2AEscDA/EYSSwUxETRlF8uFVgxCOGe
oQTYVgiZlM0hd1aHiXk+koZLFjPukrV2vy/1k5wA/Xwp5RMjrma9ibUd9HFzoWCGiWMcl2F0JStp
eMLua/zQC759dct5Q/rlHuVxwtiM14cdFu3WWeNckVecx/czl1Hv8CLv8MftHBGHGTMxtoB4ygBW
p+8CP4VUyaF6i/oXWMu0POiMRtWyk5wRWuY2tvAS/mVC6vi3GGq5QFfBgnV6KjxTRDpojvxJOth3
lVanAqIBDhnT+JUt4lVaEsVyOD31w9Sae5s6fdevEpXRHvc4Q8tafaLEjsYVz5hTCv4o+OR+M6GQ
mdlTRPiU0Gasx8+CTO+L9mOcKARKPn42q1hk1KmWqbbcUteSmAs62UkHutksIqz3k9vt+94a9xUz
U1JcHUrrzOtGiJsAB2uExJUDvZKFFuC+7/SM1iq9IE1N7sF1llEC8z7jAsFeFWO5tI5aTDtOBd7x
DI3Q4IV9hL3thpmmbHBKTM1Mk4BcfrgeMagHTVF1KU6T0r7IJ/MnLKrG8f12Hjpj/cbWZqsPmcgz
Z1fr5aJWkfJLwZzU7rw8QSTHcOOs2Ndbd/sbEmgJABZ4yiDGZQONWa7m2GzDv8YSD8BMuBWDOryZ
R0BvulJub6PBKuV6LXilrxKGSZ3tZ9JubCi/VdVipyoCFj2cT9a4gSypwmJdXAcUdtjRbDUoR7PO
Smyz4PtwMxOz0JaMM03sm04iv9QGhyvABQsfJ+v7SPLWUwPDiV2rKZNoWCLQ0pZymkPPTUo6MQbG
y5O9RkXkNTwmyUPQWrBXXP7ZRE7jlltVJr5LdJ3pLwRFQVXKej9hpaa3994Ibl6Y6Y7vqyIj4jIl
Urk66fgLwoK96OKUXvscFDGwZ5azBUA1JC8d+RqmUwPOtpLUn2lQ4iN/SqQqTF0uTFXsA4xiVLnf
A8P9Y1ySafO/bXp2CqsFZ/Zbo3HOW4UobZ5BHEredgEqWJw+FcJdzhE9KDqWNS2OWMMRWA/xpfyP
TZo1CwXCBFWbs+ZqzUqaFy8f+9Hx8yayL9FJ6CScEAxjwq5ORAQZALQLx5AjJ+HRoP3dcfXDpfYW
o3Zs4AJDltuxrdn8TLmv3cbl4c6Z37dLN7RvddJQQRhEYRSWyOJysjhhIbupQPom9/c2fNw8TDrG
GDegqCDiYyWO+5LgYFQWsxJBwHRHp5dNxrwstI6eSVnEY3RT7MTcejyTLtf4dNRkO4r8/p+4Lc7w
Em3jWjXku3aDcq1kIoFBH5FDoQeEIJSY9TTLFe7ZvlKe1KALsR8aTMHJIcDL2ZoN2W1tlWhkaY3J
veaXemjQO5xkNnzO3d7TVGD8mLmTKQqWUP8pS9UQEjuGQ8AAahi6SY5IjVQ6GMc714Oi3CXWoAt/
971mN9/m2jJ52T9D3wdrAnH5Y7GKtHl8n4oy7n42xPsdNwTVZFsfQEsxhWsRRAKCllKLOJweCimg
rxiVb4CbOn/CPfRA3Wm5NfSe8TD9Sba6GJV8NHLXtI0LRMd+iOMXHJ6EyQKUD2eW/s1WzSlJ+9sK
oo4d70kNzl8jy3hp5K9Vsqa1mH17Epv4hqpa5v732gOUnNMcBowQHGMEWmd35Z4XWluKGo2zy0x8
awIihoCrNOIMELF5bC6mxcywgHZXNdQW2musDz6uCiCaJS8YFhE1SAcuJPmM5eBPFVWDFWTw4zFZ
SIW7PlVDIW2XK89fF/AWTckHIEH9siU0DJeW85rRPkjIWrxdtLox4naDYy69oei+HyEURUx1J7pQ
cht2YQ6irQDJCxGgKl1dMj/H6ApCCCoEVjQEVB2wumaM+wahHn+bX7GxN//KwUitQGGmMgu8fw31
AtMgSOECSEONKwB7tUxxgE+Ez8+IRc4HXd+b4nrVuZsuS107LUqRoIv/GYbF5pAIdc98zEZ+FN5W
6BZWrL3SVnIJw8j6ishFVIkH2DWY0H9i3pHIpqRu/Am+ybwy05f1oHh7aaZzlauNAGzh/ObbdSvL
aIZid0ltW+c+Dg9YXcuB+qdFHIArd+463TmOs14F2GDJT+DkpOYcWsb+lXIjzhLNXWDBjcxL2FMk
tExIedfRfsaN+6pW2uqjHxYIp2u8uOJKomH9qCVO/QNxi6k6e3AB8JFNloXVOBH5vV7X7fM1kg3Z
G4Uw0mej6Gt8a1dryEmdhHsNQ75piG6XXd5VyxMN5/MSK7SjQwzDUukO2qHd3RYJEEurNtV426u8
+HNu7F9R1LSVuIsvgjqXuEWyGpZ2HakNPLjkrgS222T/ybTITIsr6mn+uLtatq6W6RS35P9nBsub
doPC/7umIwR8newvmVHkw6nVG9KukZDQWda8YJsUevv012EMczY2tNTZzs6rDX5Y60sDJT2yqHx2
gr5bXfO/AqreLkqjaUZZc1h+7QkOa4RCIZeataleghOz7Gvx3L9hSTH976GDospNdn+faJWbz+kE
Kd4uywpoPxeneKYyOVuhUIhj5NvWEllauZ4o+RR06Dow1sciaffgiSIPjhtkok4wZLb+IfTVHh78
FHKebJlpOfs8VzVUGtbTDQp8rVsDwh87mXfiNcpBM/cw+4FIK6CO4yXTKOQa0hJDE4KrZ39uNLx1
iZH1BtCxA02prIscQDWI6ifbX89d6D6yKu/iFEubAoTJ+XUeOvAYsUr5CWnldA1S5CioScDsLB9/
NN2sj8vJhtEJ7FlfhtQblYQqWmuhdlmjFLEVhmAAj+5DYGsxkS1CzOyTw9/pP2bUnIRoRTaXIgYU
EpG/i14Rxq+lKdxduTjSGLwPvFWx3vOa2H/4zo//SCTV+O4MBLauHIjnNGoYXcMriquT+SPguPer
XtND4/jITd9A94/q5cR1z/W1KzEqhcoeTWaZPy/q8pDRwMDSuD2E01Jn/4TFl7VGvxedyM3XZt4+
4+DfqHlqIgSwWZ/rYBkGb9FxwJJfOk2/4iLHhvHARTqyceGfci23UxqCSikQV2arJeNTl6kTfR+n
JASmX2vG1IySL1nju2rQwKnpc5R6qxipf4UE8BsluuG8tYhTVsOMF8eE4bA+UiiO5l97j2r8R7+U
KL6xdiSJTe94LEiQRkGVXyNDJj/TQ7Gj791ZL1WHA7sOrdQBamVw39YXbdZ/A/TBrZECB+eYdJL5
myznvyXeX4UN3U6AJ3T33jojDQaMe9mbjmn0OHk1z4H2UH6KhornUMklQy8jOCH2IO+IcM51ncBl
EuRqoXc8QS8kgAtXDVEsvz90iMJL123BoUDvTNu4icqDFBdi2eLjm9MdphNgZiCEM/xN4EVjG7wm
cYSpAcLtB+OEgcsV4WYsTn3AerZZk0sok/JzRyt4FJPehHwREk45u+UBWv9ZpoleGpnxj5VNx3fr
LHKs+QRli4+/q80c0sLXllBDUJ0oxs1YTRjLIE73KtvdZMot8tpQyDcCm0Yi+Pc3h8mpuLEiXjhp
5meo2nMNHKt7GoY4Td/8UYDWdzOjj1CtbGcXTvdDIicj7NshhGNYj9vwGzx/BeALQ46IloJlBxlc
LNDtzS0q7rhQyzccER8n6xqHv1rH/oOS1emDUwwpb8ndMGzerAJW1HMMT+89OlaVFpROb4tGGKIR
QevoUhLvGNjYLkKmy6kEtNAzj7Y7Att0nj9oABoFSJifW888+O+86Jnuwz6sVe7qRdZSG7JFNaEd
dmc6DFsKjR4l9M9EkU67TdcfEPb7btZvyqu6Q3An1sdWwUKCBww+iTRuDiFVg5oEWgbEnBj9nTTy
Duk7CRnZBDGYVekheEPmyu8NX6v/sBACj42xkKCUpRxq5ud6OSMdPHSJwhsEaavdFHOYyb7b4ull
DOxHhy4A3RVEAw5YiGOFn4H19nLh5D/WJA/2lxnU3Io62NsKROnvY+VdfwleQokG/3nz5ntVy5Is
ITclJZmHJyGPrrYDXg2wyMRe9Fvrdp0OAuDhufTPW8JQfFeT6wFut6gKpdZfTd9S8RMKeM7RdfD4
rJuXPrshu6bjmTP+UfS+dbfmU3lz2iiK+DZRlKfJdq0RDzZQBLZmHBnXSWZHyQx2YFuoPnbxUYYt
eBK1aLiNSeYw7rHFGXoLU9NELEDHbYrw+awWEPNVqnWVbyIdKvS6YhzWD/DnuH+A3DGuYMNWgyRC
ZlKL2PEhqVDJwYHDkppozlJkNk6kX7YOD0xbXmmm3Cgvn7rzNg5qTFpWYSijyU3tMo0H1jgJlY6x
Yh8wNhLGpRD96erInLekumXxdKJDP4HpTu1Y3jPzHk15nmEbtx+h2FJ7FqJzzsN6j9GACo/xe2LK
l+VwbQhs63vIQuE7Mmfin+xN3NS6BaX2rZs8ZJk2sg57R4U2aRAFQpJx/UZ7iyklHgET1T0XSXpX
MreK8VFSaG6cpoqkwNjOeUbxoHiVrfsjm0c77YZBl4IPh1uk6B+o4GF/joeNrxuwsH1Iek6kXzwM
zUghao6xg0dL65apeasoIcktNABT4Owwz2j9Ol9TtyBWYQoy32UPBkOL4BR9gX+q4Wa4AlWqDH4U
ywWhwAA9UpBpYas/pSGMmWeexUpPyxzA8Zm9J1fkq1cUa3hBv8IwLMc3USqO6y96FUtoOp+gKmIT
hUKdRKAV+HW6h7gykIC9eLw0ylnkz0eTZ/Hq5ehs5rq958svJQQ9x94y1mbYn5Ll5tGCkpcD8OKr
iGPhQAhWPhRpCuKfpv67DnEuVStfFGHhJ063u4bchOW8P+q19FkUHoZKhVxxOxUmwe5OR+20To/Q
jfKPyBtO/5mbzilwEj2lofc7OXhXTROJF4AX32M9G7WV9KBO/0d3sLfzY1hNfpzcM4nhUN8XLux1
McJjYfEDmmsyoNbp7nx7SYhsCi7jsyMqskPajsixEnBNQ9T0sr+Vjv0GFMtbj4ivqhasUQEzS+AV
iK4smrjAt2Kq8z1/bm9EydZjsMHTYWEJ8sNq+x63CUOxXxxm8LT7itQzVHfzwjaM++m6rj9W3Vq5
o7IZQIRMDw2W/TjwzpIEQn0QXkjJbF1Ke8lOF66qK6CQeuyJAW2rnK4n/IrgYffAyIW94UqUEi99
14smcf4jtsWuQzJnJODJhdMywSWbxWCG9eBfKNQmZqdqd4/rqgjcpffCW8KAb5yq9MzkC4KEmSBn
MgV18XAbxXtK300DYH+Z5Ct/GUfw0/sYTssS4GKOIHS1YSTcDdJS/VM03AHQWQhOuUYifQz5WyTY
RYRbOVhe/6goSvuztuaYB4hYWuOHWqLZ7ii0Stcs/+5wO7T2OPEK0ZKsEDbE4rf2wrEfV/WH6BcB
+1CrNySdH+qhAi1xtlWOajRKTifSN74VwdfQtFW3FKuwoWrXfs/Gu1lpDr1/IrhafJ+i2e49qBiY
srZw0BUkqHqZAZl8w9/wrNMv8qKj21JyjQdgQUytxmGXn641M3NicC3aQETyVMN60g8ztRWq3diB
OMMR1tVt33GBqzEkHFoOQ8EUH0+/Wf7NLcYRit1fZ3pu0XkYF+QsLgDJ2uOZenSoydiTxUlqsO/A
izxPTsdEu5x9imW/XzsWwEurMnNDDtpBLytH7wyiJNJe3ZZ5FfFADGkSvIqSIyWdu0hCGr4b6hup
EgwZYL21M2GakIiHVSWCxQaOltu4QFGcDwmbCEfQrv7XB2fQY8Jjp0BhWnPRBvEvWPS9QxtQuo0l
N8kDqAo++pB+xILO21a8wUVLToMc3zrC4JvNOwFOkvkmFS5K81TIuW0yysn5uFeWZB5FOzG0v7G2
JqEMXMKDpMtIUQHbh9YGPaynUnCJQyqX6Q+P5pQszAEf7a+JI6OP5WAVPeQFDL/zvSr1h8A4utBo
2JCrngFREndZ6vlxS3fNfK4P1MPyIsk8IHm3eX+6iBoLE/d6qutKdLc7NiJfpZsYYOI/TlSH+gh9
iJTwZqYiECDh8dQpKELF0o0bee7XLkZ0lRzT8qDGmKh+GQeiGPFXzVDmoywl98WFeDQjhrPDCp9E
Frc+klIMB4FeVqBYvKtIdbrT3iWW6IihKHgJfEj0NvSyrtZnIHQR4VdFd+OE4BnbJG5zsD5gNRh8
sagYyERf59sWNfB2dGYMPuvlI52ZdQk7Z5baHLb/OnNWSWcZ3UyFRYNTjm8u9tUv+/LKfVDGgrjq
qmjH/4VCCQTFJT0XB7CbKUFC51Ww5wV52rfXYMBd4gf2Dtfm1Fgf/obeziH1jE9nBhFQJp/2AyQ0
Hr6Ev8VrLbm8oXR/GV6mi5gszWDgpZz1xCoqJPT90gcrrZGzP+q/k7cbAUac2K7tUxkbKlU7kbIy
VdsrUmJQyp9AeSzgOm/h88LuoLCFKvAWj//I7NjQo1FmZ1nrr5IaPVMFQpSnSMjUKcS21NCFpi2H
VmhyYjWey5kPGETz3+xyAhQmpyEmQ6q9lDtvM+yo3C4hUsQVk/YrBN4Xcxc6AlY+Jf0DdLr1Dmyd
xklIIWk9xnlOf2+UPZmK2nSXfwdyNUlTyZhS+86nRsvybUYUlHJGEtQFamw35zXPT3eN3HUNG3mp
udwQY7NI7COmSJveKFnYURweRWENWb6rgqmNiXGoFkYQMWT5pfeS9f4LdcwwoI/sjtBF2Xs9/pfx
b3aJBELXuWG+7EFNj2oaV8fqZkUTDpZzLTGQaOTY9Ss7Y0DwP8t/PYcFZTJ/R8BylMTVJblQ2pTM
uUabHody2xWbgVBe7b4RxCL33yc8ePC6biz3rrPKUc4rqMhQQMYRc6AIlHP12u0V/uA32HThUmes
q/RYBHaisIVGajD+dXPpoht0QJ23ISvHo/LcfnzbhaQ7cdh1xgAaikOrf1YwcoeYVlfaXUjfLa5F
wjmi3zTDwVKtbxSAqemJ2coOIeeE4QHLJHSz5uNg1+EOZbjfKoe1huUFqtyYoUAAiZEyemk1TK0N
Ch4Vd27O+/I1sKk/A2iq8H7246JijLMD1+jpuvy2WuWttWkO4kujT4dZd7FL1PYg79Y2Ph/cseb4
IsRw/ErGAaFD+tXEosNdfphTVEl42kZFPVG1CuQ1/dFcgHkV+/Db2VXUnxzmk61rfAraiwSEdkAh
1ENpvCvNVppz9QKpi6LGDRUfweCoajxEilH5qmqNgoN2/HIR/IkmHFQgtf2OAYRm+BTh8rdfQpVz
gbk4Oa7EvzBQVNde13xVzrVP4bMbZZYbAkOaF6cTZmXlGJkWT1kbrXzcGyhC9CZ/MxkNYMemJpQm
IF4KUmN9I7NxepAPZuymrfu1j2zPJJnBGpFMeUktF8LLq2ncLnQ71WaaVqucPTLlHlpXA86Bkiyq
7uSmGJPT/MZw8c0guxcibig3b3XhZsptuk9aHFEj7PFOJG2B6JY/tv0RUG++7Pz+y8CdpcMfzBEa
wLJZFj8bJF9CtGkCa0o7nk506R/c8ecky0fXj0yWv8CzWNNdXxPbPhYDwfzCZfB/ViJJob34fHYy
WMv2nnmroIQF7en7ratS9oXqBJSmIXxWzNkybt0zwGP/lVJ0jX3Jpuq12/mRG7LiwDGes9c/HYiY
jmBNUID5r48W8TILiZQpRgxMSyewhXTaN+qFd8bVkbRflGgw5kA3c94biqGRYPH23TzBSWGmbD/8
t//SDURu24mY+k7drhmMNGM/xy7kNbhtdL+CanDkJjeshz3sZo7kBSpIvqUWm7llq31Q3Y2TEbem
syBpWCHqkdD0HDH5kb5eVn2H3kDb7++YN/bIs+0CmNqqJsURJpB4l2y5DpOK6+mfLFAFb0SXoxGg
8RC7gZ7HhG9Uc0DkzSIe2vNoTZh25HR0dIuvj1O2YN2u5Vt745V6GUYSDGDutkIf2mk7hQ+GHBTv
9M0YRrgtrnyVdLyCnuWqYQ4KsKq3eEQTtevKh+ULnGFFVhEwzNBc8Ms57xYVDMnCkcFsRERWA+sj
WYdOsKxsjRqM3HYdaWqGvlP+N/6D2CVoAupES4jI0AUH/nzKs7JAbsHOiRU3CxS+a3FQThfB5l7x
8YDNeIgUU2NI9PheQbdWvn+3ujZ0koK9pR4g9PgdqrVqAztgu9jSoW7JFtV9D3Y/ukmv+/p/GO2P
PRugAvKOyoc25L86i5iom4PeCVm5mkYIXhI/H3i2mF4+GLVLtf0BLA85ry+79XxIZTLNEfNEctTq
1mlvStG5PaA69Gyf8xKLHvWz58wkiH7RX89y22kbjlQEhvL3g2vXLE/g6p7h9OaADydqThvIVoVg
Ukd5mRhM1kpG+4M3acf54AX/ABGOC+MoA/053X9yvVKlRYxXGgpyLAlyX4BEnBd30LuEcRb0iTso
oTFiba15STDExaKmSTH4EV/pBfAmqtpwY9M/Hs1GoMZdzqAu81SqbGnsbfQz814N88mbrunaBb9k
g9Iovj4vrpZJ8rQgsOtjlMmrIRfSYBFh1YShQon4ZMen2r8Xotd/5td1pM3sxdAIDiHuiKXa50o0
iqBWS0zIvg2mFN9KSwaF05h77n4Du4j9LunalDXEvnoqaVDBOs/MBLLlE37IRB/IlSeTluvdPgVk
FjJI+frP5T3CKt6a5r+5Kyj2nNY3n1ggsU1LQUpDqu/L2zDoJJa8rgjKgaLTauNHgoN2N5oTAdie
P52qbb1+tyrvS8ORiOZrkCwwweSux2dsSzSFE1gLJ6AZxAA13jh7P7ixMD51ZEumb8dH5G+j7qN9
XPlVRPSYDYrdezulKCNRrWksbybE2v3ijhcjAWPi/WOqp1n8wKtGvAfpBrT1iZCVbnDVOIvXTgf+
O4SS397YoxFYVikxGTEZIqL/4TYhISKUK3GwB4tz09IGKn+Mg+noveqwZfTi7qt2sz9cRnbc8sPL
5Me9vG4n+bpeHGrYWXW+uOKRjEdqL1igpTbfkrUN5mv13/EYpMmk9hsgJwV4LyxYFghCthMVV7G2
lNwAHcAFnP0nBpsKvTkZGTiLtwZw64PsbYVMPMfCdhhOUX3AKNjGzT0ZOrZGF6H3XM9VdC+9eVAr
bpaVA/47JikkpjdVOgXfOM/+YPseDfFL4jV0AGQrFsFEsZIylQLyJyLvP87OLiktYEx5YOyObNZw
blxUAeSAeXaI+YC83ZeQmG19PAm0O/vmnQDjdAyGak9j2JaKyX0HrzDkL86h39xs0h3GNIHAM9LX
5c7OdzA4RGW7v8FH5M9wzIZuEXiomHvq4lqZAZHZfDnC0U0FUkXnYk0QB6rlH8ea7QOkw051Kie/
MpnnIhUyBGc5HLmUfB0lWANssBa8XbBAHRvcKFJ8KMl62JKXJaLq1XSMcmpx4aK2gtPSUqRQ5ruq
ganC8ueX1M8VmU0WiRWedUKx2wMGVjcvCWdubeAa89E9cNHjCe2+nI72smcwfkIgDaXzT4DdXs4L
+BU2i5ZLOam8khGGnurZ0NXi652nOODdTm+i46sFtJoOWY7RC9qN1JE2UJdCxaP062F/n/Xy+DJU
n/0FalkEKOLGubJhSPw7pk211qIm33ymLNs7SjHwnaeruvRcoS7RhFetMsdNWfx1F2w+o9AEWhWE
HQ4vIZvrc+/+aBS6x67F9aEpeJlCL3QTrAkg+87z7FLpTLy5hybZWV8qVC6pzI/BgJ77tpicG2K+
KRLFUdvqixYjjLoXBukF4uNn4f10BfmTIvdFSp+aEmxsq2JRBOEUbmZaQKu5rWSgDlA47q8geewk
O++rwLqPg60SFmqERepGPXPVGdo3T7SOJHEVy4MJW/sm70TI7y0feXJOgMfdHtfca+AF7YhhambT
S1l3RyKVXv7X8QjDqYUnohxfwtHiMWJLxaRZ1v7EoqMSVxaTX8DU5YqX5zHftuyZ+LsFg7Ss53ZZ
vSwqNsHaGwn2ZaWI6er1I0edH2LxvUpIsHkRPMW0zsoWomAIGoRayMpiICcZfUr2b6Gp58s4xJ1a
VGQDOhUyxycbmvo/oWJJS10sN/d1JnuhvGaaVrqxY90xsif8tRh6M1mTTFnSo0Cr+LXJFhVgVELS
zv3EGBhmP+FNrt5khJapdxCn9hNCIxb2aJyPxW3efTZoLd9AaWT0hwSEyBAeVgKi7EGk/h9E6hfv
Y6gL4fgocvsb1tV55W+dl8F5iuNJVlY5iBFwv5pHHWWhOucMYeUMyhCBwN8qk7pd+t5gqyXxeSbt
/VUzne3tgVPN9m8Q8GTFI84JdRydCNUjgfOicVuDRRFwk/5IV6Bod/J7IfA+oTw8zFEx75kW7DrC
nUr95Bmy5SpdfxL414w0cO16R/3t2w89rLXW6dRZQ4sbnNCU+uSvWrWzf3cQN9Yh4cJm5adFg47l
/TCuCCGHy1lYvi6/DnhlguQvR/uVMf5LDghWaNb5WRQPtFXuxh+eWpSyU5/TN4CB5VPkg//VbG1a
k8UnKym/KyVK7ea+G2iBPm4GieqVasRuDCdZo+OilV/HAULO9sSvCILt1lry9rKMMAx4dYRUWuHS
98OBioOQQ9q6pCibJc3xB0LLYKMkD3pEPgim0FBZLWuWxkBW71GC/ekJPWmfrF5X4N/BPM7JOV+k
QH8KcBhN4d9MU/FbzXFc0d8umWSnnLaKIDa95idmKO0U4JbDxuGj1dWMa0zF4Vtp+8tzizH3RnsF
vBukInD0eDDzmubvdFs+BCTfFHTAvdLZGVdGk22zlVAa7FcyS6qtSafEoDbh7Ri55GuiHrZgDqB8
AvLwuc0srvNErBpWfdYNF6O1MUvD+DbMgkLcRnthdySXfirQx2l6EED/dgIeT2bxoGF50yZloHt2
0suaEidYS1q4nQEYCCykFxrx2tD3H0yMnHEQ6ewEojhcZp5Ei/uqAHjO9MnbLHtf7e12AeUlcpBB
O3L8Pc/GRVtxBYWVkUJW7T47nwCIz7cLT7n4wyWQw//UXW4IFgzv77cS4eDnQh8WD68vFd3o9844
+efLjR2KX8c7NNSd04uwHrG9nrSSUPh5ecJg39DhEjGNLexHPuowDSl+jfC0od/R+WVk+iRpsW+l
hu5/SDZFaYQ58oMM7KhN/Bz2uTeGfdARXmsX8Dwpy1NZog2vJ+GC7kQhxFwGN8HxNQRKtvSgLPWV
7KNCiS4Kzep8Ay3Va8j4tFzHt7vvK0WT5xAF8/b8QnJDPFuVcH6CE4XuMnXvEDHQr8ER+KrcMacx
oioWZvmIJmcAl/CA+bce3fLwC+lHvW0wMcOzFb/ghcQaspfBS0ZeYS7HngcF2N6t80wJLOLFm7IV
BABTV6Smj5WuDE2/n6RXzTwSAyqHTXFztRgW/Ns98iMuNS/0+2KujhKMc45ZiFfq2QkJwJic2SXX
GTDmIs0W0G2gv9yRsU3zUPRMRo4dFNMLsO4OPTag1Mx9rBhy9qskBtEQkapgb74ofeiqMyDjCkug
PREzUKCuM4fJDLsQZ+0HOgossXlOFrdntYEuTCMTox+wNtJMmHtp1rsN4zIi3+YBdiccPLAtTARx
Ad919ZfuMV1gwJ24kx4ApbUul1JZpB3SO+MO4uip+PEkUGQs3nhj/KpUq0gAinvzkwTM+ouOeGTU
At/sGNlhDJruaN8irKxqBxpgt3MkpMLvyafPC+OgAVvcEgZ3zC4vlH7C1vHXO8tZ0gYK05A3tib/
ECgokZFOfROwMCKn0X6VHyhvBFUGgPF4O0VW0LDOvDnS77J/h+789vCRRQmHSGKIHeuo6hcOXKJc
awYcxFazTrSDmds7fHTI5xUS481GcziFNeErIbhK5EihsDOw8SMrgpMlDOS7SjmJuDb5QfXNey9Q
hzSbnZ/Faeywpiqj6iEvUtjgHSn4/M5L2k892GrKwEzQTo/olK8yZRkn4cntzgSpiy5/QAIx/1ec
FwfCweYwEyiaOOonDZJhl0oYAWdJLZsYqsoWnjPunrMDlSernRVlSKh1/ePti+eEeTSS4Eh3NYdx
NmPwFZF8rk1mPABSjoUBHAnKtrIY2A2hb0yVQIyr9ZDphO7n1KDc/DiOQhjjZMTf3PKazZkjZZcv
b07GDkqW8VcwEp4f8cS+COoI2Oh3MsmLtYOX4K4G2qifKLh4r1BWCtSQDNkIztj5u/9D9tZO9eMt
BJJsdD3DsB/gOd98lnRhPbvPEqLl+AN/Cr2RRktb1PlnpdfvHF3+T7F/RuqVGe793cx0g4bPEazx
i9VsNScJRGw2MKmowOR2aM1oIsZF3pJtyZ147wEhpMuXcU7RGH3+DBKyyNV+0RYzxIJuGB3Zl1Wq
ofpXfQzb7xCmh/ZnD+6Gd4RCTwFZtlaCTppQNuQwWjsIE/n9/wqF4kOIz4Hs223mg7N6uvu8DCQ7
U8U6WDeBf8CP+Pz/h33t/uz/PVpmmHHfPmeFrGBroShizkSXOyZsN5VDNqyqP/NwviQmVXMI+Znr
aBigbwffGHF+eMzAzac2X7/39VZec0HBVa7eLAT7+sDpHKj91GD2DjLEckScRTxRa28ecH2DS4tx
pplE7uG22bQIwXGmW0xFzT6BTJH91FDAQkaTXvU8OkaIl1JF95C3D140NY60ix5tBDy8zho+/nq8
xOeoklx5qbhKi8KS6SqeVL2n2+dNsbsgaVd7M7leEnF9OsSzIOy2Sl+lPAzLm+F/gLkyOoujd2h3
r/F7C1dWizdKH8qBPREQaXkGUO/1kYyvJutA266i0dv60gYKhushcm+flHM5n0RLuSQbgaQntAjb
D0CvTkAUkuwcLbogJRiFJvErXBKlosqkQg0rncKrYiFBLCuD32u19Zg2BZDhBHWf4LC0fRCy72RG
6JrlsvBP4H2ett3Qhf12K2PmcN3+7HcLOWhWG0fZlD3kw1zmyDiCGjKAe9AJHQPf72gSONstICDf
AS3VfY3hTqXtVR9mVp9Fq/ZIWg+gr6FnWDw6LH0JeHAzKK1OsElhsqi8nf6gDwxvLNxtqPkjyFoA
MA7O9GtQWQutcC0aH9szNX6lPMHzt4Pq51WiCQD5a1503pxSM+ALLQio5uRV0hZt8VaR+0AWB8MG
QcnXKrrPDtULgFxC6cxFAKERbQ7PJzBTRzLpP9cp+cgSSxqEJ7lSEtG34Ar4voENRr4YgJO6nPsh
7z055oR0Cedw4tRrOoA9SvWbf2aDfLTAXhdYTYkJZ99TFDdxr4HvMA7DHLFHqMaSZzSh3BO2XFEs
8Dpvujy/8sxDje24AlNu4EiJ5Y8abOpSe/F5oGB6I3NmR07Ftw4ByL5Tugpn6qxhBxGsVkhR24w2
qpaTakdljFIhUDTUw/xGpANtTvJBhKi8jj6YqMNpjjMkp0a3RYQ8sn146Hh552YKu+ZhLCCCzdP5
pN69ojhj1cnBnPQ6KH3TE93eMshBEELIxvo8uagn3nObAPixNoRojNhf8hKLOPeW8kDOUtz3MKjP
sEOK15mBSfqwsD/cYFTM16xskPLohH5KxS7ozdrNXmmTAgn303RR/qKVB5+0C2l6SJv/upcRwh2l
1PoEQe3oJ68u32eO3phM7AppWHhTHp2lKrcL4hkXOroAPvyI26hHgV/jl8dzcg5wwRtCen3Bvegi
I/jQW/TdAA4p7Ue2CrVvLzoaABVI6Ik06VUvwlOfQ1logiU4Sy1udfgW/V7BEtHQOT8YPoY7kvPF
1hWCn/m28tDOJtWmkrviy3LhNIwYMPapuWL+rX7A1xr2W/NUti3xCdMhUZHE7sCHDK2QFko827Lo
igr6F7Id40zomt3zE57hy1bSJaHK+4VFQLWrpqjanV7rDxJoJBtKZQu06bQAbtQr30k4wjKiPK5q
CwmPMHyMcJ2iWh16opD2AjmQI0W+V91W5hMPnxBaEjTzM2i/OZoySCKuOmZwXNFcCmXdBUO5oM4b
n6IgTw/I//UrwlqwprFzubTEjmywfA4K81iWDm3pNjqLLIBt+P0LeaOCUIffUxtaOoEAcpLejqKZ
61tCsjZ0Mqkn4raJ+hJSwVHlJjv3eDxEUziNDkGhLao5H0LvC5gPOn4ks1PJ61zAKMAPWk7xDvXz
3gRofGHQb0X41+PkYTymIj0XYF5+PIu8CltKPEYSgtc1QAuU1JKFfoxqLu3xYbR163f0ZgZYhILu
BEsr88Sfmi6isL37gxcawLhimMoA0Chw2k38CrmnAtgfM0G9NchwN3ZuX4R0CI8pve6tsgBcaDAy
63CUwA3aTr7zgbE3guqS2yCWoA2XQHjExu9tOFe2GMLnw60MXIw1L0I1vlGtMXRKShuS+DVDObQj
KBhmHdi39nPE3oIoomnx7HQF7Cu4rDVG9V+tnlQCHnB1gKGJWsXKOkRuhD+stW4LYpytXhLXXCoe
ZHABxtwmKpBP852j6Vjp+ddCT3LbP509lJeknbhN3m300KCjfK5mEiZRGlDn5FmLoCxU4PP1yf5X
P9FKs34Uygc1aWFoho8XtV1AhMdaryINokYYVJI33bmRqO+9awkcRYGHEd7dcGP8sDX5OprfT0PI
Wgo1sDAR+DaxFl8sJXooC2NMnXNMa/FDF0CC7TtbIlyDkgzZMPh0fnXtFhCco+LwuTPbIdSy3mAH
gqG/ZpjbVuZ9yxdpd5MgTIcDO7vstGWUwzy+hXSkKFkQv7e3iLN7HXi2+WufAxq3Nu2i+2BT+Ifo
J2sVYBrYd9flEyhix4UfHEyGB/qiXFv5updDoJ+21EG1kUqci1dPJ1eM0BQKclxUSpEFtEsbmZEJ
MySYoaJKgua0YlJ+jgM7HB9uQy5RWTE0TVLiWl3ju1JZteCdrnJzkXxT9zN01u4hnQLGOKr1aHfs
b99VBsBk50oe3WnZxt612JD0TL/RSPSh42l6/1k0aLObjQLNXsL/WKjFh+y8B8DOhQ62mKArevht
zaGaw+W07HYs5dnA0EDT57L1iYioFOqmbkIK6BA3WsNzUlyRcMJ6l18Jb8EOTeziMgQAGbN5gMst
l+N123FC/wS7YRst8uEePPRoVvjSelxCdHPCUdl/3KjOPzzcl1h73pShfvTq9rN/EXz8DQUTdtyQ
I+ns2Z03d8OzBWv/4kzsijGKvWrca74eGrB5kGbUP2pFphgEAlUre54nI6LOocTzpZLeq2dUjBjC
gb+N3f5cmjN1NB8wS7iY8tIi6b4Z6VoVGdMoNc6A8Y11dkh5/tT7iX35vckJ6zeWWHYZ6NOy9YQe
BH+MG6vKsVgNusV23d7GKXPMTwInLoGiVadBP7ybenEIUyX5Z/UxmfR2IDn/vIJVHBeZtYEcRoEg
X6rYQCjnWYYYhn4GAdZWgzSCfSLWZHNANr1BEzO/Q7ItAZZWUbxiO5PtYlQBa4pTUFzGh4ZLjEmp
YLQ4bWDudR7DlRNhuVSR+8dd1TfHQYGPx7sjDWSGKpNOT5xPiw8DxcLn8UmR8a31/T3VoLEiUcwZ
X3LEEDKrQOEhf2gO5rpn0AsBGqRdamhW58qpgIWkwwcLjjdv//mrVwrb52jphe6Jlu1dA3UF1jvU
mONbL4NOvPlW0ngWs6UTQ9txHChpFLwERHMDbF8faxCwE//nlydsXXIDlh77OY+KNfC/x2k1Ftnp
ovi8Cl1jpg6WYlbmdMtk2BppWD5EffSqx/lWqlp2kpuNzB2gE+Zph4yt5tFfhG8qjA/p0w2DqPUx
YLZH7ApUl2S9MiwW37MqJRhj6bfloJ/dM5mszLlT9iItzeJP1OItiJVbf9puK/mFxjDvCird8/sH
AKArOI+tkBm2Muf16LKyJqxv71nTm0hgyMgwOFrhBh244NxxYwLj7Xb1Y5ahIbuvZVbtvTxozL74
Rd1p0se8ph+wO29Y5zLLeTW3CV3RfbJGgWi4xpRzUBpdehYclyQmNAP4ePDishbMZbsjFDJ2EWi8
0e66N1JjiZs+At8LWo6wVYOM7q3M4O0DNKzRlCXcet/chnco5QqTQd0vCvEPWNAdaXROzwZJb1ol
V/otGOTrEQfTtPm9P6ZYqVtj3byAupLAMasf89uOAHVS+1trmuDy5/plTo6FsFKZNlYcZ0C+1AXo
YTQ8xupPmUWEXUfh16kifptwGHwUp2XNMzITeMbAnUDPVMa6B92sHoqQZEv9p2P1t1TVR+dtdCTs
HcFbeHLKnFW7pcvTsbYlnxXJxF9I/YQ6KeDL+2h8FDSrvIQ9LwMAn11fyxJKni0VD2Y8Qpijzrlc
EFL2DO+bdlHgkDZcjdCEMtMaX+kfhA84FEzLqHQPPyZ/u+hmQ6Sh2WImCnBXi2SZFheuHTrV/KMw
p6TZNJP+F5He6XOYcgeNtdpS10MATd5xZPdtzRjskOrgqmtKsVyZ9L9rIxsP3vMx6I8IOkZg7BC1
8U+rSI6/BRsEvTTX1JcbSW3m2CK7cTIcFmsIsza3UOgERcjYj9q7jdT5sVB993JJb424ttreO7h5
mNON3i3hoOa4S8ZkSOkfvGBqbT5BWbsKpm/47X258gbJbxPyPUrcAo2TICtm/9m4xng7mI1G6qK8
yo7gyWFbuGG1UBgaM9Y3LHyGPT/G/bJX6vvK/Co9R/AT18+dHZNFQDR30ZFnUaBQhmB3HH78EMKf
PmhD+JKzVin5+EamvbLCTdEsnZDRz1zXpvN0PxJxbLReO1fvCl50OiUMfIOJYycJHHyyMaQHq0Lo
q38gY1ZZkFXzpcgL4ZeRQY3ds8TWA98q/w52s1SVxc8hUvYfX9XME9HCRoWt1in52+IJ0HiWRnLr
Wil8RhysVuykMlm1Vr16vRT99VjggW714Uy1O9c9pWB3hKasVJKF8XuxmJUzGPqVHrcwWstX7faW
RvzEcg6s77aTsNbRxPCyBEhlkt/yWGEMTROQEnc/3g6UM6NcKYzZHhdgZDVJRf0ONQhSDYYmYyEa
niDgRYYkQUpnu3VasdRS7EsKuiBTcHf+cRbCsLdYSi6J+9vy6NETkIDZgjbQCDRSOTv/RMfUdDGK
f8P6sqYvNlX24aFEVe/TuXyT5GIWdqkgUDww1HBQW4bRMY9XAeafAzNrQPBIEcGWgIc/b1wAQPi2
fUKxLnezRoNih8Pji2hiwwg7R2xnkIm90CVGk2HdvhwI6TIU9V0pi3HwKRFStcdeDGzQNegvSxr6
4XBOVpWIbWYH5SolaPX/ZV0j8ySxk2d7TTI4ViF5D86l1w7OxCJmIT/xGnXsTqR3YQLHXbmSn341
whtOdeMzjodss2pJdOp58ccJ/vS+ucNbotcWP4DiasUDUGtB0LP6JRCofRGfcVemJ8kLC2C6UKUb
wlHK4SwP0mEEzkJA1yUScaZ99BpUSvaeSsZHoQk8OQvimJT2z6CXLGQ5K1Xfe9ymzATTWlti7rUw
n8JIWzSPM4tNfHMgvBOm/3NqZamRGE2FTHJJp5N796QEOaDjTGIT+tpUitizNXdn7s7l0ZStgD0U
e0lanYPLjigKjGdocQapXi0fWoCuCx4RO1rmBlnzS8FZeCi0/4OSwUv6tPCKR/UjNePRaghgFWoV
GaILeI4zuK29f3okOPBvR0dicCkXIHxDHWJWawAqohki5+v31bbXgAPlgCFEjXX47rvOGx9wONb3
oA4RsRB56g+cfQyPU3NbQdxxF0xzqNq86zdMvzm3RshD3UpFLtafRcC22udjxJ2O+rxEAUUAQ+AL
adhl2vMVgvAH76VbD7fMfW6b+K2f2JCK+OY9dmry6clRf49XSeE/nRResO7W4IV0N1W+kYOT3Wl+
xhgm+5rSfKORkl+TN8vyBDG0wWtnVw7J6GzHCqjcY3DjJ1+Mmw98Kp8iSkQKB4HEEysYLFLHv9wg
FeKF9v5C62iJx2MtvFpIe4FgdXGTi4Nr6WEl97rtWXdadbvgbggoGMgDYSgPohHLeKqVZzYHL4kJ
CwjmOK1al1p99m9LuM6TkEQnN4xdRkXBf1u2FR2TZJ15WRiX+gkvpWtqJPtMvqX4qvBnaMD5+Pdh
GDWzhApKwwNUovoEh2cDtFM4+dCeA1VRpubcfBNNuA+cTsLToFrKCM6knN0Bedu6eqv43Cxflni9
pSKHJxx2bJ2rDRiBk2MwxQlUzCJ/T1I6BLJ+afTxjVJzeIV7yEtaLMdM0ODNKGLu5TZe9iuJVrN0
sOctTMfL/q2MPOdlafuLcIAypI7IUOHdykfVZqUHEWehfvokFId3trlydr1RWGDqPtYQdgOYgATL
SZFSFAt8gC0sOYSeShd11yu5caKZGH/MHQR4C2yFP3RBpJjeh7DuBHqxydZykG22t3c708dc/dIg
Y91loklkJc9IrvYPNgq9NXMKTt2jLA1ZCQT2qLXoe/ID44qAh5sibLsaBSo64CjiKkTGLiBehBgQ
ZpE6158eY5ClYv0rNhdrvaXZVtB+YcagSfwRbnKfm0IsghiJdAI8p4Hod1U3yazkNcNBnnByvjei
pRhicJe1uHTakglOwnRt8XDwbIiT3tcBXxbkmv6battsEHG4zWENbpQMIKI5xdTOqPls60inUaaL
en4qRvco/yNGu0XKC3tmFE6yVv/0hzgsG7Keq/ft8EWwzWeU2pIwoC/k8Fo2ofU8KjXofqZQ/kY3
VI0dmDRy8Vtf1GSn7wBzgk1/tcrZBLp0iv9PtrgM6A1pGnWZx2eLgzsjGh6DFqZzoTQEpPJ+quxD
e35fl+G3of0DK0HJpEnxyQpuZyI+QSckBeUWLVA3xIGwPJfvu5suSwyE7ySkX0QR5D13n5xZcBJj
9mPfuQNqL+/qggQV52bQoz98FhGTr+6aVsJWsXpYHeWhSonzUi1AWpUYHAJd7HFCy/GjcfJjGSlR
m83EpqevTu4XqzjahyyNT7EOicXzWOuhMN6MzysFInnxiyNzaex9R/0yO+d2e8gvuR+KYZZNJDrK
OCBEUQlC9z/PHSgEfM66ZpkFlVqqAtvGmIPbpsET3G2aJjGsgxzkaZwdl7oAyRiIf8BDab2sISz+
Qt4Sdz0gi2b481EZcohlb6uA+r0/kAl+c+yEQty1QWNHt7ZXNsBYhkSKeadDnuwkxjUu4puEdxn4
ViVZaTzsOB4fxbRDWyWAjlZdakhN/LWnDxqXWkNBXzdz6oa2b8udsLU+6IDmpUKtjvnBKMUtfbbm
EYtl+WhG+Bbdaow6IgmcGutMxZiLpDBGxPTkg8U9HSVNVKlqiHUDJ3HUehgj1DBh4XnXixrZfTck
8qnYPU/BV1xIM1nuuQCVghJ7Z7QcbNKOfykok4NvJEsIPE6nrJdLk7Kb0LQwpjZfIdWtv7pQWkzu
Okcb70B1cGVktEGy+O4gasy4mEJe+d54CTzkpimj/qS1UsXpNglvr9xVZgcOcKc24Nxa3B+7LKvo
ZeUQhLr7rrdGGxvJlVBzJgnJDd2Q4DQjtWftuKTO7lEQEnszkf3IvAOMi49E2wCUbUG4Bz18vwve
l4HdlyQsIjY+FF5wtaZs99PG6qZ1DCIFAZHZ3nxySc3Cxc5VWp23uC+WSA8YXp1GqHiOG+IxQ9ct
ucKeBMZRKh3UF+GwfTx//5XKgBPoI3/l/jnOjUwSytKPzfAndzShMI56eETBaGeTUFvMdqNR4tbR
G5Y3/CmIU6F/aPH0fRQHA3W/OVbzVflpIRGmzfkoiM45i0L0zR6jOaQAkXV2VHCQg3qyX1X2EvjK
4QvgwSeIoVDkCNdX0OkkQzxtub4sZdohm14j1eHFZ2a0eGq7kA0Xs5Vs43KNQPThnCnZGtVglbZ3
6mX77gG5MC0R8ZpKo12ecca+M0ix32QSBDR2MPADz6DMGPA4zrDej4R3fQgrxabtn3Bkt8BVpqWt
0S3ArQtHX2WuocyP6JejK7pbgEsIpoc0wH5AwiCJazZkI6yQvy+yndpSBQ3RpRPE5bMNLkuVSmmG
lRRxEpil30VZXascpdz2/agmiLjBBrbU9uQnDddjrXGxZ80in408xwSmnkGZu25fAVSPPSgeq5JP
4h88LX+ySovQTOEXl9Orpntf1I8gSLETus5iEy+KtkEM3GDy/dcGtJwvM1Ivf3psL1BQOxSHCaF/
VqAduJtap/LgjueS8BtCBeIAuvCGN+3u/zRVLnnppuV5whU/WjvgpB02o22+A9D1UUjswzlMQAqu
g6lCBulhZI+eQ5NRarSTfHg3FJRn1atxUK3D5xZtgn87nlxbRKHnlXDEjkytHzu0IPOJvZ+KzPC8
zJRw75gGr4wjZYOfWl5jXAcWDGtgfdq5V778FpxrAwVLtGFFO23zYIQNQ5BxglyF5BRDBog5DwMw
XoyS6ZEeECEK209a2w84Vl98/6mEOjErLJh3L9kcdAATgGPzrLGRU39jE7hkJy5yX04k6gTqv/35
J8NhIPNn3xQvkZtoLZ+Z1tYJevGN/meNCKt2B8JppIH0NVyaEDF0jiZvJg80C1U+5NlcuyeQfbmz
wiftFi18at68wQ+r4QQL3KmsiW1K3Kx3dEpSP+oJeoWgfv6TpzoGJgTYlyvfDnOF+yYdyDF095PP
7mrXnqRdS9XX/DWWoubs2uG6Olbc1AnxDKWs7TJtrbRcea5QadzeB6kBK9ImfgE0CBUMdiXZCxgk
ydfF/1SP1JClRpy0+aIZIqQDjpVV3Nmezl9zC4QIpuckB9duBelM2h4SaVm77QCS76IK3KXx49yO
2HzP4EFpGu57xuHdMoaSmjaBwIMYXqsHPtXOihfl6k7Be/l7Br592wMol/htrwALc0NpEQ2mrfuL
baIsiZbEQRPBsrMfqJEVDpd4b4u/WbYKOj21CXxIvUPXC3o5sGD3Qn+q5R1/EvvwhRF7wDaB1fg4
6Qc2TIDatE2yExQo26112Y+IXGoynyefcjN06UqDAXJx6BW2A/UltZPe1B160Lb7N5K8aqldlnRG
VSiZJtXTq1Y20lwkH0ZmMPStXsPjvhLlE1wQgX/vKR15NI3g/Nk4IlAH1JeuqLgE6ky3Cy+8Smxr
bg92QmmCOFmjfiuvqidLIzUH0xusPYAH4V8NYBe19krrw/gX7y5ug1rPYGRqevfNOBLbTK1O3B1T
b29UkTnuLkuOXcTdA6B14QZhboF1k125S9MR463eO5IqKBRWgeiuV10RGhqMXDkyK03UJda2kBNw
Ho7rbtPe7O+Rum3M4AOXzkeX22fA+SlzNYtdK61DAc4u+gjNDAXvpgBcxAkopydnWmnquCwvjJ2y
Gz2wB5+NSdCprbHN8d8yjvfCYmeB38GszN+BlCvJPV/gz2mDoeibwDSjrRWgTrq5c2ZPlwrK/f1A
lYcGql1lE7ZigGs09/uohxZL69WHZmqchE8RKuPeAVzvPHN22DeicsVCXjmLDMJb6X9C1hrW1FIX
G9v2iDOQRGIguwTIaAm9RGtyA9WOf7B2x4s8m9wUNfJIHhmKndRHLqWIpdwIvSpmDiOEsC4lzfVd
HNkeSW/LgnsfpMMUFBoyp70t1tqIQxmFywv1W7iugFcMad2/7vuWgrCcXBvISp8B/I54s1WP3L4c
I3k54FmAtai4RK4iSg4h5JoIOqqq+MberRGzBQzt2OgwoOeOtiYxKRKAkhCZ/K20v4y66as31M2N
o3qiBUdHffTV8ApdgiojrGZJLRullwdiiIhKw9jw1iyQiWVq5LAsEKIqm1m7D4J8GeImlDO1hX6p
58iAa8HRxXssos6XIJToecdLVmywMIaV7se+P6GChTj9K/jrgaF+yF9Ofz9xi3kAnuvNMaaVx1EI
OhY2i6K+QbFb0h8x7T68QreGn4Rryt9W3egXOHpUsCJAhGmW/m4OOEAe4Km6zZYWiMwj9OFrQvfL
BDq3ODbpsRjEx6x66CImPqC4Qx3CAN4NvYgMcGVqAUH39tIisS+/rKWIYSLnVDvrrWU5M2iWGZ+e
qmfqtCSWmQZjH3X3tiy6zNCdfQlbfS4boql0GgGMxZe4jHhnQilZCHHOl4Pv7PvX03D7aCskiiw3
mmEc8TqfDmFs7UZvoDCVvevLTwJd/hliP6s2Iff6aG33rS2OGUmM6xV/8Wu2OgGipldxAqs2seT1
carEgzGqrFikNRAHLsT1Mw8v+eKZGDI1HQerm6796P8YKHqzEN5lMPsgKrzTqNLEJffkiwkmEjfF
xT6I6aNzmQ1JNZsja9I32/6sJA4OajrKc4QlbRpOKaDGxQg9MwQW3/w7hZ7TAo2tPhP97h8hVudM
w3PbICVaJB/KSkIddCNruXfYvvb80Rzhevg2YmAdrTlegyxHbN+AGGrM7glxOXbo1+s1HtvYXLTS
cVGdiBHDD//84j/UQ16P8SB6b8qhA6slTCcd6AAkdR+sRKScEf6b6krceZZle6Crxn6nUknyR+kH
g0LU9W591Rl0fk+B7oNv4oVGymaP8xOe/52yYL/dPNOM3Bdqou5rna3ER8ydt1HGEp+fHxg+XS47
HkDnXWxWbOdfg1Vnxr2cvVLwkz/l81u/CkoPeuFeQOn+jGTU9WpLavPQEzxSs+9q0Uw1XrOjJfml
ZQNBFFmUOroT2pF55PbBV5z40opwJbJSqXYAjd5sa3Afd3W1F9pjIyUpZVL/fyqmtH+nwD8TA9Tl
1FghpiUOI3SZ5+1FQ7dBSr6lN8qHqKL8ybzSmlk0Q/6+gU0tugtrlk0ILXLXY6eEgdBfsppQgvY9
Ix/C82MSq0rbayG4O3haNniQrEcga4eOMbnltQwDVaSnZ0L6KekgtCe/OBhIplzN0UjnzQbkI0zL
ph6hhjqH5QJizuDRWrmDOYv+Ws7mimYK7rCjvAyIGZkDJv5zZXFhfj5xTzJJZirtK1Pv4z+Eadfu
Z60pfJ+XMTUUAF4o0fa6Z0OoXNeFE+lUMwFLqGoX3FbCAi7WvoHnHEn99bYvKxdNXKHHHh6+HPTl
DMwF2x9J21NKpnFZvjYpichBWowtB2ZavL0QJDCd4Ig2WYZL1HmtyHWscQV37pRwUY3MahP0gKK6
A/T+aZEU6dL0ovFCTihrceMs2ZZ/Z0GVI++4dfMNMdPjMKoenNQbfG/tlSD/0J2rdYlPUs/+RNeL
Mn7s/vfqn3uicqIO9LVTutZvr2Qegw3crsqifxekis3hXA82yl0lek8cm699VI+JvST+TIpE10vX
zXd7DPm+NjXJEBW28PQ7mbhq9vZvDdbOtZ5SCnWW33EMYAxRSlHT2i7qHv736TN8RC0LMDITfP4u
8f1N2LbqC8tArMv6QDdFdygNxHLRPGuq5tv4zuJ1FfY28/W1z8xBPaLImWcs3UszO2NL5/JirNq3
i9o4jZBDsykJoCCFSlPyX8TDZzDau2YAbftDzuN9S+btzNtssyiNTaRMe9Wexny37G/6aCJIahOg
+tExf+SOU3urOouyfuNZ4M13WktnDOuckTPcuBQgk04J1aOrtjN3DCL8IN+S+cW7jhWqWsdJv8wD
87U/7HPB+I4y/saxvJhgDxU6g4tEuraSOGEIGeeTX0sgEAWfU9wlkBLk21Kqt6U7ONv5PbENEa/9
l5lOvPURccjBdkM/tq1HXjAGmCWkPvEvzq4uOD/iLgQ7BFO1/cj538GwA1+c/s4XcClqnEatLbm1
RNwSqC/YyqT7+UXFt4W3IlNASvcvmf6XFpxrU9gjaKcc3AaFdELuU/sk9b4G6WdRYhIr6TiAWRT3
3hldNMFdGvTFzD9vqt2Xg0aoNwxw8wR+7n4kTv3lJSymZ+MyH00Wf2tlBrFlENg+ay3YlO+UPQXV
Lm6zTHjOYqmuhPUkX+Wd3Y2JShEkOhDFS2Tus5TxY5zHh1ALypRT046bj1RL/rOyngwgp/tKAg/N
L6fMEPOuaOZHIgE7gHNxy6HKZ0LtuB9P11cRTG0JQDm/P/GBBpxaQnF3hu8HA+gsW3CENLmd3p/p
kSO4XW6vfoWreINYYqJVHL38aP66vMoM2jeAUMPGDFWoy/xZDBSqQGJRDGlSUZCFHL6iNBHF8pRC
3yLhG+C67YQYMq6Bq+us2ty4YCrlplaQsUopGixNxj205eZcOt6eZHsMv7Lw3DWDqd7L+cbNAv88
oHGx5ZRqDtMkCGuKvhEA+wuKW1Y86VTms9x7KutVWoJzReY/ZpKB78PPX8/ra2ZnayRnufq507pS
CZSB9rnv3JJOxL0K+MIeS8fqs8+Dfjp0Zpx3G+1QRQggTeSiXk5U8cSo5z0ybr1OzUWAeg32fPXz
QlfGoKrFpRDkhzNW0F3d8sfIuvZSY4DNcQOT65L6ddmmhyWDd3SsHMd2JJ8WX4LtCD+OQkw6qCv4
X427G45NtZ+7ZoXVxfGRnl1rEAE3HTIOKIvVZfwpUPwKk2JxP3KmLAAxhVp452NFb9qUAInk3l+w
aakCe018KmfQd9gzro00v4L1MlFiqosLe2b3FAZgpT+WA48tt5xQCZ+S4c6lX60btIgWbjOkN0y3
iefYFodzGFvwcXvRhCXO/WIQmtRBguJdr6n8gTbIbfsTOPhu/13lVjcjtnjn0nRlZnaca3ko8l2T
jkEwbqZ3tLLcJcEFtNG1K3CkXCRiUQ9NnuSkyCUKQ2GEzzA2df25/OwIk+fiUhcVRKUzTEVaGqdR
I7MuuaYLG9t/gNJzaWgV57KAQRF8HuPDCUH3TsG3en3zfeisXrUdoCbtHec240gSGjTxiK4rXUMr
VAIzc80KNDmh7opM4O5QdCU4GKrXs3vKhoESD2sP8Www+SDwHVRhJFt83rRJAgClOVkp/2Off/T/
a4DS9/+/HGnd4r3ZtiDwK3G23g275daCcIKe5+2ymoSaicLlIwhnJY7tvwHsETxhxaL471xXU5TG
o4/lnNIBFFxBaPHS9Vvp+cT9NmNLdLNGLkGMV7V5WZEnTlWNSGhOrADAKgVcrctm+vnr8zSoXrGD
798Q49ECIcyqjqnRKZQxrcj4Yoe549/VS7YyCzLkUpYdEfqINaHM5RVPYXpTOHjurRL81uNsV0JT
dzef5Esfh8SFN2gLOtctOKXVAJI/xA0J3qoVii83x+JLOHfmOt2z85VjcCJo86rtN+O3ZkRgmWb1
VJ3EthNhp6fgUJytU/e0x3dM6nLRomDtzx8eP901q7aes3y+Yk8OAdnGO6ivJ87fRVtpoKkytsT+
CR3WPt1IxkeM7AHDfLmj56b2yfoIHBwXaHTIxiZVQ5MPzBEgmk6CX9pO2KY46jfnQmcLZaArQEW6
TEBeL/kILlvi+RmL6v6z9h6G/QsopXEqSxCcH5oBJ+HWGeXY8QLjpl/ueLN6KzoEFGM0uzXLzbmh
3C0UYqj+xkifPBmbvAELkyhAFdmf26zfUnJa1NoDjk8bqQJMHJrOpY5aDuXi9sdO6YcXrUyD0m0S
DrNKqm+NgoatHRSvu6RLwHxVwEdSD0gfOn7A6KJ8f2wN6Yh7zdmrQpO0EL7SpnZdGarf+N0Ok9rJ
NuF9UNkcUc/Dx47CEsGlOqHzpUbmY3EVxiflVRxFm6rldSJEoXu/kFmzZ2JyYUi6FqszH85lPbO+
UcSrk/VSJRg+WRw/nJq+kjw92eREdb9c0K29ECi8ym96zLCCa8VBavpUvMSMGPXPkXfZg3bjkXGm
2ltS3MAexaMdQVu46umYly9CKCxzYHWUO0NfOhxGMo2wfbX7C75scEEPuMz6HiNeKG8Hi63lKmtZ
OT7e6Y02o+9xiiiSuRWnn33GDkns9e4SHj788P6w6yTRg8CcyVSXXfMli9/FIxlysP6JV4RPve4T
YPPFpAqQOTy3RaQ+gPUVxwt5uwW2TuoAlwGJnae5rKM2yezgOA6VvZI3dEuX7r7sT0bjSYveMhIC
bu5ofQi9+Jva3romRuGyruotTIqUEMNQtKaO3uNy//FPs0Emf4p58YXKj6uKC5iDsWFnaXVl//Au
20apmzoxuf/OAfAIkpxZY+GfNVZNnwuHQIZgiPOoAeflIjsyCZEpq9JCr9g5Iqhx1vybjOPGsRph
w8PD/yxdoNd3TZeV7AIL1cCvDfxEOmxrmriuRFaqFqWyXH8praVNkjHUcBJU4G2GK3PhGuAt1Ujn
ctvmyWDzLrSz3hU8sfIsK1XlewsaRPgBS1LHG7jTv16CsN4AyjL4uEpEU4l0CLsQMyd9Gtr5ycQ1
cwcrvYWr1NDATlIs6NBiIU5O62g2kZKhS/6NoII+swc5jax9BnKV7lkgrXmpG2uevMZ08ZboGHz5
oSv+s7zeQ0s5d9m/PygqQSP3yDFG68iJ8eCbk7Fy4Kfuw4meYrz2a7IKi5yvEbpZdRnytRmrIGbC
Ki5dIBOe0x8VTCUuhHP6TUfyF/yQ8oKoO374pvu+5hzGooXa2yiZBZ4aE28hhLTeGqa5lQUm8489
3KEnsHIDk3hbnz0422AD2BlggO9IZEM/Is7RN1HZRjp1U4m+pNO5tK2l1fmLAp5HTBKyFVez49UF
qcN/ctdWADpiAn50P/9GKKZBUPwtuNXkcOUkD8s9a5SZ9RcPcjDmZSySJ3MBOHYcq8NPw2Dl47rC
Q8nR8W76Dwfx6ru6hBQlDR2FRABnBr64QcNQ3NqrAa5GISpqRzDe7t/lgLkDBHSH+0UMsA/EZ/9y
FRL9tt5O8/w9Ur0arjWbEQi2EzCmDevajieRf/P5RbRlp+8l7cLwboD5hHacXyEyVBxXO0bFXV+k
lAZpjooV31pD0cMGfvYAX8pVeUHbaVaBGj+ySUjz96tm+iSZDfvqTN4C89TdFWw9NsMP7Jz4+YdQ
eP5kr/JsKZ5JgpQv7E71LoQ/ZdQZC7c40LD5svhPhoHOWj6aYJ+AJZzlCtVhtmHLwyw/6qg9W59L
CbE8baqqhm5mvDxQ8UvVJ7Knmwy4NzY64LKomva+DWafMWq2EPfNJBukXtnvDC8d6E3VEyMjhZq/
egIdGM7BICKbEOMvienRDGJwcJfl4xl+ykAKnX3TCp/p1MDznlOnw5EozF5A8scRcNtraDv/E+8s
LdkM5pWb+wq/5UbDmJdDJ92L4CMz5cAs4ncMR+LTqbmnNc459mfLiGHjNLBnZPIVQ8I6jcBjnCoT
tEWd4rSiTFY7hBLcFpg/uVuOW9Wzwm9dcvC2XvWlUTd1q+byC/A32E7f8VlmTFzJYnEfkuBvSvxH
9XFrV3OCM0UEdDMxqnbvUrQMQUhH8xhtI8gJNyatUpI5BCCwdsJw6hOjZIBFo5hlcFwl8iKg5LoK
8SPcfmEB4hnuQwF9QFZEdgkWJ7QadL0FvXk2fLh/Jibvczf92u9I9I7hWkMt+Muvcl4aUT7CIuXy
o7JKtb9mUYOASFy0mQVBB8FTYdSoAjsC1ErHfckE/nAuMcFix5x0SQi87rF8bgUMwt4Ic2G+ouU7
H+XHQp1G7usLS9P2RQjVC2V+lGha0ri6mQkAxdn6xeKrSHQQNVOSnkSIaIBSVhaF8ldiCv5cm3tT
F0a7PxmAEw0GVMHdhIHErl6OIbbuNR/ggvGZj+PrlMPWwZDGgUeNXY1+QTfiXiwo+ijyoeQRb8eB
jHiEZf+xN9icaxC/7Mt8Svq/46yGPJ5ppum126XnPwm2zvClVVp/PisJ7L++DKXJojbGYTUsDj9W
KQXrTdIIFbi8aru7CIFvrghtvqewQOVFLn7rW1yjiAslcR0qn1nQoNTiGa5rq2Aj30IgBSXo3MiS
q8rryqumVIiZ0xJENc+ypuBwaCoaImt+nIpkRgarZT0F+LgSgCTCwCduj63XKpcqSQUqKDBYVVhs
LEVImRHm1zsjwhPTJ/EejrDXKkcNoI4L59WIdCSLFYdCyPgKx7/tjrnFr8Sl89ElLQAyacu4A5t0
XQJ9q5ttaJTfNxBl0b1fbKjckIERF+advasRiYStzqwxXnPCNUIQ9hqvQmF++VTCHKYZliarReEd
d5YH0HG6OPrQLNZLMqPXAXqApe8hhWd1Z/vHE1intCcMQ7kN0ydzQS4dqMRuOYkbB3Dtl5GLNSNo
nDqqSUV94Gx+5ENhIt9MFfCMcdcTLCY9o1wvY9fEzIXd5pkqpG/kEe3UVWceQV7GbDfR7U8q4pln
q9A3QFaVwVI4AqYOtzSdU53r5thVsm6zo5epXEqv8T0vEzKLXGJ5Wf2mANjVS9lNbCT+nOLD4yYA
CUrDUyCvM9M+LYxph+4O7dXKQdXjrmgGMNgm4DMcEgS25d5sWk8FB4a7RBRYJSVVBzdXQS2ckiOJ
jABD9LtTy2xszH1/DtZe3jXEV/2Y8uO3owQ7E2n/q61GgYFRLMK85J19vpiNPvidZxNo3hCLs+XB
NoaAR0p7A/UcpbDqYoSdY3mfWlt7LD0lG+9fpYQzbVWEr2YJJ7aMnB0V8OmcsdPBi8fCxNXJP5UQ
NQRMM42FyAxi22brBlgBPSfrmA0vF9r7kqROz3F+QAJEsCLzbDcsZN2CtJmx/pBI8/j+gYKMJ8ce
alhr3vr4cD3wbzT/6dIyR0SjU3bBWFucN4b0BrfvOIxHB9pwN6SQf64FN0D9kbxcZiukoYmfrW1i
7fnrs9pHMS8MxIp8Bt5i51iO+gn1tOIyZ05uG9JwOGMCWCB+9KIqQ8WUPA7OyjJfQ1w0wsa2kXbs
LNTNlHaZ1XpqcA+C3Tum97dqGH0Y9z1Ve5T9NES0Hq0fTWRBLBdglCFjZ7Os8rGypAHZZXKG6Rkq
571TrmcFCvBB2tmzae/XNIOpQUagg9Pve1sORhECf8FBhWh8ZAOFFn5OKyOmVdo20Ik7PQXkz1mE
qiZFU4RUT+nmcrjpPaZCKHWU/LHCkJZRUKWNRIym0xMFIur7A17xezH74CNUQIbtbI7ap+qSkxYk
8u52BGfBFmBApB6J0tyRnxYi55EFkwrSJQMd7XVEIdGThcxRRwINogb2lzHnzI1sK0WqSBhHzQT1
nc5WePWgJXyQtts5V6gjiBWOOY9aDz05HmCNy97A55BUeIOomz8RRfI8uccADt5qNzXGovTnkzxT
VczKSbji0+YJDuCZtm+/9ibCmacDaPcRdt+az2TDZ/NcL7BBdyZWhxT7DGmWFrLuG4H5iPYqyhQ3
Kr0J2y/r2+a77vE932uWyxdkHhQcYQCUA3HhfcOLpl+efbyiDKvxHhEHAUnZhbgZOTfAKGamEgrZ
/MIn8DDapaTE3cMLjih6QbYJgqQ0Q6a9HCmYAoOFOa+ea2wgcQRH2xltzIV4KNxQ48Mrk9GeBQPV
3jdSU9Y06PVDLCF/pyPabN2ieD0KMtz32aUo7wYkP5+nw+HlAwJJ/2grXOMHm9EM9bTZtB35bJvm
zpapmil3E3SwcdAMnF7uSkvU6eFlH7qyUU8BFodiPetAKZFYFxItIp9ZvNi6Rs2GDlaLRFGqqH9Z
7VNg8/E6dUM14bQ8S+Snlh4KMuAY8uJy9cjsxYog759fDzt6upRvDVs/Gn8YcifFT1mLw0yfQqoa
/S3e4nzicB0dSYsraHgrZRTH26+m0XoBgo00srpC/ZLsctHzhUdXfkKAR8aiA+F7fFiFgpIoeS+s
B9jMLKjPEv/uLiSITzq7t55KN/Zfu6k4mWZLVzCiiIaf97isfz6xpvAioRufnAoxSqMab/72wyQW
O7xdQhGv1VM+iGwpn9kxEKigLE4dPImAfJ4vcBkBH168U6so6pbq7Vqrwp7aZSJ1o9YIueER6SDZ
z58Oqyv0SWkuhjlid5u5guK9n7SgLlvlbVJQJZbHk/3YTevVLEfS0CC3H7QiXIMoPzlydcDwcprm
VJPKcHoLWY39YvEgTMFARR2dfOECqaDrh57FiqxlHA529oS1oM7Co/O6IjZdSjKecJ0SH7t3F3Wa
iJ9BSyFReeayR5DoOA1C/Ejqifdpc6v87CuIRdYogfoJ+PvxrSQtks6uq0TL53RiyiQYl6JkccRy
0jyASCFDDsNohjg2xtotHmKNC3d7OPKvS702g3uBHfZP2xNbSX3SnzuCjjkCDcSL77jz09QrzIoN
f11ueyi9YYbD6FRrRnBINxgzlaGCnc04TfBufDP+4o1rgHAolcQxhDpLrZ7zSVXiHrNuTjUSXaIe
bPBqbranYaaf1rSBiOLeje0bn2wjvPCbpkCj8DRdRx+wCLocC5ItrVLQxpy8YXE1ffR0I11P1uPM
iYhfCn30s96fInICDpDCDEysiwnzQIoN2nmRahrlzbsNlbuZc3ewHaKqv0BNqS6vtnJF89cyA1s+
Xm0Z02L8Aa7pLZtw45z9s8werCUsfp9+l1XlnSrd/8luvkeyiiB+eJTmiuagvbTyNqWFIWZxBI4T
EtRYkdLSUM4bdZIJCMBPmDN11TbUlhnuUbR3RV/cC1a/msNdcZNuTVpkEkh/RqSwuz3ph2KZ594G
Szqh4ukB1sQSfLjNDzKNvnYy8fyg5N/2C76/PEa/NAEhU2mdclo5JePIhTwMcB2xmg0apXE8Rc95
CD3EDdN/4Bht3bUbRhfMPBPvylsWkwH8sBhgUowenGNdk4xhJXGefYJlp3YbiixOVcniHzKycR+9
kouQCzKUh347aMZIm/Z7qTO7ek5aIKEb8Du8UX1MNPy3RAvFOM5IIpik4ck7UrjjoUu16zdvdRd4
kM4VT/YXa6ek8zh6LOplWAjCDJ8lAOcTOm8o6bdVaZUpNVc1gmlR9ITXefpdNJkGenmwqMp/fCRc
MCSeaWuJgGpv+WJvw92y/LTDeIoDFq+ApVedcEzZAeaUfF6GpFWpnJNKMjxGrMMZkwqAzcybjMdS
FbibcysSF0zt4+SFJtt/ujo7HolP0BeubOFFCcGEJY6w4MYrgU2Wywl/Eom42FdxZA5/sy/CU4Cw
5z7H3UzyVMnoakQdLXh0Fopz3n/QjRobRTIjWcvS2lvfVEwVKWFuvK9R8fbr+KBlFU+Jk4pewz++
qoEFRbNMb2IIjb3irizkJR1dfDbG9gUQH5dNnL0te393dNUKm8R2QeITD4Kt3m3xNFB4LK4kFeV5
wHuQgPXK7xDzBRotXBk/NCTjWL5ExmL/GGXhrqkt8R38lHS8cbJcqxU0aErqC39R9coUybw86a2x
QtGmrNu/HgBP6xhqN7qOby6fOZc1YDkkf+Z25y6ngpvm0P2JQnNfUTaxjv6OvRE+noV+eGlp8KiO
m+ksSlnATPCcf3LGBJJoCtHUEpkYNM7grz5Vx0pTLPpeBsh5j+mTD0qWPM/N7Mt/+gDCBf7s3rbD
ToBCRpOljXb477f/kpddaOpiqR/RtteLtUjRldLXDSKiQJ75kDJ33hQtmZKBsSw9vICUK7U7dYXl
Mqqrp0zFGfX5wqkNsDMYL8tjF49XBaOPLENqCJ8m6SXU3nZlVR/pDoWtunUNfrY9ZX3zjpnULTmV
6gq2AVBFRxkDPqVRXizO6V5ZSYFv29t2luUgRwvHx3jrT4vIvsYD8bdS1OaY3OLEssdzd0cZkeVs
BNhg/ipcqgQl+XygjrvwSZ3SzJ6SY48GVFIny9ES3tNPkYibJ2soWjEtf5piHVj+g2Q+JtktR0z9
kE3PGtwnW7aLrpLohVeHnWUkT1pfl4PNFsdVgf+Z0TM07yumxeZbZ98OJUmSmaXnAHuZxNo7JcoS
7qeqqwGFL0+Cnsa3gRAeddkGos9ctJt8bancDMv4vzYGo2kGXrpFTCLlxWZhwO6kBRD64xsIAhDq
P5zYqI7n8nU6jAeesZPiwUbVwvvy91mG9EU78WUUC8lt5bTulNe8HVEXjHFqQEcbzBtp1DpaHo9H
NcbnnsL+7RgctqSel1lzEmsduB8wQTmL/8L4XN+n80BBRsU6j/FkoBmBxmBdVI9Ra69v4m7v/ZI1
7bKfKvxpYcQ7aCbUY7P2ze5R5dTlGfpTuDFdH52Am6Ha52i/Qh7VWPvzGEtU4uNQqKa3zgAf9MTY
+e6ht1my6lfT7B7oxiAZAqlwaMnEPhXgRjfFT3OD0YzhVFsIedoiSZRUbM+IZWj8xhXetxZ+gTYM
hLPNOhMJsnjr7Yen+LOQxGcRGTsXdIoFCyEJZf6NXUYeyAtnS3wG+ruCBiYlCfOxyk74fUnKFY4I
m4/ATWvm0Ot11VZg9CE1hx0TsS5jPPkzX4YF0JXb9Rp5vkxLvdQIl5o6n9Wa1whhC9Lkwf73MVNB
eTxZEiRbs7aon+aPDw/Cz5PLVevkFzN6Wx/OiCrXDyfUxH6xzjRsp+UX4AZnoAR6S/pag+EFlwmT
w2Nubc3HL59bMuVHiVHLafFqhJxRpm1112IZj/WxEeSmg/ccls9qOlxhnGBciUJI4vq4uzQC/n4f
6WsbYhFLe4eyzDTyHPQ8ASTUHk4YMRsfWqFkMDfEsytTAxogldBsejRl+g6ODDSctSPy7Vq0svc/
dmKQCeSiywPBvt8RHI8rSR7ABIPHL5KRs90D7+Rrj5sWK6b1kxVbkcGzYwY6ai+SKPxpIaZCIt95
/Pim+WrQ7/WJfWjVs51nURSfizFUWNY1nMh6/sqMiV79rPM53iutUYG5Ufkx/FEsqxmaxUxWeMcA
7RvmqNumMhgw3rNLDf/U29G6jsKckqJTO2YH5rNhWHXCn4fIv1xgUo4GTfJxuah1wEFGA4RTAaS5
zZ1hMSQTcloq2WbIAxj5/BnQK6/5RhTm3xNkzbJMy13+D3LHi7AbT/Tr2CO3gLld+ftJoIteJRFP
+hrY3H3EXIxFEWGRqG8DAlVvpFGdi6LI++zdAl2j1VKpUbCk9sJp2KMDLPna7JJXCjoI73l+cIbf
byk/7TsYBLKBsI6Gzt798cpFcr5423E2mSeFd6PPZn5wGJcQ2aAb0wQjfgf2uV+Y7Xw6udfSv8rJ
OizGx7kX3Kh5IWLzKeT/FdQKaSjyo9jQNhtZtNl8BHDSm4FIyMIYMoajc7fOMQIrBBHwiHDxF5VK
bhisyMOBZpAdBFZCjdhMTHoYVjQsueEN39SoWPJUjcNoQLz+ADKPna9lBdn3lu0wR5JMq9AcJr9h
zuzrcQwVDR5Fxdz+bHVcAQywl8gAhW6LIyfj38YSqDYm8aeWVf1QPH1LcxUUmL8Dtk3cTDNbP3zk
utssUCE1a22DliOJakrz1lcLAQ7ajmanHAOM6PusxOoj88/0wZg63ijhPyNdwDPyqxW0+/SHCjtT
McpvkA2cz5i58PfrOtdR6EkdfR6a6R8puWuqugj4t6Qinzz7Zl1HDJfbuqZ3tt3Tj10Tk78dNvBr
LIFb3+XroPJYrUt0vW886C9vPK34Kfh9fzqbibP4dwcslYRD5sOvHunmnmNq51lcS9XabQ3rGeKP
vtHB1scd0pgp2bZNYoCn6qexl+mivGlWG9nlYqJYPepsUqOQRs4gsQ7NyFeCfnej5V1ibksVp9z7
5+MzfarxpuC17rLuxEf7CgiwJ5yxRPbkSG1MTciI+0PstzOp2u05cWpzlHZkmkwjXhLp4IEjfHrz
Iq7AemMTeIbtyGJkJEpwoebBt5f6J25uQAH/ETmCNzSjLubXz3hbu83CBupOtG+6SSDT/205Sg6O
502yCZem9jD9lXsQd/utqHQrWDGEQ1gsXbDXd/cO/9gDH2wiOC6yLdhjECkY249xqgeabWebzKNS
1YDJzZxdqHMKYWGkh+reEUSdixkf0fsXGFZlvw5EkeuO6Mwj9U/mCp2Fd1veEEn3nyvYRupeHnIH
tSW/TiMhdpw8zwqTgjo5LkiiqzynoieZ3L0601rRbpR3aWvyuFexhUT2dKqfdC4rw28ca1MLOI24
GkkCFCeChJiHPImgNpE0bDqAVlY4OA25snVyBrN7mx9d4XdjpCMLx8FVR0NguUUl05Yh3snkDaXn
dA2oCEjYDXVZSsf6X039KCV5UxlUPD8AzFn7kSrL4cLcuX98Z1mRDCVQqlDww3mN9lwdNNvu7mGW
RI9wzXQqWSwkWufLKsoqg83+nswl3HXY2HoNZXrbnFqZm5mCRXffChYGt3DGB2dg7F0GRPp0KRol
YekdzzC57zdDhCbCi3a5pN7cC1Hr8HEXmslztquFJsOetBjDE36hibGldDtt2gZE/pvu/DdSf/J9
e0vxAeNiYds5JVFKZPMDSjfHWBU33l/1pDaoI6r09YvYya6kXs/ZBrJMzMnfKUsEtbUfITSMwDAv
f3aXMxCDARW/g1qJM6N/+UovBu/FIg63oGb1uZ7IQlFlP8ey2VsTYf0OPpBSDSrl63C55TfAQ2El
HOWmc6i2kFEKDJli+F7HpjaXzrBu4QnA92+tVDCpkeUig6+/YpBIoUr34A1kP3vypIKP4h2gyYJU
o9ZBWuG3FUjxv9SCAl7+cHi8grzxK/QNnsmy8ACSIJsuPOHNZB7TXZnrstwuR2ra+ijORMeRwS08
8HRe1bWmcZgCGTSFBQr1JV8bCwAS4R711hjVx4EsSmSs0fTpmto9jBCEtWvQAb78GScwH1BrOpQj
STmhBpzAKm8D4LExEjdEavrAV6YqB5zFHF6NVagcaXWQDx1rGkaFtB1qH/2FAGTqSD2ZQRl6zHow
98JJGzfokxUffEgFN/9fP5W75gmBFv2o0Xnw2J/2bpmeqA9l7/WxlGrHfmTMZ5Th+oz1/fbNrJfj
ZojN9PLhQg63XM3i5lOQrQ2hqy03x7i5hwytF59x2NdR7OF0qubtAzRj0LTLmixMg2nE+NDf2vOy
mEQUbf1Njy8g0HDYOLt+pZmaVCDHoeIOJm/3rFpV+ccmReTaXJtBKiKyh6XsgNnqmdbzccEDX1eA
vY8gLtKh3zFskkDehdSJ+WmVEeo7QxiVTgoUS45fdrfoRjOzY1RT6iMK+VwpOXV6Zg+FMFeAdBHt
PWW0wOhuV5ssmriJFb2Uudg36VZ00EhdI5AmeMy8T69hS7tBFEUyiqpfnGSCdG7cEu59wetaM4zi
pjVkSQnH8GjQlLO7BPdGpYG54BEo1IJ+Jue5YYn5slE678UQend8eWbJKytQtFBHxPM9yxBSYms6
pRFN52sPI492TVODa2DyC8vUF63NqtChIsj5tgY4MfEjqID6I1iucXz4TNS4DghmD0r9VeBsNuRI
kT5Go4ZYoHOHPQOyOSR4vrO9Y9zqipFWLJcP53veAaC9VQq7cgPD7zpacAZNlxsXzgx0K/V+c/dp
ZyCHA/yeesbBfdteog28+o2Vf1IR2JgYuE6NxSfkmnLa7Vz8FgZms96y0Nt1J0oRUASbtFWxyYl4
KDU/hPm80n7sfhC5yvtTj2nmenF52oYtxgdepoQ5ixgi6e1vhg/Ny+7sg88Y+uQ4zoPFZBi1XlG7
AOkBvnxO6xO7c7Detx/6vJiijrwMb7/+hxexfjpOudl6AMwWcBgTXfTkxGAf9gTkXMVTgG5mk8gJ
zrzWN0D7ak/UrCw3iPeGruy55Dw0NCq0rzxLO8J+QyJ65HQDPdIB+fgpk7QI6ueLLE6ynXwHpE0z
x2FK6L8WgAlnuSAcPTUzLWmgX8AdxRkXhfjvlQ4COsTm52OFX3Pyqjs2VSPxS49zRH5rIN3SOPFx
IxKnEi90qAy3Zr1tx2i8W52ywsGSU2ynG10QULjscSCfRhJkbx8/0MTM+LkeN2l5oGuO2OAcP3Qy
T0F9WFWT90zn7zcOEaKdaRbn3bOspo+92AK+L5M3zK1IbAybQ6K/DWLclZ7EZn8LHNkY0nFskjB1
i8IAUc5ed9cIc8btoRR57pHYcgYR6hAanzPjNjOEH7y7vF82ovCFWU1YlftzmCgaQbSFiR+xXY+M
5+NhXWNV6TVdZSlNjMk3nm47AxZob4+kwltDoH/0v0vmCZqWqSsVKGMeWJSY+NuyyCzDuAB+VdKK
6v1FpAo/lV9gnNRcXiy+wecEPfGa4wiXYxx7YFxffdX5a3gY7rQQggDbYbe9PVx21eBiJdrN91Ir
ViN+wKKM8w6F9apIYBEHzvsaRV3yTLRk51FNgv06r41gOJpXzMy62WDPk50IkScUWAMeb0LycQPD
tPdEORyGQg9gaahb8fv6WeVRmAf//aQYFly314/ygbzfba91W2Qfz+VarEs2hbCYOPTZcxkbuFdG
WkRQE5pm7d8NJb4+SsvIc687+pKklCFoSYisMN+pCvQQsF64aC92emKzGcx1yDFcy+OEiDfX1rvq
llUkAgG1y/+JXSLWIYfUVI1Iotwu1XCW7ROhWnW+nsDqPr1K06pHOKIRYclJHeT9zwc73OvGuUQK
pQQXQXobXyakSoS/n0rJeB5LJq7on2HGwDq+SQUcWn6Y8+QdGtzuqnXjzD+5cd3rnRrdsPxjP4Mn
S2pT+4dKhexgucw0heiDtQWKbn875N8HQv+MMCsCJmtGUnqNwdMBUW9fIfy6+ffDUKTUoMW53ULQ
szA05STMg2kZiLdCkN6hq6iy2i2wMk0DgGNQt8UOHmy9x7+69SZJUb4oZuie9UH1TchAs3Y2a8LQ
E6+9ct7HPcH1gLuVp5vHKn62+LNYoHbDq/OS3Qky2VFo16UGP3ewz0CGRgWI6sQv//fH+VrDyWtl
MKjScnq4ZetTWGIOgUJEJFi3RwFG9QZq6Ppi1UyYW4tHCgXCn/URAcT+LDX8I/ZniVQDNJ91MXkJ
CbZ1H+8iRB65U/9V6/7Z7r5EIWekYMVRgcxNBJIXwK6bjHVC1MlyjzhyqSJ1n44akNjQC9WrIWeW
X9neZDMl9KYvkz2QOewoDSH4tfZrsc1CmQdnfLLUV9PAQApoxYFutYc5Eb4gG1/l0EalW4BGbqrc
1hEU9V/SNbDCiY25MxeWNCpikeB26y7WKfGSN8S/g1ibc0l2s1PMYPGlg0+pHc3Te0ufOf2kfPzi
IVXymLJLFcUaOS7WHJOBLUZrSCgutTg6Pz1D0nNapJPd8/Pk731ywj3DLEKmnxqO0Awjv6HdAcIr
X1AWTeMy4LDipnGn5Av7dsAzcYjSYeG8ROGG2QnQbGMFJeNWMJMLmfdvAI/t7q6ipBsL02lys9FA
g1XmrVmPMEm8GGVRQ+6BB9q8l7BRSS1kOjjEPdIgG8PR/RuscN1VIFPQqtS4nlZw0vHDOMM//iZy
UobV5Kvgk4IDIKsWR7X22nNWqn7delLikqTf7aBPMjxPcoPClKMZ6x4hbMdnvPorLHDG1hEPzzlC
T5pHnzwtQwaM4l5Nx0dlfByEFqHZLLsxZDnPawNnrwZcHVKQKyNp7J2goMYDMoz3xdcQsBxlvnIL
5SoUbkbEk/cAuLIorIS5Eq8JQjys4k6vfl9WkUApUeu/Q+E/OyNrI7RCavJmdDVP6vykyDPoMqL3
oTbaUQ0C+fehrjDV+P0kly93+mcb9yZ7dnTFRCNafuaj0Z2rOCcZsmJwkntAxkK3DXRey3RUMMp/
+YoGt1ns//OJFoM0mHclyWerAwv98Bn/UQ9FNcl4EOG8YNa7f/DbHsLQu/u/0q4jibbxSW/aP+Wg
ybdI8rImruCJgXYT++g8Gq9eEG4/PKMoK3s0Afwd+c6Y/REBbedf4VEdKYbgQFns6faKZRaMxaKn
G9lRK7ZwGGKLuyOjuxNPaRI5/Ppqh1sgnQcizM2q2qup/kVPan8gTHEaMHRtAJgrAqUq+bdKYZ1p
n1iiCPRpamahwIFLRDjcWnB0GDL+aSVOXipY9tdhtuWP62xt0sRCxGv2+K4AyywfSTqJpGTLavHy
V9udyFGl4IsBJSGjbNuPRqSGmYnrKTN9jQ3YBjXb1nNPJDRIjDGU3ptmZNvQDkmdJ5WwNFJ7r0HN
gCvx3cbF54PZyV8+gT2fFBOdV0/NsZxuNU+0fotD/1w3ahI3iYdBfqQfSICoebHl8ghLHVH+NgBb
209OuDTKEQ2I/IqIzP3g0IYqH2zWeXx+PzZGIFT/b66rrtigCHn4uQ5+wF9X8koSnJ6DCml/vCNv
E5g2N6ydJIaMwtgHj8TXz2kIhWTLqgzLz3OJToU1pIyp3dYQgggAP6BAm6WOm6R22BJ438YfxQLo
CuXdjO8VvWxd/BAvJ15a8sI7fNFfgpZUQcwKP4gxifoiCaGKBjQFnpz8kbZVcnhwu0OJO0vvWLzN
PBhFHCQiep6xtb+TxVct1c3cLWEPrA4nvtyLva97qvO9oBPW+zKPWsPYs4QYPe2TXuJbAg1y9Drb
kyRWPISmS7FDbJleb9riIgM6XctcVNyfYA1bOdQClXwe8N6PeFsSiIat7/mVshWkgXvTJtD2DTq9
ER2exqhG/td/EH57fjdpTvUu1J3Ue9eFighMAz8QSwjdtyg+oB1ZfSTDAcJqMqfGRAKMjnAwzrdA
QHtYdmTJMpiMs2z57bWG2LSOtjnVxIq8X5pdoiJcXa0YguIDWh563/9NHeBgLXzD+dpYBYVdmpPF
FBh01YThnaC31C5NeR/EyNcB7Wjwsgb+Ry8VIa8ig+QB+9uEBbV2XIHKTEkrCcl/gtaBuKXQAGsR
TLyLMqnhvZu/grxLF01ukmLXSP/ZcOJ/vwhY1oy22rnTPq7no1Ky3o4HANLwao/cwxNEB2xNKXH9
3d5ggWiXOV7mUdGv6Vw4RCYBZrzH32cTd6scNoEqBbyCEsGmEr9rp3JvAkfuqPPUPHw6N9YF+Ml9
m+2uwQQevgs3Ja+b/ck5SLfD7bHObDyNYVmpkM/ZYHazPzOSJMb3v1iFaxL0IVtusJXLwf2sn01g
dqdBZm6KLDEQh8mENOlkWwYIjo97+7NP5rRHoymkNSNEp+vswb3DHk1VvJSoFyTLD2eIUUHOhIS0
nmDr1kjLcHyLEUe55lt5lLPn5ivFU6XoKYVRDyro1kGkddwf8KWutjqw82iIUYbmG2JXFaqvp3su
rPr2/tN6W+PqUFFjTvGbxnksp1z/mDLwOqQcGDW/Zar5Q/Izx7HLQKZM18kF++XAUs9PQ3+jeWRk
jfUPolW2o6aLaNf3oYCpOokxgJ80ibfAQw7Vs95uTeBe13x2e7oUGK9hCv17uT0stevE5LAsT6eJ
h1dB1kY4woo7VmWixx4OyH/ylJ/F7NrJQBxb7CNpqBQuu+f5KexylJckXmqK8Uu9Afvm3A0BB/lR
NFScxfAau4M0xauYEPqIZGyVoD8ONkbkRdEWNuv/YikYVTtosVCQNygkRon/i13IWJvPyZnipM1c
mKynGf0Nbe1jjB0xpA8ZT6gy4B/2CBRMyIxxfKowRUxUQ1eY6Rbtgv5JgvODitovKR24ZU01wb4e
D+6CU4iVKSd45sXBMgY57OY26Xu4chrJAgaxr4MPSuTkXHFVDplT+vgL1WPDPQweD5e8aGFdollZ
jnh5gCLt5JG/pKzRz2Dtv457zy166waolnUSoDZARQtpd6LkwVwyF4kn+sT6HjEGBpwHbsyqSEFa
u4Wk3i8Ss1Yp1NBBli0GDhmMS1eX9mCaT60kzbdnvxYszPPQ4GE6Cl9dpTzyskoihSPp04EQJpf9
FNvZT2gUjYGwB0lgMzSK2/Unk+O134mr4eBalltFKU1+nBNr2P2Es9kXFlW8G08UWCvDIIEA/a7h
qsp17cE3rdDZWRdAAbXHLd423YG4BdJEEcG6l18HEAg05qVXUZF1QKM7vpAOnuTFMKU9ug905kGk
BXDmo5usmfWu79n4lBDKBQUrhZoFI4M5vzFHpEVwA80fKJNIidOK3BslXtVUytf13bf8u+pK1IG0
Ay8uWJf/fuZAIHp0VBUh76FLrez46sIPjowmdMnxuA6lv4NC2SQYKOcb9xa7N4K2k4OPfEdAbJVa
M0iCGvlAC3wz5vLb0Tg1kJSu3KOkIPs5Zr2JbaR0IjK3TTka7EVaqApnxRYJqvS9JEtAFbaZj8y2
EZRbSv/sCsnUkLVyRpDwrBzYqyETquL6WzdDGX6F7AKeTXWThwwAabOxx1gr4ZXe8jRHbCJ//A4w
HWPUYIluk/WzfiriMAtJdq/0ovDVcZ9UhSGicuia4rWKgP1e5uEwZtxgzVxe9Gz2UEwr2KfQToXZ
wReqaELWB2WdaROlMu3LWese4tl8MuMq1fAmPwh0Wa0jZkTh560dx8nEdNYECbpJclo2qwCRAeeL
NWgYwX2sWmhpfxVLSNU6h175eg8Q9Nt3ohNLasRHzh14scD4h2YtiDYfXtgX8d997FTA3HDkjW2/
ybQU00Z++20Ja53mLV2S6Gl45/o7qQvrAzccmAf6+Q27w4sqAiejriUQ/0pO0dzPDqDeUAPHpi3K
ZxBiJn5RVxSXC6tYT+bD9zXfYutrm7Z6Zcz2exlEEiL+BP56kXvHkv8V3f0BJ0YXRriC22Iuob3j
GrFK7SCcjqqy9dyszTEGQl1Jq52CT7wqjUJbNfTViDGkYKuhAa/fG/SgECQE2zXwxlae9Rdl/Osl
VmO+6/eBjnQakIr8sLH2n9H7xfvHFqc2OTxaVLMU5AOZSTWlSKpM3L/C7HZSwkNnvyOn2bhAbwFN
Kb6no7+Q2Jl5jLDq1FJz0zJBlZbmmZDHb20kBos6Vcr4x5f8HNvOkjUUntxh70fHb7F87LCBPobw
n1wmrG4F9kxwPhbzY6SQxcgXXKS+uVrsVN99lotWnC49KTesw9A8bRDzpJO0icSPZ6M+Ff8+Wibq
Dl9dyjY0Lesu03Obm5TQJspbW+13TsbMlWrZ5NSV5H4OE3EEgWhkD945vEBF2UdQdYxKPw0yDUN+
0Nrzco4hNqi2EoSP5Ci0FWuCj5nX96W0Sf0jCnXi6XeDpiRVAAmzPP/aiB7Q07hOZygiEiejqvrC
sK0B2Fp+yAzBEP01q7z2KD/l3rIuNxkbintMQPbAhpihCfMEsOIQYOJvje7ntXH0KAd4jKUVwFzO
7AzKtbx8eVjVIPfWOh9SzNOASTjx6QSQzoUt5R27d5kngUa4IqKm2j1YyLO+gkLdoKaghjFx0pGe
1A5YXLLlC5K8fWhpqL+vDO/y3t/xAMmkIG0jLUFTDRI5A+4MKc7JSNCZPFrfUw+NFoyzlH1Q+jIq
a29iqzKk2mruuo/vunuGZLI1LnF2BrJcR/ve+ga5G4+Ae9w8ENBAToy3zA5bbtSGXkGO5MRWmSVH
8HKeNCRZf6G9wrAlebTYOPCUD1RRbsNy0r6QUGmdoabZyay+YF2CU8UmghyCd+3CJaw3Cj7yQGoX
loM2xUgNzhx+5IFKJzXc3XxBnR8VnvHIoQ+P8JDwjQnX0Q8QVekpYzgWPKvx5lpxCwtP2KsLwKmC
vdNT3g8Q8S4yOD2p2UqtvKIA9saliI6qnQqe+AiqbkFCriFi7xUPi2Gos6Ajqh1QkaEDoYH9KGct
yBDDjqth3v8YrCj8N4DBjHBbWoSBd/AOJ4jmkV/hyG6/PCggPd9O3r8pVC0GFH5C15jM3YzUCbA/
P/vtQAAM3FDvvJSBWk6fWKiKUE8UD7dlyNcqPMXhYO/kRBQX4JQHhfNHHaDOvbe5ya/S2xGHs3WU
rMG2N4ttN1h1eW7t02EyQyfyJUUoGWdnj2orj/HXqqc7Nw7q7oZdXWPupgCA6lwOFxtY8DZ8bfHK
MAzoFun3mG0xnCc37p6jGfYyKk2NZ0okBLniBStciyZ2JvV/K2gE7PzsLAwt7YdTAPnNWrczWGjA
rFlnPUKR7+UAwfbUuTWiMYRZkaP4SFabAt5yulKJgIOPs3e/0rm/8xm3SIveEs1NhG4UpHZvX4EY
uVwvrtBdXV1oI37G7JAiASU1s9WSH+gK5hW/HTOKL9YGbLPakULvxsUQ5BtIdmh95mk2V17/2BY6
ZPQSEqIFWX9iOoHsZWz/ZbJo9EGb2VAT04jrSrPcZ5fvFVa8XQFJldwZxwM0oDuUoNPRgS6TLnQq
oVsw8KslU2TvOWOFpYJzGdDQdBZlx+F7yzlhO8X4cgkq1v62IanJgh2MRL79Vl+kFxrUUhJQBdEB
S2zRDNd/aBb7E8AHJldh6oq8K8tNuxBQEzoMzbMNWaN1hLBdto6WxTkMeCY7pU3RX3AiiXmYLD7L
KJBWOPcDw5xOI526kV9ZkmYLaFFaUnGbGP2uDftazDBvD3+NsqiJwrCgiaA7YEq/468ZcHmVsnJx
6apYYvHEPVZlENSgz5fjMTPFaE1cAkiukKineQ9ZD6vezC/fRu9nsye5e+QMjQfKrbnUNncqnYqe
mdozvWxazJlhOE2ryk26580sDKr/Ed1siM/AgiUMMwyiRaM9FNIqEqPr0WMDfD6268XAJB/zn9fr
e0KE8L4gKEWB5InduNeBLxmTtAfs5Dw5RviZl1PjPo+edCtym3dN6oyq/721xPjm6u6Nt+QLFQzk
a9SEbFHxRGHRp6i4mdglg3ZDxro1v1dW9sBbXvJsibVHaCjp0G2DVOd0BYITWofPA7N60MsWuRAb
lSBdfacZ9ehGKBUMXcg9W2MxsdtwkKvE9HwqjZN8ORbJUR1c8m0yE00wMW5i50H44w+VjqfejtIP
the4OE1t6tAJm3diNXUI/+HYnwe+OipwQ4+gFTQZ8uur9Y42ad9vojgLJT5pRCwqwZI0K0TanUDF
wQzpfqTCrDb/foJw65ABM5dPBFjWdv42ZRYgC3/7vMThY9CIOlPNFY7MKvkZPPAXdWelLtIfySeG
wDUZQEEPQd0gpmAPZb0zBhV3+jRhB1o0rIJZFhFy9QVdHAOI+ZJVTn65KaEjCwi/pI92jWjRN59G
jG2tDbdflsybUWJ/hWZUHKkpdvLc22DOOpW79ZDiQp0WI1qGMpRqDTMizMG6lP3MS+bA4cf/jvha
8nW6f02bdLHk9VT/VKHm2cL7fRfOfMuGu2PFNNAe0rd8eLm3KLXMnq6rhAigHT3Tft6/8TNXLE2e
B6TXAjBzu7yDd7eGuZIY5aBNZ7p2+BOpEMKvVKtxAsNQNSpRpAuDk5O1BIMgeixj/5A4qkFdnbR1
D7248zIfUyYsCUdQ7Qw/mWzf5ZKeHyn+ME/Xtmr+FKR1hQcoLSljgERv35XVd6Wikrj+EeqFnVQp
p/uqAUUVJKSS/03pk9AoIE1Kx8AmH5/XIr9egtZ1iWhV7SrOC4gNdKJsxwuvHEJ5WoWWF1PfhjUs
hUaaahhVIVAYCj7SE3Bzfd4oCR9k3v0X7ionAnBuIhJEJBx99SPh1Pgt00c5G/BWJsogc0TCqEem
ToPXdGs7g4MsyA8a6KHkMTy6QPfmkjlp15ZSGTJsca9fpe3gmaUxMCuC9W7Tkkhbjw1SUEbYgoCe
V08x3GQvK6nNuzBSRy2uoAdTYWSbAzw5HSdwNDpw+uY/o1KpvC6QtPyaFh+0YRQDR1or+s9uN3xw
PWfd2h8F2LiaKT30Sz7EappaPMK9Q5zVToSyWK65aGtZALyhCDK6fn74ORSXE0LOtS9kgl8j7OEC
wf7Y1bzw0aicZJIP+qrdvrZFw3nBOjpUBS6cn7Zn7EhuOY1INCa6JM9RK0fziVsD23VyELwQ8K3/
Wh9uAX+n4BPZXUvhJ8ytfcAp+nUOniFieV226Dc9Qv4bOmstpmWE9eUaGj26Rp8SkhkPSOqJwB6i
KHvr6/S7lF8VOMHhDZ7emD3fG31gk/1E4uR67S4UiGApzhVYuvglpTfYZe5fNFgxHHXnolFInHP0
IjOq0HCxzwDv7h6iFpCEakZETVl9TKxsvwy8U1MATYS6z1egZDqtksogWBtR6ZuPwySVijBOSEs5
S9vioEJ+bAYks3x8S0xk7l709c77nyDUwQ/dbgAlUtjKuRuDwgJBkdnVfb5zR0AeiXswo2UNFnlw
3nUOx6/JAlyIPuezN+cRCZWIHrbUVmTXa/T2n8oR+QoqwuttaXGS9giMcGAMChZn3vWQg4SuYCY3
TRa1byFeVQuniHDSdABwHfvpERN1/PacFTSpEVm5nki8Exu5V1ZN4PQAaS4Nro4MG3UfcEpP1Z4x
QaKPtVNJjm2HwFcMJLeOby3SttmR4hd4iMuhQSc6rHfwZqgvbdvan9d4JUKhjDnLbPz/ryKZxRaj
tzYmApS8K7Xe2JpbOeoEPNQd+JrG9rVT5igkZwyLl5NVJWzR9RxRUKMQRkSv4nz9Mb16u16p/Ssn
Ie6B7UIQV5MnxrT8HVMlXqDGBtFWkAeZPOPxdPwpYojukSOTStfR43pdnIXy7Ct4Ejh23E6q/jx5
U1OdrFskNAp32ouH4mR4UExKrExvMOovwa7t8ckdj2v31AKdWLTwUtyjxfdlanmhPl5iMzvXN1AY
25pYxbzWyjzLOqYaZEmnLPbBy/k7Rxo6ZEtp6Nrp9c117d9c2C2T8gA+sKN7/ixJ4HpC9pdQtizp
dkbuhWbThf8h2UxpxcKYWGX8Y9/AXtQ9Gt9hSMoFGgJ1wjyZMLJlRah3in7frA0cQMVaSzl7IfHR
yArhMc67j/P99Y9M8owEt8lgzkgwOz5lxIDj8IJnKvscY+WudxivooS+him9/PR13qgN7QiNld4t
Tz4A7yNbvokRuPjGvjOsVnHjH5v02rIUyX0JWiRVm5T2LyCz0V+lOOtzJkcP/Z9msIWb9MND7tEk
63ni6Lfbx1AJc+Mjg6n7jjcx7p8AHpOJt6Mh4/lN1QBJ2cukXQfOcnH8QKqe2DhChdin3CfOzeW6
9d5tzw2nLcBfP2KjLSZvcpDN0yvAF0EY/CsJRXipFXkgMPLFB91h+2gJK3Oc+AosNRaBjoWvBVKZ
gssm7zlNhNYQGGd7cYIiQKjh6D2WlZQMbHw5GCRBKH5lYEHmhX+dAhr70Jt0y0FkLL6g2HWg/I0M
4Zic7T7d5vBqBLbHUGVE08f02kWpvF9Ve8GgicjaCb/trOKXPNWh6x7E6sZgAJJIu1IBbz+npDp0
+g47CfSi4qnMfO7sIun5X91wcQsoZOroN28UGeyWEZhHIPzbvxfOdK4OJiXxthDIb7VdiPqowXyt
nTs91UC2jHiJTDlPkX47099Uyiw0UdGTM0AcWXByD6TQsSgJD6vO72TGleFSBVosFAylue5UrSlk
qQWBHiRZVCoIchvl2HiyP4HGNwU1EDI7sHo+0o4pq8XR3Av0m4RHtK3BxaOS/aFyyIpqainVY3Yj
umLKSsv/VTCiRhTAKeh/69BhS7ggUXPwOF5KtM+1L0NFUSWVlzk05HO12fcVgqa0+8qHf6ujFHUk
is/hlmtu+axohHVCZfODX7HeStLQAItVGeSLQHAmDkTVlsfHWSKVO1293MRHrsK/Kp9aH8DrNuCo
1fwmblyxH+YEojlHyBv4EPaErb9uByv30mMTgLmVsINSAWBoPPYONfqpcsUkkWnypb92KG/A6Ajj
0ow+KgutjaGQc+IV426fJz/cQl7oUcdKWlrSooVJUA10qSwy9/kBuuybiWd7OLzgvb3/Kkli5ksY
Hz4GbZJwo6qOv1fnuPE6FxB3mbngNIkuETCNR0wus4n5qZink82HGKvlCuQ1Ry0JlouIm6Vh08g1
D4iNopeeheoWimn/eufBmX5MqQw+hjQqBwC1QzQEAeL1MgVqYfEYZjX6zy61yffLkFxPn+Uy+rK9
pfdBfO8a22ej70MEXIhrONg0Fb6FCoKDw6bKqXjDdDni7Xrva9yO9ij8gLBv169mOTmCfLBGNK0D
j1Jj2vAfpdBYkfNODMvkslnxi+6DmnGnakSEdHHwD+LTMifo1zmYFgy5Zy6jOuGfePsbqdaHwzge
o6w8qJycOsarF2HwdwKmYkRhrp/ARcezlm2huv9EZDEGm5HA4F+MGnJNJfvWi6cIU7Qv0vrdT38m
b7oIm634igEuwVPb+NyrElVbmRMMNtm0e2K+1IaHhLmEEd7hYYEjDixLeXvlkzNb804MOB1YiC41
13/JuyZ/ptU8WPoUd0pbJM8MJogTG4AXzaLkSbgGtVsxKKp89ihiOxvbMlngx7HFsDXVGWqiGCpk
8W8EHU5WipAjWWG0aycQSmjw4VTTwSEoIXN6l6XXtyPPn8/7Ngz22YWPfdIR0uCc1quaIEEUmqEJ
BgB+gFJlBXc1DyxCPdirBVEOR9tMF8tIT7WFLGKVncjZ3hPrdDzCkVQHyG+3HknGfdOUhcaNFUBy
yT1WcX7b6qzTCNRhYMW8QnG/UT3zPrC5cyKZrRbhnkkdcaRLWIqaT4mWV40gGuHpBbMu8aViHn1X
gusPvY2/JHh/Yvy0nG/yLXk68puQL3iikMVxxIr4y24DyVJ5kmO9K7tUBo8oXuJ14koaPdEqp6Rm
wMiIn01nsp7vhoE1ouq11zUGkxauJWSwNG+pFlq/2xxdTafYBpsFjHkHuUxYGl/3U9PY1NL5J/fj
MlWqNkqWglbdCOL0rnPPrOq6jYDu+Dk1fJojEaGYxXiXEO1k60egsJs0KuNOwP3kKvZ0MKz9p7gn
rI2xYa8UnHGubftHdQ3XWm3ZAEOK/QJFqicbCr5RqP3Wl/FXSq28B2guO4akhYI99LMu9jBt19j2
n2c7TCLzo4b2Mpyfka3mqSyitO3KsJQskIQ3ThvIVQnM3miMglAA29lQ5M4NfCG0XaobPb1pWpyv
XcRuuOFFkrru5ODeHB4JwIsMxU1/Az3VEeJA2da67bbUyyNsa20FgaL/bce8psLu04IE/3ZI1Yi2
NRrluyAlC6AlXeEpC74apTlMwh0KsBqKcsrK+WvQYWxWu58kiaA2M+c1+7LKiomhlvA6P7MDp6sT
V3smDwlR0pXbTgEjy0pqZ1rStjwf5r6lkw6caszVIF6yFZMhBt2X7Xc+24xkpmg4tbm7UY2nod6V
PmbUJ8ewyuRwl8TIe2fCKuQ3KYhCeofbjolw8jAz3kDjkBdFSuA5VM3BT1T0JrC8wo426gnvSwlc
7L0GeSQh1qmzIrDXEvuUTnElkIjcS/Bl64VzXqni1lEG9J6g/BRlJCw9MfVp8silkq42M2LdKBUp
C0zlMrgl4MQjh8NxuZS0QhsM++1HTGBmCmEmirtXX07E/2tmMOw5O/5VnIryHxKchzxLcBy1gsyS
jSrL4qVnLm9+Lt+b+ZcWs39Rx+99CGpCuWyR4Ogw4DuMMzwEJxgg4PNphJXNf9QtAkd4XTr2nlU1
2VQES83YJ/E5pUZjLMglRgXiAi/V0o8UjVZAmgY2v4P56/0tewfYIXfxsUD3dJ12d+tLDXn5n8Rj
m1P4+V95EIDJyHUxypfmzh4YEwvjePNR/zOX//oRTWkLYW7Fn3iM3QUmI92Rol37AWwhGhfKHdiV
oKK6bZhcBL4BQktSYLOZux9s8dVf46LJTJ5SzaJEbf6zOy+nRWH97zwhoGUuFCHmlnRr7XUTY4jO
pA48ASIpbbbe8QrsI+7JP3TKs5cwzUsSA2VynrJwpi13i1AU6GNk+3nid+EgA6wmSfCVWaIrj6vQ
68s5ZfVIFqAJr99avwRB8gklaArNSlBxrfaAHcWgQwly0hhyXvyzxzIUD1HK6grQZBy8dr7SYEU+
i1eMX+iK3z9A3A1cACDwx8LR5GIyEXlSp6+YuuFQd2imDDZohAh5NER4hDFI6CTMKSTdN/Yj93cY
XfXhEqOAb0faQ1a2YxF4yzWALTMfOPyQq5Rjlb4V8eXCINmYZnpsazPOfQ8E0ZXKlIHtXlPF0tU9
ezLuXNk5nLBtqmgq4ARU5d8bGVVGXWOzctKeAeOLgM5xPNAkrSS0pZtKjRXMZhBiwdG3UMpQIYn8
vrDWBPdg2C9BFLW2KYO6Iwm+12XJJ1dL8zP15ziA0IeyA+ytrV+ZWyYKf1P2e5moSYvwEryuC1gy
o24/8IylNxYf9LZcQe4hvZ8cmBf1hMUYPt2LdEOEE3e8EbscU4Jb/fSAYxYxWjavhC4te3sGe5SV
uLRLfUsI6i4Bp8HK9WJ0QSfUwYEg/7bhkk4Dl8r/epKNKZnZ2NmrLjtRlMBiwkKorAcHN29KzCI8
PysxXc260/Z+mhxtMB3vhAq3BvGZZ7IQtE501Q1P/bPHWsYNfYieUh+FBPlCPTSClNAYHvOztXc2
QgsliXkPkjf1GErJOgv2APSzKoEct1xJwb/lKVdW0wwruxXI669AK8tP3jn9pZdjn52opzmjpsgX
Ui/3TjEKrjfMGhpVTBdkFToP1qkXlZcIUB1aK6fF0WVBChE+LTBULknOLfHSJcMnnXiPta5JGWf8
yplYETFLBVRaJLo3hndj3lso5XdjPgExu69ijDtuEcUJDW5fJRjwOtW8DdktQBBo8+zr8imC4Lvg
Gc9ym2UHSJxsN4QUtf7b2obW3TcEmXFWQ3suiM5fd7uj5yXYoRYbN9/dDzWSYXiWz1ltjaoagLhF
QJKFCnvQMVbiZFevDoxPi2dELtXZ0A2agleSyuvyan55ZyNIRZyaBZ4qfCOMwoN2it9szAfuU3ok
4zroemHdL0oVAMAcuiOAY5s18wRADH67ho+TEAQkJwUQrJA5af2J6kInp2P2U2YcP5PjMCsCnBSW
8pVkrB1PZaqCBcJhq/Nw2cQAhbmfXQZs3Z31ZWeYUAIh6BLtTNmt8/AFLksChmT2SZHMxhsR7a62
S+ODyJxIeAXqDQFGUc2wxCG9VIlNDJ1JX4NfPvo/8SvU+aHi6UgWw+22Kq1zJdzRZj5gaTVktp7j
G+rpvT33tPDtgkVatnMejQpYCfXMg9TmokuyQVdjR8VZg5JS/q/YP/FIZa7EMhYGeQtM1D968DgM
teZ2RiZzvoluvGcqAVMRCD389vVGvwRhNAuLumTrV3b86U6mTFWdw0oLyHYkiI6PKeWKPcTXZxRx
3SRnm5IZa+GEApQs7b1UcTHpyvDvV1+mlnLTembL3y3xW8mZ/2hO2IAs5NA9FlLOoWlHnDsf7p2F
TusC6ASiyIODZo+SSJbSa/+U+75ICWNk9rdckXpqlQGzGvwOiBVNDrzoNiYB2B8/nGOGc1KnKyou
C1tn8AULEw8EmiQsaIiMKOjs8afR6UdpXo/iXKPMbAZP4oVK7EJYD9LW4F1DPo6yXJKIODw1mRMq
OwL2ZY2HHVMDiIvozrLrtCfNNbGhdU32SCszdhFExrQV6MaWFmWukHzslDh4Q+IjmyvdYu7sFZdr
IOFuf+FF7puBCTtjtHBdI3xcXfjEZtuv+mxF4wNjdtZ/zhdM16dQsn5xSlmvy/PvLk/4PeCiwMom
RGvL7zcnHyKyhGpXXk78Sfu9ltmDoZ7w9diMH5yqCD9L5dm99umkG19qThftkC+AzOuYjwwu7i0f
6hAhSMm/No4Tzkk5UP2km16gJyWBj8plhy/cE8bDm/roVHXuI574NxR8gIqfVRXVRnrGT9uF2RZC
Mn+Y3wLnVxFHpifFtJfTpPXxcmNtQo7f4hHQF9+nfekZQJk+Noe48cRCGOLBOwO+8xHHnH6dJ80p
DQeb59jitcdFryfwA8whmwzGVFqlSkJSucE9kCKXIR6K5GmRvcz01eYzyDbhZcUZVL4dXrkDWfvz
T1vqvxICgUJa2FX2uQ78nsJwB7611vXr0geRyYGb014hkqCnB5FEkQ3nfG4Wbsy7XaM+Y+RFMB/R
rzfZH+tsyOy7frOJJS53BaHhyZed5aU4qwcOEfdpwXuD4CmfPXZZDl5ZAsYwg2RP+ebnauKZmZBN
WfeDFP1KtlilCwAzBx/DxcamGrmnsdLOOpLEy4O/oR+ZcFLnlLX8qbW5ypdBJVG8huNFwbPt1sCu
ixSEC+mTBc5Gd2bcPq91wqFKvwQPVV9fPOcI2jobvjO56bRpYpHiNmMz19yupTNb6O8vYPs2kFcG
XdQwXtQQq2xJYhMe6BBqBvUUH/VRBXl9iOxI1A0ST4KFGLzGjRgWU4CkpGTziAYx9Z9wvwUXoPry
h2kNg1otko2vsPpaKOqUlqVsCXtJkBTDy6tP7oZ5p/kXuWOlXDr1kagko6vzFHiDyb9GNHrn12gA
KlyIXw8G1UhE8nGtoYvJC1WBjlvsLM+R+RxOpv70WZQTV7lhhT2WdVKJIA/5/hblLnaB/jjvAd0/
Lp/2sdhI1O3yRnuFRe8S6TRQdMPPEU/FF+KZTJ58w8HPyTMf/HwMf6ZyOm2qM3M97n41iioxKUAm
k8VF6rEbMTk7suacSSJ5nkz+QkcqcU+mOry83BDS8xY/f7Ux+fYQoQh2UVa8XGbMYZmUCffNuOEt
a294VmhnxntlNkxQPK0he8Zg1N4iLPijs0DVup/nc4G5YYfSvs5dHMf8NanN7UfVGi7DqxtfoB+Z
N0TTdEETusHuqxnQYk3TcyAM3ET+zW2RKBLUwqrp6x5YspfUJzMQHin5ehUU91vPZPbTXi9Nssdd
KyNRnMU8Z6TOdTPDRtfUhEZVv1r3w5h6NNQZQRrbRbr9tBw/rEAhvUqGCiOBJGOY3Jiz5vdbOGrV
I5sgWeuFTMvt1MBfWk9j8cDbF5cXBg126M8qnxzlA2ZEqGWDWW7dcj1aWDubS6jUVxVvgFDlN6mt
4Qsup/UvJwD0m2oKhHeL3zoZ+1li7bkLY27XxSq5eCLLvDbHt5DGYjcKXAcRzLm/RiG+ERUSS5l4
GTL9PXBpTLfm+ohJdNBqsjSntOFtW03hBZmQD9u6Q+mQQ9GBap3lLOEDV+BydCcZzdddha4n7+ih
N2pqMplvAv2Ac7PW5PHBKoGmfRVE/BcvnMlShLSuLgKRT4W8hXhwndpfBBtBPTrfBzG+7rhWCfhK
71ocZzwpCPTvigCNUY/eCYqws/af5wNLhPrMIG51dXySdBlGJDV6N40xCpO5m1eQlVIUFtVif8dY
qCDT4+qDlp9dCTDwfZLRiWy4ho5PljFTEJ69yMt9jhms3cx4jVlSvjVF975iX6jVFrn5aKksCVYf
DFsqi7DgtjJ24enhdn8TiPMM+v/FIk/I07cJDkdD8RAch6q3UuxaiC2UszY9IoycWtStcDo0OYn3
1YHN5JXIJZRr6Jbj+gBByVPgLsdr7d6NDfFIQ6h3EJ1P9ObWMPiqGnlbZRWFByXKro7plQQWJm/u
gBjPdE0ubjwEqTqGN0IEPY8j89GJY1AiH1ee2WvVKca9TEV37pi0o8XF6pk/BRwbjfPpNp0+AKIA
sMEx47aFip0A/SDUO/BYxG+DZHRdIpDeCZcnoEVpaOZN/BfXiTmQTLBq8syBtmeP9oUa2Qm6fYYB
z1Wdkuw6QcNKjp0HofBZQt7HKcjSPHc8OTrukzHYD/F9z0/o53cbpqewMaem4ynf65K4LP0QlwYp
41q2QVmvUFsBjgpkNbQBAp1oxHU1zZspDAIm/PnMvmtzgNinuLcQy6hUp3quuQcmwDLdyaGV0wwj
V0rHLiA/8QABX+tSKq5wsz+wHVeT4BfDxw40pR4kBUjftAFxtr8Ra8X8j5c1vvcbAodcOnrsi9yi
aGzJe2AmVcavdmar4Iwj0bk3bmbCXzOL8/I4pEH+LX1UTE7ErRiJUiCg1aaHjvqaU1dJCNa6POmf
YPdEM4ioRknU7/wy1YxGIkWslPY5rFKGIcuBIzQUb6YnqE1f6cxh5v74r7ogdHX8qWcF2dCPuVVi
rn/UXjgd/GdmiaqR47/P5Tk6Y+4FGziUiJEh+/i+RE+nOdKFc9u8c0w4YsK7t2Ikw//j5DUPaq0T
YTZSEu/x2HokfoSvXHsBiJQmN0PscqN0twJJAZCrVEMFWrOS/jRj1uoOPbu6cZxXzv3bqzC9b2oK
lhEy5R7dKKLpwbR1Zzf3kj7c/QPveepqN56LzabdmSbB03ZIoBKyt6uTsiMgbyKmQFpbLmtsu2v2
5Trkn0T7WKXTVsdW4d1AKrGTR1wAUVWvHnKmH+02AxSe0PGvBw6ldTpeQoCUkI9R3EF8NLltySIA
nzMfh82Wufr+blTxvfXYtq2KtHimKRMrla1+MFFmNh6cLTdw4YR5aA3vhau0nq14OyTdfKG60R0L
PFFwcSs1yJj9apnSDiOaPUnsNwzMH4+kJY/sJ41svC5aHgpYlQvcm5dBeEiNEmnsr/EFkWkKEaB9
XZCSQnFtjFGBoSvtE8ArX0fM660xHAetNn6pvGw3HvQ60sY6Y4Y4Lq2bGfC6J4Te0xsH++QqmY4A
MU/wBIOWKoNlNTYLUpfRP8D8EdNU3KODD79SIzddXhdPxJQllV69P+sNRRIkOgAdBchtUTXe+o4g
2wkiYzJBBwmavosHPSukynX3ZRBcch0kPQ7KwzZAKV1PV9RCOaZkhD13jpERqLduygqeNiOBNDGM
j0Q0y8MMSM1TzeQbGMO1r/YhgTFn072gTC9eKmVRssZVvnK0rwnwLj+SxoDCdJJjKhr2o0ndSczi
rB7K12IzEMm7XVjBV9Xvt4pV3N348Ik90Ctiqqpt8AvsBZjlNo+v0FTIVvBXnn5EaSzNdgKXLg62
18LhAam8JdOON/QKA7yfG+yUyAkQlbVddKhhQhzrozNyIR89wCiLS18p/4OFwmwZC4mXYLP0gPeL
opYJNOKV3i52u/p1jxj89vSE5sEMe2bojWuFuvfSvhT3P9CyhPo17BcDpTPEWoCCnEqVSm1oXbK2
0HvglHZR164BHgWSZ84dKnREdxvixPqRY1aPP1x4UCYiClsfby20+fQB/+b8E0iJOSN4M1YAuPqb
3I9rqKrLkjncPq80jCIr4hBqcOTlfo6QbFijUwhFv/PMbQ5lfLfkbDB0zHYGLoEiawLjzCe1vDkm
kV1W6Wo08hwBYugLZ5uV1rLqcjq0+3gkv8kFCS+vgVws96gToBt0wqiCTh4J83ysbCJHrCe9f+FD
mCiB5qHxS7DdSHLSTV8XDwD88hmIsn/jLsA7WED+K0CK0xdOovvvXI25sTOI2SyHLDgbd14yLeci
pfoKPcluc0eWa1/s46xqpM4mKlLk/LW8a4b2Nc+h54tOayOy4uJwd/m9KfA/OdQOczHg5W+zi2yW
68s6gBwiW1voAeCdoWH8CQH/f+BF9oahSJhEqVybRinOAXNwtNERHmu+Z6IN3O4h7OXVInLEYpP2
p0CoEBcFbQxZWowPdl11h41SyhLz8R/jLfPD5XX0S6dBClkWpOEOd9cTPNYgUiu0mnFtK0ZobNHL
QIWIyJzOcN47dxhTQbhwIoKAVQT4FkZQ0BVGsTizwGG5Fv9h67/2St5W9NMO5j7n0hM5RjGhl3kM
MTR+H7YJaUWqi1KNhQ60QOhXt0YcKDiOY9C6eyBPxuA7Y80C1Z68ax+z1dGkh9RnnSHlwCdE4Ch4
oizGaMxHmw91q136jg2c8yX12nm95iSAhV3xbDbUXzuYWUlx7zu1XYpBilSF1q4eguvOaiqM9HDL
87+XBHaTT/zr01GLtpsKPHMmRhTSyQHxdvi04zb0UBkLI8akv4Sp9NdsZKWlC93pH/zN8je4Aaku
JIn/nGh5ehkAqJseI26+4U20iXudo4myDif3H7O0bbptNYTPvpZECYV0761TCfSfapnPDqyNmm8Q
rYXobz9AUnjIEx2wyjb3zv3yR0VysIleuNmxWlMLNJOycsTnnIX5aje/BmjRA7a3cCWIvifuDw9a
i0goqzf9M8kUWHgWeL+iSWtjDwR1vO3E34iYx8goG1qaxcyuQs3dVcZlBS2RohyyQMNWozSMJaH7
rnB+tCx84wKnnyU34GJ+mGAcEUYX7j3MXFjhZlTPRjanAQhlwpmLd8LHouBMHAFjhSdYaoel9sHs
jLT8LptWWmInMyEoIlzx8Ka9qoePDuEO8vxeVivomYjgM7xYW9Rgu21YE3VbAUpyz8wSFzMC+kCT
fcK/Isfjl+ThZMxyXJsC7CbufdCvnN5FkNoLhfVs4K8SZ6NmqBW3yUc3WHBEv0hZhUrv+NpebdQU
4mYtJFo4/rs6GOkEIPccMWr6qY7vwI7fmulVYKkNg+it6UfYF98CXsa94pqt3/61+2Efd4ukIC1/
PkK4nDhIuZhRRcIA33OwKZw0JnxS8ZTxwaNMfPy1WAO1/a5RIOf7D4xXJNzMvGP7slevfJFm5OGT
bhOY6hFvzAwOMaREKCxds53rVCPWY1XF3fkWqVtWZ2tIfAGkMiMsFtTsxThfgUKsIbfp48BaNReE
XEIIIGKjgebYzqfGF7LcM1CHt7DXUWc/82inhkUaHMfDLTH5F8Wm3vmBcX9FNKLY98R033zJ3t+K
LAxSyTDJ5r4pmo0OBlLbBOzlla/2wn94YSlKHcuUPCAP8Ih7X/Z3PMRD0e3Lp4uYO+/S+RChuLqH
WuxHGf49bX0l0wmfEB+7o4h0qwW1dmi6G4d75VT3sjQNwOdl4MT3KWVRI9TKlT+Bs91CS5AhHRBA
Cuju+fWEBxm6iw647NctHHO1aUi1T9ag90deyrK65xPCY8ObRr3Txb7oT4qjnYdfLztRlPmW+kLp
MVSJ88GaiT2Fq4h4KcfqmpdMQuyECVmTlKpGKcoeXPU2DBhjTjLz1Xihn4BdW5n2atFfZxabNgzV
uq4jUjXaEg0pcH9BO9skHoaR4Um0+swoGDO5mneYzvm/Ldr8cRmCKf0gEnR205/VcSvATizIKhDI
oChZBkTMLxiplDOr65uDIq45MNnlFxv9c//jKdOMIfU3PxX0pSpyaJolHHeqY3bVPnNPGy7qP1dJ
1IdDoE1Zyl8GWGwAwfWAssolmZYYv4jEA9TAmiv3yNlQVItZ4aWYD1hzUL8Fa9LkKVlrt0gx1PEx
hiMk3/0poENMmJWR7EHfpDwx00nvVgecFJT/jFGYsF6KFTY7Wmsms5IhSFaGlmEhfnlcEycbg+b3
0tolx05KkkK25DN2KDqWW4HCwaIOyD2UbBFmpvXMvUqr29gmf2Xzcfmm0Ikn6/mSGf1qWViu8iAm
JXZuwr+bLXcVmiP5TUShvfgxdRqaRYjRIec5QPspgQzV69XsS48kmTq90zsnnFwusS6J6y1tN845
6ktqB2+6YH12CZRwfXIbrlZwTZQoKAqJO9Z9VEUGOxJbBRpMOxzHwn3PbA2xz4M6Qo+grluFg3F9
6AaG5Qg+m1aGo2TkELqgaKGD9DIBi6pszToIU+cEit8JbSSLfDiKD0YGYULKDL9BVFFXlyRqjoiG
0cK5sPPXnfnCershIH5NIoal96zHVtsZslhnNH9VetuEgUfGPEvhnmuoOVU5KK1c2r9E8O1bZwcQ
I2I4quHHIhYJ6mqacNoWwFYt1B8b5qnhmPnWoR5AziaElhJvwZZEqQOUR4RA7bzWqF7So4UYON+9
KOA8Tfy8/+rFBmd4lU5ANhaNDFxiabbTQdmlyepyhMDG+g1N8nqZqIbOQwcYRaFeJJR3QitarGm5
H7fpcedpSXQGskkSpb41Q07X9UgpblWboTanJHdHfMcfu4cCBaYxULCFQaiUKO0KBJFoesGkOa+B
erVagSofDXrVJhqhiFgtaJ8rXG1jbohebVqAmosaezjARuk2AeBA3u1qgETNxyHuHsupKtOVCqNF
suIYVDQ/iEd11edrLkg0P/VhRHzm5ztW21F2YnAwElcN5arJBOPUoGcbEkloGs+ZEZE0v8KUJqVX
giz0VXDhkT0BoCsnCr14yEIFerz96jI5tGtWMv/d339f4U+7gdRaHsbpqdM6TkcSAB8o3udXebgm
EII1VruTNG2V+Auy1rTeaeak/nDKSHjy+zYcOAyVFJJ81zEtPTFt9YTbi3O/XSsUA48RY42wj0db
NJsd4ErbS+79++cafdMoCRnTUtA3JciqAfxf24i6WMVXFvpzzHJV79OVDO7k9Y4aqQ5bZ494B+t+
GNg2jvHIIDxqU204JYGLFGpGg0shYJRAYqVRVXOC2udfGTHmgxL2Nu04ZusB46JP/ETsOnYJb0FF
8XgCCjohOo0jtF8Dmo62m91TGSqqFE9PJkSLAHBc1MivLs8K/cdUfj9PcwSWH/YFKDC4h7VMbxGO
dojDnF0Ibe9zmcihWPoMVSGroVaaP61g5cs49eL9gbbMJyxeNyb8/FBpA0uiyxRpj5xHt6Kvvs+D
Yp2ujZNe8khSroZZRZM7247CF3YXPAZpl+37bj5J3Z0T8M3vvQAtekLVQunKjKjFSYeNuOVL9ufW
dKtfKbcjhDmlJw1QSREpgqbafY2v92ej2VU6bbG2VMknP5TEoMLGgbNrDiAvQIslSlk9SSwgEmQK
xFTgPY65XP6uR1llNfx/nPOY/zsCzdOjqvhg03t5UiAl/THNmgT307Q3cuRTddTokymRtI5VEnP+
94AXqbbczEWMv0sLqRrcFhhGr2WpB/aHjZbubGj1nhQIQ7FjYJ2O6698TzYykJM7dC3inJuect5E
dB4Nid7QQq0IE7Kdp1qfEEjqjE/gWFhJ1AICMqJfRVJnBvF8MuAdKDrZLF6LePYAjae6baGVX8GV
76CsWj1zjKw6GHR1zgQL/+cGgYX4E1ZAiaBcjqKa5LZdsevUfBRIapf562/3aNiScZJCfPhtQ+mz
hxE3z4ACPeql0KKpwAaH1Gl3PIs3lkumcfz3wtA3NBRvl/RY1dt4EuhDGaIsSQvc+XnPaF/X0nw0
/mdEMP8paddVmamt/kXvgBAa/3cCyULk0s0GJEjAmxx4LKVst/pL7Py41EHmxbix/q9Jyt99Jdur
IGrurLDp2LfNyWbU26w5/fOD1BagVujaNh70RSTtS/WhUNctBi5KX4GmIyw07ZDOumHZIWBjOFlL
bbpNSZW81Sb7YT7hNSzqFFKo/5JQxT9MPHarI0cVU3FZ94Mo4Q6S8d9+J9lbPIj5MgPApH/X97Bn
ULwut5URjsKdYmHIhAXNr5c50fckywHM4fe2oDD6tb+qqWFJBeeHTLSgPpQpMfC6cI44J7Qulcni
RNB5FiVRUc69lcL/JnHkorSbKSfBCVTO/IvFUW9k4wne76P5MrDULYzZA4YmFCR7eE+Lan/OWvHd
U++7RFYXsoxFw0hauXFe5ZTTcOWS/cWVrTDlWXtETiBNk+BZfef8iVEA8oAEnHeOTpyXfzn4PsVv
5Uixv9+GQS0+Nozn5YWN0jn5I1l4LazqGhBiimEjR7tRzbX8PNFekTIPGapFw45FkQIKkqj8jctO
6+GK8ivifAYim4/9IL9sf+SmFdqC3VEHA1rwXPL2v7EKLA6M6WAGIE98O/PifXDqVtMLT9icoZcn
Cii+eapzZ0Lc1yCKG38FPLwcBe7Z9O3UE6t4Dgi4VdaOO/MtLMa8ALvkp+2xSleFrP65Tft+5Mf3
qsedfqJ8I8OU5W6reOACpPL7C7FHedVigSnJ6U4h7dQ+aCj1Ua7zoMLKqsPwd2danB8mfOZQBUAZ
ksPw/6Laodb+I9wDWRfN3W5RVGsB97e14HuF+TIVe5k517+rW9oB64BPlhlEfE0UlqvjhUuZvm9N
rqKHMoEGqgjfPKFZU7SXsYmPxfwlZzBVC1AqpVcNRF/yhLSUNlOdkbPNnDj25l3ArOX9skfBY/Hy
mrJTQCV4ha3Ye7OvmpWWJpoNxLnJVVpJjCtC/VSGU8qZhahOgPPs/6BKU/KJTI3dNljUU2g0IUjB
bNTPfoV7vfGHR/Q0y4Ito1v0JtmZ1E9iMD8ZOZHYRhQuP2oR/XSsrgdu1j4inqj2xor1RjN2t9yR
fCBo8xUyH2nsq0jTcjVPvLfVHoO5XqLH5jIhyujrDmNLz6OJGtZ3RvaRQoYLmapZyeQQOOKjbQ+8
U8Gu6DQteVvxrpWvAysf9GZmHhjGO0BrahOfqkbp4Ik2bcLWFe6XsyfNhvODjsLua4krzDPBBqsr
useK4iaKSVkzjLrryorePz90aLCf5LYEHXCntRI9ymw+eZZJF/J93LH1pPr8Y4/ErpFHXZsLvBLt
XrdM6IlbbLnUMag1EswgtVZJw6G+AP8VJ5dVYXCnJbJv4HihMMPfc5/X1+9FwDvPiVlpkPO9+y79
j6qCptowagq8N25NRRDNoWTKxnrxCF6d3p3bC/4WnefVgqx3Zrg7XuHnXQ1RgOH+awE0qZJ8uRTP
HuCcOgEcG2gRDzA6M2DSo7ZmWzVMvJrlLq3HAXv/WoMcy08pLdk0XQ9cf75nxjxW8JRlqOK28oP3
XmJWG5O10OFa7045ghAhzsLqdTEzRcQ790vBWmgPZ1zDfxhKy8mqcoaM5FbT7cTrMM/dpKHc1g0t
9BgNulEd303y1k2q6QucHohhbjy4UbKm/YxwYCy2b5U2DCuP+OJv/xpJtpSmFtzEEySvhFjcFukw
jLFKQM7RKFQMlgDnjouNVsrKSAlttmjm3sJxxusRpokdrOKUoIx1Hj1/pxgbh9KEUTrUCXpy70/y
lUjU7lJMW6qy/Hh3md0yE2Kr5SlskawW8/G3uHdC/m0E93tnhV2OmHiosOJ4g9fGL1mRNHE/Pw/4
2uLFIF/ceiQnEi6KQ2FF89lgPwvf3J/r21U5jE2b9TrTqQZh0fta8yEfevyCUgZzdfo2vF5RIbeq
dScphWvY7VpUFS8UzCLtbvS8Jdh1c3eT3Q1g1D+GOszWfanARCM/mXW06svvbpmHfvRCGgCmyNwE
h+TZIOfLXm+HTeTW8N9KXlbzA9uyulJiA9AkecoTEFeauKZtihJnm4E3r41qOW4OB3aZHUX+x3Kd
jDT0ABzqTjPfqrypekdo75yL8r9fZcu1F/BOWpoZd4sM6VtMPSAmywZUUIQ/m/eb93w9qJYGOY9n
hhfWhOBPjqDTlCvcXXvd8+ZBnmMT95Kou21sYmaW12XjApaRJw4B77EkjvzcUdePc55aIDExjQhS
6Ltgajf79d5XmFcBmQHGETgXGTWAusZDdCWtyyN82a3nb1+tPdjTQtVnET8w7PRSynWYLbMvTnwg
pEHRJmHDWd8A/JFFvNOJ/3HLGNfAEe1Z3yR93lrr+wOZ2jb7jej2WzJPO1Egsqxqlv4fVUC1m6SF
Sx0ucEtMFyUUSo7hj5Bea68TLyHZUdcdjIT3AhJoVipBkLn1THuKIlRMWW3y1KGljzqOHdiR3B1C
9h2u6B25qcODiBze9ksY3qyCLOKiXKmbVrw6MctegLiFGmDsMRuEzkVAg63gMPmeA/nhBRY3SHXK
3gWNMd4LMZ9rueYvWyfZy8l/ZwbatpV+3sCoIaC8IB6CmTEmvb6ApR+h+KzflWJSxhJmepL2y1eD
F4RP/JxmMSSzq+uoXjxZ1/H3s19nSei5uWXHV+Ec8hhthb4jmSM8xMMqiY3Jm4k85y8eZgBXhDfk
82DWdrh3zqXwRVUHlYlEqbwXmBb92kHEzIUzD93b9SKf1LNbEUJqo+g1HIDD5aGIm8Bi9gYVAS0C
hCjTxUEEOXyIouW8XC2gKT92fNHpD5F6452MAoVWzZ+mDFZH+qKVYFr/05PtWprWoktPvrJdtA6k
oq3Rvvosge0dXmWR4/SqnIhBVnNK44m5v+A6dQAobOSyWsc0gKKfdV05uWvHEcIqx9UciKyjgbXS
RDHyruFeexKl01JdAJPBbM+d2wYSK33maoVd3H5Dev7Mp13hrbPhghVVsJK44ymu8tWCksVauTwx
YHDvhzu4Zj/nHILPKBcE37A9H4GSQAdGqSocHqJF/b+uEB13r5bvWpkHJo5AxKcK8Z6T6+NPW1xf
P8YEubLuWihl+w5HD1dQ2g0M7AH+xuf+4XEU39+TtuyWZqtndlr/fsA4u2ka5PBDLzurMk0qQ6Nw
sf6dcpDXbz5aY7G31+7RaSgkwoiJmRixXuJLCQzCBjyBg+Hjm08kzMJ4qeTmWg8FGhQyX/gPbAjZ
E9EOabdmr8REZsrXSo+l2SE9J7SqG63Dp1h9UgGtmfbZtDemiRBIF8M2pXZNYTNX0XTXRMP+s4vH
M/tulbScvRklqhR7N81zRU+yGWod4l69MlDS5R+FPphQnoCkwenblkJfmF1Z0x66hZWy16DlnaL6
liM+dsAAgWl9vGzuE8K2XTCZAcIprlIr/Nx0hQuGKN4bhBquq2cIxgCLj6WTqGa0xeYyNFkWkFsp
DIeLkhpMMsMUQp+2VhEeGWxcjyUINJ/dttG98hdZQAF4bLmILvcMwMZVynG1ZI6ey3WQzJjK+40K
Dz3fA1NAVSgF+lQvr5poNsAYIPtJpLzfsdKlpsGz1WUtq86KqvfB+NtOh6vdhG4WUf0AvK3AW7RC
d8ZtA2zxQYDs7nNtKT5oACI2o3d30Fm7V1pBntg+RRe+fiobwI4BMMO8D+6eQjZaqbwIm1yZ3Ts5
oIkOtBhYOBUK1hPPOML0Y2FzXAbEF1gTSaZHxhRRzyxMmBaaNSDjpmIF/IS0A7n4SG94Sgg2OBjU
ClW+Byn0KcVUCNop8xBAI2j7yNqNIBkKaat/mfFAnZPqEo7jXsF4300HY8g68Rp7m2zRCIEsIZ9E
poORckz9nbYxIa/QzSbk99OY93SpBkAl0htwBXChFxujf2ymQoBCbVXmkWYGTEXTpevAna2Jvy2I
+rZK34lFE/+tu2wDcte01KILfsFuRFcLzybAPXx6YdLLYMQS3Z6y+4mk+S3Yo2afzjf+Z2lw9ykS
WfywYMyA/vMiZCY80qNGU1DlnEZ4c3GP2yEl6Y9MMyEe+gM4qQ0QIDuAQp6mIZFFigW/0VnAVlJo
gb3XXQuMxxaxtkzDYa0lRGvGKMmVIzkrlCZKME+C7XnZZBmEFcMgEJBjL8IVpuU5OMyw4ogl/Qd4
SAM0sOvBNjbLxHczhM3pnyEyVhEqJdYjF8GVF/bS6zpMZpveYNU3zlsfG8r8pi1Frm4bF1c+E4ZD
Ufvj/DP1KULF37ZxRYOEnuC9Nx5nCFcDCDgxpUVkcw5uiTwz/xz3A586M2OSWH2/EI66rQM1kMxZ
TjKBm8lgy0OUpcRtLMzHYpf+A149Zl4t+sAaQ3ytZ8oIqRpvpDyIC/5ka5VLhZZzgAGwHfEzVSg5
QBXeY2ePfEHg7UB9XG3mMYDpKHgV1TR0f/sfQM2UrKAfopmBeYIGZJym85AY3J1GID3ZYKRXg4IT
XOoZ+sfkGMI76nxaavfoO89uqOWIcC9qW6RyGw3kEAdhnlYFTiXJbmEqLCR4eRq9zDYjKqZqAEuC
7jSHWNutVc5PHU/bfRlq7JQaHRpZtDaeTMhbpoG5APYoVnAEbegWFbl7d72YBh5obfSGFOE5PGXi
i+C6133kflTawfH1fW3nIJJCopDJRUhjwrL20mVzmazF9T48h83EV7ov88fOH0gkPQYultnar9JL
kAtVMRVq4DI6bQuKMMMkSTz7jDH2krDvM2Qa2YwqaD0G/8iLFvH1kJpty5VwkcyL7oQeJY2CJDHs
EwVV6izuXnZvcGOb1CiYJBWScVYqoSuZFJZGkDfuLV/ONwP2nJ8Cacz+wIKUSyAXnYTz0N2rHK0X
/7tH/odrmNPy5PhNSCyLzsLw4NNE1ZcvQj0GGWDLaEi0ODo/ThyOXxZa0pjtF9KDmm0+50GhbPUB
IeTJ7o+0/T56chR5/bnatxXTWNqW6gsQn8e4G71SH+eXwWKFBzzNaHhhH1a2SkyAVkYc9CMWBpHp
IYwGu71eJFojFpAZVxGTdGL+IcZLsde0X09OLtQ3BpYwR5WO9U08dVEZplqfoy0xrrboQY4uYptM
tylwhXutr4YUi/ZyaMHjiZKdr2J8yIIto/SQvvBpyfQjqa/woAb/koQY3DSCyfdAJiCiSK+rIE++
K5yH+Z7u0D8FPNlBiyeCWN+VIZk6KIZeR0FS9/BNE/eDZ70g+KfVkOEdzZer2H/zQsBeRCxxeTzh
+G5x6PlX7uxh8FrN6Ja9+jBAtLI7Ug5WQHx6B2/mXZXqhMf/E+2Jjz0PnLDgdBFttAiWkVqz4qYw
CE7LHJWydaEAnCoMyOsNmGzjzSNiao51Vd6Qdwr/gY+G9OZgHD6HQHn9OIObhQkUW8ugHF1eVRO7
D0X8TNXmhshynB6jSb90kAw9z+VDthl1AMOk+u+2yMUAisSm9SYuNwsu6cBYKRJg9pRtSmjtOqa9
aDXdS61ENqhxpLpomOZ1Ea/IuXLyOWaFVKA0kHVShV6w5TTuMCpN+Fh/9Mc6yhgg2MiNz6n9huUt
sv7IYbLKL6qGiMmNERq4YnfqDp/OeQA3gvQ48ky3BoeCmiqEkpZqEpl43rLRMqoP504J7rgPCbQi
2PFd/iri3Q0Jcp9xY/TlYdcKhv6mYR2ntWATXOtln39TxSdJQLdf8J6tE4kXc/vS66E0mRSuFQi9
T/VdadCP0+Zu4tA53yfkouDKCz3l12A1ouNXmKnC8qRbyxgsaAjM/wHw7z7vTwwUnx5v/WN+WNkT
q/5LblCc65cVpgGfYrAfPfMNPEJQNDPw+a99iF9djXA38LGEYSAKJocgNTBIxtG9drFzcSeFGGd+
AHJMYRRlwlHQ6hRCyjXD7w5gNK/ovgQ5LdpBStLXqPhSrENeBle74bVzWgiCtgNzPqKhjKW5HPht
co6f74nqRQRnQA/dCNOPLBUPV2DR8scYWSGdjE7uc+U9tbUdIq7t7vz8QW/dfDUz+ePlJgSaXmXp
AUd6yqnFMxMMCSKRMPqajyyyZHlfn2fry/TVsdxbl4AvNubaz9DTchHEvhJzGvREWHDVJ2wSGpZH
mPUw8bq0vsmZVFAtJTnPFFuuZhPXQxZTsnEFQIIzWGITloav+Ib22HymxG1mpsVWmoM9QoxL0JoM
QLBYzUn9YZg+MdonpjoILdHtxdwMGMzOPbavnbMeOJG/8dJjojlc4OoapoQBsStLoejC8A7nqCl0
ceSlOXcEjp49nGkNQ/S6YKPYomKOuSHMWpfEcIC5kvn5bJsikTTkzSZ7nM377ePeVQZMCMN4OYPa
8+8LnMS7DX6snegD86g/0fp5BMM1xaKc5bh2amD5Lf0i8XPDLJr1kOEQjud3b/K6R4pZh2onWWED
fA8JmOiBokhmKpEQw8IkpSCOWdjm/zNbA7ylKhBfGR3UgyV126P0yfle4XqsGcEhqE6lDZS0x0wV
NdHlF5ZgnEyoRcliwssWF50psVQcBmUmsFicTCBM3hjpEl80cHBv5CxlURZvfTYdPdsUzzHNGvZj
bUGYs/4/uS6PB9NUrfWzyRvsenT1i3SgkEl0kQ0JOOwGIu0U/s/6yhvT+UcGlfd0vS0ZmYdF9SHN
kENVTH6ywkcK1L4vem+8vlJhaSfhfCvC2+r2vAQFVS0QLWoC0bNyNrDAnF5//9WKvR4wF5RMWL9G
Zlv9YDdYZNwoy8+CpQKIHPU6EVVkOXznLPejcEMt84Aih55zJNJe6P5pF3q+QmPMJid6g1Lq+z/L
tz0BctnR+2aHXMVTGB55K9AIEDd3bEse6tnn3tpvn53qKFHTj5aRCNJMvwCGiZiVpzQDCcDL0Y1O
WOVAX3eRLtVIbLRESChup+sktXrkV/XtpASjuNkqjIlEOYf9AQ4Uw4qNk0+3XygWmdQ7bOoaai0v
cUqXSXP2xWb7OY3bHkPCiRJMYvS1pcCWgDmeB2+Z/1+WS7gHAsu1t8NZ3UK9KNgzRWAzQpt4QKz9
PHlNGnx8LLhThVsDxC6dTB0nTM70hRaTzazBiZKffAQnjVYKv4W23T8WpX8yqnziuNQdSN4J7toX
mlEiPqRYHlrlkVrJ53CIB40sRb5QM/bOFXQ4ahl+fayfbFz18I0ce/OHfjZRePhz60Jm/HhkBXiB
JWT4IG4W9voVL8Q0dcZS5+UFBC6mP2eSFWm8tQItUUfnw6yn0JcJaa/CcLpW4t15ZUHwRV5dF3/B
CmMBfGOOrEOmZDARNLrdsQI5ZIU5C6vreb0XM7XNDTwsW41NPjPBd3rYv5liFAHnsEv/garzLB2D
Q8ulvPND862WUWU/ji6RuwSvheGli4hpDcmxruK8YSl7ecks2JZaBNAFElM56t7JJvtYIDy25DF7
o5qbHUobGF2CkZdo1gzzwGUnqWpSOhI85t4Hl+hHZ6ZjZC4bMu+JVuDWV38bWJLiAQzWXjfSvEZ2
jDlVCZoV+CySxnTUuqDiIZDjCEFLzK8i998YoimY3pFEd1l9AyXNdNPhJ7aUnwskeC7mezQfMoe4
VJP6XlRN0MAJ8+kozwDWjDugU7zJITYR5Ne1eooliz3xCllUr+Nt4rCUEDgwYiKV+qVFki9FBq94
gOsq0xBAIznAxX5QRmVIEtXoBIHf1zAzRAR85b1vM8U8gAMLfLy4l9hD2HWuAuclXhhIEKuHTaQD
KP9pPAz5K1iCBQrfIZcE7sAB1rO5tB0XuaJIarGQcsfWPxX39xH5X2VlW6zOTWhJX6ssPYQnOcnp
CZ6f7N7VBebnev22y67fRdfCqfy08qJG+BW08/ibvlPWW5I94r0AVcmD7TXjz3/J5egqIrB6YV7h
Tdy8VWs7SKgjfgg3GDfplX8yJlgzypp7QHkNu2ZzJJX7JRjWNt+GPj7ovxXXT3chu4zQS8TqyRMo
VMjlDc8G0ACye9YXdFVumI+muWGYtKP+ONx9HoTDWl1VfLAIYe3QfvDZOZqctwNm/bF8/iI50HqJ
vcQh5L3lenxy7lCMOx8AX4gOqlh08f7ijCRFf2gM2QVE03vu29iv/scRI98ryNT+0iqo/aO2RUbC
XXYff/lv5iM3s1olUuF3ip93pH4UbG+x8r8fw6xn6KltgTKHKD2It+BSMDGpGo9CDZf6UIvtgWIi
loYTf8rGw0EX/aY/tBMt/MORxM4SHq8pzmJ7vRppVxkp/4gtH+UFAe0dC+F4Ccwb06mph92gWJYK
OuF4rqJ4dV/CU8K4PC6DP5u0bZ/ROtHecb9vbZ7iCUUKCEzCbNaII+SkVDKlRQdZs0rHaBauCrio
Oo70hMaLFEatU3bLx8PiEvIgriBdrtvSbcY0RP3l7UqV6C115svmaPe+CRcB1fh1+IyGN/cbk9jR
/NPgZABF+LmFde42W3Dvg1S76VdgzCS9PnTuYmc40iLonq1Tg0Xe+E9GzYl3Q1n06iHDNiQ9Wv6c
aASSAqiAVud2qDUiGGprxY32FFIp9/lEwi6IhRHdio25bXQhT2rzRgf5OgyHzF/AyOGfyj/bB0e2
8anTIRQRZMkiM1uiKD3zDoEKljoF/F5K++hZpWTWXPe9sOW6AhZDX7+0/NVO5WTmRAcGJAZ4jSTw
LO4sLQ89USkWOQYBmN1tQZzqK4O/EwTq5m/tNOrdkrgWFxPDoePWyLX9eGVFCZqm9DiLNEk9Rx5Z
nGyPb2+mDsqMA1vrHOgNI31OQI3WhFHh+1MvGlIX99AjL2kiYFiSWBXk/XXmHeHVLw97bji71uRB
6SmW6CxM8Hl0xUkYio24P3ay1Ew1y0nrgJHRBMdAPpMAT85dlt7OfsXyw5AxNaEgGpQOIvHzoJTm
J7n+x/n1PV50N24+lMe7fJe68genGT4bBvf64L3P0diIBwWsrlT7Y/1/Ud3sk8ZSGgGDL/c+ZgmE
GZfTvHLSPbx33LQlCcckLYyvbPCOFFbxOArriqMIBxjspTx5yrUjEGMBjgQ9iRW08yXOpZWRoMzn
eeagjjj/Xos4lksa+hqd926ibjyFUbQzXfyWV9G6B/fAegrlVl0wyAsAKlgWQVCz1ZYEJbGi0LY6
8LG/pGPqXin5ON/+NMf9yJjepk9CSxjf4q0w4T+ObQ2FCVjHWlkzIsvKWuTFUaeZ1h4XUgwn9kcY
13np4eE/o2Aq5AWgVcfJGiiw81K94tiroiH3z5nE3TyAG0SIk0GoKRq5XluNai7QkOTxK2WbiNGe
Q37fLgXs/RN+uAK20QNWCROEZ3m7WkuSPYf9FXtnmvHAQF8nXxe2Xfg9jA+Y3/qDc3xkLUGaXxto
j7tBeGJS2TQbJ/KnrlEQAnsLPMhtc3/Kpg7Ul6jBZ2NFLrWz4/NamHbj/Q4VYo5UzktxMxjH+efi
x3iXftKck1wMb+qMugBfi9OoDxw3w4xMUb/JSDjKXNLbycmfk+aRFqXSiimQgLaC3MXH0b8PBvUV
g5wkp52SZvBXpvg3pJunof0A2qt9XRBOgfOHHsCt/hb6lazl4e1WCdoW7NNqXup8UOKRMN4R9CbK
t8eP8MTZkjJEuc+WtxkXLsFceP5plVhcgu22IVAsWn0w2DeG3XBzJp7xrBhWyLUefkkAMxwYEpzt
uh0fQfVlZiKZ5ecq6U1IUudG/8cJPk6vBOFKfKhbXDJ4XTa3LgXY943rCbIwYS3hpuWy1O7y0L2g
GLyWEQby/W7JkUj5N+dJFtjjzBvOaJV00NPFpzybP0tFxvxGWZghArMXV3SzbgPbnWcs4O6bzsvA
630YKpQ/sPs8Frd052d/zsotq+xYdVPvPV1h9k8oOfsIpftwP/L3T6D3E1TFnp3/sp0nPYeHHyLm
WVwjlauMd5+qMpWMaZxdgIOeOpcXXrUjboapVwzZxhjHv31/xYvmTy5FX0oDV1VCutNcKD0r2g7c
BIfKXX1y7itGw1xHGrcrr8KttqIM+Hlv7i79U9KKyfRJ1VamQIER1b1TAR9DrJXtBJfmuy1KaWv1
Iet3oSDsc3FGg09ka3Atbt8v0zh9m0RGhKrshDngaMiZ2epiETLvnYUwpT39Q/LynhVv7w2GtUlg
hORu541mZ5lLeCrzS+k+nMyrhmKl84dO/muFiYcbW1xE6esF7WPtvrUXuK/W5BPxAXks3TKYwmI9
GjkakUSuXEZTuH/kdzqpBXB+cC0YUe+Ynp+D+UOeStt3TD25bWRhfahBUH7foQrenzibuc6w0p77
BAQTcD2pDyyzTwpD8Nw+fBr61wJ386LGuu+6u643HRXk++tZV1b7UJVwwFHh3tj24EyhN3R+eji0
Jisw7Cc1KZgzzFn+e2rnzH4Xlk8Fg8j2YyQdWtSuF88CHjMK8x7POo4gX1WtiAvTYdFTChsNSJp2
eApjMG1wnunF4WMBpMHXnI8mFrY8YmgBDSoyq4xlTD238NwobTpiK3T+cXT4FpBjomihIpLnstc9
93sEPMiLBMz2kdctHOFsJpNbXaZVRFT2BoDGaNCdqpz2qAHba8B7gqIkP1C6tkt/T7Jmoobm8hS2
zlw3a6tEqaQmqDcI5INRx923sctxIAthCLZUiCsFsJ9Okw1vie4ySO7DTvRGYbI1yswMJPq1EIx8
DvjayLXATNfRm7xR03ZaITY/WwIsZouUakXy4shvjboUoNK6H4YI3hk+T7PZkr3K0v44dXIul35j
vbrlAnQwVTSJ0+uyamXEIDfF9eeIl2yLuEu1yEonfecnhmIymkjqbc6sui3e9UspLSebM02xd7Ea
XqmFqlstCBnHPdY8SQYJc9iBkx1pqYwp0abUk8gmJgz9YHyRf+0sCL6zIACO2TeixYjjq/op121g
XjouR2oCgom3/hYLZtOUiNVr63eKVHwBzOyiSYaPkDaHumMKCu332/ygSb+U5KQV3MHUNpwCcPNL
9UvscfKXoXP4TEO851Z52QB8tzzXGzB1G8x1Ty7Ft/opO113D7+jGe3SPEguoT/Op1prcPJ4wuQs
xZepWte7hSBnkdqEFsdH/C0Mpgs7MNSgDzAWsDSr58oMg8XiABaGuWPQQIT1wLj2ZdCIW+N/5d/q
yHOJGWsXHm3n4oB7WDezzxCpZ3nOZxDaUnTs7PirNPBQyy/CMs25WFnyDkn7Jwm9xG6U4mvi/EZU
k8ir6n2yoGFKMbF2A8eT7w5pGWrbMh2osq2eQ5UQLkQVujzQDigZ9oztXvRmVbd1/wPYpu2XVBfZ
ErX4ofopG+Gj3frxRUXJF7tI9crwiL8S4CWQ2RYlsrrix+ULbrzgO74We2J0jA4ABouY2KulH0PX
469Q7u5aZfra/ywXDUpuQVlQvbfVWxTfWp548JSiIcKuIRxlZcXNE0dqXi88MV+ZL5tz9ktA8SFK
Z3mUn76G2czAAsmWYoO1yqnpVD8fRmLhoVF5z70sBYCAUe21unbcBYAV7dIKVW8CoB088k/bCTvd
CKuWgTcfrfW/09pEXPpkHBkYWjfKq+KMb87EpyWWyXRGaA3XsJICu7J6L0z+DW4WW1u3qnq3cQ7t
YAad3a06FtuKB+NXTExhPKMHXT682k1GPNsJmnVuFWVUJmpt94Mg7az+6X8Hi3xTvWTX8XyHTmB8
LzroGObSl80y+XKzF19LjO04orpGyt4irtE4CYSPeGOnRAu+YE+r/hUXOFnbd/BkyYpOKi0gZRA0
4vf6YHQWvcwd3gvXbwLaeuoWNxbEpW1dyzsjXdl9EnXcqMjqI8kJC9ENg6uqdXfOoKrG1FY5+uCe
UcrcYwgO/eEv5vyQIde60+yRHyi2cV7DThBi/qxBLxfUujxp1ee+b4XMrHXiiQ/t1bzEbWRZQmZ1
zeWV9REIDxo1B7fGJrHxTg1pRMxULv3EJNrZPtJo7N0w8+wucnrcmRYpLzjeE5OgFVj05Q0han06
c94bb6usHLAtuPhMVk+zGTCF83f3delvilMan4b9w9vPN0b3Ha5fHpO7aPrAplLqzhDQCnHK+UKe
Tgm2ucbY9uJCyvk3AQbC0K1895k2CGv2DLWaEDVfASfeeJWOh4qC2wk+FPZsJoZwCrdOaUGAbg2g
i57HOkesnT646MYSKp+su45l9NOoTEIweJ3y1gp950Hw4dK1x7oW+JvWC3vHef5a41ZCu+caRrUD
qYqIQvresYs11xuJ+6bvhcpApx/7qmaJFfkhiesdOTNLZBcMEy6BDr/u9MZ/zaxozLFMeqKWBqF/
pS/FgIMi1Wf1AnFc2cZX5DYp4ZGqh7/R+ChENZKJJ+J2GAWssSONB4fK8A2q/avmk4MUFGgDRbCo
1NPzxvxX9HEGX1B+pIGXkT5roHvVNuFA5AIwG0OB+s8iOsygkDfVHvfjus5MzCoVjDNPrNHcphsh
SeknJN1gC6Veu+JnL9qwup9Sf1L7VtpgFbkHkmhZ0FtSOP1GqzoB3DeH3c7R5wAVzwjPdjpNDWgY
f9+t2lhDa2cdfqjqFLG0BPCWep/+E2aWV5nxrybad75bEBhuYrd60SJG+nXXygnFhF8SNEPPhq9K
cuzDGowFyXya2lIQ3HnYfDODkHVx80CItWPnQlJODd0ZJaA2QY/6yODjgKLxveZ6/b/sktvEHvcz
JLTO4nKJnwpXR5zcbiEg7myYKbCKaWSmuEXoGlL6blyPkzaBUsH5ya81RQB1oIflmrttE3me8U6K
UC6jEhX/scHgReh1tya0QpZzxULRPbwQNn55JFQ/PTzeFoE5+Fzf4IRH7yNgbDXwUPDfe039grDI
snD0Vzh/1moQI2x57l+1BdQ8+6L2rpM+rqYdnHhN+NLIlSMKboIFIKx6pT31aQp+DcGnWynxfqv7
1Ll3HhxDiMGyhfsHzJxn7E8ApyI2wvb6Y1pJGN80ScA65cbds2jthqLIUjwzTVZzAzc5RezygzWL
Ran6H/Kxe3XKWPbyC8k4C4dvsy/ENr+/uzyObHwEA8DE/dtCcVk1wO4kTQaGwUlHtBr55MZ/o/hQ
zM+sXqn/n7Dq4FZXWyvGZ27LhNe0AswIcL9769mkYRXsnkNwkb7J5i4iT7OPn1dlhSEBdPNH7xVr
reoYc539wtIVxDbTsD/M8r3IQx/cuh7ky0FuKVRjlUMy59PEnloHgdcP20Hf9rayLveGD51QG15q
oKo6FIhwdHycdt5bGUDy8BahFsVeN8wd0q3lleztwnWuOi9GXZPxM33BAyylr4KAQLrbTDOekN/B
k2Fa7Um/yQ2jlYNKCkx4tYovOI/CbKCS9InAWnCmBqJdelAZ82e7PXg1z4LJcqsRipA88+paXT/O
pFFU/4BiCWT4ELIA8hxqrb90m8a4VAJrZNYbNtMBjCtfBErsuYtcbQdIzwaM58tm8tKKYAdTPDpT
T0+uDWUvjsff4H2p4ByNaWAHYDegWIea5IvBXIL84UsNKSGEC5HKgi3aQw5f151TBhoJeHzA0vK8
xpJ1qmXd8QeU4Io0zhLsrx1+WeXEYx+OOAjowpjSRjwhHJsVnJlu6JHGD26kOftZ8GsgGPIYZl4J
RVFywTWhQfBF30uN6pb3DdnFCMhV0ccDVl+Nn6fvYTi/7BTCLVryr8Uhv0uXE8/1O1GTWdXNGSM+
eDXK+8oV9oc2Pmoe+5kC/WXSvugEMCW7x9G+6pFHBX+Et173uC1KQSn9Sg0ooUT4U3hxPlbQ1uV5
oEGdIx7rIDhGRHYtidmWS7j4h5Ha15JyR5qbEXKkYQTYLiNW5UKb4lID2CN/O+n0uOI8WETOURmP
6d+U45YqUZ6o8rSxlp6jHa2GPi/+1A/jZRGqIsstGrzI+DdtPLI40ufr/6FK1miObVb0UPXZ+G1M
UK+9PBizzkCznxVpAWBiSHmGVZQuLkiZmwc1T5Amszb+ffI41imZ/RAFzVkZ41ayxbBO293Ybd7x
AMMa4pdOopKv1YHghnWWChGcTEpeihsB1nnWczU64brOPobYrv1C3dub44iYiMlfimrApykqv/53
IM6xim20XmHxKrIEW4NIw99N18rDKydkdftawuwFlSwGsKcVJj+5ND501ddSCKpQJ/GN157I4MRD
ENmoj29F1PPCNl4642uIUGRSN5p8dmCA0d1m5D4HoqZVL38mZIfm8ucSEnmJM0m6uzP0AstjDlrg
vez4L29a946FOwhv9ozMCbMuqsQENOp3jFOfU7KgnF3KBklJ2EoOPhMG1imqAKmCHsYKfNMFAdNr
GT0qvcjcVxtqzI+QxAtUSzH5InKVWMoY8Z1K1gvFTM+ZGzn3upoui2Q0k911gjpjhtXKHbAsRVTT
QUrFJMJbqqEisXJP2qmFdXArZjBU9M/scqC7M9U6lnfE/PILQS93W3bUhqyiPwJ+icvXpJn2SxXC
uAIMRej02LrYHcM8ZZzx2AD65ELyAbftZsPtrpwYko51Ic3Px706/B60fHMusWK39J0syjP8bHxh
JM0VkCqQQFvfefoOt1BQZpOvlIRuIKHDVWcbbpxmc4y86SksnYJ/w/Ks9+QKAnUxFy4xLyP78I5J
JBxWwo425rpejcG0mWlQw/j3DC/6GymQPeTyiSmfAm/OVHZz4paROy/9ST43hHGC0995eKcW/9Bu
0aQe7cCibQN32VrmE7syWqCKhAQ60qMeUL8tRGGE7d6HPHTYz2wBVyfdNniI7935dE1w342MuPP+
dWVGeWKW2tXbSSIfFCHRV29kWdJRtDFoebMmR1dbPX1CaP1MLoyoWGzn0gP2ugBy4vhJFCTCbo+c
QrCH6mvBi5KNIoD2OgbYBB5oefFM32z/7tXxKT4u4ovUX/D/cZrbGVEEaww4zlkyi1dpcx4rPUQP
3WDPAP+vjSZQY/1DH8jmETzL3YyzIHZFLVmwLPBNcbN68iT4FhcyWaK1cYtKk4c8fAFu/8LS8T7S
oM7XXdjdoRIvkx/wW32DXsrkZ14CIxjD6rxOMvSic9aKNwTSraPeA2IjIZGuAxfpkmAqyMbP0UOM
eglmld6CY4gWgMg7kKjg9M8cErtABf01bOtj5O0eaAJZWznsYeTFnjaCOSDHEJ0O8FVGIPVWqw+l
8rYOcJfHV5lBKsplJg8n35KAySXEz94z5BqpunH7CBoVLFKYD/UKxTWHA49W6sT9xTCtXVChMEkE
5sMfHvat2bWSNlzWxBPAp7YeML9Ewdb9ARQI/+rU+U5u+On3NTXNQB/9hQL4s4DnDgbw/1pxoktk
qh3bkgqvZj65YIkajdFyD7Bptf+9OGdtvCyOy+IkLorqMBk5oDRSdKsJVIn0/Vyv7O9Y8yGmNbrd
UtflB1hBLdOi8t91m5BIIQaCDzwSfqEenXG+GLq3bToSHBMgW1Jwoz3DBR1YQETI9xzMUHW9Xb/O
osQabn8Cys9hxV1NhovxfM6LQXjjtcMM+9TsKg4P006mFzO3/9PWi8Us7gVfmO76FIKx7qU4mGo4
2XePPO11H5nKlOoCqLfuEK8G9MfbGt2XUbB5DP75LM/lgmaiOtw6vaXJJYTspAZW2HJZPRxHb1bW
9g0uPTJQAi2wnyHld1uS4rSECdVL0ZoYgg7/jkoBnNDOt+8pj7qrnK0iKqM0vIpbeHJ757qNk0JH
k64zOluhhiait7SqU/3i1vPJOPcg70q0YPhBLZFjWcT91pZ7UI+8y7fFI12Pqx1VbnIVHdQg52Ee
t7zt6ZiS8IDRzUwv3yrhX/wJDfTbKC8NWkKfgJMJTRpMnFcMHstFJ8H82rFG0fjjXu4j7jq9GqM6
mh8bPFA2o9Q3gtkN0x+VUYKPZVOryu7G4ru6wNoukx6Y6a4xrKW8sdS1h5uPfk0NJzhyh465/meL
I2MN8Hx8hKt0SIWwmNeQjX4d+n9Fjzv81/P32iZTHAro8aJ6NMPFEzu9JGulXGkTfrr6K1Zs8Y5+
PXivnFB9dvl1gR9mtqrBiU2P+ZIdSaV5GFRPTfHiSA0qR+5i0RXjrXHNV6SSW42GwnhahsHdD2vy
6ZTEc51LLnAlwhyz1/MiDaYR5UNsOFZQHKq4XJv1+EgR6FgJenVvlBX3Z8Cb7K01MnqjKZWoSwsM
ZB1CLJrRQE2QhxWIRRpOyvBTXHGy1O5Sgu8/zixBxvt0vwtH4sl7n/Jw9t0ZsyJzIk7LP+IyVmdX
VsI3z0/Ad6EWAUSLvYNl3o5GYHlrf9dWLxLEWtVrMaLAolb4585hwyKrwUViGqx3uOpeNIPrlf16
q4IK4MU3am3zcPaKX6hoxkL5fpNNvb5GNK5pqicb2tEzYQGfwhMiv0CwDoO1qIaJCm2hb816ZHCe
7eEbwehwn8pWbdU00AQoYTc9FNi1lvvZUkIBZv6qijPvUh5nbo6GUgd5vtUgcApiRcwuf4mpx/1B
0iZnYizFZw/tGbEYBZJro0X9AfrR/KawomJ6NTArwfHfJQtiBd0yi+bFRMtEPHU4EDklcy5zfclp
hpaM03Gsl4XWCr1LNRdyXNXb2iUIH236fQyoYvwDqpeJhnkkBb4Vbl+Cha65tGpXdOphQaEV/rI1
9XpovTVL3TLHlFUPtpz0wKp/nr7xP0Di2gsFp8M+yaJYR/0XJSRjA2TKLON6CNj+unSzNTIHG1+0
x9lNh+bTPPY7ShJE2WZYcHb2ASiyVPOhNlVvBKpLVB6ta5P2JfbWJO/VZqZ9t50mnMkzUh1WAEBA
U4t+lK7Q0qK1lho4mo+uWp+ZAPkWxSSsOg+2oMGyTLWX3T9RIaz8AB5dHfTnQebw2pd5CgcosPoj
wTmbIHaWZzSuv7efVtCozfUc/RsTEn8jtP/GDnR8pA0rXwzHyqpEuRs5PIiuusDPbK37wAar4aUI
5MX7r8UUvctQ++0QzZQNuFjexsNv0kq7/1An5L/cMK8HxOiOT7XmewWofsgup7V2hrke0NqtR/ad
PJTNW/SPL5mj049IgCxHRcwE1rsd2kMq2iB8zAbp9N6oZgkixPtMyurcKxoszLEenYIsPduQlcaZ
34mlBbjABb9U6HU5Tg2vj30vcpwQzSEtDM40VX8i+cZ1MQ0wYxZKbAKmj7/BVIPo5v5G+FrcTGsZ
WcMY+EfaZnycIyf8acho9wEyg17a3s4u1oaQ1BVjRIJZtmkzMnbXDS4q3uvKNR8NmhvB5gsSCbt+
gNTb/tsBnqS9yW9uXMOZDAFCvN6vUUkt7SgJsxNYe4JkYzAY4QurJVcjrejhLsxvAioeAO6FDFC+
PvV5XnO2aymAmIC9QJa/II9q+KuoRFSKI+5MDFpKn6i4uPXQ8UUmzIll64CY9kzEmu2XiXx+f1kc
yHbzhpdyol5XGvvWMXNAbTNjY49GxZSCf7E3xPP/bugTLtokGV4yZf/M+ZorjF9fDRHewnUOjnfG
OJH04qzqxeEy7YsZ3jMBqnp2MfUoYFlwypIjJvAeDRlyf51PzrVtpuRdqJErXCigj2Nnz6rjnvxJ
V7+HEPaa21S7VjQQM1muzt7JMyHdEHkPrmqO1TXeEj4TMuiCtCNPC5ftKip7Xmgx518WYfo/uFrz
dAQElUYgdbOGeZ+voPZ/HzHCEZ0WljnGN2cRuYKcbQOzKOu40nhcpBrzO2cL00cK5EdhsRd0rX6P
stLyNuoXg2DZHBdJCP1Rt3ctiruI70wEwZKKY8Mtb+Uuw6vHU+JwkPrKlxxQhhDrZZLu87Eiwmp6
8yLYE9/0KVtX2SRwt/y4ccWS5300Z7Y4Jpaz+Pzvl4ygWCbKiRxXsVfgkIjYbNBH0OKXYfkzMyAD
On4Ndj0Gd/ZImMi43wAFgnNxOD90C8BPK8LFti1sQwamVtBXZA/X7og+JXtdriuWP1gS/YRFXpFR
U9a8Rgh7eNxFS4a9WXJNQormcU8O6IFIEBtoYsMchlgH2LZCRqGNYGj+CdLX0IU5vvHqtpyq/OW4
6gMFiDnmJ05+MwV6i7FMczxezJPOTESGiEB0Yviasr2OD09eZwqZ81iSkP+nIUnS/l+JDp79o2J1
lOuAX91lYvXLasM6SKMy+s6DJOz473uLW43l8Ag49U18l23iErLZk+a0W+TikadNTK/HN5Pe9Dmt
OFkl81htGskTbNYxeWnfYiNB16WfBd8N40Ru5ihJN4tPj8P4ZyhFe5pnN0Pl/b2ZvZpRm/feqvBl
irjw/i6sCcfyEw6+5r54FgWcaHAvWoN8cMARC+DqUKLbDJ8Os9KfBGYGyfdzigZZ7LClo9O4vBMm
ITcAc0geZ3qB5lKeG2vOkpPTj+F7/B7Nmq9vpaSTmW/j2+QAH88htAJ8wBtpvVk38P2MCnx3UhUG
807d+wc/FFfGnw1zm6nWFFpW5cIcHSHiB06XmPMaGpq5NPIEmUl1qbl4luh5LdTvTmW0FGB2gOSK
aeRPH5fwX8YT1ifA4YJKuWJk3vps4IY2EEKbzs4kRLc/Bbyx2OaN9He+bhiHnpST2fGHBBZeLn1R
f46F/4Tof2aD1OC081kFlhEUsq9cQuvZ+GonDIdDzNeBiAWRbfgtaGD5tDW1uJNT6fLe3ayH9paj
FsmZSkxtYydIrn6Fy0OGDwN/nFTrPr1PLY71TY8xwxguaadVuKHVIqBYDCpZ7v4I2ptBVhy82gcx
2R4vY5nKjdM5NHGO6+cJsubCeVCI1NqnSzETybwKCLVaQKjE0tDGPSPDP7eP6K2WQZN5YMiwpnfp
SfCOHf7r/IZD58nDAxD14tQXErC6xlj2KjGYQCQuQBqY8ZPaEsr1fkbaPW6xTApj1I0ep12Y8w6W
q1XkSpYvZBGMOiE/h87qWgX7K/YfbcxfOwQS+OsXBpWJf06A/M32va/0+GhS6ZIuGlUSCV0KKiCn
4NsqyAnPKr1V6zQqvdEfnbIKRK6MTA6eV1xXLCK6jyLe94zsER1syZIiLnb8BQnRNXw7QdI940kR
mebjqoLPd7OtDv1H58qgys+JhszIAJDGsvscNPyRxlCkLmG6UkUDz+52ooSL8p5qOj3opOIAM+xF
JDQAhGrrlk4LFAx1TYdyCIardprkOjGiOxlXQDHeq+5nXJ7FolVEocXgMfwhJRdDGwDF3eEBk9Ix
yxPoIXR4vHFqsUWQEts21joqNZ8Oj96MMGk9B5HFOH2Z72cXTlQk8+SNjOiZwgjvW1RKtEfN1mpl
ikdYhs8eup8YVk4Y3dJs+8oOzGPSYTeY/Hp7CI/IxfqGDSw23CXzG4cbiDGlw3YHoq1xEge1B1s5
EX/rHfKVsV4j/KLdhv76iDUUbyJkT5/guQfEmWg0M2ZGX+Uv7dW7XTUFe10pdMvKpFWdUNFu5Nac
u6jjhP2/KtstZhdL5riUE4eFIWhvFy4H7SHOQ3TsRUDVEYCdLdhIQ4TS/3G0JP7Ls1SPuPevAwdZ
xnn0oCfU1dRdkjqKgEFx4JJhPA/wq14JSBAaFGgIDV6Sn1Wv1qc8dBPFZ5+1oLSVvU5n2hEpeXDU
wtU2NAFBE3GRSRFnW442XJw1iicao6E2lYj5ZIeR6YeVDYm4a5aTdQWNHhnfvEKS+Dsc2dFIYfq8
wOC1CTjNX8PE9NaLpTp7YZtwhLk3y6+pSG6qmWMAHKiTUuAlLosifHgzemXtGJdZw8lom8T2B6Bh
KGjWSnP3wuO0VO8U9iM9ldVQUyzWqxidYR7wi9f1wP9lFO/wVuGcvHzMB/jD8PD2Dgpf9rj8Bid7
W5AZOWo4sVma4K+P2beOR/zMHimlALlZXeSJTumy7bKMoClMEyrsC/FjH0UhZRpMaHjA6bjz4G8L
ZfjUWzemUgCH+afGYcA1mt2BklbS/HJlLyL5+yNsBuPX3VtYUhjjyKPO6QAb0LNFNZiT0L70O4YF
Ug3Eckrw/KuTXYbqnWDlBJ8+OcfsLOqnavKvuBN6Jt0ydLZ7BEKDwvn4o3CiwfMcFv65dYGKTVCm
Ba8L/IMy4ieMyULigIA0Qe+qoaNy3xx3SDxA2BDccFag+WiAqC7S0uDIsdG7Guse79pofFPpLp80
4uVUz72Wit5an51JUXMByu78of5MJs40XLvMZeGUCoPeflX355BxBMCEBF+OkBlmbxOddfKhSu55
2J5v2/Frn6w0HcwechcmaVtDo2buf6fcw46eSdGoSLlzKjl2oBqg1cpDc/WxhljgK5x/xZukObOV
kzK1QDez01L6lvKWoL+SX4ueWCDJlwDJiyRWG/s/rKdjZ59nmh+S4HOn7FVPsmJ3AUyIKWzE+qh2
7XU5+qzhEwuWs10VlOUD9T8ftqSR+HXNR4OGANfZZPa4Bq4HwPF7T31lVQqtBxEurjmvsWqN9rAK
I4YT7TIA0pmp3EdFZpwNSWgx6AJmzNAqu3um1CLeGEfxgzi8twuKkHqS0EiLoRb9nggrvlqWJRRC
JEmNFHO/125/3t0Sa1aX5LyQ8/+oyE6LXd5t/PzLOngsZs6f6uipnQzlTUwgaQmYlAckwLATyT6E
Pj0+EjgmKWk0vd/yCc7vaT0bJzH+8idlbxrfncmcHCdpVD/3s4flxe6HYzBZ/eUGo/pb8NzOTo6z
OD3ZTPoNDl3fznE9vjmxalxZsUmW6pOaLoggjKLiCGCLZbBs/0Fgj3C1Ggq8j6b/Ol7M4VnXuFgr
Q5INrreNJ1lrpH25aomE9VQxfZx+yhqjjRh45FSVmT+lmpC0lPAm67vO1jDJ+sK98ruir1xlMgUa
o0yNJ7EZNYubJ+1QUztIONd8TSrZ5DWae02YLltNcUXY2gIj3OWevpblWr3JZCiPcUK2AbmvrnTA
MxBYRzDuJZNLSc/15brhSsra8O/kZlFsAKfrzekwiNkrPZYxanITMMZuNdP3tbhhz5nJfVZYQk1U
bmCfmVcW4Emg/G7Ueq9pXYg+7E/88S6q9zbRQhkZave/0tWoSc2HzQIIwHzRVIyArcB77x3ndO07
ckM4XD4mxEx7JPK8MUg/XhOWAEaKapWV1ieOQIDTb3yjkuXiR0V88aG139bqoX2E5v/SaT7XVrJk
PW69LYI7L6kjM7OH3ToIC2fAOF2/5R5hu5RB5b/WqQFB3PEMJ6NN5fRJjY0gPitJI1iJSZdGZIIw
vwa5YqAc7IMmV9Bm+cz/4sYo2/5wUrGMrqcdZkPBMGa4ajcwpJUyE/M70pxGKQBkUaHX8jZA06eA
v0qro1RcXoRVjIUqhEyRHqKLnnxMVIG+1g2DqQXuPSIDgShIaM76IB73sSsQ+cvWmRtROl2HrECT
LD1o0lPYSWda4+n5gcsCd23VZ4VAPHtKKsbkM3RJNlI+q4jzrb2xS3+z5YkALFK6ZGiVtuZS06Vg
TnClsYUxUTTIA8WfHQEXVh2PNaquHP1TeOTZi1/6rpEwHgARRT5/h7nBVW8bZ0vWqBlSq+mAkSsK
Z5yZ8YgBoW+mosBsqIpQwvGC5OcxXgzZYPHz20Uq/DyhXNiv3fjDhfERXEgcIqKXYilvHjZPIG4e
KyVzwgORpQvGNpHrft6Y7rqXPERYZDJ0wMt+XJ6Nwk/2zP3yl2MPRKnTqOWLRkWBMRBC3vu0/O2Y
I3ntjDm/jAQDe4ohFcFIxlqtW9I/mQ4m48aoathG6CGD2NcWtMO5Rg9f681bIghhzW0Nv4hutQiJ
XVDdfXZcwSaeM7U1uGxjss8gO7mmYPhq2xDuKSYRqM6YMjQQA4rdMIbSnYY9i+3VNF06tpSckLG6
O6S+1FRLUUpsIoum1puxJcjzPFFtiXlitViiZNoV/QK/hGZ7DxX1Qo3rOOEa55JjBkrijy8Omb5u
nGL7EmjUmfssvS7GdaVuSba0JBn/cGxNkLbUJf7ydCnheTc6+oqFEqBixiNqXLfYug3jAu6ERVlT
RjrRQULlx/4XaVZ3CjOi35W44CcP4M27Bzty+OD1Pvv197M1/X8c6DcXa6/JVfQ+enM3PtMK11l4
GWYLQzmu8aknYrxX2U70ujqmcUO4DHaqM+iSK9SJSh7RjSxfU36/1WeT7rhgHjtxamGlKqlsASWU
fJ1C/yv9HEh6+A2MzxMUjLzUV4PzMgU6WdlYRj3/B36wY1Xc2NClIMd5uk6LzhG1ssekuMTc3SL1
VcOVK8TYhbYHEzuehQLBAn9fdmHipckLwfLTZLa1todQkn73lTK2aI8X+PVi9a4AQbNiPoOx/2AA
KPkLN1fpJxcjco9u5+ZGoqzu4vDSzx85Ozpl6H1y6P4xSF5k3a3TEa/3YMS6zdOpjeMUTDlkwH2X
Xa6LK9SOwjmphyU+xz/ZyWD+MMDfn8UTRjLEgMIzy1Zanyu4eP1LYmYCCUpGxWgDcRdQyW5Zvj1T
UtPzHiQpLII9OGihYrYWS4mncAX4wqhqj+lDlTaMLJrS4QPkOrzJClQysrFNF0dC/eNoGbHd10rp
SMF+YsawwGGXr8EymVJ8fwiuqNpbFsdYQ9vn+Y3crdYc2DEVJRk5sDSFv5VfGye9fINkQjOzUNMu
xBrFf5zuc9c3cdqGC3ogRqWe1EKUkwuXf7VAlRgazS21WPCfVJ8VSspExNepH+B29sbU3Q8Nc0/u
kuyxM3TLNnu9zid/Wg8tgOpm1Hdk1sBbZ9RJeh4gs5yds4ds0pEepx3uW4epNPBRZGOOS1M4ZXhO
Al59zr7CHPxu6p6n0iRg8KPPJRgyRZQ7AmHzk0JgyF6TvuVv5GPW6XZTfXtiBq1fsBzQXxYo9UxC
qqcIsckAKiqgQvEdmJ0uMIn5/w+Vn9imNfYjCgzF6U6IkEC5HGZJpOsfEGstgAHzu2BkgpAMJ4Nl
snZaJiysQkGoGJnCHMh6GZQGZnYkWnaVhAMSDJTuI8rc/RXIbj0ESxFZPKNHtQPuCrzwBNhFwG51
jg0O4m9HpvKCFGYLwbfFXaRxXfUCPKtpPnHdgCd5GqrqrYXcrzsfYCntk14xZ5rw5hYTmzAmc2Uj
01C755V+z5Zcg6nYtqrisVHnzEk0zkTzoe+wUL+v684mWSMDOXZcUMtNgIoFbpRA/VqDfHSfwwaA
mSrlxfR/Ooka8srfh64DSkLSdts3Vtq2o1zFb/AxSHDElf8JAi1KFtifjWZuc++pEBitoXtUvqDm
5t6A4CHk4CIK5QMaBolhGHOShMjU4P1/0ytFG7VYlK2uQJwZqgWq3GGI5VNhH+oywMpladcBOQYX
1rkj17WEPYKiVIw3NuV9SxONQxWRrmDyTsX9DODDsy9tUqjngyOmP8ZBli67OYb5KoewNpGuscui
Xh1i7FwGxXYCk4Fst6zDcx7xU9SjRrU7LtFnQHqd0wZiJ9rc5k+IVOprsblwCyBZcpLKL7IHzU9C
+wC4fdObKGN+GZ7tDjlOp9OH0tKlCLDh1kkeWjozTstYewq1uYCLAi3XS0ZNPlAgy1Lw0aNJapyq
YTGD2QzXK3HOmtr4e3gCCrGVBjDpwGElF9YYtSwtBfJ4se1iLZ8OE/5LHcBcFye2BeJE/AaqhNt+
zykq0jG87Jo6DjsS+668lJqvUC7QHxrByuK4EaomXsVPsSoET3TJ3aWl43H23PIDtTa9LVQLYbv+
a2rdTc+gtct0dZgGgSi+FeXfVgWVRXsZAZPl+LqDox9ySe3orXshDVJzVJe7eyBYkZRu6eZ3J5mF
9ZwKKIjoYGy0NdOE9QnJDEoPzLPfLug9F27ViFXr2fe/vgM6w/3JCFZ17tspNT/6eqjMw+HmmKJb
qhTx3JnlDHzEXdWQSZ5mz0tBMrzq19A8Xagq5P1I8H8Va6h+E+Z5nCttkxtrJCe8ciAz1F7WQd0S
y5/lJeNfwWEQ5tI18OzPriRS8jUUj8sQJdxd7iXxhSCBMIPB49EKCKH3vqgc+1OZN7C0M2jLG4zR
IEZTtQ/kSKL24e/5XSiDmQjwxgx8/KrWPJbOqDTVE4bysARKw9sSnfrOgq6kElZnLajY9w2hXNP9
YAHhTv10oeL8Ge2/zubJZzi52pz+o4qtcegdVTvEvFDXn0Chx/Kx2hHlCgo8DbGrPSFAaMlAPPCc
H/IpTywuq118/MTjKW/Qmmo0dx69Nv7l4Tf91ehKTvWd6aM54o2xcnUEiyaaNCzUZDC9BE8YOQMM
h2M5BMPHw/iLUGYWbvpNx/tpXLn0hcKHKDYwBNL21YT+yQJEu0K8IOsxAdGR+a/zza91taGITcgH
fZSV32Mcl8f42nhpTdaBy6moVpvO5Avo4zpL6jMAWVj9oQjMiFYOq9fblHSE3ok5vAM+IJ1kalCD
p24ZQI+zQdN+XvY+EshmYZpy76wHxnn/+OefnBdGzYTczYLG0JEM2lnza1c1ziTtNbaPAXmwoSDX
2DrWWmsEVkNcaKk2afJcS2STy1cW3uhsxhiqHylW9EoGExACMXeEAminSAaEdHScPxj2WI2DzuNV
mGtOjx1+4gVxARoyhsmiefqEpZ+a/dO/F50b4shAXo4kSDYmFW/xaKEEAxGlXYq+7+3wSVGtUUjr
wzZbJV2l7N/NBFSEOV6pcONvzmmK39fsPqQUFyHkDHZIso08Kz4cmrRhe41GtWNebabFr9BO0rEV
r1UAsx2JyAUqtSdDBhGQz0cIce9VHszRREPWHjOvmFtLq7QnLaKFlOAtscT/UG3wOHRKAfHdV1nm
sdUBdQYMaR24/NFODzB1lGgrIyYioWg5KOGWwQQCxqcU2LrWU0Toiqjbn9GT7BkPUvjxViXWesbA
eNLk4t8ZcAemYHPaOf3L+yEkLikqufsiv4ATWFn9V+///ecDTL/clxOO1yx1asW0sR7MfSwgjsPY
jAJaWqlUEFmmmN9sW9snZy8LSLKIIi16FdzzE7k6HapmW09d7BwrpiCVNmQjzGbK5YNt5YqL2WHy
nir/hsmKL6oSbLoodzxsQqSy9JCiPVroOIWwUHUFvrexaa5uekOU9WBeeXQVCDCWOgsuYrGEROZJ
OjFsdfipmph9nUeTYSpHyj7n+c15nrwm/j8x8hI0u6kWQhXvFZV0x+L/CrCHZ0tc08mgcmkl5gsk
lL5SpXrB/oGWl5r2CEI5b2SYwHUY9arv+zpcTGJKmOxYU0AAYHdj5IVLuawan0liYDUHq+m6zQXR
TVyy4N3urBJqBDaon1mBskQq+gAEAIg71HeQGOpnnJC3QTD6hEnfyAym6Dg+S85YuEhZzM27u801
MIuxMiP04qV04kbmSAoueX2vS75j8Rct1uzLH+BJD/JwyuDgpLe+0aTfxDE3T/7QrTPU+gZUNw00
JfhsxrOIFhXxnVJGP53YowmEkH4wY5NpZ7jBJdplfo+ZoAfb+3UdEVqSQSwgEnXvYZUGrUHStMdr
uHDfYm1SGKUCHMyF7L3Dk1OiXv3v8cgs87uyuMgtmrmsfQabihku4I0Aw2XOv75vTmnYHbzLlo+g
rSkbAyJSKTj6yg1h4azBFkqYAPIsfwfTAjqkgEC8QocHsXVgq0MH5jmBqm2cSQJdygJ2I+ZqT+PH
Cvf7bEGr9ZyS5aHc+v30/UOB8clJujOsjtFONXWfoxbauJVVVKxDd4L6FRSOaZyDzdNVYOAe1b3W
aKmwufCDw0ENLoPQEpKVkUwyA0BUy7hvU14l0EWU/Z8AtujD4M0qooJpp+88/XmAj9t7RaJgYThf
F1nAk+awDpD2rWTcELQTSfLzOGnaqMOaUO05XnRswmEJrLIBJ6gtuzcCquPBLC1F3+dYlwufR3He
cyyYQ57KHZniMYjIUV+ZEluFE2tW4DIO3GUCUIGWcGWcDvk3PzjNVlqg+5n9cQH1YiD3i7h3RaHt
/siSAR0rf3dkvN8rdkxMc/rKUEtXx1OjkkkwPWmuwFCfvgHtHe9zeJ/m2Hxrv8l5fXzIiDr+OJv5
SBEuRdML1Zp4S0IXWpDcVglX/ikLD/RYYNQqZkLA+kQJdTk8YG3Y4uosZd9PDiR7To2xQXErFlDa
vKlfHDWOIdt8BJTkwPNSMsdnaYEeoaHzgYbrCCPZqmuXHyC85qrOVIJHpTF753N3DjoW0w/6LafQ
bubibBXCpLNXffu5koQbGhTFGF5Lqikb19/nDkIy9h7AOaWojrQ2odeRKAiZXlaWw92IE3keQCTm
1hjB0poMOqgrsrsGAvTlbf2OrWi9WIWupfMNXjjMpCfHlz+U67QJ0VuZRb/b6p7SCiae8OGuvlaM
QkXlaNov2+5ntD936T5oWKNwClJx33IEwQh2IJjKbtYZ8/RD8oJpZG4musTZFqBJppdRrSejJa9U
FsGRME2n/5/dIQNTmiCnS5xZOXbUwG52U1NMasWKiAY+11XtWULYNpqZz4B4uV9BtjwGSDHJvItr
YojG/WDnv96fxCViep3APMfNyQbRQ11ZiwoFu7Asflgl//ZZhD0xixDMLYGrBJi9xMRW+8dp+9kX
v4XQpw1PLwh63BWVZBFuQ9SU9IXjXUT1VIOBtS06cFJom3dK13vE7cbzWAwwgwn1gqL3njtNe3bM
0vYIkhPAp86i7y5JQK/VM9Xllcdy4nkwvfqZGOgsR01fpi1irPogHnwPKrer6mzuA5/k45I7AOgH
jI4WN5KRevklRTrkPDnoV+vmpeWI07UVy0/ueg/PORJCTSM+hyU2AD5ZaXkjRYKAGuLFL0nbIGNg
J2P8lfYBAYa5vekZbNRAW8ARuTFNtki4aYjUsNhjZarK7tpW3msFVBFizIFlgLgrArw7mUl6/4MV
tm2hwdxvqa0P3ycJ8eYe9Z0Sun2lAr+bjpjlDlYRyj3mzWxU7hAmnpYcHs+IZpHsYjiaPzCWT2e3
UANyBQJwn26vVnHME5bLUvC84/UCtbVTWJqy9xWFQWlFdvtxvD70wTxddWCAIbJiEJpKnkpktjRJ
OJ1aK7cnlhWVW0rUWZEW+6cZLpJAO6sJzFcs0EkXNNP1r8te7qPB6oiEqrxt69HByntjQJuKKGkI
+W1vyApMJ9TpNrgnE8uyovf3aK+LB9+H4o/KEVbBk43AMJCwp4zGJO5YzS3YN/i8YqO8dOZWVIZp
6TYTvHRLM4umtx6FCCWHTy7IL0EbQYZevm6wEgJukoBTJi3L8392XxzfIf/zCfqny151gQ8sicP9
UzR/q9Lsko2VtLUmFD36gdf1eoLU7Iw2rd4er3e5zuPSLB1dDrmECjB3gtIyupNOEaGBveiFDAXN
1mgbi6Gt8ztg/LIt/iHSSVbbjIK6NTvXy4m7sznOOkeU39/oKCdH5Nb7RuZsXkcFiE1L1K/rAg1e
JzA+Qgwo8Piz+R4fAurHLPKTPmeGVajQ1RTwvP5/i5Ve6L1RZIjCUKOmQ3pQtdvsdIjlqb9YEbWJ
AMft2G4A78Jr39PmdrK7wWBXeMRB0zcZgfOjwdlu+aBCnoqY6YmAI3UxgL1zvyMXmdL3C7qQ/OfL
mjtcgWcujVXzGO2iINr0IPavuZMm2kXID5gHShbxw2V3D+sxMPIvjRt20uJYnMDpIA4+vEvDcz0c
Md8ftH5kd9bYlHBEjXqU4jWJeS+u/fXwzFp+nBspPSSdfnCte3Z/hfQFGpzI+Hxg0Dutsarl9rzO
qZIEJIELfFJIHNhkK2s8JiURjqla9Ha3DWBHP8acRFs8Sxzmxi3xSXz3hVsAsO5AdRvtkWyPd16+
nXVFEt6HIhTaUz8SOYyZALY4kGIw+o+rOGBTVNS8bakkEcJj2cxWg3uck9o04mAv8wwybFjdctwn
98d4KrHMDpQj9a6z3cvzjbGxB1k8gCHyP6vo3Fg6j+IjAmgkNEtlGpZhURLotTBgaHqPY05Dxu1i
8QR+ZBuK2SlMlDJhIVHawtuUvWtm3KnU5yAmUpWetFEfH5FSdYGe0PiT2tZGSV5bvsJLJ+P4gEig
fQVR0Vg3oWn1wO5JW2uDbUtnKDxRBdU70bRg9huYglIo6MARNXTdbhktdps2cyQQRytypW5EOf+2
6XWk8X4DKn1/ZRymcZoij1tft4VTyiwOEvfEACwCvaoNZ+1s0RvpX6VJRxsbfelCZAhdqJ1LeWqY
oMwm/jbPc2qPtDTpjKS/bMvw9Q/W92XFJA8j83tEx4fw11GzMr0gbZ/epdbK+CTv6NA/jGzg/Pxx
uulBMZQJCmy7trw4/AdGv6NutAQ6//I7OTPGFc3Gkdr9LMznL6GlCB+VBo0opi6im3yKuUoCDpEU
JXGJRLAVHjEoJY7GXsop2yE5fEC/T++ZB97GKjawK66LXSXkrJD5RUnvnDkRAANCP0MJxtI9jqBY
0rexfA48+Vahrju/MKQWVWYnZ7EtDPKdJ41Lzj6XG9H54xfND2SJju8h7Q+7xl2sJ6uq/IBpjIXn
iI50kTAwGhUFpqU+lEqyIDbv2+Zj+EXugLeFCklRsQWdrQgeYCUQFA8O2i9p+8ZxBphgJ/6LgSvW
3hZjAPwrVQaeCxIilPWLbxudGUx2D35o/6SisYfUX64MQQnQgZI+CHIZ62RzyFJZ8vDyAugG/Zi0
VPW5exVrgDf0giBpZ/2SrPQYIc6CzhzHhUzgwif0D2ppxNxt4hyDlH3vVTTsU8NZZho+6pkxmuqP
uuvxVjHt/oSNz6Rd1xYd56GpX/mUhKZ/HzIagGb78vmnfDTdcUQ/ktrLsEOctWJzBeXofKYPSeqq
Y8bjHZq91SxRLBlxuUk7G+NG1ZJZeXMxlbJPMhTnc0j1k6F1l2YYHn0WiEhHvWF5xbRKaGjd/dYp
f5qBbD96hFRKamCKQpEqRnzPT07+dMAi/ql84S45MUBzfS92McO0o5MjNR8+qBl42IY9b3Xe2/xd
NkTfnWNVbP7fyP/ibHoobmzfsA7ZFt6weNpoOBR+u0Urbh89nF//zJjhYmoCmQjiXgsxkpa7bC1v
gXj+vHvlDtSMryDIS8E6p3MwKkTAIa1ZhQ818o1pQxsVdL4V8EBu6PAIBZQ/6jvZrqxfT7buKO/l
yC0AzWieonip1kELbhERGSOgzPhgehxaZ6V0vd6C5NmQXUmiEF3CYpb3Tl/iZHYsV3lGkNdIaMbt
wIObLi78Rh0kI9t+zStcQlpzQnyl4EEt1pG6hDqittQ8MoA+nqL8rR2VlWNvXN5/+rrGlB0tE00p
Xtig1BRfnLcp0bZIwQL9kh7Tc3ec1MoO8o3h2LjLR4vfW7OIBlUttDTK5Xhp4pr1G1HXbtAT8Ddu
mRIzmp5qX+nclG59/Ff17WLFFwa3UpreTh8LHSxwP42QC2HmvV1+RZNLUeJjsazy7EjIsHVcDq8Y
oT3PL1i0Pf7fsoSwy7R9sY+BEk29OJLOEyikTbt1m9Jk7gVGd0uzMMuoemlq5m8BSmcbfHZXi5Vv
PVD7C/hobcME3u/bMeFVG4NANPlkylOofXAaoqs3+SyfOC+/K1SdXdWlApXdALbgcaUbuCcAtnGl
9DFBRFtwCRyrnKXjRnEESw9oKRebGSa9JBVtFdK/Ct/0Skd99g1T9Tm9FmB3jezCu+jGbskGW7Fd
qZZJuIg/tRxmHmKehJhkHz1JKEr9kmMIgnWgTsU9cj5JCl9KCQ/OGKdbGHG52r41tK3qTef5wTy7
UAtFOTw6hhk1BJBwUxd6LXCEIzwFnrre+eETmtiyL+eVvRcl++RygT5rO6x62qTctFP3HiRSRgod
ypQH497xDtsnlu5MiQ6wEJh9DLtFr18dTB9qAkfg/u39vWt7tWAYPkDeVaXJ4LxMjceMZcqYd0GK
H1bjcOSKOU/YNuLWMiAIBZFt5qUNzqLwlPrM+26G24fVyh+FWMpwJIe4SSiEzomvRwo1FZE/K90O
Nec3Q+3AzzJU87iueSxiwpzNWo/9heTM1oYYykumW3zRn3XMX0vA2eWsroQR/E7qE30Kk98yDUl3
5MsHBKzV8ziGX+un3m+7QuJ+bEfP5Xg8zAivlZt4yE2ARfWv1hheHPJu2YI3rsBu4/27/feI717Q
a07caJtyWZWmEmFaq6AseU4CA6bxCx4snJhva/WPKf8+QXk06D3jCYL4kmwtrhlHnXpc7Xw8VAV+
gdmuWuFFkWWIBF0UKdeZSNYRVBcNVnVOgvnF/cY7lwFESyBTJSB1kdvlcdJmw2jeC5LjuQM5qiKM
LqumSuC8cqCfhQBdhm1dX1/V/rgATa66mS/xYy0csePhtyQKNpyUWyYJ5LW2rgAEk/gwBhPWrXkA
8fwkK6u/D1T/fHTCLWEZZ4Q0xR6MEfOmiwoZa5My7WSZJ95QM/xi7txxm73F3P2riYvrfPu4rBnm
A+uPgomk1JA6xhbDqOnAPRXgx11Qv3+GurvUMHyzQq9EziYZyl+jScGH660r3UDfspJRsU3ipM1S
9B9pxTQI73Js0CWN9B+w4BiR3QxuPELwk9zCyVu1ZwJGv6zXMQ7gxVHG4QIe/sdahNp9WbEXD97p
Y0WZRKtK4V0Gf4kQQSPDxr3h7divrOb2pJcbWgMBLAyLqP9XMkiDi6c4CxQcP+2EH08+ogrE5mHW
yjniba9p+6ZxzjTVZPs4OKWLKfSAXv65BRTxs4H7No0iOZEHtWPAcNo4i0WtNAQszTmEEQJUN/BT
ebE35E2//8fulAlGSQqyHZ1oeLOf6md53VrSD9dXxmZ6F9UoIuhd33NiDA2VJoCIhDarsU15mPPw
onFSzQCy+wszh6LExkGHPHS62aWroJHDI2Cblz2uOc2coovtD9yve1xUowMPWZ3sOUTemFrpIjt/
pkKs/8Dep5XX0qt9Hc/mD1D2W1KX6huEDKyWD0WLZzYx0fHTbP9nJPgSXEK85wyE6lhrqCBQc5wZ
ATDqX/77gt8fLOLFUTvMvSmN8palBWI45ZEGlb0kYEBbY6Z+7041G5/e80uNFgEtg+RWSiXki80v
lqfYkHMQM54QXLvlLoZl/LSoBT1Vw2Ja94A1HFi/3p2b/4SmxCNs/OoRgqgy7XWA5g/FzxmQvNau
ad6heTTnPu8o1eLC9L/NejhS3lrmMx9JwzrAT95iqLxdCHCnJePVUC9ymM4ztlKxoOcSQTfX5V+R
74fjuUSZS9rlYt35Y+B87vcQ3rJmniqYIiD9vAs3di7HFjns58qLcvj03am8Gsl924adxcHzFY8B
CMEEQiyBEYtavjhpC0O/eoAmRjE+7rEsMtGq6N5Zd6k/lmKGFMFkyBlv7D4MtyBEJfE2/YbCsrT4
VChW18nCUaweKJEgK5fGXj/9yo2gcxcrm10HDSQw2Sf0HxidUtimy9p7JG8TnuGxLQMMtOg4egRp
N/kINnxPk4T1W5J5DSzMPfuS1U2iBHsojEciSD4Ft87F/kJnuWvYHAhUjhdIw1etKOpjldQQSAor
z5NQ5sMdJqp0ELBKlCqJdV1/kV9v1s/3xu7rhNiTQdC9/w0SP3TQdZhervpyul2d1LgglQcJ3icS
zJkIYdDabut9iKtk+lI70J8YmvqBBXdToWvMZ2keYlzJSZcmGNMVPccRHlBH5cH9TkgGrtCqS074
W9WqP4WnOk8+HRLeSQDVYLHuYFsJ2ZWFAvhsJJ+oB5qOW6zOlrGksWoMlKGP0HhccbdMEjGcy1f2
TNhwcwkLSLh6ibUaoqHxQMkMO/kQ/S4Y/Xgaw6SU9hb1CsJ7L3vp/U636B5wwpreSSvcw4NxsBX/
lEGziGQJrqroJNgpEPgfkrtdlwaCuBGYVODybr/qA9UjCalqYrKKPlLhM63jg/Pu+uZA1kdM40Y9
ps1BEpEHFAiGv9OQObC7AsvXy/VlPr9fShgjmirpl15K6cYs/aSRTlW20IAWs1fX6DW74PCEznLp
LO7FXbafScO5FZ0jQa1G0VgfruE4HXJNoiFK3fP06SgjACpH7Po4ve5YxsIXA5HLvsTrhNXVKECo
6aP0Sy61WSeMUSpvkggyzpqyTlaTBBQGeShkfHCK4+DG4p2b8GHVJfURF7o8hYT4ENPVD4/d/iN+
xREGfPrEIJDbyQf6SBlUkcDua7yqLSAxrIRqcYx3/NuIOTXCkqaAuaH0JZ9CE9oBfzy4dYChvFuN
+Qs/fV+qzMkcBDHHgEeBLVyWzCUmpe//Z27GBg6NFlQsM40UtRwdVaM6CGWiOgpRBI63QAfzPubX
u8MptPlDvt0jBT6ndsoWkNV39UBFn9asOEGfKe1fa4ZEwS+92+Ow7A/wFtzS5SdT1W3Uph8SwUZB
wzBhy3dxQiFvbYB/trH1CHCRroI3e0SxUn16aLSMjGjdvkw5NVAKo7G1DEroY0ro6KQOgbxYULfN
upqodRoKmL+KvApSASHEm+wSIW6ZMBb/Kfqn29NDM/g5xkX5N5YHqKXWJM4mE+/xQuav9BjjiIGN
aQtkk5mBM6YXbP1lHOjv/imoBWQ0Dmcl8brOxYB15USIPUtvOQ5oYLZMWyjFdj9MzDy8JuMpQ0nE
heXz2grUx11sDKEReFrR5KC1/jrdnMIGLy4SoqkKJgOfFVq4WoECW5NPvU91xzcM8tH/CGwIDoLh
sDPuntlokoaODofIeRspDZ8Wmp6jeimDGVrf39/urcAF1+TY+camPtzLjwIsuIRyrpTrCgM07sl/
UBpZzT1fOvNbSBdMA0wklGe8MoWn8rC7kjiPEkNiRQqxbPPZ+qJ2csBKxqpq0ULjE5mKh98Wc1Pk
aT9qPeD8YHHD32MCRzyGCZCWt0zL19YgQ8v7zPwHZSAxe66gLjc/jYrU4nzHwTk40cD4Tmf577/a
9/04L3j79xOSYVV6dtkQBeEMz1INnctOYjmL+ovPxbOBPkLqNoul+FoEyM9wFwQp5Qn9LQIf+C4C
qq/4OA8plD7KXEgX9NTzWYfYwuFH36++MAi10k8uf8cDWRi//8bPA0OdL4ur0u5j5SNwzRa1Tx4v
JYFzvBiJ4kmz49Xbux4GUCs1slEjJ9wVbAcZgfdQUKLF70wceppAkaTpMCAls9ebls52HruQn0Z7
ze4st1crocPLei7QZ/A3ZcdNycc64DyQRrRP1bd6PqKPFU9OwQa/SbM+Wwg7gJkoNkMSSyHQ/b/v
MxM/J7Ok550Y9oVjePbGoLLmzUDGbK8vmZDeOtAPRnTxnKgjK1ySNEAus/dp8GL5MJHhdnNMP9vn
3YEvhGUGswIbqApTOUwSd9tNrIOWWsXcF81b2BqkOHJR5JWF9rToed3zOfeNg6CCF4rOs2ndbekv
8v/ACQ1w2BY7zhkVJug+QnrbtcEf2cFWT/Y1fooX+laGI8BaRIvr/9it4OFdymvDKseSzDiA5CYt
gKgbIUsTU+RcjvVZgeTMk4XNdoIZOPV8t1chbc4iLJHhk6f4ZLCUeBKvFwxoaP1uehrIV2lBsYki
z3N15GJpXxEOlnF2l1hea2M+wr8k0l5tt+th8p8VZCIAJgQqnBYXunS4pJFeIgklbsQd7Fk+q1vd
8Th+jc2cHYDH9h+BkZ6Fgvj9jHyF/rgLC18RyTR9UvnBQPtzbMCuxfxSTtdU14BHBHMxb+lfvrpz
q5WtenhVKEip//+aRtstT4oPAVkK0QtkFhNBjMYEKb0JDiB5806zs5zgUMSRgOkSjNOWq8McP59h
THoJPlAGk8QKPIthY1T+N+u3cGAgkC8mqN0Ha4x+11NKaOo8D8XbfuBLng3y42lb/JCdxRt/3Rfr
yQcyYIvOorrlRHOcb4Z6gxA1b5Yk6KbfQtLdgPqrBxevBDIy1AbVGhdksVNQNjBL1n0SJ7/G+c5l
GcbryHYUZQ//BaW7tg4NjtcWViw166HZ2rhzJ0zlsENQCtCm+iYcr2JWqpvyJEuSV9DIY+wJZoxp
mje/M0Tf6OXIBN4AqPsK+uGavg0gneKmLwIRB4ZyT+rAmixlYCImT9zNDAjG8c/qy0MOwIsRUEdO
c8iNVVVJb2kCCQhPCNYuv8/XHA8VK6Vdm/ElnbRTo/khY6maxW4x24Q4OzvoQCtX8MHRTqtIbOB5
/SzMhpmFcDFy97pzB7s+vO5H/V9oQbxmaqhJ6RruiPFa8hIdVZWJsZ8U8hDVVsqSW4KNbvphZukp
lLJkIICl95uYQF0wm1cSAmmbAWhhN6HMH6XN5oisssni5H+B+CHPktn5OFZ+rPCdPGmGKgbfujBv
jQVgvvXl6G5cZ/hwh8P5TEKSzyFYArGoSGgJQX1ez25/8ZGC3B6T51ZIi3sWSNRl3XTlquPEcupt
ij14l3rhVTBvsl6i+JkTkOL0pTTSrl1m6bWgJp8l3PNBr2OcDqku44XQKeiWrCAx8B7lhKgA1TeI
9vgQYrrQ8CuxISb6XvtXCxM0TZEgTRM3i9rkMB24JXiNZWC65uF9k+xAMFWWQvxnui9DhYMlt3bs
5AcGfoIlkB/iIZY4ry0aP5G+KxvPYVVJ+Yy/QXuAc5ArOFMBXpvGMCQtCU+W4WrM7qCnd5GAl2I+
fhOg1fH0FftsMpoupouG3Aq9MvAr511pcGAKbNFGt0KzeHnylwcxzyK8k9IO5q9gnHfIFi4iEAWO
CxUOHCwhRE1JuRCmiZwO2EAAULfLv/Fh5sPDz2e0y+JePld6uzS/J21SXmeyoAYcqjcr0D58srMb
SW6JTmSoNP1Cbi8BFdLpY5fF3ScrfwihaB45/EgxpLzX8+FUZkm5jthZSQQbT70BgcJrnrdUuDYf
Lrhw6YfhPtYxEboeteekTBNX0MFj+IGKyswC/Z78cQTMtrO5NcnF+Bcct354oSf4mNPXPodNs1T4
En0PxytjOJC/Ko7u81ms2ol01ieOZvmUrqDQ0f413ifyVe+vye1exVih9if4ntoMGU1ubKjlp9HD
zmf2HLUY3sAsmX5nLTj977nYmYL6QPrp7WfRHsAOqU81lvX9pG9quXbmFRqs1gJ/eP8QsAM1EMxw
ucElkLg+knSDCFvA4mHKBTwIjne2xvxnc0OJCAi3G42fcfFnz9CoZjYzqhBRqRlM0GuXRg6RHEhg
ttnOtUjeGDP6P4LdRB0etHrz8r0qObUJqYr0yuw1h1aSGc7WLH76HYkxs6ZeSvHrNoMLnxQy58bj
J2mXmqsq5PaNfppWRsgXiYak9z/MHSTbx5fzRWQ89DDxsX/9YkUOHBrdoA60WztrOYhMLN9ZxdAD
rZ/F/Aq23HSDf1NtV8gtcChHGxNXZDjgaaw29uwQ7ds93AUDGbCDdZV8k1/0RtlfS/dx5uAUhLy+
hWetcwGNAMb1DiirsEujMV/h9xxWXLw//R2wnr9Nx34MgsGKTwo3yWqPOvkSwUaKDa/tV6fpktwN
urjDUJT/zV1k1qZ+WJFH7XWBJOV2NGLDCZiAmtDg3od4UeQG8usmHSGay6hyYi76CelMEU/Ioc9w
Ca9+5NdFZRAPq2GDg5cOgqrreO7nXRGCSjiJIBaYJJMOfS76XHNYWmJt9uZI7fE3OCkiTPKyXWe9
0e+p0ruPE8SyVOLMfLZ6nali8i6JVqxJbsgt1VuYyPoyDuUijqyfyX+QMUWuglu9xaDieajjjI/V
JyCI+wdgE9DzqfdPSzPRox8CLIVti1phP82X5Us2pr38UJkoq7v0YZD5mi/tRHppu5NGB+qpQTOC
GzlGSZ2oYWFkRENcKOfva6VxshO/w11/DLrC1YbVx19G1QkqCk7S4PJVBSMF4ZVYVPDCf4R4BlVR
+mC4EMZmY1l15pP/EH+kHbobPPmj0LV84qoE8VXNhHGNSrp9rV1cOiKTFp8AheIs/cqk4KxvVQKe
Y6wwJFu1KrCateREN3DpJ4TFGbidh8/gLQnyjIDvApF+kOfRdG4TOI2Nn8VWD1vDJDfNuys3rTCn
0w2ufI/Y7qDQHsw4ctGC3Kfr4RpP95CSEZiu3ywge+GlnLMiQs1iEpiK+KR2vdMvHASfalELQrLf
nLyUDbDVgkRwLnZLtYKiPbnFbgXA8NtLnrDJLMKrIBnaiHjJTvZoiz69uHdei8XDrUUToHmuEjVj
21GHwwht91pieFxWpzPeAAqvp3qCfTlDLoNzsn4lUdFYKPrjd3S5yd3p7/+0ejXT50Sf1ZLu2/sB
ytFeUtbTMVBkKyBP+zJirpPVAejl7ZnjszKH1KtktPciXF2IlnV9gFWvkOQuPBmXPnmu2zjK0I8b
0cFm/fv427Um6MN1NYAKueQL+IQmZBtGdW0KFXX3bvGZzBEOOEkPkbfuLRms1WJn6qYnPOlTyUOa
DOy0P9FuFAmVI4IpSxRt3t25Q1IVzL9XdbaQ7FhAd7s0UhfY0lc+Rxzwsk0Yv5xKoJGAr9o4EJYR
sOoCWtvGHbdaQqGHTIUw9iGzhjDlia+8mReuE6yYtT5IrbFoAKRIWFBOU/l3z5CB+yWIX06l0jx2
p8Rh0oqpt4dDNgvgioarRd3XCqDVuoaH4hWGrMtmEeI0XcIaIAG5PpkzJgsECwZ/6EKJd+fvpGNu
9MZ5TQkOl3W2O9HRHfO2U7tEXkgsqJGVIN4XhYeGNxRJBdx49nJH+lVbDqVhv7x0QHTQyuoMrh2K
gT0L8UvKjMTMsTxvEA5HULyB8Raf0NPnYmmwP4aguQNenO0NDyOnCeLAHKssh4vUPPR3v3nDCOMr
rETh878Oa3QWUR6UxCHIX4q9h6l+BWgOO1ce02MSqwbMkFn2Ggvg/mHKuvG1IvNh/FwvGbmQLzU1
QemgRLdeSJUTjy/oFmSTPbfEvEWK5+hZl2gjb/C3HOJ+gJAAbztcLidOtRPt9M9i79DllZ5NTfax
AqekZrAvnUua0bGfqXUnxzoTRf53KkUW5YgxzaCLwOVldEUV6fXVIMTYNAblEjP5zHdis4PfRItE
qfFG7X7VWnMQGpC/El9/7BQ78dsI0Jo8dvT1hTBNtnSRkx5vlZgx8riu8+5j2veIm0ltwaoc3u3n
Foozy6f32iA6C7ZG1Kbr+iarG37fctXk0jp41HKa3FEcZI0SXU9AmCPeL5z0ja6gx3KSD78jQWWu
mgAZZtKAc7xJYiuGKA/clS4U3NG7zobNph4al1H1kg6VgUJ6DS3ahRsKVzBWgUnEfyOQwwktGYXg
RK2gU+lwT8WxMkNe9I1B1h9iz25O8Yc4jm9uCgDRWo5Pda4JhnvRe6p91VVn7SXbrj08fykZ0K6h
js5A16R8n+gpt+NzTjKLMKki/Fp91r0BURLatGj1MmV7QevLHiYvjfjl+YYgkHMTLqekXzzkC/l3
RICMLdqj+D1vz6N8zEQRw0iqj9kZ19SgWHF+x6xzfYwcbwFrBLVlef0bNxmp/5/mLdlK3BcuUk+5
iEqsspPKBww8T4cZnkhY3rCVTW7BDBTGDKQBAtHOk5bLgS3fzhAGefXkfCkR3GjTdQd8d8uFbeEX
8Idq7cw4OKGxQhUNFKI4WH4teFYhRi7B3IHMDRkCaRPDmUhTL7fY495G6XSkCQZjm/G3NtJQM2y6
tzU9DQu0yp2gyCN+fEip7QTNYLGTg3biFE8Tj/puIsNAd9tqJAGyjuofjvBfYpNu2UXdeMFkGTRh
aX7m31uuV9ZmRTIm0UEhZRBq56ZvoufC2xUrcryIVv/wPlfYOhm0y+r/NlqQ/J09Ml2Bo9CvgDuU
5VAs9x3fTH/1E6gUJWdI7JGEuqYjKq13VmyQfR2FAaFdZvOKg33oQMy9EXJ3Zh8l2Hl4VhBKoOhf
If7oyVTb/Hwpy1wGFrPDG1V9Xz0r2L0UiJWTKFWfUX+XuqDCm9O/hAgV3axch1NTK/YJgNfzbZUB
8GOKnkiZYt0DxLJQnQiZLocTY4xgJn2Iv3dWmvf49VzJ4T/g3iSxrgSsqJ0ZepLZHewchdp56IC1
5H7a7QpPFpMn+2xXbeJhjZ9/COKDfwxAqiX5T7yTnFGb1kxnbIGkyw/y8Qdt+QW6C+n71ZgGB/P/
LdxTGK/vc2S6cPOcfff0KGBytoCvp+H7abuHW/JPkPPbdY7bsdS6r6jhcvP2IUGes0ygxOB0iT8j
J7IXY2WftLtx9u2341gZnoQ85GdR39MZdtFuT7CQ7OcBMjD0DbbSJAqyEkTUjnplMexuj4oXiTS1
5Fv3Q1BCWb9SbLaDND4gcD6vC2B7MmaRctniMBTb1wH5wcsR5QtsdIfQC/Rb7N3VlvUJ8zSQlfso
zmC/QFWGe5qlJClzIr8TP3BbQjW5Lj0fx9GIIza2rOO2p/G0zjGRatMPSNXryhpl8oXYw56PdbNu
WXaT/WbqACBo+4U6TlSdGPK9cwOcVIfAnHmqDdQgQF1lEeu9aGQpb6tdzI+qZ0+rG2UKa0oj/hPM
KOqP+mW5cnBHu+igdWAE2UXGkWL8UfHqf8e5k7LvFTsa/4eWj25NtOI8Wj+91IkegpjHP4s6Spvo
fgf0MnjIZBKe68HmtutUp/5WYkpMwo6YTAQ2CXWQui010gNC7PcJ0rZfNRdpCQQeYh3/ovW5CKI6
oGGBVnYnw2sEBS/oAwR09umMc1g3TbN8GRrwpxnhIZzSNER8g8BTR5CqTKMljuyazKXJNjP5Vh6D
zzZ9Ff9IEuX8Cu3FmsLbhX5o/XJ1YK8mCijjvGCdUrPNDSXvX+WD1WWQnipJ7NvJttznupj/6t8e
yY2e5i9fjtPV2yAyQrCeFN8UpvRBa8dpLK/V6HiI+8ofRZiKtjZFL17jNADMi7bSZhJrEQD0W03+
uqWUhWmScI5qK6FMsYitlrtVtxDdLR1natfVmrgb7FOJtfz1SdsQglhhRrUK1bgt4If6QwA7574P
9S1yWQIyqX8M1dLUWuBwLbl+JyY6ohkDnatdeQlTToF/lbyKJH1bDeZkLdFPaBPfcVXRpK7jBU3H
hc5YVWujvt2sDTueyahUdu/quPnJOlJSFM941u97W+oaAw5leOXkEXr0dJFOif2OkRmV2rOTxncm
wiMOYN6HVywrGDIjVU70r9+YbV9CxziNrVmhjFyi0PTf7UTM3tlCMbozDEk1JZ+QyaBlkn6v5Exg
/tb5zLfCC0mchLaaFPZKJm96HxMBUwXSQuODLqyho/himecv6A0Mw4yiEXAsouDpoy2X8FcvRKYG
ZWWHCXxkFFMd4fFIFnwJkTAW/ttqo9uvq3Fl8IXyENz3iy+luc0+LzZOB053f+/kfo7yGO3TDwTr
w5KUVIRHWDGumamcBhVv6EWPh2go9pZqhUe04OR8WkKtL1YhkqxPWy3ztZDtyeCxWxdc9Efv8gHM
XU17mCZ5qz1GZ1cL5QRcinslBzwtPnsitBSoxy1GVTqz/3g4MtOTnVNEjr4cclwbua7ODJjuxq6n
JNZBZNI/8tYd+g8Wzve3HbspVfLyy9eqIIh9cP9AJFnfju0Z6/z9C7Ua3/db3YiGOvvN2ptcOSEM
lPUBy8T97HW0vJdLCFXhjkNtNEcDVFI0umOnAY32B/+nZX9LIdM7S6HWpgZUyz/ezVXVF8YAQkxK
3zq4pYNGUyDfJFXGM1bQ0JK6XBY+mk1TBG7WbrMJTLVT00PPro/4v0civ4duMOBgjziWuXhrV+1j
W6fml3z0KKeljbrxHVLbcaqOmoW/TUTd3Y7ADpwxYOH5GhQZlCqob1n73ostfIphJA//iApLdnix
d1QksWZR+f0RA13hI9DudQ4DlbE0Vmf8gDbGaNm6JoisuT5Dlg8JD9tKERLDET85ssNZTaYh+Hzm
/C2R0KMoWU40IEw1zVVq3JPcjgmNLcJp7LQihYByX3zkpLgBBWG6xcy54ssxrctwGlcRS9ofDveA
x42oRxQZDehVN6AqdhpmACFo9MeipH2gftsMRlYjikOlvw52gcF13VGHv6nFtRoRXkrwEGyt7363
KLBWXlhq/pLvSdtgb2JAFFcmRw4wjO3woAb8WbOtStTQCKeHLjqdaVVLwEKXnTjQeRfhkhL+eHVH
T5fbolsjlDlUmMUxgr78oVcHg5GxHeKN1zhj/nGrB/qiR01D1Z7sWgEvD4l+osE+25rkTAB/00qe
aFQLwUonLH9Am0SzCwmWshynag0HcKqQeTDxKzi/qT1mcVn7/t/HdvBp5hB36w85OZahzoddZMX9
UyKK97v7PdPn02lPxGru/ZVyeeAGEaTtcN6A77NhPlasll9UhLqLVSzRR8xx1TfUop8aA8RDuZ7N
CMO+/x2fdBuTNieadwl5U9d7VENn5iZRAKLv0yrfTevVmfF7jhlnNXuCgcYxrOOcyytEp31Rwxf7
fVct0bD3yra2xWQu1fa5GhPyCxSBSaUXMCDvPxZuBksATplX8iZX0oCe8zZ41C0ByvGWpxMtZV02
PVCiY6Nk4OqLfYjIQQaX5paW/fyGRTUSTQ3lXZFFAvclj4r5x/0BZMskA4uzdAyH+9oXo6YSrTGF
5kfylzEOqTe2SfhFZJ4X5kQTWlzwLsBd/GgcqqZ3ORFkHNBXQD1BDvn05gNjYze/2KWyFkDku4cA
XRsiuXc8FezZLNqq/b+yo4TL+l1k70cI7AIGAMiHXyY6SJdoImOQvy/l1r12KQJWndcwCASK656M
tIyhoXyEeCN/jMrISHyZ8arty5dBujlVG7g/Lsj/W4Rw/dHAQQrwDKLJ/q3foWf4jCCzA9AuSQ4M
YQnhrMArz1WdkpEbw7uLPQ+z9usBB9sZwheXyluhblxEY0Pf5Y1vVzhck14ptFR7vQ46ZBlvhyeu
ehgixENJps75ERf+cQIuWjPx9i+nkWqpl7e7PJCKvP1fYsK8sBCNqFl29f5IGa79Fi1GZo2y4Usu
fi5YYgq3wYeR7IDMSIRYPhhIse8bfi/rwq9itaTPL+q8ooB6ybRYg5nJQ1cLYXA98YmFtKQz+Gf2
SCrKtp++zo5IankJx0SeuLSM3WdoMcNiRHTjOKIaLkoMpAdxy+Zdz4LMkUw9+LtdttErlALmSSew
Wr0DgeAi6HmnqL3juPJ6it3o837SIYLXTffLOEqL+9osAshfhoGT+cQIWtVJTdIij2kCeiUXiEgs
38vN4FJl0zPgKsHfrcqx8XYzXWPgN1RcixuWwSUrbzmaRrftQtJpfT/6UgjFRAy6MotzYM8OECJJ
juBApStCT0z8VRTJh+NzPTQdXwp/+iDGIQznc1PFQZqTx702jX9cOO0D90TtZKbVUq9ACnNIzLG5
o/xxPJ2HWOtcEam6Sgdmd/DqEqo1M6z3qfLVurJOIWzaA1BW4178XFZQp8F/thNz1XBM5Uc7jn4V
yyZDbIQq0Dhf+DdsazwKMHEcar0v/YoNeJ/IxauLX+hPAgla9wnECRRLsBpXUSSwNOdgZJ19R1yV
ZLmgq7gR/7yBZ3MkkM7WBfUZEKEzWT4FvVDp6qF2I6mIhcbWEQKce1Z1BfoElWA8pc54cqTOOIQF
qM3pnCFoECBeFebMeHTfzqyzJ/xrLuxAGr4aZeSyQSaaWwZZyjKn0uOYssOdWySbyEzkceind+DR
wiT6Gt94hl7rB3s5FFMcBIhZsj0kkoBgVJzTiisqq8nIjCSIo/A49jiRIDr9W5stw0QArm6DGre7
zLHv3Y5EjX77PUEWJOH+0+BXSI/RtZ/w1rGSN6ZOfi64eJ6qoQqn0hluhNwtY56zPZtyVWRvD8tq
FFSa9syVxxVGhALA4AUcWAwNmVQHJPPxxV9d7MeFIrGrZLL1XV16VnCsdFLDZqleOugClr8ffjZs
TtyruTMn+vyjzK8N78DF6tTnwn3RgLZm/zfvkrfYFwkotggwHpB+TdGI6dWDloidwg4qzNzTfYnu
Sw6vkye1CC+rclu3MzCF8W/XqKzTZCoKy+dZ0FkE+GJMD5Kuq13hsiLA3ipmGnBI4IjAmcS5UUa8
tikyF4zKYmol7BY2IjQKAnkeDRIEtoY5CrLj8Dbfo7AJdzAAqynsquo2bwZumR4aQEPGkpC2TicC
TVGA+YRP6d9JZIuhmY2VfNOVcmyUEUWV/YnsvMrL/cHHJjnqYL4HUfLsjmsVtgi85odCmunIjQ3S
+QITlUY+rJHECtNSmcIr17aSzJNaxSG0vGlZVbhM/nsc0SdF4MNLHKuNlu1O8uQeiisnHivVvneE
kIuH02t0dxbjt173+CJD9FKVnGH9/5sfFwABnhzNT2P+MO3EEvFhpX6YGwIZeHDCVNZ1U/8whUt8
7xEd5Fd5KI74GCYfOOasuERUAszoeSRmxL5PoATaIrK1XxzIUorZMQ/bpkdlZ/Ubiza/o27c1WAd
CIZXNWdb/ULMNKJ09ZyPTgpbrEOz3h1O+2xdEwj58vL78rohICrQmJQDGz4PxLL+eqS8418Dg6PS
dItH8oPBEVQ8Vpo07XZ/lDQcbtujPOBKjAN97QQ5WwY+SmrF1KFiornosld01+SpBbRLwH3xn1Dq
D/CY+ycTunvdHGtGMGsFm6Lb+zfNwIVUz32r7ZjYzwPUFnzj+sNDeD+H3+fbQX/zmW83HmhS1rH2
Kw3G4WJOX8ATr1ZpIVh9PUNCSoZmrwrGO/af5LfdQty7OKu5evoA3Fs/jjUXUY6X8gEgq5H28d2u
nHsrvM1SxiB8iaXbn4Be4F0Onsk5LUkvQJcHKTTVSlAVQ8WqqVEorwU2NyHUJ+En7cEcK47sP/Kv
nrNnczQxGeCp692LKU78QwF0/YlMrHGLkB9bUQE5KPmRHoXcGDYDNLno4Mb8zZgqHLSi1/yd6/y3
XY9eHwNsQWLb4RCy/szMIxOkar6Aznc9X06Id/CgzRsIGv9mqKZ+blgN3MvTdirX4Cq+j+AFukVd
OxCWX9CbKPbHmYr0iqgPIPLPyo2q+JAr3w++ipNs1aXooMZcviFakpkbbxLJgOEyoBq28mHx31HN
WkZb6/NEcWqogOKowd+MEk9cYLZz+q6vpZIOxiTEYOf9HQlGnwPnMJVL1Bgn/W9LEKfyeW6GE34v
pF7BxqwexWZ457ktfDssoghcCfYxAAkmuPpIG47O/D0vJkAx8JUE1YF8Y7zpJG3DPk53DUSy6Z0U
Q3ASN0kfIE1VY5kn6zMqtDfJ/L1QwWVeDwvBpCoLYnu3m6XNE0pcHabPcUVbKrtke+2BbcWnSl5b
AkKGdnAWv7fmf+gGEbtBx45mzZgIsbovvK2HuX1nuLt7frgooNz3Oq5GTaBDwYUY2VEYe8jkvZ2o
fvgmqynAQ+XPOVYRN6+KhHs51P0+EHjfS5p7RfzK3PSoeJNxyPGdr+O2NZVnRCH8qPsr63bcckCI
/n+kMXYBcfV8G9WbYF8FvNsDae5MgUG5xCqNV0op7G0+8fP7mdeTf4qSk/23ijOcL+I4Xzq09Oza
RLGrZCAmsXTnS11cjNIAEN6N1oUykx3EbgZIfIt0n9JrPALp//mLM1uulxn2TEzNi0P/Za3b6VP7
QsCAryFhZGJ0+xcOIPAEXZNHoRw6D5IOCdQN+EfDM5KU3fyoL8drPDaPBa2kkdx23ZP4BH8ikiSj
WxVAWQ+9ujUbHlJKhkT9wSlvgArFV3rxg98gAGEyUd+fO2LQSeQM7EoRGnx1+0dsRBZFJOZKvnC0
GwFpx58W9chsullRVWgE6qwAW1BWwdNfSaDijsUlEDzZVu4OeJ29Vz/8e1ZGj2ku4Tq8DllPPnLg
BCI6kXT27yqQCovJfFIZ+OigtxDXu8J/O5bgZ3Hy5lgMQCuGjTFzrUse7JGTKLCA81bVzfKpYMyp
UX8z4SzfT3lDK8zS51/Ru3A+3XRBsK4voWSleinFqkQEHE0Bc4ckt9a5bzUfH3rVdieB2+9/bz55
BTNK9JFhRKd2sz4G/c7cHtVjmHSM0oxb85kh1kq0Eu4e5x1k5L63YU8/7s5JHwE4REGSriwKgF7/
upVLuee6BVmU6u85GikplXLhckITcfQAZAC4IaIbHbvd+PNefmXdpnD4P+wE8/LvQ4m3y/qzK+OG
8jJwLo+/LKAmL5Cjhz5hrXFwP9d5mkdGmepWQbP3u1uKfIE2xCRdQi6dXyiAcHkFxhY6n9ac/ITO
3xgFeGKVTFqOqZhl2mb3+Zy1UNn8HvOzY+/zXGdf+q974CWeM6QsRABXYDGm0x/dXcOELi9mto0K
W4rdh0pOdGYQOHQ7zrgfDDHriJ2nyXp44V/rVnLuZHTzwH66YqubTKz7+QLsG/m3qQZEhRtQbbB9
mpFly+iVBs62u8+xk4c+eep7qcydiK3IMjwWbEynwg+M7CkdOoGLF8BHO46Ms+qQjrngMZxHmDCy
xgfxLKX+OAKpFtHeDPOx443DW6HVZtFNdZmEXJLXMC/vzOPUMTTHu4IbRtphoabIZIzuXOA7TY+t
S3IPqvzWrGxzyUO+k2ppFIdd/lNR4OpytGki1fxT7jyIF6tvp9/lUzl6bL6HkqD7/Ju3V4ZbSicP
7g0h2fEvswRuqLcXNNpVRaKO0459EtXwrKamTcLHcamY0+jIvvZqLTY2AYt8jw9e82IQXxd2LHtx
DkJLS6jBtj5BvJ0R0eXkHgy7F2sbsrOxXV6R/vuUt9vgA3osR4PbeAt1J8hOAGelhnE6S3oCUKT3
xo+0s+/R7tQdiYSfMhrHR7rX3QCyjHMp4NuZ9w5OMUXm+DKgSPRWgKQaZw7gwTw9KOY1EuGdIRRm
M66yt+43KESr9RJwOEEwky15thjkvtZ395RO/grAJem1GKf8DE6yT+olxyScDuJDCpBC+hmFZDnj
hzgiWjX6g6RE2gwG7fkgI6GXe0Ds+EHSUQpm5jLRhHKO8VGQFLsRdSGAq619fc4Xrma5Vxf9OOeM
3zfY4p9NA+DDpzjfGyMEMuq8WtH6B38D0G6S105MAbfr85ILB376Vg9u9hxlnD+fCG2LSwh7f1vL
qlrNQiQM5zY7wT7xEmX8gq1iBDDm8vjvdB15HjNCcSW05jeFvrWhxU56G2RqHcSePyh6GsABz6cm
u5wkLh/g1H8onFyV414J8ENu+RAgsxo8F6uX8QdZ2Kxf0TQEkPy0UwnIArMfDLEXhSPG+tf9dRKP
nI2JRvvMJDdrWiv3/6pdN7FTsngg+NEA04kRtsTqH0pog8AJEf1UXLM8i/fpNpbcvO8jiRj21DNI
evw6r7bDr1oICPxXE9iW84knSS8I/8G7khgTrHo/qrLUmZZ9VPfGBA6ft+MnHHeRwwz+KaEkJ3nE
9GSHdmadCUyluaMnzJX1GVBck6YseBFEhB/MGxxT4+u13w9HFiI+4r6dnUDbfB+84PDrFJVfWW2i
rgIv+5rAHZUAnhYmqg3Og8Q52PB0yEIfGMUawREMS0ffvlkKGz8ATYR1QkUbiu3mZ+ngoqJlBnRo
VpUAi9pYe1YYp8vmQaOmXWjBpqerxpCaZTgf/l7RTab+YGs8VsUzMVwIaHNdN4FlK47fKQV97RHc
RZ1lDilysvaQ2zENa4CWYUMkHYyS5Bpaf06GxsPlNgojdyu9h9PzmmiCCXzsJG4ZxZC31f8gXylG
sDeo4tfFR2FxtE9aRmfXztyya2dBCLA+7ohQCYPAMZ1+uPLKZQKruhywtJNBcwOl9Gt8PuYMki/L
Ye32Xso9jJ/zPSo0tGwZFTRkaeZRCjzOg7kngVy4mX4QOJIUpBV6Kq3u3Xa7jbx9ppTXwtQkJhp5
qNxgIRYUvQ+3IhRMBi+0DO9XWIEssxZMA3ngSMD14X2RwnXhdQm9kPlUQ/t70lDidlZNZv3uUfXE
zfvFOieqox4fT2CM4UndJRqxPy2YT5soZLWyB+kPZqUDNjgxrUfM9Leor2UBLrf8chnhcJbH0bw6
ANkV+l4bswDB4Z8S6jrNFUQyBrPUhiQ7POJTHy2VeAOF9B8DAnD7jAAsDGMrXv5qULTHk3sofBe0
mqM/yDuWm+SX/XJHxie89Eb48iKDoSRo7RV+pLVCwlFpUDFaE251bWpCHKYgADHcJP+HF8yZGN7E
QA31bbpuulF/HynmXHzhf+sEUaMSF0HuTdP+sKbMq/5it/AHvbKLAyG+mf5LjAScK3kRivWpvUBJ
1uB5aKxL/m2GI1vu/owh9y7rjlOVUGFPXDLeI9gfXXUKcUAHPr72AjkvHYV0iLiojGw3kwlk/qgc
PIj7K/Zj5ell1otVt1G8OeVUmz962yTTbdGwRFEWB0+EzO3QppV8wBeMJYMu/gLuxjrMeMXA5eQg
Hw6NurZiWs3oRQuWHB2/fRBImw/ISrZvXfzy9z8kKOSLHTU24OKwmR+d4hMC5HOgrYSOR6k5dHQL
7qI/1lA+ft0njvzupvB2Pra/xDy7davScShsBFO22b2LHNrzcd9J327Hx/xsEU+YeY4k0q9/TUOZ
Pp9Pg9BWkhGRs1MvkrIf+A4jl/96JCwP33b553JxU8dre3Lfj6NGSBKqw0/6g+625oKWzgq6H+Y3
OmEgJtWMP56zQUJwiSdElbbIfM9j3wUU41c5Z7FtxNxcdpzk5e37avz5GkiFpWDK+iw/h4dgNRIZ
WgVXqiWVimz2qb1FfyZ+tZ1YN0oxzWmc438x4pR+KPyxOBBQlza87wi1vvVbbHUQBwOYLtTwn7+M
G5hotLJZ5/zfYeUCPmjKIWldIFHMv0tQ88ssxh+OJRkkQfvi34ie7CvjqqYzCWkGPhWZHJQ52jIb
guav3ygrnsz0QO6loV1GnF1UtEZW0iIRfjIoLQ0pAntJRPss7oHjA9Eg6v6TCU0ooMiAjDQ1HNwB
VXueGdlWyx7DUFtRjRXan8x7M9f+94adtS2kbQT0RkFAIEBPdK3m2GFaZRZjQlrZb14YRRRldG69
NKHHPpRAIWEiZ+/su2wNAPR/B1dTv5Z9m8xxe0YlJyRNvRxt4RP10WpbVmqpvMRTXHJUfa8QQw+C
MUobCJIqv86BpnWqdPAOmE7V6pp8DFF9fF1Mclorr0cwpNe5siCLyL1bw/bpG0Uaz6GmExKBBg8i
NUPXM9tR0RjcyxBvqz2OWSjddef453rJZkl/GioQoK3UO1TO7iyrxxMvcdnXgOoAalnLWl/hx5tD
kXkBhpDOv1Zpx0dzQc244IATgqGDml+53G3FjdIRee1W17aq95ZUkTsiueEdEYsyDAlnDJe4oceM
ClWrCDeDDU+KEaJTvolHyBhK/rbhYquW3QV/lpIsjG8K5Gg2dHxuw2WaO6+PRl7Iw/hlH7NlDrpr
/uIYN/G6RtdhuUSFeqPNut+rB8ykN8bikTUVStKF8QgLm2+3uRmWHrdm8Ou000iHoR6a8taKwLCL
g4RIKFoXHdofrYtTTG0RBmkvShoEbFHqtXZ3B7W93IFdyeJinH4O4OWtLdHDz7jawtvQ2TnBCOWU
5LU3r2ZkMsLZoqb/gM7jfS5ZvNCrSDsHTLMR4Axytv77FwoynFZ5KYAL9vbw6Tj1mwSeK7VgfJRR
tPylZAehXlAEh0BANYLTe5yO/zRSzR/g25bZe5i2gYMOYPcdQZquCkbHhm19AeaiqtbcLXep9pAK
GvIKIWft3SddCKQrDhiH5wLRqs9OU3yW4d1wtQTb1K4KyJrO6Un8IfvB7kEElLRe7mQqKJPwmDW/
6ME/i5ntjZaeU/7C9NL159mqDTOJIQYmC+uVgNl3pZ2dZPKT6nMGaFEInOko7iNf1YGOJzpiz8T4
Df38Gw0OZIm5tw2PDtHPNurUl1QaD2bGWhQW+2TuyT7/Nj2t2Ut7ih0mzbx+6xOWGXE/IVdOXwFm
Mo7SiAfIjDvQpBvZiKCDQ1QcimYeTC7FpVQtk9VBTNV0I+lGRNNKRP4CNyGWcvJVBljEg11WGP/w
LtwxxBMJGfqgjQJ4QvS17F9VXESzqURAJEZhthYMQSmoViLgmkTpCCE9XgosvMy6p32H+WjdDF2o
R3Rc2rquhqHJFPojvIhJhkbqug9W/QkZg3QAnW9ygLVZL5f1jrTsMQjvoGTlbn4O2L67yupGZD4V
Cvp/oCUzNVBCvjOveGdgEOK6gnQjhQt2+pVDww5TDKsWrj44DuHPA/70gq2ZK23uZ21cbaufYc5Z
9Bsk5gGtUV51g9psP8X9nOvH+x4lOaDUwZolleg9EAvRuUuMgUrFokwu9TNoCtj/D6uhmTQm8fce
186EMkKdFPIgBdtnFnZG5oc1WXhVZHic3q3WNJiRG+WAagm8J2nqV9fcqdhFveaoBzGJtcSmeoun
2bJPAaItNhXY5tBgL5RUcqmI5X9B+Rn7hYeM3jM3AYTqBwmJBF8rt11v2b/EM09FlPKYnadsYWks
9Y31cLXXjdICmEcKo8/eSckJqAt7wmjeT37gt9hVooKFR4n/NIVv94Ew2SlFDrwDi7ieT0AMoZmA
OMC3bCNp/qgSJrUAfy1sHhzdcCsOSACP6zrlpT0i4BxICqlHjloW5gybw5vzeZZ7LQXFj1ujBrU2
zt4Tz14He/m+UaPLsNK1szOOKoJT6n6s0StWDb4Ps1wdUSNN6gky6TaxmYW3HOR1bAARWejmwXuU
AbLGsuDdtlwtTVVvTc0JRuAoHzGrk2FK5tBu0wYhbSue7Q8JB0YjnVoUCM/XJQWqIYE6IKpca6Sl
O/XgrsaIqbu+NBkaIHCVbVBvJS4e8tIJ3GaiouedOMusASBQkyJV1ZX3NXghNJkCzQE+UBsF4YSx
mX29n8oBM8MX0yMs6ZpWS6YXeMCywSvlloBJPPILnCdxNAmYSki4wntqQKvJzXTxT+WLd3OOqXey
ULXD5YQpmM8XKFBCGZdgvUWW4Zd/s/nhZm3iPJVpZU3sihi8GTE4s+o1C9W7hCdX6fIE/oQjItEZ
jm55pjnDBV5yCCJDS7zB5uSznmUZsc/6IJYw1ZY9GcDUdePsoBQXnawtlnXxtyKefbR3KY2zih3a
iHvME9TYI6bIjn4lxDU3B99b/IjFZ3Mp0lwvijSedjuz0jc+67TWnbhSNb+CjEiqKb1YkyfEQeEw
OgGSLbsxS9pEqaxI6XJFavqgYH0nIcvhGvq1nC+JIKS8Fpgtdx/1vyCyK7E0Yf+VEKPFzzWTzTBN
gcNUCMdV34SkBht6bVC3P2MbWOGZ9RNTEChusKyUSh612HHN58gWAMkH6r7kfX46WkzGrDVxG15b
PHsnTOvotdjP6qjzBVn2GZSCv+jL4joq+Qayl6bRHGV3buzPOHC6CH7XFlN1qa5oiVtVBWU5KnA1
ysYNC63qin1dCgv/5yMfNc2VT2qYtx+sCtoNksMbgEXtfH/cVth45/NCatqMyIZSUosHpKcVEC3v
3wD3rZAGTxZny95ebo/ci9yFRQNfsHbvvKymDESlfuJhtz9iHDnxEOWQtBq0rRp2CeDymZM7/MqV
17Mzt3LNQEtZJB154WM9U9MFOq7bzOR3k1gv7g4Y/CifUtiY9EOkDRi7SnvRo4Bs8iVzlVXypSBs
ebKAyvpHxDIBckRBV4ziEwpfzpBQBvzMRg1PbrEQ2KoLZigKjZaC27uiq7URJ0RSXJywt7CT6kzg
IhJoVf0/TPR+d8kOxliFlqqp807l/aChR6TAzs4GqcEFIk+rVWdXyAp2P46O1kYd6MN4Oa9YVivW
89VOF5ORMWP+ex5275xrF2qcREDDqVwDFfQDi0Uq3h03kof0BzanJBkm7VS2x3YrGZYO0elhsj28
zOj3AkYzcMroRcvlkkiRwLUeA02I3ABmh9h7FJBpBeFd+AFVGyikBIDtMn35cWKKFGAes78Qu9xL
dYX2kWKKIjSwk6Ed85N2AcuB1yK9FW3Wj1b/ClyK5Pu+znvnK9jBQjlhaAoCumbvSAPaM9/RcU3H
FZWLHbAnGBM2cEcL4DdTAgS1BD5afKL+joNDDx10IDU6bW4xEJlQoWn/p/zz91doBdBmaVcSqZjy
a/NMWqjzDkN6IySUEp8qyT21Pr/NwEOV6I0uovOschHW3fdZ64/M20Ij/biwUFta7fkiYMFzalWt
spv7t6o2Ga9KkEkSwk/ak+xWe/O4nERM7BNDVe+aepOR4zn0QUL0QsHIVAbkys3UvGglhHOLpHJw
ktv2Srf5Tt8dGS5pa15GK2+5UgqVzM/DmD0cHMESzLMstiNQTgEz73CTZ3CNKd1WZ0VG3Ew6ylp8
WqQ8lqFaGB2B4C4qJD/vbY89tg1MlE5AyrqRKSnEBV5BzBUHw8vNAa1Oa9moEmMJ7V48N4fGm8qA
bShI07ABiB1ssY6E+P1hWd4QdiYIMjSb1TA64DUC1asc0Zb2IMIH2IyrvgejWn0sX1c+hRlco57h
Z0RWXBeW8WVvrVujFJnqzs60gZQmYiA8YKH0TZlOu/hQpq8Gh8YK8C+DDKuTprvUvV39c01V+FFa
Q0KocG9QWxTyCrga5e3hVH13ph272dSmhP5Ls2eilqIxdZmhQBG0czboho44aSuxoRAc8bo2cS81
q7PBAyAysb1+rc2ptlo9EK9qxGMD7RcrC4z9AtGmRNsRX7my1Avy0z1mH1xViJhQLWb1vwzJyLJP
tLrUI99JiOyuphSVrAVoHNTZ9IdkwJL/+FH86VztgykZGFI87tcQ/Wl16JYOTu5ylhpKrdIuCfpY
weXvmH+Zq6mtD1Af4Q0ctPyYzRixlB/jlt5cOVzsQUvPnqfY6GN04VGpxPLrcqGRb/ORl1hOMTZE
ZYtVdt+F5cXNt+8gE8R8d4ch+MY3eyx2kqMLi1zgwyHHbbWXaiNHWCl8xqxHT895CzRGeFxcpIIz
HV+JX/Q5LyzMwU6v+FaP++asoEQqj4WvDyf+wCWNKpVxKLBa43TrisOXqnecKqRSRkXfV6E5ZmWc
inUeJknzFdHagSXbsv5KRKwpTMBoqaigiD2RVW6HbGoXZeX0qyQHbQjoqFcPvRk6wB27ewJ+mZki
1Kdea/Pa1eDCf4Q8dzWAk5Ux2+6JUPh/e1sw42mdfY18VY1FewfTUJAh/dlxNm664/oyjDjeszmh
XnMw2wsgEi4U54UvkN2y0G6yDcZkh4RJIVDh65QC6qHE7iHVDc6qFfm0Zu/0xqC6BgYJTNj/EvMx
phsUoCDlny8X32NwqzCs9+Y1C99MtX2LWlk6Vm3Dhq2SI5s1W2TT1OVTdWDXhFm4/1QE7xDmSsCq
0yaagFCG8Q7J3xzDbG+3W4exrIdXeFmMUhuNrq8gRBy1v2ZsQcEqyJ342Rd88s/KY0YwN9vNhlqe
YjVHfZZkunkhf8Uz+f9AIPAgAv+RXRKoWDyPZpTv0AjFZ6eHrWHh1fKhreRey8UvjhAWPLIx3GkD
oFCIbhrFKLjQIdzUPw57BteMjXo+JjESROGKZlJBjdChgnY91YI2y9Mck81iCFoSJo8jne6QNtGG
C/x1f7roTuvT5AUyKhFP12rBf369eftD+2gzk0WG9/8A75AxLxHCh9X+lKy+l+MghQKBibYYaugc
M6LHy4KB+D5zDDvrpCcrvsKhetcxL1pJ9XhDEfU+YMhg2saAumRsUbo83Du04lTAqHjpMMcDIbXr
EEvp/r+gNbuQJUOseI2VgC41Sp5OICGcUzLX68KigycIhbV8/osK2EpmA/XZdh6J6fWoD87aJPUB
8pPpgwfloeyO5kMGKl85AtPp309Y9gMzABSFvEuVyWIZW/nX6XyGVoUJK1JP67e3kaP3gXvxN5uJ
wJNlC4gRV2i0ynkV/pA5dtYEcTUwK6by3aweRD8XlJcjKJD0ImxyaRZWqKOKBFxaYTVGxmP0K7MV
nb4lM1y5zz9XbrZGfF9688/yoS7nNYlm+uaFVVn0aAlpigFI6A0p6tGOD/DS86TyA4nMlbZiOsEz
4VLgYAQi+2bwX/4XFUW9wrNEMM3gEebKJCqa0qWiiBLcllmsBpgOsB/pHVO7YgUpgNKWOKZIPp4w
RNwag5ika3gSMhbbwGVJa93UzmMJTynhqGsrpxQNJGwQs6Uee+rhfu8GRIzdAoSbqlD3yofLzH/L
QcSvL3qtZdjG/txXJFLGpdmSQkUUS9ieTfe+cl3x3S4FIcS89OSmgliv8A7R83ZoNYxsrsI6ik+I
mFfx3IoJyXjo59qERzs1HZIMpouZ0r0fW0O8eB14TF5tQmnVjP7H6O+oorXGIQEOmZ0btS0FY/QE
5CZxM5cIDOyAWJYGT1hHKJi6JWr2CGS0TRMppIKuh3CrDYQTshnWV+KuTGg2jBSsnzj2avOR2VpN
KqSxUv560mAmWLF4qZ2i2tHZT0A4npEDAV7N7pQusOzuHhtAFcgExarlfFhMjLpu4hsM5UFwKiLP
xLrvCvVr0eXk7xDskVKqdZGIKKKmrCx/jPvFMcavuXDnP/i/IuBmM+nqH8EY/fWcNZNUUv0p4DaH
csS+sd55wY/wJWkpi1P+o/O8tWJdE/KRNCo9YaeD7DGs9BxEt782niEw/zVoigFsAk6wlDkUbirw
YfDV8TZPH4LZqLRi9/uVMw6NWo05xesk5Q0A4hh0Nb3pGhph8r2ss8IULYNBjn5ioiHXMmPxYz6C
cZzIH+CvZBEjaV9U+jOg+++MsIHRODPfr8lmNzEa/Cz/vMABweo6tuL9hj9atlTFdktyIRwkyC1R
XIV+aNLFu/6elkY+1tF2wMFwYdPuS+m6Oh7uqvKj1N0BytX5edzkIWLXSwgwfYZ2Xq4dOwm1Q8Dh
xMTR88xcSRHCC3oXEbu7t1x8Lqzx2sDucFUkahRFGNsPsX5jFHxuc7VLXcuZsoVRZvZA0I7mjNll
Obuz/9GXKfg/BqVa5NtkHKzY+W90A7dnsXFQZTg0q7ZcGUcOdWzkQR+NZBG1xfOzC6IwijSzSoW3
zfdLmHccSzb9b0rjBgAShyLWLkv/QE+Pq1UfjgAQ8iNaKYUnIdirKvtEUHGZotGF9K2FgEyfLdgi
zRXnpw9ZHU6EC4U2d0Vqm/vZfs5G00DE2fMGCmFzxSgXC2qgQeBLGy3qP0joRE6e8MYaAGJs3PEA
FjKOJ8TwCx0yeJsh2xNmlMhnfYlrYx80kLywI8/lWBzTYvEV8yfFnU2VYh15YNjthJ3MR+xG5q4z
SqyMrXs/FPfBpGp2dXYoLpFoViBeuEZtyJph77giT9GBQepqKd9csTxvyDSp/2RkDA701I6dsW3D
PC2euVxwUz77g4R5KybGzRgM7NHq41TXpZmYvRMBWPOMcZ2V8D2CpTzAnFUB3UGvBGg/BUBwjML6
SZrvp06aDUH85XDZsIjVt6oo/6JLOoAEYBb9ZrDs/EpH0eflRJdHjJ1nbL8Mb9KiITSXf4VDdFZF
ltY+6hNUeN/n4RoidqDr3rnpKyqx6ttcYTBqw0MaYLFS0ioLAG+fDjDlrjzasBKgRHIyqgyr+vqk
ZRRVhWK6djmMabG68uYL4aNWDceXzhUnz9c5AvaNuctWMPUxGFGeDK+vD+HaU0HiC/vY/2hfnuFO
zqlZGWz9NR1TdWYGpFQTSZ3h8crQH/xQQh0qYGoqiUP58oxjgYXvEgiR/hsXZ2J8RQGLonJCZym+
Was5PRsEMq83Rg8FUtzvw7bpT36JSLFW2aO2T1G1EhCmKEc36X5ncrxyXS+NPiGFVLJQZwEBjhYJ
oANJo1F9HAJPdqZ7wjcDbU2EsIKUEvpngec7CfquVsZSph3px7caPYFRx2CLA6Viu9FW+LVd2kP0
tCmCPzP301euoZJRcz9oZu5HOWzq0W7FY3075gzmPjfGFdU7wCKoYvffeNP5rDC1tdiwolCmZn8e
wMrKY23G94DngltS4jQ5/0zJqGxLiuH34jze6ecKgDAd40rIjxG3xaImipPIPVlGepUj28rw1j1w
wZToA34xc/sLt3ZU2+QWlyVPAORfY1JYzA6dMTW5w5yg+OQck1ZPKvvIIoBUETo3d8m9HBhrv0NC
O+sIuGd82FM9eQTn37if7bvPCtgBdqY18Dbu+XD0pJlE5hqn6nqanA6AQrq6nyzxweT3MMeVxjp2
lTNJ6LGKhNze4JV8taKV2uEU4Kgv8G5h7iLTOHZ0GykvHv88CMnjjnFFhTbAZ79zfW/bpwkQriQc
zaJ2Y6DE7e5F1vVwndYAvwwuZsUSTLvOHf/R4/3Ke8lcFyUehEvpFeUpJS8mNajF+MC/xx07C6ll
e1+GTLAl/0Eodn4lfZX/wJA2SSxxDoNdoF4qXlytxyM/KTzVZbsfv6MErDFmXlF25QzLPB3MCvMB
szBpco1U5ANbZ/j9NIXo7dVOds2EaFVs/p9XvySnji1R0tkOlcSpbTx/Tu1fnAwWOkO1ZqX0TP7/
SfCaEJt4uhUh4eowumcmvOuTSLbDqD95ab6ONmaRZIc1XgVvQ45nWwZzj5misjmCEQ8OotE9ieT6
kF/dLgknLClNTTNUlAsU2piUl8Ze6sybzuxsYW0ztbMWXp9K28Z4RoSAthmlC6OoC7jU5XqXMrzs
MwudBimxzW/tgYjOWiQ6ifhGiAeSj7RKmN5+jTptrPcSTWy02Vtm3aEBs3gz1KAgaWLwa79Yel7A
cfTAi7hK4HoXhpbwBHZonRMwIesEuwq7MHMAVBI8NfqZFbVVyCNwEuUIxPQD80i6Ask7QYRFdf98
ZpN6V5bQKBpd6dLHkz02r2JTbX5pI/fT7d0F6bzM6izApD8g0kVdnPqIPgl/SHB1fxlIpBiFbP0B
uMOs2NxBUfeUBdAwh4RqIz9IoS0/U9FAElDLZK2y0dXQ4BjlJ5IyPhnJVU0JQ5zjJawdR7RqsONo
WAoHSSns/eX3HeU7nPIcTmHPYQRceKb8FRx/FBCxELqTtwFORwyT6DYGTK/S0/1Y/9MMkfd5dF+1
ikApDM7QAQYYdh1dlBvJXYvweXMsDuGpP0mChyeje6RQ4gDmQkfSYpGcR2GZFvK708Vdg+tG1ibe
7yA/9IOZa19Zj7vEdXwfbm/3UGxhSp3fJsDgi02ntPEv+zDePF2Hq/Aogwb4OUSvd01hCo77GuF9
pt7hVFg8a/fFDzxAJvCsdNJeKddSsbl73eShMTfkOhk+waUkjoWHVEoI8vrePjxnjSysgIIpYLGS
cRkpYP/oBuDIkRtD8JGwS19NvTfQAftnTDKQeTVF/dkwqq1Irl8mhWk0daL+EvMsfqb8Xl2bHJEN
OptiJ1EFOG3tZyCab//1gXfVnkbgryURoKsp344Ceu3KGgkPj6M+JotBqnof2XK6dgmrgsynji8L
GWKsGEThoxu8zfL+sLj8kg/MWYh2fQjlj+sdB5DrQ4SSfyFC4vdnzXPij1ORRLnrsVaFPAGkYipw
eaKyIQUzdXodw7Ee1+Gq6xpQuVfOWvatnomrbU4tS5a1QrnV8p8x5ZHn1dYp1697orXg2eAFKPC2
z4mp91ibBRuIH0aO7VgsLELYN71+8ok95NON4N/Busfy4FhiC8JCy0vJ4mJV0URP74hUojCbq775
ENqJTT9T4KR+RgMIoDq5LJVD5vf1GxdeTm8r6otKZCFm85zBDIeCdv6ZW6yIKKySzS0HMEkemkwp
dnFzeSob9qWXxl+n+736vCK+wCh0HWCE3OOzQUwIX6hL3S6fBrXRYyY8miSFlxVHUQiTOn0q6RP4
2Y1WmXPYNIkgaDRrUMN16NlX8dn1gyYwWbDapk9UcMzr4UNNNiZVTAhUhcotKS6ObkeohdokOfJg
HKlglvOw3CZBGJNTZBpqvb3/dlF7kO4IFxxWWIvcmxm/w3qW5poPhf0glA8IriCOo7kTu53v64JR
1VE6h0ARRSQVzx2W+UStyoDQevoG74Z7SRU3T3QghaPx68jR7yBAsl8cw4wkzNr+y/ZVW+5ab1Xc
Kzwb1yhMnhf6v5WcqN0Feiu/fEzF55nMBq0aS3JePDgQ0Z/YHtvPMwUNv3eFaf93rtoc+QgQmufL
kFQ8g2To+1byarar27X9sZAffneS/hWtCikqRPDrjJNJ4AChBEhsXOYq/6Qr4UAjrkVfZTQxZgaF
wa3prwTKP6O4dGQkFVIqwFyWWZEGirIErbqCvVC7ibvV1Zgh4yG+qUHo51KBDkU0aKeLUA8MziXC
7285hww2mp1BCSdhgva3u+5JdQ3YzxskbO0vbIk+unU2vX4UqmxZywhG7qYalAepWNyn5dwS0ydH
POJj8dgiDoT9i1MAJ3NbvFwuSK/Qoh/mkq9Ku74muwW8bVuy40/u4jhS6qt5XLqnwLK1hIIzeOAT
myF1tIoL8NEzvhWdTtYVp4gkINstiAhvzE/K3xtvzjA3e9UmXzGMzLqTV6mELr9rl5pHnVxrdmUi
V3htth0KcTJh35xIgqG4B3gTD+6APAfg9R21+hOz2BrzIWmNs3OmdWSO+EZo8SUClU293+Fbqj9b
TOkc5PaGDcR0zNMQkZP6xIVDenjJOzrb5BQZ8pqeW6eXJvWraa5zEuUtCzxjV1kMnMv89dsl5sM1
6ckh/H+jtU9RTiGBdUSNW5pNi/616BrcCsW8mPZ1qqUxsYxQKViBj9hVw+2rSNJCjjINian6ZqB7
4lue2VfcT0jbcn+JEQD56zYXWOwoO8xl+2vPOB4Cvp/ftUyDwy7WbpU8kXYvELc1UrruVaIHOuEX
8asMoIuTVaaKx6wuqY+JbwT/dx3OKK+VCx1fDSa3czrCmFNBIxu4Hxrine+i5X66s4X6Cy8tfMS9
p3f75tqKfuP7DsX9WY3ZiBqCLBL+h+zRBlDZnaNPshRQ0gUGm3xxv9tkezGn3dawPnwg1DjOeEDe
SsJEcgbzTFqxWQrGGltmJMdWGYzCrdz3Xmc0cUi2USAWrED7dAV0EzCudzHpnPrL5HYnYsBHV9s3
LByh7tbv2uV8AWHn7sIYb4cpqHfgVpq0IxiGsA6XhQpmDQZNgDYKpdH8agxVxbogSusmz9GPX2Ur
/hejrAIL+1IhLFhi3IiBB0vMquoJwGaPa2eMUFc53ih7CzeL/JbHZJMSkJm4Bz5QWnukSBsa5+gN
sQ5QuBYKNbz+TRVcaPlwA8YRY5u2ReQxYVfEICqM9ig+7E3WeGCRKYZDyoOM/TsxjvQqI2EIxm7R
jbXlP5UiuL0FDwXVws0dTS5pubMeDla+M0zJLMyeoljz+hBVN/IapZhZ1M+CLBqGAf084Y2kQ360
1BHAN0Oj3NHXOGJCgdiT4dcVWZnjFdsDX5vMFTn6JSP/05tqOp5jB+b3iQ/8lYHFzOQcaiN5lkII
jrqiNro3ToEYG/VmsIgAVN/HTqmEOiyrH+Jk0/0xQMdKiUbvSj5ubShlVHEQQEyXT04nLVtDliqo
OWb9YSW8MgZNFYN6DnpvwPSIDr/3OBmUEJnXFlJ3zp/mJiMemX/PPwSeMnG5YXR2qOu3wFsR3OQD
6VaPntJT1FTLsPRg4Nd65Q112qD+Wcm8QEFPg3pXRvbVKmhkefQJMgxd99Ged95CZ4xVGAl/Yd9v
lBuJJPcpRrv3Nv7U8NYSTjVBg/cQs0a1widdY/0/S1PrYbpI3QHo9+ITZ6cL99D5zv2K+Q4CMMe+
F3/47PQja4mSkOtXZpf/4qbf7pLdKUkm0zIvN6zaXH8wmBuGqeHtAnJOCj7/ZQQQXQls88N9jzBf
x/T8BGN936/Hwpl1eDERspJ3T2su7rBGl7TSIspcemzmJjhzjHIea2Va7vSDKfuzadvCci6W0iar
gP5f8AblwwIFggqCiy7u1/8OawdFLjye2L1zHdlM6scW0jKDlpH1iiCOKCFjEiYeVYXlJdz9fi36
hFnYHjrH+BfnKTHWUmpTMH6/EbNq1ABTnwf7JZVGVdF6zvChCGmeTQLKfks2tvKtslIVkb4KBe2k
HT4MnzzZzj0qo2J8BOqwWSWlM2+xJ4oySS6myRVOUvmPeOvyn8vqrEBtedO0LeEMa8XNmFigMtOz
pM6XYZvmJT/Pc8kmuRNTTIBP1pjsWEhSP45x+/uMW6Dm8yCVanE5bNPBgubbItzWZNHz6X62NFul
R1uZls0MFiDDQokFzP3RUSHj9o6ySlSRJ1RiMrH/OCHCW1LzDU1zcT9+5gzinwHRpliml9FjwwA9
AW0IQIIZAk6Xd8ErDJWX0uZGShaU9ZTkcbqKeCT4g6SEhardzH4ukfNAk27qofp4Vs84Ef7T4AEn
mkEsDV+X06b4/igxa9aQgO+0TMvj8NigVstl9JLMIhmHjn5TsvXiCGixDVndFB0EG79fobEAQfPz
RT9lLwXG25e1qIezYRIjZqVPn0/JkP1d13k+RZRr38NQhJoQRlxQNDQZQzyclZBEIgEFvaIy1Q1Q
bm2Fu133T8SCA6ABuigP9LPIDU3UILogvqGu7ScToQUrcnURvKaKNMSk5Ihsvipc+L7fQGUS1ow1
QQxM+Mb3JSOa2hJ5p1ImoWnYCxgSF2YkD+nBwfOIEuQsb6gSQP5PXIyH/7cF3MRIzpwi9FftihGf
YbFDmn248tA43kpbZLxEi1js3dTgoT8ciQh5XuIiCtdrEmdbZbUY1BPAtq8moppFbR4N4cu4lGI5
P/MWejTdKwH8KfbewWOHDIar7gnQqkMWXJOU/HwqAH4DlKmDcoePCN/1YjVVo1u8UOJ1gYfegmyy
5sOU/3135xsAu9GDr2V81CdPsTMK+niRKfR13pyqz1maDhHFrZ7HUWvdoNSsPrpPoS7f3hN5CjWg
KozFCMrlw3h3Q8Pfr3g1h34Y1OhCzkou7zKqIPYZ5UcmKKEcmFKpjjwsKGq0CH0JxnO3e9sYLHYP
Fbm9F5sItAmCAB9xYsBeiHVcSbPckQeD4fBzdp294tKs4vKsge3naLWUYcMElTBsDe8Xvn+QE05y
kNio8JvocAkFjc7Gx3DGqZht7tH49kfz/RLPAZX75nAtKPUCAEQ3rRi3g2y+LMwO8tccm4iftTrC
35U32rMUJUnkBTA3l4eKJXi+ImPMb0GLYYnPMGHAHts5hTLKxCZt82xbnCwZ3Vy5XWVGC9C7vcXq
aL6H56hxqrESApoweT2puYLpFEgwSS7odjHXdyV+OuzvjKlbTQfhFC+OKDs+d5MbW0SYDDmbe3ui
1YdvmjoX+pLYpQ1PmYvYgyg+8eD5lxnPdJNrp1kOS5ohGtt/x+/uJCx91xORDvlsYM8VC7aI7tiI
igay9Ef4SPQj7x6B2O058oKeIH0YtIpPerpC116nf5DPRsVSTiryz+NIhloVBmU4O4u12oyFps6O
k4gJzyhg+DC5Z0nXEioTao8Zg5GXdHRGC9l7hs1KyWXkyyfkSabOvlJRgyHNcCjZJpJgByGB18D3
5OFNRQTSi9VG9QkbkafsSYueaF9XKDtID9/LB28dmCZg9TCCrh+7J1577ZnggVYtsdRJu6jkF1Q3
KRQOJdFoJcpuzz7NFm56WCSlrplMYZO3CuSiWB1YVJMAXS0AYHPJSEjZDNiUzR89YgHrLYPWpmAc
yGEMwGd+onbuicbJ3KMHH/6Ox1+pyTWY5tZxSMYtEKHZGjvHfT7n1nPltuTdHB9QfwQ39KGgYWuy
2Ha/Wt1jWrd2LjU5IYHJAdMnC385Ib0TJIKOKgaXrMVaZjdBszeiOmwkFdLd1d72EepfRkaKmO6e
0y0UDSEruk+F+iICxKFVP+7XKObJkmOOHLt9LRxboSg5wSASb2ykotJaLerpauFdplxjGH7b5ysb
e/OOmRVUKCiW37fPuee5g/uS/LQmSYPUWf9VPK9ntUaCVc2q0hi0YWLFH79aC8l9/tsd/uDr+roJ
014772IjqqJogyJEaSiH5k6y8JewYgzlJoBIYJFkFGQ0C3ut/Y56l3sOVtSc1Esyt1lmVJtNj3D6
i8jN34A6zeiLMYrfHRkpxOJjtzlLem7QS3kHziZA5RYtpg99KAnB86MNcaVOroJfK/JPg8ESFIX0
7wgIysoionKk8KcG90gMdUMVn3tuI9oLzkTs9FiIw4Qdkbh/qdbtevdhqPnhcca1qzvM/A9NZCIl
LupWTvdWa7DFUwxwlM/k0av1tDmmptz5Ffs9lTOr6MMYeuh6higCVivt3OC9bLNJZXnl9V+7JGKW
qMhxmd/No1ScIF1UFbgOselKamOuTbM2xbpCYeCpqyoXPanztkuCFz0M9+ekanytmahBLG08q5AK
5VfBpM/i6kit7p91t1MTDScqM8VtZmvHnumXyYmEENxlHmtGQkW3a7P4FOynTOD57IKK4RALQvVX
tBwSOKobsoOuqd2lAvtM+P3sSPL6zvT6gRGyRFzSnIZmjHDqDHum+pOAZTDRteZJhK0dC7O5TlSH
Vrc+kuP/W6oU+fU4VoZYPF2sVwdaAMikAqqvTFfjOyBy0U1Iy9w3CRsegYBVWOUuCa+u5I5FWGdT
mrAm7+SLLSUqeUfNleZ/VGrweXDz7R4+/LiIxBD95MeGMXa3Kcgvv1kVu0m1UZ455o0sALA7LoR8
0D1BvaP4LVTMgcocFP737mqktAPoUImeTP4LIx3dj3mrQnK6FMtqrTXeJHC4PU+6pZv2nmGbU5Pg
NLuSZau5uwIisTrocI4pbrV1aN96Dchx81K0TQKKJmnKIGZd29OGeQQ+tnysvWRpkb3qbEYeouN3
DRS2E5DY6M8T5hS3cZZvPTWPIhB5UVSP3cXPRWm0Hz/knyD8OODxRjYFz7e/tBrcVPJKvHCVaW1q
IZaK/iwMi/p459B9RlvLANTrrrSqYMScPMNtkpgJXqxwq5WMtZA6jb1W45ziLpEoCpkcyYizCaPD
beULmoxV/Q3dNWk6mCHWHG5EQaQk8D7BPrAGIc7ahkbUft358V3YnKTzJp08Afgvlv+R2YvtT26s
SIu6BC1afGvmncTvqXtSQts4JLzBI1ruwrPwMmjXQgQuJ6dhnetSI2CywyIUd/v3t/HLAYyHzTto
5VpTlkqMIZ5zg4yhVjTSlUG6M9grCY+YZ7BH5Ih7KLlds/E1o0Yzac344vkXe0cPYFnOGIgE5qK5
Is2GLwspXn7DpEDL42Nte0rXLZ6KQxvUwdGcpJY4iGU7Shykw2BYjXLtDh/8QSGlJYQvQR3H+4mS
O75Dw4uUvhpz49Mv2M6CdI8Irb9zytN/Pg3MZLx/S/eZVZAnrqCFFiIgnXFHWF34HCeypHnQG6TE
0Du/omxWDmBmQ4fQYIckU6HhRv8AO4k6TWoOV5k/w3ujHDCiI3/bVASRoDrMQvYrqOLpt9o0M9bJ
iIP9M3w0IjOI+AVrgmLb7NH3PGw8+WirNkOFLsHdnXHTp7EAjYA6eSUEEkxDek7Q9Td2NFdBiS4H
pltB5QuF0Xo/1AGSB9qTsAjDAeOhVed00lFt7oZ5+5as9cV9aV/fDB+8PY/PaSV2IFwfN7muUmU+
tNjY+SxTd174I2LQqQCJKpS9un+794e0aDU88287RIx2ajpVGevUy6HitLojz7tOSxsVIfURDLut
DfGL1GyjbT1Yu4xzos6Ckiibj6bgtrlnuDvwnRLmxYvf13KicXI2TMdTVN1oA6w0Lgu6Y1BmHZRk
6om9rQ9U9POsv3iiBd+gOaEwR2yUETAVaCzHdkekIWNZr7MjALzsIO9PUswqgq9uKkhYY5Udda97
gzTM/HsjnnZnyLHLbR6kIbNIk87V76dcAWnMfHUmJz+2uTEFK2LPrPyx0WylWlbjgxT0dgESkR1E
ryrNlMgK2z+fMuWbkvViRaZmfKM9Qv5twtj924CtzvK+pccW0iwqEQxsUGhQpnlgB1+Acrxwx6B3
Xr45GgRFR67Q1yM3XIQgGbJdW7dLmzSHNOFJydMuvVc//DvAUzwj6vUL5bjhoBzEyFsG6ctca1ak
geltUTIkE/fJ5MN81Jwoxo+1GcKs7+zVh3xZGr8gtypAMG7f1ssq0mNj3o8GyoUSQd99OJ4YSYSI
mh3NE0VRLx7U2I7AlEMpsHldBPExoBFByeeDFRZ+doa5ryb/9jVk0ClfpDKZFbqvtm3hTGQ5gA4A
Kz1XXTYOGkDGRMPd/8TUeuZRtl0T+dSUwfj+w4nfVwz2CpqWjaB3gsxBSQJJZFWwgnAPtiShvM+M
5peuwhoT19JyID04WmZ45DhbChWyizSVsohOAfl4X0uvC731NDoF6CLPrtbXbx+2Q9ssq2alejgP
VsFNLvJ9aK8UPnUq/LyYcuIPjlo3+G7IU+5GPqSjELsPQ/59Sf3YaO+I3JkqG53oO4wf1WtzhuF9
QST17OTNGBR4KB+uBFgGKGuA30Zg44QNCTFOxoI8W4zwlms7UxPpwO9oa7U2hrxEtGjwHm1d3gNi
UfylZJQpAwt+2XcILAtKkNzjJSV/IK4CT7OfmVY1P1kFIINQlSlfpR/9zUmFSmTtXeWbALZDcLVB
1UM4Qa3cdzCPODnJqReiPvyNM3nzv1E+5kJIXJ7TUMhV/G1YUdktSlehMMS82KAdQMFKd1UPuwlg
dqNjWVWQVQi211ibuLZmCmGbyo5f4aEcdWx61ABkgS9O4YIJAhid15DKTslR0+ZOwc6xN3C+UMIv
F/v4POLWqmhIoNR3vxjt17ngdssBWr4EfPadpUxaNgF7We39ddP0g88OyjGZhO4u1CKOwaaPWtCV
WOFixl+1fEd+UIyS3exaoyXlAebO/zet1vdtki/SzP7jUBhWUcMYvL21K727eYQnMDKnTGQGvTBv
3T0qEsgD4jZE8W2aChr3SdIuYUctuhQfcMA+0Da2z7ecVaqDt4IHCNPMssyaiW7PDCAjeqUGnEDz
EuSfngfH7PN333MoZUjp0U5FIWvt57Uw355DAk2jBhf0ALn64zVpvBWlxXImJfV/HKLGMcS210x9
631pn7dvIgx8oUT1iq7CWSfnfzPZxG26Ng2Y9x8gGAVeM6mgrRW0Yy8H0Nj8kYgUm7z97gyPrxra
Y1ZVMfuy0GDih/9GlPKUzm2RZ9jyggMMWDje/6a0TF3FM/++/7uvORQQsFgAuG6qwvAEYx92Ae5L
zO9Jn/AjNjGSuF1ZhT8V+cupkHFV46tmNLvEDRZucQvadNwYcgclt5x01HRe3h+SUVif/QlGpo6Y
5URdUtq1fXJuSIKRJSEKcxWxEF3/Mkf7mLjmwaaQsdTQxOGThzVAJLwlmKzCg73yYDMdpz0ErB9u
cG//n4d7OzlfCujIYSA8DDGDB3UvrcdKc5EDVK8zkcS72EDFbCpPZ+76h6SpQr5Tk2FI0AI1ZqRa
voAdFNsuIsyOig7Ov8XNJzR0/xWV4FP3gUxn1BDxYt3V/yvn2kSXHV+CXYqumZN6SoXGVSO20+u9
NJs12pPkib3q5vnN6XgrJatQ0sd3rH+sFARoMWlnyVVd7q/PhZPq7ICYtDCVUqzxwc98wzI0XSZZ
gkn3q2/Ye7FYN1YWudUKpu8LDkRauJZUT0S760g09UUZd4xol33QPtUuwT8DmKV/HUO1NYkqR9F/
tg1ha7MPPAdZopVNYJw80E79SzVRQX0KWAFj+KWRZ/cpYTi2CpP8Z1d2MbPlRxBfyakOPTbW+qil
YDnxFn+Qw66w7BAQYOEytK/X1tNnE/QwMTIFEvj3wxVSIyDkhkP3ZFvDTTrBsjq2HvP4NlWAOalI
dMnxSSstBKwVeTAIYwZNSle4jA3pKLzS9L/hTanmEvV2jK4sUsN7LOLnjIrKv6wCWWLZNrmh1iIX
2k2ElWOaDvFZwbBldqT4lT7m6Vb6561J2JqhftGUGVuJPzzHFeFEqPMvXyCRaMJOyp7v3YSLJtAI
Yt8Q5m2t4WTOHP8nGM583Ns1j8MjGq+pRepYbl6P+VPDmJOqrJyssaEwC0B4IIqqgtY0S4rKqev1
OjcQ5izbCM5YtSuo7DrypbtJPP+bYb9ioxvANvzAJpTFQhncdDAQ2B4+R0Am0pRxMYydICLLeSTk
DRC8AxlsO80LePKWxdgyOLKO1Wu0tdYw83bpO3OS7xzNLe4QO+6DNqmv4mkzJRWf0uZiCCmW1pyK
Yl6npl+DrkH25q9wYai9BVTy0mnqP4A/IKCKEnMZp4qhw0ZOIN/njoXd8UVHgOYQGLi+bPOozJUM
UXw4CyNKv5mtWXykioRJMGWvDLnPHretML57FLi5kzUMnbwtnso3C73/Ora3/q/iTRNfC/0IEi3X
WzVzqKptwdqcqfQs0OO8lNDqVFMtxiiIcfeH4M+lssoc5CqpPw3o8goOdznuu/CS4E4gdj8WukwD
l12u5+JuZ/yLOB6A9YbJ75JhxUBRJ62bsc66KJ+YtHDQhj62bz4VbYVjJagbw/kBihZ4HrzrFhB8
E3WhW+9ch+Di7+gGjhFIU8sf2C1i6m5QCS858flkL0O91Y4/5n/8mZTkHjAANvq0k4EeGBrqlU03
Maq8OccPFAtv+yL2LEf4PXOhEFX5gdFvx1CY5izHGuxjNcsmYkvYQXpI/5n0SIeP50K9P6C+0WCe
nu70QoVW72dfYgRdldv5z+4sGzeRC/JfMPDUHT8R1hklvEQWmTTzWVeji5KXkJfJGp/k3dsnmlM7
he51nVmqT7Vp4iuoA2lk9r5/x0MZY3J+K6gb7ob4mKuJTr09OE7WduZGhWaCBxzA0y5d0n9RQ+DS
AScbNw1XT2/k21VenFAENRsRDQ8dvkqJo4/yyTOj15oTCZoJSsrIeTck14nh0/ZiMjqyiIc4XtfD
IsqvQu6MMMbkNukhlbOQ8lak+MnU2SYqejhVFK7DJC2gnAhMnAOMJEm1JwlGpZew6QH4u9jAX+at
3PiyH9K+0Uob7RqV8dA+iH2+rwO75I/U1AJqwz+rzi0cJRsANs/n4Hq1FQbAuwpMyx8lRn1H8toB
m6I3Wr+Msd6GJdIzs48s4XFujoTnSmkPjGuZnN+/7Tet1yJyZWn4H2aq85D0Sz5ZUjqdxwGxNHB9
ZIR2kbGP6Ctemu3AItoB77N2lhgmCkfaD5u4r7KjXCA//D5JOpUiMihVwGBJHgsXXYgP4x1Q/iSb
ps+UrXBz6NxXQnKPH6mWHouaVAwP7lQVpB95eoyaBMc40l+RR1nseSclm7YEM3e5RaV7li41APZx
W+SmmHgrG2ppJBmT+wF2Ry3ZUzvIUyVGTZ9pb1xv2HF5mJaUzNlcFYK2WUjB17xkF1tO1liuqRja
aKQbNwpU6hKIj5oCRoM7Jx33WuPlIgwF/BCWPrgHfP4xD43s925WG8r0PObSTWDSu30/tG6uJ8Fs
SjcIl3oeKSOUVQ8KNZrPSg8XWTy4fsyXOXPxN5Haj8X8qMXghv55pOTVyNpUTkWnr9XZq/RvNgNp
uWGDqQLYa+p5Jfez70jA/cl2DwgXSUp2KaxsIaaxsxoZRPAwdlhQPcTddT26/70hIS8tWuCSoZQG
VjqqPsM+/BnQDWXjbqak0FAMvh0SloJzIrEoh1pPWc7Fjsj9T768Q4CmgZ3Oj1AnkP3GoXzuIQZa
AFMljtAfI9qlu3iQlxRrZMmR+BxZK9QPsulxM3TA9BMzRS0ZVtM/9vf0AAFnt1C/8T7pgQiz9ZsU
nY6gjePN4neuM/b4WmA/uepvJJRcgek6sLp6X1/YqczMa5TPxY1Rwdstf/waJP7Gm+Nfej77Pa9S
Dt4ZhA+bYHFFHjjqPEXQ7KR49iJZt/Z4t+T0dpUu6eU6n8fASTNUzFk229KJ/Hm/5icHx+nD1+ze
Pb+Id8eL4aJqj3kwHCMFzocMB26Q/mp6FrJZtTAmDKeN1yextc2McGjF0VCZIdY5NlPlsQGFXEvT
pQKIxKRa9FBdwmNYdN1bW7J3X5lirgTuw7YNlXQ9uyrhiIRufXxUh3SZdTNVTP3obBdmixiehdgk
TcdWophsM9ZM77X/y/2C0q3jQOhJMPO5Qltc5moNBNbFz2evPagyVjoMHsWLb9DbFyYViWUp9F6g
6f2/DJgBVWv/5eLpK/sJdRQqp+/LXa8x+lInOWx8XyLcUGmCgCcQLbK2FxxOUkxq0KE7nPnk45uj
I9fICW/Woo7S/A//qh62U2F3K6/Y5+0NVnoaZ3RW7PMfXyl3ylVGa+fg1OUr2EEfNMgjocMN6/BS
Bx7UXgFsQaVQ+CVvPoOvX8Mxc32/qDTS93shsL3m14tUtMad/F1V2xEDt+uEFzYdJezClisa5wC5
OTHXQIv26Dqk9Y3kyPFq+2SsEc467w0htOdB+XARwOgGGHIYGA6Ylj4khumhyLm80fFQicVWu2u2
zR+Lj/CNyuQaInWnWKA58OYb0wUG3xJ5H806Y9JHpkKOdFy6ToLNgqQibWn0kMd0fU8eZM6OjRVe
5RVlVdVxkRPpqyoEMVVmN9/nfuT3a2eAGl9ZRiIGAN9UldexsTQoQDUXjuBt/lCaf/5+NTYrGvtY
zeG+OK6+sQT3Jfi7J5LeYWOMDlBLgjJTpqnqeY24sxPP4o7gl+gxZFoy5v9HuNrr9Fe0R3tz8Y1r
rs4Rfqv4oF6hEHz9LRqYgKZt9CxuOjKBDIJ7caCQZm/MYWJdD/P6fP6LFdu+JcqQRknm/0ngJs0J
/HOVEPexsEJM+WuWHwR7Tcbz9U8fVbCEXYSbzhjci56KKfWx4XWgnDu8MGCAsDaFtdpaw7epHDAx
SOIUwTo7d6HZlEp0IcxzqDz6dURTtLiO2Y67Gdn61o7p7kf+E1cwv4u46b/A5I3qTNBz12ehg1uK
7MMXC88V+8gGaweQ8Clweyd/XTQE/gGwfGjgv+ODB7/+0oUPN2eaRweA6vkcCXaLAKgQYRMdh+yQ
MmvCZbtgT8jkNVJoq4ghS6WcMr+SqOOKa3KzqNzaWWWlHNmAoSZqubzGSt6FPjxJrkLtFLSSJg/t
m7xzbvYsSrSXvh+QZ3ybaxHN43/U10x7Jad54f3odHmZ/L8Kx30AqRneJUGc78Sra1474dJpmPu5
Bd0P8pTJT8E0GdNfrIdI87bUEAzUsy7M3zNkR1LCzMGu2Cb2ssX5eayNJoYZ27t5mAzymJ5LzIVb
/4T6+9dVguomMXX4SvUhZAuLSfbnEHqcZmezegVpazhwXIeu0a22g2prIfSTBcmSSA7CzRQwDvc5
I8j2a0urCW34/ALZo3Helf+QvcqMOWN4TKvn2s1L7gjRhrMSzNKRmPIZI+u6CwYDy/hYkCMSoZtT
QWILMX4ht2V8sb8G34+cJ5fJMNCOJTDXLLexpcbZ0ddhF7Wx++APrJvKY3SEpaRzpHSkuikEDyqj
MyB9cYE1n/YhYkoX52S3emVW/K4QFCaBrKJm/AxUR02AyyxLwnLlOioBw6VCmrypctTNnbi8y7Cz
OgxR00qYjmCaUbEcGXNwIUkdWhLrpOlhQUpki6RzBAxizxF/JuBBeCdH7gkeaWG4ZeGZdsUxqKgk
Vi4iO0NkKb8afNHbxxK0Zeh3+Iui7MhJNzP2ifcU8Zh3iyfBle/FPWg5+GfIqbph2D4TPnV3DE92
fZ47deE2uUzd5vMOrfDCSh8uqH78f2qUcgf/g9qihZoJRGb9vjKISG4SpXF7mQ0u/bB1FI057bVN
zuqRD/5iPfpAvEwmiZjGdKx/bvo4WmMM5ykAHnQaIEABaWQbzeA39M9z0g/EI71g7aHY08kRtQ+h
2xjKjgAWgxSsY7zTVCYRisSZ9+wJz4XOAk1AQAdkCbOxb4jLhjx8l3ZpZ058GkHwUc0vZiBx+DvK
Sd8BQxQYC2mVU17mMpGUpWOHQugS9NLYlPFa57a7rH6BRIudrW8PAMe9WqeNoAYOmaM3pIeLc/Y9
5oY1CeJuogkdIMJ8a7tuXNcEXFEqLQ87bJK7ASTva+pTxHUzt+rT8Ww1p3MW6s2jwCBnnRl+tPWL
mIUBOTOhHjwFTU9FJUWYU/aIsOYksrRS4IUT7JBybsR0GXV0VZPhje9FcI4+HSsv5nhox3r8rm0A
kkBhCaAVFTEa20F+cEi123dmC4de3BTZOFDYPjMSI74BXzmWjKOQO0PCBxw9gWKMuEtAIZkyf4xd
+GAiS3I0FjKykj7h4z4Agbvgp3IPSAckZmtAq/shtyuCyi/MMEDPDf+ahB67jjqAsJ4aD7MkXn3L
y2YrmBcJesZCdjaMCCgVIeLR9C0GzkuMmnvC8xLEQYcnAQ0GTh3zaKbHMlygzVy5HtiSu/RyiffK
DWEaxaoH3u4goR99CMglWOmLOfECWY57qYb1fopyu8I+bf52Xy3C8gj59jhCRW74GBST50LQryaS
/tKaMFjchcRMZtKC4gRNazFYw4QSZvoJ0w7MpoojPRILYMGrjpj51YX3RlFHPVotUq5gB7bVM/9t
AT7bLKqAXm4sdgGG+tidM0q9xFkIDJOy01ngIqpusrmOhEIUZt6u28H5DxMZcmN3X6DOqn+rkV63
Eb1M5gPA+sJeJWFGr8u6IWs+kRxc3jgSNB6U1Edsod5iplhDNBZLTtq+uZ8wA+KindNhUQtHGUGS
pIm52MzF0+AcrtGT62hv7RHdReMwQHoYhYu85cqXAUBok1ZNNsL/wUoKX8D5P5b/upSn0yhkQ1sf
C9ogfzcbEMdqtZabbcfQevUhrKsvZ6UZn4DvmDmWq+Z3062t/m25hjQCIfi50GJ+LrpG+qZTl0RW
Wpye9LUquQbBy6lPOSN9yw3FpKYgJkC1LjUIsXX45aB+K3QnGlNlQTfUdWtfVyRSl3+p2wQUUy01
f12LhRlPy9aU+lwX4/DWMs979pLwUGN4CE7OZxxYN72kE3sOId993VD0d4zUvMOajHPBkHlAYfI4
kXD06QX5L9btY9T0I1J/7t5F7SoTcs1sWuS9f7B86hml7nAu67ZEygN6Kgggfzg+ei++ccZOlODm
SU6gUZnwUGajbgxP7QqutwXbOydvYr/hvjYy5IdZvF61I/CD3oXXahzsb9UOvuTySfiRup7uAXb9
xA2fpaQNAAQ534renNWTpRPd37/LW8n05nKoab63L/r0fcbg4wLQT7rH+4zoqZze4H4SDPUv2IPQ
SHiOfrHTKSBdOg/1gzfbv8JV4yhlb0Kcc3YY+Ab5gsaCgu07yxcFDkuslr/ti7chw6Nnjx+zKkwt
58MOVY//s5/jSDB6c5R+SI3Oo+U9FyI16NlMTndAV66r4sJq+heNXUpSCHj4TUtS+9oLejGbgKPq
2A67JyC5ZnwrDfXjXjMTgf7bKBAzfhBV1BwVxZIpgorUbj0jgh09diXLj9LDoee1bpDizymzbPED
WJcrihmhwfNbY7isQCHLGUYyP5DPEOmms247sIcR9/Ijsq/XqAac5IwKJMt80NyG+CAmFAks9Aty
oXXQydMCVRhGhgLrm0yRLk57hCnEOYIAy9Efedqed9US1HOAzkfk3ZIL2zPAkpyL3anTRB6mJ9Hp
gHmMcm8Lsvo9b0btGeDNpnq6c2+OmeQnHWXcX/sa62J0mpvAVl+cwD9zeQQXyg3uJqAE+bZ4rgo/
xtOtAV8G4LUM2ETLk6+8sd3q9HPgKiN8yh0BH2aPsPnKcc+bd0akgnC3KvkRXPiVgtL0SI1A4vLT
VpmkW4BN0B/dqlK6NDVPZ2VNXlMw4aembDTn5wEWj9amGUbBtWmVzL0iz6A5RY0j8T//1DXUTz3q
ysx3TXbiZZR+Yp5Yl9UlDyz+5HqfARN9//99Vr978Nsrcwu6nzVpn6XbDvtknej6w2O5r1xZmR4r
oDby/Q0lex9OgGp6JeLRu/lAbgobnmQbyBISQ36sdpqbv6KMQq+wLVQIjKcHFPHJEEkEHtwuXMxd
ZeEDlllnDMwr71cdMFgWj9kEiYOGfmW1EGlYrJ5l9V1MEXUNh0lFnVoTZCjxGrrW4HUz+NjRLS56
+weOGiUNHfxyz/yS0dwsrNKXaNjB1E7S9CoPNzkkDfan1lIKguJTEG8PTrAXKlwV4FYOk/GdPoNe
DwAVCNe0Lo645dPR0KaamDVfkXe/T90pAxj7u327zfCfY7PLPVJmv0olzvZus/3BEVMij+MGDwXK
5i+pICq86hGNmBoHeLogCCW0xDw9aVI8Tns4d6wreCXMyuXO3I5d0wrLC0g7yAyMPTl3CYRQiEfi
GNicPloDH8rKdWtM462SjDqF+XrPkAWnxc4Rdkvq499RJUL2wJantI1xeKUYUzycHblDM0ikKSig
vqT261LDut6b/jZhKah7uihHBLTMmBRSVqzic7JBeeKoaOUO6lMVC2CWfBp/JlwhKg0eQsiTt+zX
JGjC2Yd9SRVgAjtOLI+bXlk02wEJIJK6RQGXWjIJBqoJsZVfKQr5jxUtnKrPnfUpUsSoYcue8e+y
DJi+5gHc7EwsIMqA99ies1ChY5GyBhQ+YGGmJIn/4Hb7EiHcIhi0PYsUjGecJ6/wfx2tyejPc2da
BpQmvOI4zitrp3VWj4HUZggWb13CFa6oueoEQ8Hj59D5Vqp26jc/c7Jkl0gUeFvxGeaHHvj+v2wu
hN3iCBuD3YZ8xB66KnSCoya0W1SxoZhgsGV6wA4S4LOH3n7CXZHt0sAaI9iK3+R508mNfQlPHeKB
NYKvk3+/PsV2bw/B8vqn3MXS0SSJql6Wvde2D3FSJEjWYy+DDZHAf2+08++W4LBrzxcaPk4xqscA
v2IqnPEvYGaoebpP7nz2viY7UonlE0FE+fjMscbrxZcRp7ljowBUmlQwCOFCtSFdaaAPqARtvrVD
IJ9ECbyuN/OjNytPZHsT2CXN+Wvjy8PnHjWWtigvw4lEojvlJiS5f94t4zsPER5XZL9eW0nGhWzx
YkKE3/18BUXZLyJlrBoypVA8TtophrQHtp5qekNkSvZwOp3GD3iGcokVrJDWUevG6pdE1zNE0v2N
VfeJ0dbx5d/AFjpN3Im7s2h67uIJmW+LkZzhvwnVQ0c8Leg/xZkODb+bmo1NF5/qz9BW9GaHjMK0
8cfJ8Jixf8eoy8YjGwG3zxPJI1RYz0wxEeeB08ZC67UIuHIT6s/tGtvYz/thbGUPuAvxABp/Ildu
9TJqhdYicfUvz3Dyaa51gbsuDOuVD0f+ztqiTjsx2pPRG0hjaga80nTBh/AgxHbkDtE9BGJI8qrv
MQSPKd7vdoOGb7cfrRI7e+kpxKTE6W6+My5M00DVEtlM0JVpvVAJzwZ9ROb8umXY6ni3NvONJMwW
Rm3cld5mVyLZvUibV8MuvLaRNKEeHrQHVQXF4sylNR6G3Y6JZQWPpBvYFC7V4rJ9s89QTWqpMVgs
bxrqdw9UmYP2AXSBLMuG6W5aF2Xi3Drq9XeRfIOh8KHXd5xsny4i8ZTA2D+FaCpgAQRt2cIENZk4
/UXorEuwXkJkZfHg6j0CzAT8wO9KcfQor9uzMZ588ZYXrEqMXb35EYplLFTfptqrN3CmE5jvqumh
rFoa44n5H2GX8f854BTqtShmLgx5K3/mNY5NCOf488NzGakGH3INCgbFQZlzHwH2fP6FEshTy8VF
0i1WryHsoc3DOg1HjKyH/Z0IS8iFezjed8X0wJ8dNlcfSE77zzXffRl6s0CXI/DweAvp2omznhe7
AUBMi2f98iwWkUk4aTv5bUfP0IGxJOUqRZL7kHmb35mvq30apf5dm6MlSB3BFJNy31NLS24+fj9T
sAWi/41OCJAun/2RKgCcGXz6peV3coxv0GZ+sm8yol54DT3Ri+PfsEC4+modGDWTy1PJPblkOmCn
cGQDEwt8+AQqWOHvOthTh48Ipd3teIpyr/n5xwEz1Dt3rkM82iMtKuQnfNregU2jXTmfrBP2poKS
kq5oUbhQu5BPwK7VnSDCJqPJ7d/LuXqixxVTyxm5P2aMEuaImKniI6wtg7HioX5JoA/7419NNsYB
tSbUplSqWm6FUTtkxKTXcoCl9FfMYXjTInu0orAWN4saVxhmRMJDR1uzxD/zSwQPNEyuWOFPWJhr
S5TxJKDlwBrtvp/27LMXRxgY+oBSebySBza37r6qrFh0UrxD2QxURopOPavWcBuoqov8uKeTUk7q
9LCqB68FJNyfHox14GUPpdnuXvHgKRDNN6BiW7ZeKzyU83gOZ5Ky2wx4RUXC931p5yrcSz8bAPL8
MbcLq99SHdo8OhU19rfY1KNreqTZg6FFjbzGP/zMWXMNe7kCq3+1DOahfth2nM0rWkCIbp3HMbyQ
f2HRtV72NJtVPdkp0Asj/MEUq6UF5P1eJzFi5dWt1SipN0P3OHZDK8PGEDOIbjBBPOm6UuXsdhaC
0plRYguwz35Wztd/ndht99vEVjfL+9eMIreAgd7Lh9Z0sQidGXOPR1/3pFwrqqfLTmjJhc6IA0ze
R8DkAfRO+4IcY/CPfV9J05iqskmt+iwoXVetpSbQOUip4ZCy8S5Q5Oci4eAcF8q6Y7AJhyzEcAs+
BF4+thZzsdryexkRWkXbgwLcp+Ogsv+U+8hbsnRRb8P+GadhrhuVsYj66KbRXqXC1LY7t7VDNHdg
Ip9fDm5Jzhw9G9u+fMgRAcGhDkgl+rTBZHGBRS/l9otjZt5td1DweQgyjrVeMtAUo7zk7AD9pVen
zhff6lBth7F67ZwsKTAzzZI2IVAXOAINsI+SxUDF+esxV9cgx2WIaeOSgC5E9ZY4jsTV0D5HAYEf
I4uH3wxLP8VzT54EBpB2EHdZLl70IK+GrIAnWSkSmxWTH7FprHnNOkxZUT6l45IkWk/p2hzEEH3R
+GqQ0+Rev0ll4RtlluvaKC0JZQVvkrDsVxDL0u5v+GjDuF6ZhWMpj2ZLMMJieoseHWDj7EmHU2r/
A27pLXpsUjTgf1sC4KM3/aEff4i2Ju10InRnO2YFMZ5/sXIWfxWIOWETAASZFAMKjEg0qMZEH+RT
Cv+g4Evm2wdvrFjgFFGME5ArZn1GId16Khs2kTZW1usRCIo0PI1kqO/B+Annu9t/YEJ/bDKgf6BX
OJil7Gd86tK5G2P4tXYdQYxnA98NghYTUSWqMiJcokv1ZLhrNVRJ9fBAs3abLRDYMwbjroNLzPX+
lZhqC9LhZlQCLycecdiQpcgFgxWhbW7A9TVDdP97OtbcLnZ3lIVpRsM2aRzXe0HIyMKWy9G6yUKa
BT7M5uFU97ukToF56mOFxGthdoFiNuoy52E79i9A0Q9TO+kOG4rCgRLNFDpJtS3P5yTzfvlF5IM9
2rh5Vreq3m1qgtUYY/mEfG0HGLQf03d+nRRjZwK1aAR75GLarLyxiHm5vXDTz8/3iVMb1cXm2qsr
5U/qgMyYFeOLwRamsuYpg6/nIaT2V4I6RiL3St1dqJ8rq22c4k0Hq9dpTWjHk5ecY0upVx08MvSl
QC64l10X2gpjlj+S6DvrX0cwClDw3cmlMIgJ0C5cSnw6ZV/GO8WTiQvZJowoJqWNwSWpY3r9IowW
857eWneOk9hoaspALABkeLjjMl+ewAvzRS9jLuy+0Et7+so8HqBIjEzLMhr/19U7jLAtzr8il25H
YdV17Q2qNIQYA2hPjtPs0n6iHho8bflq3mpVSaohObSCIJai/QxdaBlP9obIHE8I6/wP4ESDDhqf
9i7+QyTmRuy75KWUcDowZv9Hl7yGqRwR0XzS0JsMDTTKuKnXguzqV6d6+OaIa0C8XD1hc3a/HEan
wK+cfQSnI3Ojz4dlfms+kxZm06bAxpzQHEGfwH+q+sdO9F4fdb7zD1uHtESX/d9P36j+xJBMfYEy
aqt4Xy7uRJV3gPq4p1BF6gBak86CzPKTdtpnH9CH6iLMDwjWt8jDjALVgnnpWmdJ69lusEChmvI1
ClVULepbMzEDff+aTjG4fr5GEM6cFe6enTrXOxFJfkIfPI4/RIXibmv+SuP5y7YxnaeuOTD80Oj+
oS1vZrhuOuQWbpU47wHkXi27tbLW1qZC9hDHKkkMuz2L7e8Aez4ZQFAyvpzmhcd+IPd4FMkgjWmY
NcQUq+x/cHpCYaRl8Uz9gNvFV1W5T7VMUTN9TIYXyG9+6IHZI50Qa+nCCEfukymKXqn+SImTYCHW
+WpZE7T8zJxUEoSiCI0Z76Y1nOTRfbp19e1S4wcRiW3SxhHkS1LOdFcpSa+dzAOks7XRxHgjM5ss
iOOih7p2ZnsVoxuOj4nBB9yughc4Gk4ZjCBiiWalmRIUqWlunZ323xtWrFkGgam8RRNMJVZbjnkG
YT6Rbt/bZFpUWwgWpTBf6we8HYsyN6SmDETjZ3XSftSvKwmCSeoR4O2TpZ50+K0JBRvNroajr9nH
oGmRk6tntRpebIeNTVLjBgXpx2XAi6aTuhOXb789SIOvOmcIQ4KPfDmQDjTsP0NbIZ/IuSt8cdMo
hLWPKDoAYcRvSXTzB+b/nrxuDK4z2+LCQFCUciGaErpVBpgI8GtQ0vTQYxQaAlnkc6Pc+pqXLLvC
FL+JSYfRK7GJgQisd0qtt2AObtsFIe0YSF0VN789bXtu3i4SaEqadkb9SIiVF+oBWkreJDpAO6Ef
Cz9x5HTjhSPdkMP+Jabq7WnGCWO6YIoJE+Av2c4oks/8UBHFpx0SQ6XZG3CGr/0QesALdpuzZZTO
rLudYjmdKRsMOuCGwaLul4YlCamzXdju2FbeE7pwab0+YDSOmXsZUm3dwMVkySTJI/R2Drf69OOJ
LaVyIBneKRhWaYjpFgCjqE6vgRsn2ObdXwIXt58/2zj+dPLOSRHvO7BBFZ97Xt6Whhx7ZR6MFnCj
T+adG6eyjAqmSOX7fh9raRhVR5FzsySLfpnirdbB89gLJ1cpWKIigFW4heDUHcmC82/0fg0Bi+ts
Z3FMC5kkFbU2b+NBqIsAKnsmO8f0ONq61d9XpqLGAPYJqBqWuLHyZvsPfLwTUDk0dskim8ybkgC+
5rqkISXbm3GXPCVsC3cDzuRA5IOm3AW+RrpZlJmqD/YSsI0ZkMg3dN0/ul+zxFZpvmZ4ffJx5hrM
t32VrbBHueDkj+Xz0fLtqOfYUmuSdvG3+zv+jxlDMPSVpt7TjIajs9hr79sOH6ei5Qw4c+tDWxQj
jNRBasFXxsPHRm7TNetWIOxrAHjFQOoCYqzXDhkf0aRIQ3pRUYmVzLGImdUVxpjapM1okxf4WbmY
HooqEx9ytrK3McsaaJ08GNkNM0MWsfuxlyZMFSBnfrZOcMsj4wc8F775jXYROJaq8NYvVEhfohV4
tjStmOar3XwxqcpReaZB29c4A4GYctRhEp+z/DHzbr3ILsU6fQdogrS4xS43c3JAmaaEti+eh6q8
pymDbkLeVnygZ4GPvrx1M25Z9Mrn+kfId61CPegYvMdIr/k9XJhB5uBsXZKfQ4RZUGQMwfr68ccV
4yrY+LLJ/bBPQEVJzEeixx4hmtSkaqDfuP1lvTAaEY5bCa9caqv5xtYcY5SS3qV9NvoJszykfyUL
TbgCjP1GfaKiF2coMpKZdiOvadR2J0GhzvqQtWa5T/jezbI6UczWLbjLZ4lkNmtr98ch4q8SQmQp
9JduguwCEuWNHv1pu6CeQ940BNuFQQ1LLhfAV7qQtpFSmmgd3W6ZfyDwtwDr/mbNy/iEP3uCAbbz
y7zoVAP+O1N0IYrcudibSSlD7yaT1fb/2CSckCjSQNFyHZ3+IjAxZ7TrMT3bGFpaN1xf+wCsZYUJ
XD0aFhsT82GC5uzfM694j0qmo2YcTjJLaJ68oLDohgu1fv1E46l3cIjzpzXwmCJ7B6orHTtUk0G6
ckWyNG0zhO3teBgsJnkgdh3CygRrLQjYtpCCUgbprQhj8OxIiV898ATEwum+ffAELeM4AjNKUyDt
lJ192mzd+Jxzgl6EF6uhLbVKmJWNfi3Y7Q3H25XdlN4o7CRiJGxtDZa1MiSisLeqGb0wGj12Px/9
r6JEGo/eQiLQtAkH+QjFbwng2G65CmjlnZy4fZwGkRCgs4crHaXjq/ulxajNBgOZv7VU2Tnam3d6
0kCnD5nIVRX8scD6E9A4Iv0oy7M5ukE+uTajJwxBL+ZPNd9rJJduGxIf7O+JM1G09n5AmYA1Y3iA
RrkeInjMzi6Wm2KGRFFfX88FuR/15fZEntZqPP8JlIfc5SAa6wdWq7VlIde04860kuODhpg9ntQe
HrmLGF7Wc44AAAqfYNKGibFPAzBqNqKzzXbcnFBgqqP1vA9dYrgIkX4KfwVozpEdQkqCbE4EtyW/
zVit+WNY5ezamCDOdJBUc5pFauhMdVBH8+d5yJe3mucjDxnNjdHRNDAukmgVoL0umwoPPYABSZoA
I26hMZRWxfKdLKdxqePhzerRfG+pK/j4i5OSJx8oS21403nMBt/Lp5w13U0SkfKbqBvbM4GGBTHJ
A8s/PVWSUJVgF2V1MGvFvgQGHCQaZa1gqYTcbggYf1p59JZKOrgCAdycWEWJbUEAHD5JoyvZ5V9t
OHQaNsQ8Gv6AcK23XOuv+W1a3UzbtvKABUZS0iT49ll3JJLAY6pM9NLQovmu2AaIQPxxSIQuIgKn
ra2vFTgzMNlHNF9aQakwmMXQwm3GbTMjY833vSDVcLnhXfa2kOw7CAzi5lMiN87cmUTxIoodxyHL
g+NgyF71Pt98lT91Z21HV4frgHwtFpxSfNjJERxwl637Du+1kKa1T6Ap/dx3UnbsORjU1NMOB581
FQ9RofBuQQzSumyvElxAa0RKHswowGqNAP8BtuUxCpctKh9DxgWUZhvgaLFqFf4qg8aFplPKHTrW
gPNHH5AEL8k0eoAzjgQPFSfIx5IxZcPs1Z6XaWagV9Uf6ayHAEyXBS5P8TdQaXjjdpmMn/9H3yQD
J4b/9/EEfFzklJrnfwrDn5tb0S72dCKpMawjQaBhRQ1fZqj2RUKb5flxpLeFSTbF8UuqoNFKLU2T
VztsNsclPz8yff4jMoGwi+ZsZ4D0mTG/w1sXWt/JOgOqMijUpqy5fv8yVdSxz1oHX1pKdUjWqAhg
8BdGnCu1eeC9AbTqQhzxZEl80HGZpmDP3RvYNwf/1MDp3tvVMIAGfhZ3udTogLNUDouCoBX4ZmSs
dftB1kFusVQJy9Lv4jiI+dPg/Un7f4/GYob9iN2S8VvK6MIhC0R9kPesHmO31AQjvHjy6PHgqQVL
mVzdVaDn1P3YEffwj2/VA2CyzmlP2Hj/fbSbuzb1AueQU+sVHbEVQmeaw/Ne/KBKWyBuhgTZwowk
DzLlng0qFN72DmWrW0Z7TxSTpgN1xfNNFU8vxDAToMXE2Xym5XBPmnBBnNkkXm+RMo/TsAwX7kFs
tyi9adhd9c7bTh2OwaTnSW94Cd+6+OJ2EnpXP0Qb3UfAH3TkW/5J+e7nqj1Yp6TxLnQQuqvbFX4o
5N8jCnzE8rH8Tgu9upGeWwtJdgIDiKxhldWcwNmKsgr1mTw7Ai5wMxxnGgSWy+jzsni2GfkGUbwG
lWcBbUejjerYkNWa5yurmCTkp4ufqrJiwp60RrFE/DrbGq4K32eQknDLzy3iufU3F6gNk+L/H6Io
2hNPE1z8dBcZ5CzOlYfEF5V1SduN65b7H3usDwjuo5KlsqrAzSggQ/hobEiVZzrYDZjyajTGrLOb
P+6aF9tYeb1ny5OHycITxhgH0QPO698e5Zqw74XDoCfKItundI9kQ1HIBCml6azIJq1CsFXPw2sD
pnk7ySCi+w+K+xeSBiaBiprMHKFEAw+vU4wK8OL8LJ1KgDaEI1vhiI2kcLF2P2yYLchd8UuRUeEY
LbICfEUpfwZzhV53FMxENqYfVQbCSiLdNVEzwvbIy3ailrrmFj1ioMIgtPFr4y+/DzWURMK84FuS
g7CLWz2NI/hHBtAcxjUPbuFIGapQM9ikn/UwOZpjmHgXgv7tM+9uv67+uE2SEspPyEnmVtQyVMrE
TCNJqJDsVWuQfdDH29AG9GSx6n46I/Y8UC2ZN/BXQDxnCMy/yhFCGSwfVMkY9qgHYvs9DJLjOSFb
MHAd7jPHeY/YlvTrBSdnX19uCQa/Qr3l6ijokbGGEX/9sdeHLzLwND6rGF3QmorXeGvPjXK/OJ4f
AkImBHv721+tSsTU0pzC1JSOat8ZHRQna2300kS02sX0ymvsOxAo/YIUuFceDo5FF460VQdybMEi
b57r5xxfaXUe9grnDlETPOoD7Isuv2UWXM1i60TUS35+lkmEvOrbXcJbw4vnsuXh6NpBCrtVECS9
jNx+qnu6670mEhBk0TKwEYTh6QteqCfHozK5Iyg4lP13RLu9DkMNKft5iK8WZZ5DglKkii+YMrcH
Q1O2xRb8xpDaecf7bElDPEQG8+JSoIlokV68u4XkthG6A1yC3+rTvDWdNgSGFE66oO36rYpuD2dm
GYIhc0nWwJVR/Bg3bcOjn8vJb2hWTufiiAYz8Et0VSHstxz7pJHU3xkwvqxgmOC6+gzxRL2qcx5d
Etpjhv5uR3KZvZEWRCl4t24nHIkCt+NwBoPQcbmBwK1Vg8YLdmHeb1puFEEAW2NYgORjOXzyzF9d
TYPx4xg3rS/Y1wHCQHBmbSFKKPyzdR4Zmrnl7NSenZ8GvLBOqKnAyDaQfwZRHT3SMn/QWkXERlEY
7B6poYKus4HZzRP6/pwtENIaRAQui0sBL7zDXIHAJhbFIT/YdHKfgSu34VZ5t7SrhsJR/Gzf/dCk
g4dRL88DUAzDTVzk++xZ7HAT8JxzFXc5tCej/tUjagBrnl0+OkyD7fDLqniQ8ZnJgOS0aozKqU6m
bkFwYL5kv+KaVzQM9lGBjnSCx/yjCBtza75XvH7x7vWvmSrYyXgxGOa3rTPW+D17nl/ITDYBRHxs
7lqEK/lRyYiv2K6V5I4UhzIUN8gK63yekb4UUfIhFWiSZFDbfBhhTBdS/Ccxe2TLnaA6RMHj6Xhl
gbBhG9hiVB9P4U1EkWCSt2FwXlZUVaHz1k51WjEzOLzsGH9fnGF3POu5KKdq8hriFSiuld9vToM+
ICbldW3of9uC13AddlQob00I6jID+ezodltdql1gIvK8kC8WrVHElhFTF3cFduGV9wrA/xDpD9B8
kPtQIqJy6sEBkigfm7+SYhv/gh8oePk07emEaK10OQHrsb2WSBL8bZL/ty9YcJKCUQuJxqOjIvaO
2s1HMcQayc5x7SbTSCFXCBy1PBtA2iQ4idWEENax8ZRj7JUWaVI/ozV85RvLVBXRhaApgeks5f5a
U245ATuJrIDw5PR4yWTly1trF8HLpLXGWpQw4EkTWODOzfPfCOupW8hIzOWNlDVdAMY4b10gAv0m
BYOqKY4KNxJ5+GatUD0DUHtScg4TN6iT8RenCvDGMuAx6ZLEFmdZfLA9rz8OxE2IUiESwTX/T4Pk
esxwFSUb8rBWmdA9uul/hV1BglmKx7kCJ6c0QKuZFq9PpNEkudrzs0zNYGvhlPKfLHZ70t+GYnkh
OgM7G5VGiBsU+f0roTVRk8SKJD6IIf4mFAKbBOGIF29WNu2xeuesN1ecIP6J5mcdINbTGsnCyBw2
fSs3ykHNG60MtJVOs/NjoYFWSoeDkrLunRr9/fgTEp10/6964ncWwRL6YfUFIwOCLqYdhC61caqq
pf+mLllR04+qM0JNwXD7iA9S9xoMd0KpHdf+WNj/P+ZM30K9vqImRBqgDerO08wuU07ULs2W4OlC
rVZLm9B8QED7aPeSpL5usFyP7Xm0WRWbj0Ua2/SnIyGX3Ks3A1QbaDMMjKYPktvZs7gwHZ+eR8rN
th7vRCoBh0yzDJ0jKLVOyG/3/1UbkUh9Dd7SyTcYaMfMwDFaVwNxuCDfZLycbNPRCDw+7jf6N0HO
YJfdibNvV4PMLq5YI5pBiBcW4OFG3WtYjLGv9ArCKxxj06EHIR76AYlZb6jB+iuM2xsTBk7lmHz8
XVt/PfbdASaIixXPYOuQIbbdDP2YoQ4tXU6GwtyfvaYpgyI8mRFRW9H1FnkQMfBXQaq2cpdYc4q1
LNsSDGFLVSFXnXQtDsZhfZL5q08nKrr9gbak52jjH8UF45h7x+rV1hvGU5fM0rHFoeZTzWe+j6sU
eTaxEBJfXGKIzAwUlxlJCcbP9z1br8sSmNdZFl8XPiGTq7/MTSYycsHC7FHCjrcy89RELyZpadrD
AHdZG/uNJbf2QcUoOA1AW5SK0Ydx6MfQ55h3tWs+8xQzXSDcPPq22ofYJJ21BsYH3wi4X71L7mTs
OnGt0W2cNeGDZSKgYJTHL1OxiDkBxxjUpTXpqs+VPKIXLB7yZKsHEspl5tPWfpVMYuLISGvnKPOS
Jxuj4VzhPaAjyPfwBDmDcgMK8PRjMyaVmZjhTPNcjXjnlUpcOUMz4n3IIgfn4F9KeDWH7HUKXb67
VN2pKc6UZBjHWkEBpR1gJ/qPiJq3kYexnBztyEEiSVn1Zr5Ht35+AXP2CT0UNzcg3RSXqhKieYIH
NJBZ27SLFQrUqD+OaT+wZpwMQRlgK+2z9inBHwbsVs1mt1m0BQ7ZxsPK53fjFNHfJI8YRCgelema
ed+WhsnKPDu4XV4AWQpmYTVIuCk1fMhjZ4LuC0XcD6J22xPLmcaL11DXWWwjjd4AqWGhobt1Lihw
odvLQEatbfQYk9qICqLJAWyr7IXqH894QbnZ5oRz10aVYM6AL1RWInwSls32WynFo/5drW0u6+ze
u0jjmDeKkm8tqXyKeolUBc2EwdnxZl7ZJV/JcbHWsvZuaytHDK7VTmhlfMgH9EEvWXMvak0m4jru
zJ877cv9ayzk/ZEEBWeN+RZ9u2Q8bPFA0/sVkvtXGR4nOq7TboYmQvv/IV/xmXqn6msIr4ORjhz6
eoICM7bnFsJ99bsrUsRBwOXYT05Uw9Vn7+P3655r2fkHIaoothN0EVe/mafrf5O/1l/+UOtncG+y
oi2bEFsSpE+iVqtj8LSaDMq57DOOWvtG6zWO0LdtY9631wiN5PDNh1QbddmV11eEOaJsgdMyKKmS
YpmszNACThPb3rlSYv1D92aZ7ygjVMjdZjlLMSMmduItnWhNRjjysQXxHXm4y58BkxlbeByfzUj8
fySixdfT2alB27090Bilf8mFtSqRhE3tvqFecgZU9NWeyAi/MaE0ozRwSCwvqnPXSevYeu3ANOK0
/kSu0Suewte0vwlTFrKLDc6/pd4X6uvI5DVzIxntYs8KVAgYYj4EalFvgB+JWZ1HcOC21ezE7YI9
eRV2sOERbHilq5SnAqYnfugX1INOWGTsxChgPDlN1xROnjo2BP8GpQTtmUNsgwMeGB7+Y1aMUyir
b/0V74FqcNT5CT7VOla9FwkLTUfU6IwlyVFC3nTo06PhAy1MFrhxYugeK54GtMopNpFsr9YbuBGA
Oxsbw60xnkdO69gc56rjyywmSpffJ8CMFgA3JzTFFsBsDLy0TzrR/qzVMIzqFAv6baCoUG7zMOsu
rcWB7BiBQiIq2AhbwSkS0ZpPAbqPsN+zaJfD3EMYnN7uEIKClTJXBxm7tmB+HyM+2KBMACdW73Fx
l1S553ZNdveSZSj8ID2RcEIj8Zb8DL7MOc7xy4k78/c6LMc6y6srOUZp+CNcCzidtRp8R+/fY+w1
iL+N9S3bbluBnsVrRq3z3S2NoDfyGPXo0KBPAUy5T8VGqIFOcWaWCU+cuvNuMV+guuLyutpM82EC
fXnqs3IRnQJs94DDVLqfdS+4C4Tb35fE5hj9gDTI/slKhq6zaWeKtCwBe55jVbgU/F6K+g71/CCL
2I4r+YqodQigwsW5+xNLQRTEToITjjoziWG5bzW34Ye88UDb2Cpl69sDXfYBRkahWDg1jK0IfHJZ
KE1XtXpjxwdaAQPAeXLDQGc5twWOe1VSCkslGJAKBPEylsjI8w25ukAHuIY6JW9zktsh7qYoMB+b
tR+nClXzIRAq/6UPfOD+bRgzUQPPriHnUUYfRPHQjtZaawPxbWYDd0/soEG4c9Qv14v94zfoLN6F
aAi1VamyNLNZt8tt/3azGx+gKTxySnNNUDAh1mjKUYsR8TGcUO4As5W9/F5IWmgIEWWIjhaeebVq
/6pVEnnEdndjJ5F+eUjdS81TQmVb8i3YlMIRcRIIzUnKD9SQ2Yx8ZPvfD3oEQWgjWbhupBMbEXWU
O/1cXM4M2QVjepEZcndfc/jlYN/eyCpQrgaQzUGUTR3fUZhbyrJ2PhUiOVuJ/Qx8rRyJ1mKJqox0
JrTxmoGjZ9WZo+vS6G47wqHhQl1SL1akexSxiXVS9EcETJbfbgLjolcqZvLkBXaUfOJSklCtA5NW
8WFNDF9oi1EIPFcEGx8VpSWFrkE5GYprNUREnLi1yRsfnqeLE1oofiWUQawXtu6+Pay8dcuz4H22
cWhnUerBWTNJW/FXAkRotofeBUrJv4zfggajEFCj3ImFH36HRA8UHj8ENzvadJ/lBp8WHOFT6Cjn
hWbcDZApC8D7HxyuxajS/rLHIFMHT+o9rAeJdEv679SXpq02WAJfr2ey3/E8hZKnx4zrgJ7Tmp93
/hjcJWNRcBTbRPcbnSTxrYinewm5BYxf/m+Xw65kh763/1rlkMbMWm/jEBz9aUVxwKc5iuZSRaLA
vqjWpDZX05RYtSblos8i83hTeNNnrF0AfKLzfBG+hmGJz4TbWFxioU0SmUs4Cs88a4TFlabdI698
95DEykLXzZ+a9SzwYsShxRPh6e4xiOwnms87BJXZFHiufK/p11g9QeLZn5Bzb8wN+Da4EUFbvN3U
O7udCUASaZmT6RYUWgb/IDvWa7tSA49rle3TV32LJYN3SwMfd5Wgn/2BqlU7uKJ6isvZVBdGW9g4
TLQL7CF1UpR3zaKOMN0r5u2d5BaaGgpphM2ydRASSMHf84f0WSKcC6DnwWsoax1mm+w/5iGvQkcX
TLg+pg1OdxOg48VHae4EeLNnFdOWiKiL6yw/QE089J9tfh8tGmG7RoJGoH80/1M6QYbdjSNiUN+t
oe0n8EcUpEsZZGIic/lXxVOYz8YfSVtCPUQ4jk+spYAxgBaGFDGaRWomjGTs1H9H4MjnziCEWN9+
vomVYu9G4H3L3y9tTd01rVG4iDxjz4WCTxl+ZoTBaYU1b9PKSGJ8w8ejrLVFYUgZXEXbsb1SQcys
jpr20bMHipYJ+129Zf2WbpO/xOxkN1xsYMTNLWS8m1mCNwAqlsF+NUegw9j4vUedejq6UP2RN+gQ
WcW0BS+FzI5Fiphhk5rQZPQZkW0YO/gPO4ivJ8xXh4bLhpGT6nmhhxQQU8nxo1KupyIl3+7EAbeg
6nT2fz3pMoMTrwMY/R52SFr5cSd3HeY7r6lVX+HpxpAj0jdBHpnk9cmEqk0L1GAS3GJQFRnOVJAQ
dLnnqdesdWpzX0rYi4DlOcx3UKt5iGLE8VH+1PGw3USDYTFMzjawkhaVzyZXEfCjSO5kCPIUTLnU
ENENwLlleL/iQajfOXDZ3gsNAp2b4fj+UpiDqgbLvdnihcslQdhrzTrRPGQNSDwoZz8J4KjHtsWy
CsDnQT6GLepWXijrydtXi1gJb20ptFqJlj1IAK0WEyvmKfO1jEUwfbYlsMIKrJqCCTs3TFlb4FL/
P200Qnp1WG860Vav5z/5e7sc2LetZY9BKUzjyBeD8eElTKNbUjtXeXEGNq6KKLrGoCNUkGdx7m/r
XPk+UoWgJSEs48PQvd2OyxEi1yfIuHp4uuCdWN74/ib4satkADvZKbWxCMCWGNfAT9ZX9EmdkyLW
SikGbvSNYBIjLlBKi6vHKRwZLeiClu9JMu95tNjdCnLKN7eNkbYpKzhA97LGyTKLzXtxgG0ieWpx
jIwkHqNcy+Hv2HUjpBxYdmCtIa6tQqQvAYC8ZPRziNhtl4V1uHQAfdHvy/VsdHboyn+g/S0zd+/y
iQlZ7sPQq2Lql6APkCF4BCfD+zJxRyxjzxdaB3QKaL1vlpP4MM0ehv4LAjy0nJEN51N8upCnwCqP
dsAqt4LyDU+xt6L8gKMKcrkRS1ooONxaU0hOaPCnVT7XewfyzbAzwMAmihZGuNJzo9IfXYnS96oB
ug4YfSwe2GxDvNOH2xcuE3YM/rbgFb7sZYYzgjlCgUy5rUtKllj2OFqaq5nmJyD1vfvAHvPGRbKi
cFtiJgVZr5XmBcqG7ptcQ32YzYtnrEnOiW9Jbl+4OAFJ8F0yV0WwkaJsnktJVFLrgR2f3e/ClcsX
rSGyaptYPSnV6ZDip3WFfPefbVEEeq/EGxAEmLI9Rw90UmkNvjda4nXbd+cKx5HiWVADes9zMZ3V
qtcvTv2nxXNtH50b11nqG/sZ8lwZu4ZMlvvrsOvmx5oKrFBRACFauBe4g3NqVe04ras2WE4LNoQq
aig0e0FeYngmJ9/GUvUaizcRKspTRJepEuhtymJmlHAjtWPhzQhXWIjBjAGYRF78iuHnA/rkrEOM
ljUBVHTo35CSN+2+NJn1TKA3k+XPfhL4Df7Uf6cFtpODUw/Ohgy0Mvj4CB9bzQL3orQ6aidij+7I
FJjLQWup8a4JmkfTO/0M4UDATqmuED9pqiMWGxvdwOXgP34v9mQb242McnqrrJ2pSGk7BU/MGWt3
ixOysJv/T0kXL4qw2y4mGFw42lANzqxS4dAkmcoZ8u3Lp3BX2gZMlW8uG6KenKBwOaCf00WtrLAU
OGNVLyTOJRUWdqcLMGoOnJ8zuBr/HQBfeMD/E4CXvl/vdjiaf679aXryaLNor5R/NauGBc90IlPY
/cico1wM66NbfZW5jCIQpehTIzjsMUP5WahU/n3btGy+ffq5HK1TlLjo6BdoDZoGGO0QWdO/0ZT4
zgMeMLxQlQIMFLMlFGZjcuJG10QQws9tO3gCZ10a/2yN3vf3Un7ZAMBngwsa9oWDEI2RL3yPAxoh
lapSu6j6YFXq1YnqshKQn23Zf6ioKBSo63NctDCCyVqHiNZVfuZal8THVshNbSVrhhKRYycDibrj
duCmlURVggcokLC6gZmjKMRKJcXJnO+Mjvy9XUfnRmVEBrrH0uRof+NHqJvnZ+r3SWLdZ0rc+a6r
ewq8Fnjwp1PgbbMIfq6XGVzF//GjY4r7kwCfaHtgkxCPja723470dPb8/wqYhuPxGETTwngjsIkk
jbHZzZsZf9NpwcDvxNPnVxYjnihgCLX9q7bmJzN6gdFL1a/ZzDPJLiBZOV8/Kz8csJbm7OFV9BGo
Cn3SwuAHqfOHYoTY44JYgKc5Ub+rX3WmobPsyboRQqmzsSVlyuMDDbBUxPapc860p+v7CKGmFZmX
rRYMVVYxFqbtbJ7IHxIS5vYBaK2TBq6iOwd5H0dDN81BKCQ9O9mEEixekSx5WvdRyhUwIuk2FTCR
b/JufgUEmrxJx2g8gWXChzbtDZi7UMrGQqGVPZATvYsbGMtXWRwDevkYLBbFm3g+5eZzuNxH/gVJ
SRAY3jRNOBZQTyaNfTjaZ5ltyfD9y7z9Z46SLPyv8v7CcqI89Z3Oas72jxOa3vx5fd5eMT0urs/o
0p97qzrubAfYKhNHw+F2aGIQXPujmH6+WH5z870jx6PrabGSEzRBsx/0mgmQ1opiAHC9nk4zLCtu
RoDuaHpSJ0Zy7xJQVgf/Fn6kJ7hOFNHuMPUMl4CKy2zQatIDGWhqww4jq64FiuAlBYSe/QZVLXpO
Rktu4jZTPCW7s8RbGn/HmQlhjJ2sTBx8XchkZueml4weZ2phkol/W4dhItr56pM3N3MyZ237OwAv
EIPwlMykqQE/ERVAYFopp8P6RmytCTyLfWGYVwaW57gJB8N+YF1SWziBTG7TjEd7tlmW7zy2ObQd
XZuZxFs02PfHXIuRLjZfuLaB8me+RUeitEqmu2ZuDbUngr5vZUkOBYupP36EXalsUB9icC5dKDxs
Y3qD7Oeh/wGJiiPqrso4p4MBbsWS9h54mTkeKIZyblSYInHLT7ZtReIN/gglwMZsx6w/mcn6qoZQ
sX28VImep9GWvC8qsyu+otQKXiQQR5jN3F1jGWuoEpazCvRmv9sJv1q8m/K9CB7n4BBAtW/TVGXo
zsRRF0lwZE6i6gQwIuEC2sJiezhZT411XDzIaeCFAUnu/tl1in5Kc/WY6l4UpZb7ae04+Mlo01fW
7neiYQVnxLpCQTUGNtHYvJRQtd60KmRDO1+RuzS0yVkWW3mvvl3H1LvBmmy6H78E1eW7lrNIxmo3
te/g3B6fMv1+NXGKiW0s27g/nzh3UFZh5VKd7H4RwSNz0dIc8oxVnshewH/ddR2PxtPgppjGYIaF
zfyAX2FZqY9qxBmkU2/dPPyCJ4/aj1XniTxfb+mwXBw2rb/R71Ui/K8agzDEetZjC31d2YdrJPnb
FOC3TcWaCrgDzZkkABXOD+S5oBprZ5rEkKqFEo4xj7FNR5YlBP6Afngf3Ep9NZ1Jkx1Qu+m/4Otn
Fztwr0MqVVnyg8uUknPCxcU5LEbnsMFvQnK+pU0qAuUTw03fXe4v5O+dZ6WycpGnoveqsh8jlF/m
uecnz4gxHJE1x0hlw43D57qR2YlueA5GZCMOuwKt4GGzr6dGJo6VL8QL0JAvMPsRxYGCt3hY+Cj/
sX4FXcZxAtovLOyHfDa0DOEJQbTOuQBqnuiohJXccCGvnoCyFBEPbgQwsQzOFt3ixQjjUbPrxbOh
aoloo3/l+4XPAw5+O8G8wuTRxJ2JrimsZ/0iuLTglN616Q5VjIHIlvo5G4VmN/cZ2Ctk3MeEzLgE
7JBTkxD4Ek7GXHM7dB8gf932T095RklY1L3JRz02F61nMw1X8Zf5PfRyp0+xdqhPHDZoxRf3v36j
GdMH74to4jHIeRklgDey2EW1Kx0pOWOs3hUUeDqscbAw/ZsLW6zR4Rum9y7M6vptBOeC2YATsqFW
p4ZOAaXxaFJntdhTZVLkK5JuGzAGilOE4ohlK02Em10KpbJV3+c23VHi/CXFlVpQ8WuPFEe/NczT
R9ahYv7zprofaEGmF/WoA3gh6rydXwKINdKk67rGOJVrBlOPourFCJqhkNVMA5HsLqYZP2EQv1VV
utjJEFJH1HEcS+VRJ9MM7IGTWJmz9bFJ6UR6RqOFQnHRgTnldOkdCNB8uz4X1ko+g+e+38sIpCkz
VBrgwdK7MBdxjd3rNGZJgZlLs3694kJUWjs1Y9bf/BVnb1UL3vW0Aweph8P1MhD5vXfzLfL6xcMZ
F0MWOaXsDBKlTnN4RW3HvxWa2NiVNaXkce+EuInCpuKXFI4MhldWVAJT7xKFXsGj9LdwBn0/QUZQ
7Pp8dlBHpIexNb1WMd8wJywKJlfEyTBeAbG2/vFhjAY0JHfhW1aUj7yAhpFpIRWQv2fEqwrFLbom
AxoKil5W8XwC33NNAYZp8julB1sZfBMf9TfPcyu9EkxZ2orWxy1iCLI/j1sYe4T6NFiTKLtN4Lsa
xMOreFHiVqikjOkwfFWzQ9xZKxepPbAfdJauz2XUNkKxJJg02CS5ctNQwy0f/lSSEUHRamYe1suG
MIU7iPZlHe8fhwMI8olS2hMXblEQxIlPTgeDkoG0kSdBdbZ/gZUr5Xp/PmSC30Pbqm/CDXF+H9Xz
m2EkvZ4df6FoCavSARqryUBVv+cjPUojsHgs+b14AaE2okHudKyeiFxAVTu6Ux5CwYxuXx7JnDgu
LsVUk4FOXDZkv700XxD0LDjfLhKOJSMWMIwhT4+/0LxXICFFw/NvZ9Jfu1iT60Tv4LytchHavHB1
vFchFSHxCztJgRZxvS9iRro633+xOpAHN3mIngX7jsfTnzFA3edbNK6laOQFHOrHE0/iTTC+BZrY
9ZOs9uCkC9yjpStoSaeMyi9qJAKgh9B4KOCXJH7/cjbXqnsyL4fXRriX3/J3y47vLS7UNESiDuII
NSEH/jDJ+DhUqrRGjGAusiPZVHBA81Ax3kTo81eTGsYmQaGaeqJHsmNS9qnLqAI5V8PwSVo+FmK+
UtueJxuVCZ3ovucRqYV/smH1mc3YU4NmyzwYBD2ZpyaOqH08RU7BP0TsMPvNZ9uoiBNQu3T+IWZO
09WVjcQ1V3QOAXpn9tKjhiibvRqOjMJL8Ag0YXrJZCfJ8Ix/Z+PA0abzGaIaPsLJSLysvD3IcKCG
XdlMY+ldHi3PojYGk5JzrLQ/d+f0kSdtFcnX5+Yqoa5r2vJlX1FSQ2A5yN4YPVqWzUnfo00/IFK9
n09CRiDfvqTzQlGI5hxaU8slSrYUIBVoCbSPq9H8Q7O+kC6TUFe0CJJWzd++Nr5n7vlW4bjpT0jY
IdApwOLS0mYn2rM0lKZDPBmHOhHiuqnn9ForOYxGiEgfjcH38JR6Azf9Gl/EBpVpAYoCoqPi5LOq
YZkemhFgvzcWltmiAg0/XYNbDuuyKNgEFWchdHjx/aR3DRe3nI8PW2gT8kuNcXUWAWDIyg+H+foC
anXObEPZ6dsOKdCXEc8jKNIZqH32zQvtkCXJuazqjLuyLUFpjy9UvLukMp33YX2IsjXcTG5zomEQ
Zokl8xvDHHyX3V8wJX1CFER1neNNbkTkm47V/lmlE3pl1EttG5i1DU6bjmyl4d1lPNdrsAyMtP0L
p1cp/z+/gYs5Kgvt/aAH9HIY9bjb1fpjOZbqji+MMUii3Pr4gDN6TVbD24uP/nbPP6g9yDRUDQDw
4VEEeGkQZ8pf3FPFVPthlLA5aIOqzSbo0xmxrnKAmmaRN4SLt/TDxuqns9X/q4DMTyvqTwK81Foi
fRm6RZnDjRmANdvxUtk2Uv2MZ7cnmNc5hPsbAoy8IDflri0gyj4xheCaiRw5wCJWx+ikiMO+KMRR
Hax24gqtCa/d9y7ya5YbPFtw9t4TDzlkC5fIYsGr1l92xTHmaGQOQhtFiA8EwmSRAuWE/GEVnaAq
rc12+JXzaZMnflHzAeLvIyS/qFoT+mj5vyzxDQE+mdW4yYVZYDYA2zpEQoE+EGlYI5YZipr8Ykoh
V6b7AKt5dl+RjJDq09r0Ia2G0O7a+JlWIfusQJCz1LXbrpPC1jfHyka0+RDW8vJtmffqb7NiORr3
2SSY3VDm4Z9NiycLwAn6mEd7jqIH1OljEhfnqvQBvqMEeo6+k6FkhqV05zf2U3OMJs7ZzPoBZhZz
kdaXaw2QXiolc4DNbuXxXrt01HTl7ZpUCNMUqKDQ+QHVEq2HiHof9d5a3J14f33jAuwbOJud7Ns8
nJgFo/QPDM2ntDMWC2D/PcMTkpxj8jaFOvCoududJ9ZKqtV40vOSJ584956N+Xhd2oVMlk8UljC2
uVl0UW0Ss/7mKANpAeKUL9ACXCUblihZOtQMafyuydx82ySmKgY9Tw5XkDwUOgSWmYqs1csrwAef
Di8Xq5t9lVZOprFO16JNYjkeEFCsCrWjz6v60q+29GI07/SWJ0ODcd8es/LRJSv9bodoAyggWBlO
nO41jQuzCgZ/eZH3Vj/07rcFEhcFi/nfnlUe3T0lPpSV6YJJJYjQe9myJ/1zui+0KoudTyGo20PX
8LqEU9dLMOOSdwcCvy61l0+5zmR3d8NtSGO6VJT4vF2zcAsavgPRZ9BhemVBNEmbGzueiMrQWOwl
oK96PxLckiY4487ff/BMzKznbqVKYjJf+rjRMIzDO9x9UrKyB+EYqy+hiXLbg6rjQvyl5+xdulpH
2EdLCdLVEhuPRjCpuv1Fx93vkyL37A2XLMMfuLG9230+qJyI8+dphf/EZKvIm0tUqHssEqWh1j1W
bZyyGkqlJY5sBS87zEkUcaG3AsH8fehK5NUG0Ih49httJE0RyjzUWIj8x7AnEx7v5r/psRFhV5YF
jQsjGc3x6OQEMAifDc1qh2kb7duvwPwxcKmCSn9a5z29iVXDF9WbSFwmZ5S25m3mf9cAL2V97Mhs
CZS+c7Loh8DeV8ch1m1eMbbqwTAiDKlbPMSqoYBLvUXU6xnyRzDtJTIODyOjXlsuwOmtXEtZ1yvo
0WqvG3pHRERcWEf/MTvsOGMbIIWUL1JqQaN+Lwufn82IwMGyNYXiRAUycUbifvEV6P9HKQRN+/XE
kdgur0BD4ZrY+BDP4wfkWZQmFo5P3FqlEIsM4k9qc4yReKaxkEkn0s+9mLeaH7nnAptIXLcL79AF
9VOU+RkeOx+WAT979z+9cxWO3f8ocSQBnVMgYBY4AWiy0M9rm35hr9yfqMvW61gsZDOUCG/CpaNU
QstFezx3V1ZN+njxk7TqM1wQpMhGborNeQaOdFc1xBDVR0bqug+QB7Nh+m4JvuiAAM+ZNsPcFHEt
Hu1HnIy/55S2x7HcTv0XYzGBfsjVUqhH1/nB7dKmBVQc5H5qV91d5guIx04BZkI5cQJ8HuhT3VJC
THEMarzpOQdq+5ETTTRNbV37MIoWv6mqpfgsY593R102kE9zs4JOcpXPkvSM1fHl0V8JTbLEfd/z
N30RmhUii+UA9HlWSwAsvLQGl/59RHsa+JGQY0x7JRsvYRlvR8Ak5yRWBLfS032vuYMJFL57QsC1
NZmttLjf7qmoHRnaiiFZvnDIRG1lpEj0TUWFIzs5fy7pCmDxc6ssY/mq6ZCPvQ+uO2KEDFODmUSm
gNt3aU08sj3prGiwvW5KOByLeHrdT+y9cbNZk9B0tKDkzJe284CrnKkNeeWPy6hTakkBCZfx5QmP
uywhktiMJZo+/lS1xqDdifzRxQgOARufRd1SFphQyoVifpC75CjulBDZFoPHxg/wwr9RF6VNmHma
E+3kCwsJQdk+UshDattqeqGfkIeji304BenRq5BecbBtJTySoBBiYaw3BeLLdP4qbsR9bTY4T7WL
SKXO1/s2Ux3PNNSSfl7pXw5xO6FXp/KjIbVy2M+g5tdc+TjQbF8dkqVKuNLXl3LYN5wB6YkRg01i
V2KtX9590LvnyDK5dBlKX3qP2us1fDUSwKVNhkhOMSURCDt/R9O8KDKQeGmlFDkSl7DBWE2h9q6f
PVC1enJpjzWvv79d5Htc4G108naYHmrtiss5wseY/ZiOzIoBPcmRwwgp//wLqXk14CNoP2B1pw9O
vKuQ/lPjR/88cz+DZ4+Yp7VdnDsbYemxRDKrHZ5rPWHXWvUFUfZKV6B8drYwbZVG1emIei82p57H
V5sPYTMLDfVDMp+5jHLLkrSoPWbVOZsoJ43/wIr4eVrq2itz1qkHpaR8p+KMvYniA4YKxBhlJTuR
wW5rs4X3YfHmVYMx0CH1CYVgQPx5ODCkij9+2LbECfxgiUyYbXzkwW5tP1XfOaAlOYsZ4NKi/A6X
fqRdGBnrBOptbEMlkdTpiF//XTQ6TxGHOCEVzf9DLtc3uTXR+J9gYcDurtdksJToW0filc6/CHlG
D9JnSOB7W4p0ECvSs4GkbsjzD8TNEx/ND2RPJBgfoZsSndbGstoeswTNT+DokN3bx6kb5uJFksD/
bFNnTulUzhU+kcselgVdXOzSUUtcOvNqyaNm4i47P1fYJx/gN+YWA+yvuZM1Kda8zrAcDl1U3m6b
Tqv417eJ4hNnHzeJaV14/B5WTi2Tq6MOgRTP9wOVReJqxuR8qW4K2/8Nwnhk/LfaDFMH/9DM1PCL
MQVaeFTNC99CX1e1HShovyomwbgiUNqekWGj9pbMC3mL++ifmFmxrJE4588VeuPCJyAjYq7B8QdM
N04Cus4Zs1SiP6r/opiX0wR4EGnobOxSXKfqnzOkzD7PnQOQptDmozhLZZw1bMKnLRpsHDK4XomI
8M3pmDAyW1D54xS5VoYCiPWgOOkbmCRy6kbjJENLxJCL3UlPSpW42TYmaDZB3K9YOnl/GYD4K55z
vehUTNW3rcJ7o3/BtpwYa55XAsCya8whCkiLJk22OwmY6hj8hWeSsOsICsuVoiFNmAj9hRlyTh3C
QXfB/59rp2436Tm5SxLSv8Y0naHFbuipmksHkmdYZVba8DFzG+HV3rykEV+j0USxIRzuqJqViI9y
wwKhryl9dRHiYnV8LC9S8b9dI7ira38LmyVFXrTVdumFioLvFeQpdYzMFRrg3bB6M6IjewhDMUS7
WY7ytdFx4AhgvOmId08bF7t7/V/RuV3sgRxQrYhxAlnKEk1JhS2pRH3nQq1aJfYE9+DE75NSuwEK
rd+sRA8BD2/Qn4Mjmh1ineeodvqDcMukJ5t5YNVL1AlHYD7m+klsGH/OqPYwd+aj+xJnSdUhCdyr
VhRUPt7nnjiZTdy3PkaHOL94DM2DnPnfyrVxfuFqYfB/0iC73VsErM145SBnh8/iP4FVdK2vjy+L
yVU3Qs5Wj99wsHMHHY7ePFAfQI/0qtfsdmQKXFPTE/LyEksRRrtWhnk+LZqIjXByeJ1kTEZlrURm
eLQRLTDkKr7/RvhxxKN7KqpIBy9JjWsIhzE4sfbAKnBqJTVNQlZI5M8Fp+4cvS0UWq3kT9yFaR+T
UXISPAtcyeQdA4z1V14C6yhy2FLoFKVpVbwsE7DgNj+TABB6OQwS3358Ubb8gHVazppQVNYn2VV1
LV+3hH8k6iz7GfbceYND+TEsqv7/jGdaZhUq+vSZ1eeAAfkyeIAqrP3K8hh9GU3pfYuoxQWowxdk
huD8evjX/3k+gtjanDhs1YG+9MOEBz8H6LJJs70u6ktjOJioqmTv6R7hVBh4ngkb9OKai3juRC5q
tIfzmM8jmg3Y80hqcRDo0H09jSG82SneiMTCNrjwnwVudy7CDDD0F4FkRs87t6OoH4p8U8WQmXxM
bI1qwd44laDuVGtBOasQX0YSo6GZ1IjPgAKyDida9HjlQVOB1sOl/TSJ8qqadXAXsR7P5K1Uri2J
P2RHkW13G+OKCHjD0VRW231wwq7usCytuPeOHeAix9GMbN1xO90DtpoHn8SDCIwELEb5aj+gm236
NotEOvZQ17hhjjxphV49navSb05uEMWqZSdzr68r4SZn1GJjm+4zfmJ0M34FRX3BCaUN8GYdu1IM
ZLMTFfDW+1ZzkBnUhvvy+r0TePTFtYnAcLWHwdxzPXL2d5pkG5ZFsoLT17TMgFXkMEwOvcZgAPaB
32R4sLKuRnQh2oSWlhdwtOnu4MCcLOqrZkndFZBjsuYIMV1BEHB7nPaWpatCcRp8WgldNwYKXZQQ
VD1fdWZCIpSfyyPe+XTwul+A4XpQS2LVj5O6zb7nT9cu707HYS5wzEStEGM2afRo8wodISpodeY0
UsJvPwTnZYy7/C7jOF9AyXpLGbynD5CrrrC/L5OyXrxaUGwUYpdcspCNMW2UYv6LSR2ExhXfAdmd
otfN8QnzZxKUelLXk7uwfWsLtc02H/UwmXAK0xfCEhDdkbN3y5y82dl0uofuUO1abtuEeg8gLeYN
pUXpvqtx0hv5geuJvy/cABgiQ3kWPUAw0KYSK/flEJVqPCWVTB+TluP1Cy+DcYwhEXI5etzSmo+p
N6Uv6yBrI5P9szJ3hbHZE1fheXwIDLLRD/eG/zxIg39510AQkNOx4rYtWscpj2XqhQudbWwhGAMo
xCAv3BR0cUx+kPJL05419dyGba0WPXWc485nA9MfTN1LEJhcNHa7q7fgyRIyPlGp1GC6KBaCYq1n
z7JuQmWrFhnKyFIMRTKJUpGKITDRY1Lwob1TqV2vPfyNtCE+g5FVQxkLYr56zuebBWRaU3jDfmn1
cuu22LshsvcRgiwt7ovXixNjpvoq80KJFOYB6faIrIMavCsEtn1Z4C+OLevEl/yh7XqmzBYcFvXN
2bP9ooEHQc1NPCFAh1tP1I8MQy/8/ekM9Oqt6vaTWhUNoFMQn9RL5skNVNwNKtQ0p2aYQe0J6GfR
0/kVGpVNT3Z9YGOUW7XrxupKYpmVTaVLmDhqXb2gTv3gxilYsFtGEtyGTqYzcWZhMZh35VgAeI+Q
VbzcQyIuiYHo+usQs2P3T0LCco5aD6DxA93qEughQi0iSLb6dsWGl+2TRCQ9MEvzzVeGkIJi12fw
RFl3QXJrMvzg7zQoN+7ytaG5gRXBkQ2dzKXY7EjHeSUAj5Y+yQbRrNrYULhz1Jsgkm+maIlL6nan
Rrdnpdz8RUyHHgW0KureU5Q+uW5GUVOMM1J5RnzcptNx6qxH2Qh/MdDeJKIv7uBd3aFLupmzKSP5
NwukenFH1cPXS7QifAEoGW/RScqZT6DQyG1E7BMMulGFr067w/n70ue9xKwQ6/2pcuOrxYouhFXq
hLgi8stNj4u3b583s6SFEH+EN31E8O6/ZH32N9uwTMD6NBX3wisdIRLDln2zdXcE2VUiQqOs2Hy0
aaYchFVspjyxU3h/rcAcJKVtI0AZdqw5FBAZhnaNBCs4meSeTYyW/Z9M6mlQkiThm7QKUUKNL7U5
mIF6SRosNu35qcKXeYIeU1Mi4YwJeU3dFY0vpB5uk8BWd/0JhLptLW82TZV5YBT/lhsIczBSTKWh
QSFOpcMVOXWtSPEBPkIDo8Lmxx0rtvTcTOWAeFiQohlKtDtEpG0FQmCgkbpoPocQTw/SZtk/CciV
TQgFLZVyyUa+MZGZP9Vx6z7kFloTCvs6jt23d4/I7ZdSjmdZ96EJ3n1JrwGux9OWaTb1kQAKBA9D
AdcC0f/zRgC4hq6W/LQouJmgp6NV/VH5eNxZrAD84JcNMRRzUCWQ/sz141IHibfOSbAZ77FmoVKD
7tLYb0HAqUBnaOnSg71JjvVE3F6QnEmer2Ne+hDsvBl56QvMF+BL9hZJ25dpu684bbd8OFvPh2sf
2Tb1kqWlXG1m0e4M8+X8DK6aoh2bFQWGay/trLA97CxIp7+b158OAIknq9hBHyUzJ77FPidsjxX3
NxkWBDHXsDFV1Y1DQGpo/K5KluE6bkD73L1oF8znjm9Xe95IxfLzHXRFpItLeAYuUa1pCYK5+FxR
NWvscVyrRlsC7EWtZb/4XQM78Titrbi6vt1hIzMXWV7wPEliZRrmclBkDJ3LLj125kMQMy9E7o0H
josLCsGBiwqjkdCItvb0DRbuLP0BJx7CFhGsndmSy/0MLpfMwV/3KjRvLGW6ATnyswPOj79cdjR7
dASg/D/sW9C5hvccrz+X/SGPIidhOoEdS4Ax9q8YgClCoozZ+Wfv3x0+3GTW1aiicGYxd3X1F9xZ
/V4U8lpPljeJ+ij+rrewrhPTxuA//0i/SiaiTelEEaoiG7aGeJFqcfAzdm7YbuR89C72Ni6hgfsL
eLC533Wa6IJsOlVPQt4v4ACkthJOjnp5nzAjtw3/8B5MmrP+LEOtG+C/ZPQE4VYeFua7E7eesSZi
IneM7SquQ5dJbrm24hzNgYtOJeZ/e26fbqCEWP50pKZqJ5QX4akgQmSjr6xZFISdbE6QM4bPDvpu
HvwqpHR6yMz9URJnA0YBlR/9sSopde0IN4NnbcA2YKlETsaHWLMf6hjc04SEDykaVwZeN72mxHg4
QgRIu2K2A43Ju25HT2q19n6XowFGKn/aL/zsNO35A5odtFcI9cW2oJpxIdJnpdy7LCNfmc167mBH
wjQwSFK2zzn9jq21N9ylc8LUBbbx6bomfVcOV23V5gHEaqHqNMgYXHtiouexum6oHPneVsEzkjql
7desqUKfE9EPRif+MelOr7VgoYPmXB0ydF5EExBMP6kLnv5273q9A2jI5ZOnukyaFRLg9vZDFr6k
5ec60LCvh1FsoWDyB16u5a/KHIIlqq5+jUGFvbWinkRUDPkFEKOfq8you3UFF2YWzvmYY1FXfqWe
8cfzMuzdeTJwSKd486U7YowaquwkL9BBhxa/T5SGCFvfjOSu0I09q0ZsGgTWbpktVOo4NWPfiuJx
irVOVbO5Ka45BdLh3KLY+zjcIRbnf8N/4AYPl+tE0oWUYJZSw+AIfi7oDjcy5pvz6qIIAqwltwFd
yvRG/1XPBNyJ8BVi0dbfpm0on0k1j0ihPtwHRZHhAXMyg2HhoTXTe5dMPaqfj3KlhlHFZt8b1Nca
t2O5h5dnDayCA1nhAyl+MjrBvUAi+D29adoY607Sz8E1oeVv0Mje20ITKizqHfTm7it8xDFxESnY
BK8ttd2xUvO23NHgX43NXikaS50+NcyFaXqNp+AtdA9g1X7WOux9yr02lH5rjJk7IzSrxwy6OFhz
LwrCaURvPr0ETl9lb1yp6JkcVPW42e+mtZLbgUXXnthWogH+cx3a5Y/Lhi4lRVhSb39G23B3ofCZ
fX4/X8cygl9gN4i+3/4l9ciRFwsb/gYuPs6RCsW+uyECQeHlhn0L+K9nI1xNnGirLoAp0RlhfSw2
tEYoOd1GZEiIpDuqxrBFcW1hbVxCpktd/JR7ofSHTfJU9+Sexx1Infg5m4Qa9lFtNo75PvB21g6B
mvDx3Ai7B2GXvZk8Qt2M3bPU4pX+wTLXenJ4Y9jpKUSOgrARp1uVg72xPhUk6dqermBU63MiA4df
Deo1vzhPTwJf5Vdy8zjXTGBaH7UM4KkPfnm4tAJKaamYO7IrtCbFQLYlTbmRnfZ4eUpjkILMyRLl
p+XTieuC6LcWGRbiYagyj2YSJdsE2VWNnNn48m6nn9SRB0ihp1t/jaU9INVgCYAhOhlpjdYjyGga
7NxsUrH7ytl/BBaus0/FJKqENeBLUS43LhMKuCu38idLHAe4XnZBqgfNbYOwSahXNNQKXU4pUSLK
oF4oy0K3wgK+W1HB14QHoyCVEpQ/FyTwBy+W2QyD1dwkPJ0/Atc4gu5ee7pVfZj7am6w+Dkkn7EP
g6KET5+zFZRn4P0EtAImAOMKp+MsvZEakK2fsmj+14lvBLsEEHo634g/GOv29RLICJOS94sPZjId
aOAMGdcDDL64tX6JoCYfzoE0HHfPYdvgGZlA0UUT/QSXYIqHsqvenAZbx/b2847fuYNLbs/KZ52E
gDIoW78qTPfqq48PiDdZHzhMP4RPBGbgMnUhvl8KtrOP93XkVQgv5G9knY6fBu2M/V+c/Rw4oVkM
giHDXZbBKHEX8HmkDKE8M5e191kPGiK5KKmZ+AtctuTjd/ThQW3EsXNzPHywK60g2SaVsQ0HO9fE
lhUGlmk21YwZ+NQX3ujUpvdbFpVR6PE5Dl3Y9tqFUM6zknS3wB39+7anKL05GzVT3QiFqJlk4EfF
OiZ1Gon8R03loB9GvMnJZnSSszoOO0FmFQMB50ShPJ/3aUIBilRcyX1cLm+bZVEDCCoHWo0HqvFP
qB3/GrHXfs4Y93uCuF2oNlzWJg3ulMlLcIQ48MXQXfsDoDUffaik5gBY3+d8vMizvqCjN2lTLyXV
72fW6dUNmMkhRcw7Wz4/aYzSyeVL/zQPb2abhFCpcrNExqEgpTTB4WIkqq/Y2E6Mc5uX1ThpgKRr
58MkJ6vvXqOf0RUJfl76HMKgKbERbWjrTSvWt/o86B5lWn1+3LX2HnO9n670uu5C5EaSQZ7LBvQ+
1Z3X07ofU/iKuh2ZK5hldC2sZVRIU3J7ezAp15bhLMHED3LMwUWH+7t3jTe+Ra2UnZco7RPcQi5+
5VOLbxa+GYt8AuyKAUGpnRtTz+NKSxs8PEjN5ZwwAZKLKgyHKrKwc8niBBJzCqEFs/QMqBp4VCsV
tQEJ1UMT35yuhYMU7j084Qt4K2JozIBAjFLMTfdWeHm0iSDiRehXoO9Bb8DQw31QsFk0SzujEDCg
SFdLJW+7cT3IDRUwu9jb2Bw6BAnK6DGbJCTVWu8DDV3+unKjHjIAwubWJlEjoh8dYGxzAegwRYKJ
ol+3oWV5oWUrVcN7elSxnZaQ3kOU3nISC4ardsAab6dqaA93QK1DzGDlLEuOysGco726YskJlHDr
LSRcFweCXPCcUpl34rXCs9QxuZfzEqFy23HvNd6BOJ47lfYGVWB3UzKjqMcxaKSEglWlXUNgBRIp
B3wfajNPkVJthmU+BQMyyQGCCT0PInlTrtAnT5NKKgQbTAnnjO7OPrpeE/Ul7n5lUFzOG6XACYsh
hFxqY88EyLNUQdwYU6dxTvQfYzTt7akAEIx1Vaj80zTVWVNO9wL9VRTCVVGZU7om6hNHmVZQ4PZJ
y+rY+2AEwSuYdktkTIJQg7UhCJIYQQIl3mtz0x+6AdalaAz60fA/QA7iNKQbrUeURJ70hIhZyuzE
eaoljQ0jhC923nY9kg9YjDy3sc7oVyJd7OPUowSk5I5vX9+1ievoLwRs6FVaoLMj9plWQzssjzt6
HywHgzgM1rFXxFo8RzWslQ9I8K9jama0OeV1HJgbmtnYRt3qOADooc9aBTCgnhZgch4/wSOWDxzi
hpJz+5mh9If5/C9wG/+V+FO8aS7jZJ7Tj8cUB0TvSnpNAFzelBVreF9HUDy6M9oA92pvaSiePZjd
9HfDf5hQzQXMbfvn90FMxWWMWHqyBodMz2ZflSiM6oyEAh/nm6JyLR6rCYQ/IHX+PS75zq273HFq
ExKjHifhGP4bf4TvQBg0rSixVwmu+TXLxVspHCuAHKS5VsCIlfefMpzPMV8e7pUgWTnomE+r6urE
NYjRO9a1B8Y6GDqwabYV6uTG8UV7Sx7D/y3iL9ZdcNkG4EoMJZu3jmsTdTG5QSBmVjmN9LT4RKPf
5B8p20npSCJ9hq5x+rG6L9EwjFsOxWC3xuBKMsBA/hifsvTbBM+pX2FavY5afUimiWvvAkiM6UM9
dbNNJ2hrTYUEiRX+7Rk14TH7M/6Ya1w+sdO6LV3cLHOOCaGCeNEx2Thn2KENdVfMoc9KDgmzPmc5
KBHxszFdc0dUYaDL5DFeE2QU9PMf9DJnPA3CDFfbYWlc8tRc6+CXyLCOOnXSI5ySqHudMkJd6anq
bd30emD6F9d1lP53+MurjP87192lwzrW20MH+6FYhktxxZpcGBAYdUx3LU3oGZcw66owdKp6hqqa
owGTk/4dNuX2z2aKCsR/uOwrIObpfiQwX3J4TCzJdVh6tRyLXjwDYmnvx9LGgCnyYpjBkx0cSWxc
qyrzdbrNw8MkWUQt9PP9x9AeeRki/XebOlQ5GpB0gIU2V8T3L52hk+5GTIPCB18gh43O770TPMVU
MYNNeFcHYLIRsWNh9X90GeFaDcnINfYkfCQWV6QDyr3cKhMAwfj4U+nO0sx2GETQ5k5yLTrC7iyq
B8bYKkPK4Q295D3uN6bNnlpSgenYFvc2ujvphfRMRgCsOQjt2DC8U56Uy0bNrplMmtjX6x0qS+9a
3bZ1Z8SvLfrc+LfjJQDgRN2Ld2RLkFOPYNZcd+BuTY0cCeN5x4ipDhFsY3ERU10tHoSYmqKHOW9m
cAoL9x7N7dq1WizuD7mAM4O2MZlCIq5BjdCMm2tNIkJXkJoq4atL9cJce7p79rrD103v6CaGfpry
d1Zv5XJLh++CN3nny8s2nEgBXhFg1LYlOHMck3QPuTNcjgaGBaGkCNtK2KqwOvl3b/kQj+Ed5Y18
9pq046TFep5cyPut+tcM8dzfxbvqyVrgfdpzkzj/nCU9t3DHnTACJc5+8LNX6j6aJO9/fDOQxXUs
F4kW7s899OVduHYyM9Scb9qjsKorL7pEfk0EFWnyOnRnRC31Uet8EKSImzE9705Qq9H7KuOvkIqD
mqoRCte9KHFpGpkbP8/9029NJ3IyLSOupa2m37K/lDKnp0XtJiCMkXRtcWyDYDOWcvyQopBI/CoL
V1WKT/Otr2J7rw4G7m64vp73I5V2WymdpHd8urQV86W7d3yaBYmAm4SypCHiEDL/39unLcEtz4tr
nkeYUY6jG3ykmnvh7Omq2NlhqGm5WMJ4BhSoVlCIS3J39ZJBCVZ/mYD+dhQxbZtZWlHWE6MXQ0wM
Rpe4QUmeNY+xG4Yc0ebSQ1mdU+kELbZzN5BmoiwZ/QNat33dmrwKym1rPhHxK++0rHi2FS9hKSXC
vwvsa0QY8T+lpYMS9T9k9P1pkeH0YWNsY4kL9mrmO8GBXxnFMMtANBC92Fy0z1atg2exnt2Bhi6t
cSg3nn213qm1QgwihtP7fi9cn2MW5JcYtS0BbPsDdPQbDSV3S/d1RhJBMRVrp552A7+VEsKgG4Ax
NgTEoKlSIoxmooB4wWFUzmDN8Hfvaunx5sGpI6RpWcr9hQ8k2UlJovK11LFwofRJYqzxk6o6N0rW
bpLO5legZJsbqq0gjf5UsMYCZCwCxgaEOdLwgCT0sizl8WTYbQ8kuYqNypq3umm54lrvERxodAhe
ea0jXG5Mer971FGaQe6EgCNZiJE8A75MnpU1q5qPtusJ5nVH2WTL+xusgzOBneNyaVQ7E3VTEN6h
4eb0iy4I0Phe9zGpWbq1YpOS1p0v6oK2vV0YjXFk6lqnzyitKdKAOBEDw3pPp79nXAgH+P92ROe/
A2qeiaQ5sw7WSJFE4Ukgx94KF7WzJah9bJ4VWuTjzYKp1RAET58ovrhegGhLG04K+4ZjcLg/cL8a
5GOg2wHlLD69Oxlk5LrZ9IGzxsvruDmo/Ou154JACpSY7EGTVgPPN31bQybKMcJG3eSMCvSIlXdU
ELooqjRptKSQ4XX4SVMWgGb2KPIKP3h0pC5mTyRYIBwGm3nGm9zbWaApWg5R1A8Gu+R3/K1cYRs6
XSGNpiWHfT3wVVFmNwYLQoC2xEU5NUfLk441WNzeatXdJzRpC7D0dT3yn8Hla/GybwOZaiQYiuWD
nIQwi2GT5n5UM23uRDHOIutKHoxuD1cbfPiGBOXvuTaY7prOr39SQK5QxBAx3SCjMWNvucTtiWf3
5sKHr50R/4WMey0mYXaGQ+fojOXO0u81ZQf/F5PV3TL3unbKyK9JRUW3vE2mcFh58B6MXVbHcQAM
MuH2Eld6siTdiSN8z9rVXmbqew2RphLITEIIqFvAGerxp24ZFqhEFwlnDcENBpi0ebDejac0IsYT
S8et41529v50l+Gkd15+25tRlEAYCfjA7Up8YwU07e2M8kcEDVdk+BXBiG6a+UWuQjhiW5+osKxW
rCjeGuPkHbKuReyot7JuIXEL55bgWmmS1/GozuvFuc+MAXdf0ZtXBFnMwCW5lluBYkQGJa6RnM55
LQlELt8qQlyqku5LzggRczDXgFn2h2YgEPs/nJamoRc/d40ZL9lOquxMzyutoqNlHR7nP/hvLdGe
zLSLbzKp9VUEV2UV4g7TwJlx7CYn9MvIeX+iYW7yevo7alFiIqmg1Wj5YZILcKyMV65qtgo3juQL
j5lUM18v7R11/q+Guq8ahXV161QCLr/bqp7L1jdSPovTIcsUgYMxKAOsMEOeXvo/UTkB64rHdenx
bEIh/p1+mfQDEMyf9eQazGPDFosBnFYNprhzktTnPr+yh2sVPI8n4XaAhAAzf01xbZdQW5/kiqnM
hYF0R3GjtEcKa1v8l+6/dWYaKkor0x/i1dZm1Jlq/JI4lI1tsO7Uuh8fTP3CQHTjt7q8C6QAnOjk
cbmdVIQl013CKzJpLQ3prGKvZpXTZgBWYkq4vSSvEBfcMETXc8EWnM/sE9D2oPNfZU38XCg8FUnm
9+Jxn92tbuhbdCgjc/egIDTnvQ6dYrKbKNgT/SdRuzJe5XMqB14MOuPHPcRg/GfUOO+TyivM7zOB
6rXOO64NoRQN0q5YD1fNTfhU80p4IvC/HWOm+w0yAak4gUC+OSCC6CzwUUmzkoHf/r8V2Eo+Nduo
zj7moa+SIHYKGveutb8Vll+Dr1EO2m+IVrJHWjY50ua4XD43/aO502DPC5sbo9gDMvK6tg8CICB+
DoDukOJaBFLMeuyFunyJwCXj2bZehwkj3k4smMdcldsMG7uLE4IThYp4s43HqPpd/92OgV4LTLNx
U6PLEIykcd9kyDdTVUmMcWmKK9ykeA6rSC8Xk89JSK4bu/0h6oo1OLAXcObQGImiDIMdLeG5tERK
zzraNS2fx/rbpKJNCtbxr1BCTYndy6G+n4fSDoCMWDLXJtyJ0l6wwgIdmDCljBRd+QTZzkNB/STE
Nb+TWP5oYD72X6uWS9PWaMOvcmbLMK/+fkSgCOgdtpSMNtKg2MoF8HfXz1wSmPOSdzSxQz6LuA6X
LWzEOvYsjbKct3Os/ElU/Q+rYb47fQX9ZYjppstmDQtHZe/99tu66NU4/b8en7c/FIMhRVA+qFG5
lgI1WVHKtesVUgMMkhOLaLx4SWSJd541BpfKDd9lJj2NThQ+iNC3W6svDB/VUC5LE5gMh/gN1tVU
OeDIrmF7usMpEMY9n7ybDjU317YngHbTFe1uALWqUMI8sCE65+QVsHMufREJKqKWkri3uS1GbgVi
cmJsZLsdEIsizDaRXuq2HChbMm4iNuZN7nRsv+RJDDP893UlmJt6DjYg3y4ktt3RxkkKYexhsGNR
ceAUFN/FucuqQy75kBzgbTzjTVX/Zsbk1JL2epl/d4fuS5HM5HrUEYHZEgXHK0rtfQVCGO1viHZU
bCvD+eBvmkGEo7hMmyUV8SS5jtlqfSBfBZkORXiKmVx57OZtmuHtL5Ip7DJJA63/8apNj3T0/KIt
IsApZQbW7qrYyKZBPULQaHACQ0WSbfa2Ft2uw3lUgVUOoI764MCMQfRfXBOXzzyBfiSFb5lJODVW
ymj1uvBLAyr6ZbFhHL9/fQfsphEoAo/TbptW0noBBFMWg++U1k7GhRAA7k6vKrUhb9CwWpuagLdn
ClHJo7FsjRYmY0DA2k3Rx/qHnhy21pRgHS1FEzluVFZYB5c2MInPSdfrzF8Y4hHmm1RLytZFd+ip
PD8OT1iZq98QdXdDICiqC1D/+r+D05ofMBjmzqRiW5EMtE0Z3/SCzOOk+WErxvczN6Z0VsCGzibV
4s7fGqkrCkGljrZTR2lbOfkfUiqe3m8c+2RPFODz+RAE6vNi6dMLgHmM84oNlqImGvcCZ6r0uhGA
ctQeKG9nmT9sJw/Oxl/+0KONDFvJyC1hu8x04IuIJ9mg08kGAKJZ5tOkUyXQTmDkstb7Db0nsUub
DhZ/0jtvtjbG9dpzz7mmat0AYxw173Mz+dUBV2S8175j9qYinFK0ttimh4yM2WiBX+qwtqi19/qB
jUPQJnkNFzjZa3TU2k+loiFVdQCJOmsc4Jpk7Cb2g9se7z4MdncVdiNbheWEYpz+saGJy9yAosZU
b6zwrg7c5ywrZOAokl9H9JmBn+vDQdPhjnV2aPwfTds1aPsJwUuP49YPLlzuFFpjhF/GnM4zhl/Q
YlMznLTOXMlbu4p4MvQjpTT3j6mBd7ngWfvO53oA55jMgDEoeTeHIGr/YpcZV/0LLAl+Dl9RdyGy
TEkYp9OfN9Z6SuuyrLIXm5dwnayO6EYdMd3bp3/kVzI4XiFoi7o3D7XouEhv4kVWtHyQQHQnf+HN
k+ySur9Wldu8qQJyQvbxnw8oyewNA+X7e5557gUp1jxYCUCrCelujD/7iG/XYFRZs4vRHZvZDFmy
ntjbLfebQ0tX1N4ZAgG6nozO2h2wfqmjFDmOMnUmZBWFHTvB93r3UsqXxsmuyjwLEKH7SXBHa6Rn
N0ebkgSXtZxvZEyCD/uFd73ZQqxgvBTPYc1OHJ4Wx2SvPECkFCl2jaIirjSsCbmfCZ4ldHx7BXGf
2m8EksgmTsiUc7rxNL0FUMpHlbPN/XMuSe2F7Rm6qdg0ldrRf2waHu2hh2n3eIuoFMPhP4FbcvuH
g0yw6J/RxuRBFSKt/GnZViU1Tma/GiZNwhfFJrYW9iplAcw/V2lU6yB87ISA6erNgjYNnoO7TNBM
Oa2CPDNejSU4zAwiLznjqiySDAOF/Xs7TLYyyPEw0jK8vI7fluU24qhcxrOx1yZP6qRZboBf1Tfg
LMQV5GDAfruq0IT2FZRoA5YYACDkCx65VDEU6TODMMST5MR1u0xSCht3+kIR0xgr2vbuvqoRdq7m
BLVIi/Pt1kgaem+Sgx14Ctwkd2jeTxE3GT7LvKy34/YAMvEq7bIBSPjIczRwgcXYrHTVp/BV4i9g
aIi3tfZXNEOaKevBKM6z/l/OH8cVhrypAjnB/mny0RGwBjBhf0jVjlklzjgzOULG8bi+hTgeajfJ
S9vyA5mem9vJNn3NU14THSAXNeq28lcd57yv0t6/OfJo6xFAJiF1fFUB+C/inRueJzq9ge+wVP33
LnF6xR5tfxH3CWPaBLybgQ5bZ+tzbrrXaj7d49LTm7IwqTh1yGYCe/vU8NTg/nxbnx2ShUy7KwOG
N5DyWTNMsqlh24pJWqgZGhKunej6slFs4B74sj2Y7BzPMy6BFuME75xA04YkZOtBqHmGFcA4V5hT
bBtcU23+nrFr0kHSZa2jffMw6Y5RPyJ8vWvXJCznIqK1NJv5HPxybqpSHmDVufyyQGLBsvJUM5qA
yYh7RTw/vNY0pJtx6fXJOnuVnoLGaFQSHzsliX6Cr8wgbON8t3oMLY/rSJwz83gmHIMLZEYXw5as
/Tkz23dOm2QluCJf1GSH0/KLV+Hw/iuyzc/gDBn/StQfENFmadW5syOaBGCLONwjFxLZjGZx9Z4C
Ly+m8TnC0uPfo11w3Pri3KjDAFDKPMx/Sd/a8CgqCjDFJ3faK/vh2oJ5x8eFQ30qFxa64Kb3DEO2
ZOrWUJn1T/M9M0UyDk3HDC2NehtytgGGcqzK/yAPhjuMJpEXhqUecIqpY0NsNlbce4Zmt3WEoN9N
Mf7Tw/koHzChyiHJZpnOvCUmR7bia5keOX8XdYwRAtz0mQ/H7MmwIrKuzvIqtHpYqfU8OhgCsAui
NDxBOqAmgns7Z/dC24N9czz2OELw21piwmw4cl3qbU6ZqZN4/ublMnbpKMwdPA0OY34jCpMkC/un
jPSPiSseAyNyo/7KtReJqV+jWSkrIL3CghY0KRMvF9cCVpA8s4+1sxzExWORBpKztuWzBVoe5+Hg
QbYK6zIrOcOjt35mBJ5nau2xWGe+2EplEzLcT7byEFEHAakL3bHtvY3Q3EmcAlImLZadxeVNpC0i
h+VZW1z8wK2WDVoiI0SxnQQtmftuC7QcwP95rIgkLCNuVRNt5zB0cu9hqa8Wd/rZaO9vWYqqWSE8
Xxnetk2IBs+JdYyGziBPn3LgjE6XiiuvN6Aq+XynY2G8McEvVpOWRttsmM+A1iow2MdKiGswCWu3
WAj4jP3VFoaQxlW9MHyIlq4VVHq4mXf3XZRm6jUCEMUQaMtsMaVltjRKQVonqq5G5P4DkUaNoQm8
dx4OciA8RbV+xWwfhYM5dUpz/7XvzkHzadMEDM/vRWloRF2W2o7Z+wLiLZHX4mhXgAlYmQPH6ZQf
Vq76MhorgDxI5Lc28jV3YLaMhDEkwUqH8BfZ5rWaORfqGUxilTWtEdyWVpJjSu/tYJ4ONdlc0J+a
83KsS+aMziURx6+gVegbv3FFZpnBTMDhHb+kaA/wT3RRnKvFlwpnOab+mv0FYHTBxXQ4JxVCrgE5
UxhwCrsBRVi3aMP0dv9664eLT+xGqfulyte9ylyKFpyCxoVt+QQE71S3jVTTGR7eikimZIagLTAi
o9ICyE2VaPLQ/ksq/byERYFrL3aNESMmUktZzIYwUGfChhUNEolZCbxAKuWkMV5LZ+0b/9+Rc0OD
WtlBE0wg1uK5+p5bvKe9jIW/PsMJSwXqpKnE/fVNnO3eMP80cIFzv/PDNxyy20Jfv14KC7MICDBC
lR+uzAdMxly1220LuIkoWPLCMFNZFIybU0Ymqs15Rwmn7AZXsIvTIbhRNwYSHwDinT7CyyBKRlmS
zu4aFrKDuphbVGksIao3WwJltYf1DGIGGAzlx3m1Qe3PJbxivBAzu2xK9gzBqBEBq1HfTwYnBCmM
aSmih1oRzqWmoAkIQSqR0ZDYXs00O8zBAYGAQ0lqKFVKnAWh7D3bEuKeGtvv0r7PRTby57H1n7Sb
VHG31u+YkTxHfE0wZ7+XrX26fLqOJX9+/+ovg/WPXDwMNgcUWYoQhXBX3qzCziewRRaJWJ0icBXi
dodl0Xa5lEuqLII0WOUDcawNFTDSdraexX9jnYLicqW2k4OtwHuObekzvrJvRaVx/Ffih9MV3nCf
73zJlRQ/wxMaS8oYGZcuOsV/zjxrNVDHWNjyfZxY8z1IH06i7LOTWDtrh9Zcgb03RTxvcX/TKPx/
PGkIf/+GVebKNtOJVYsishI3Ty3uPbn43v5skQ67H8wCs6x9VUXFCWVkrfESX6ovDVFCSY0IN4OC
B+TpOxH9wlCDqYIQzLIn8sjAEqWYn3QAifbiwfr0QrWmiCNTGy5zMQcYteobyceXbLiL0QO8O+Py
Y9khr9k/kkb3BPcduM7EWGpYugEzo3LgCN+X1EAY5Z7RA9/4AHB4/ABP1Ff7qhsa4qvmvzUEEGMl
+Hgo+clSTgAJznDw+f+PqWlvamEDHSUeYw2t2E9aExNUQhOlafbWyN7+EVVCLeKbmercgSVF4aRh
0MA4jJCOIO/ZBZrUSLvvYmhxpYk6tpxAwpjmFVHfRmp44LC0h+LTWtR8+r07AIHiHsiARpyXe1Lx
s8z0zpqG8IpzFvH9RcQ/r+9ffvQBcssI6cfIxuyreHO0ocK/Os99yxuSd1e6GomOcv7LyQZuoU1i
ctdlAfEt7vsTY+dbbDRg+sjxoUBOf9RtIpRfhU+IHBhehJAoHhvhNQigXGwifahkh2j4edmB0kc5
CrI3qWEQLS69oCTHw6ni+LMrUWKpGnyBLslmxYMtb4bKLG7st5CiWDyiZRyGEOz3clN5sjGjaB9/
SLUPKcYlwdqiGxH5NTm6k8RiYcY/mEY0WccmrgYdC7XQ29U02yMFCqLGk2/p3zO9GRUJUDIbmXV9
SI5bPXSRqoEO6vE5icuyz2GQao4NBA/MkY2u6dnFguJwIXI5dLOEJj5z0pAfJuvurLmzWqV4kgv8
VxPjpq268g0dXOp9f27gQ6TrHLihd18thx8JJGlBaST34BpM6NHnFBsMtlbgua3WXvsTzmmyV7m7
OxXGBKYVc8yJ3Alb15yV+6IU2vep0FtY7t+rGkBOeFYT6034qP/znj0cQ7NTkuVqOr+BIB2zCS5P
DN4YF/p+dQu+wx7NX2Y4zGGzGhOTs3kHe3drpT/AdDlB7vcJ3+R1msbjkJkLhxqfr00T2IgSeOgS
tPt4C8uUsxfKvPXqY09f+3nEOytA8P/m4T1D4nIlc0P9YmFpDBIn4ncXy5XvouDCTlknEc3zw4ZM
t1pJf6+gAaPetaow1mYnxFFOl+JvETgOl30EFs6uPKl7CNzvvsXRP/VPoy6nBFmRfNqTzhHYgCwM
rlsMs8sjhUwYGm1zKGNPCnbiKVyhM+9B0NoCUUr6hqhzzG6YPKmoYCprWCRSM5Ecdke2Im5+KMNX
NEkYraVG0vQekcjwjAoDUsAV3fBjbp1PF6AtzoDG4uEKeymGTq3MH7K+KjPrCSpcuP2K7ldMnIq/
05hLDJgWPesH6BVSFWe/RdO/jsj+YMm5tiQQxu7QYkcqEkdu+5PCc85yykoR0LNID/7JfM9x0rhu
EhLWX9NTo0z3dG0PO53lo9f9RXiRghRJzWZIkQ2QJ0+Ti41z0As4JqW0ZmRTtSfyMhQ5v3xWQeIA
F9zG9DoO0xkesMO1DVKdNUhjU1idOxM+nKM11t086wNHnsiXsnQImT3qUzz20UqRiCx/OgtzHY/f
hr5UrhusrItF3jJIajKgS0gmxrFVaQBZKEgPhQUR6ibhsoxa+fihKlamLJuxXrJih362vdfhjDRA
xxkHXOv63QI3TUDs/PJKC9+/oy4RoMtZYigep0LUimOstXiLYbRQPNPMZwJhcu9brMLyw0zPFvRo
k/OKJyiiWqYglPaTAlJ+Xk0VzCZsqJ8Z+0jMXzyNizUGXY56K/p8/qGTvcYggg+pTDUbQ06R9vyg
vlSgCBqQ4Dhyk1obzCGl0hUByrlRwJDbMMciJAHJGMag2L32WF9DBv0UkqKvRYlYC5RGqWb5724B
bI1QbYP5PVpWJIbPgtgI9fuziweEAD7jA5/f+wZoz9uGq2Uq6glCKsRT/qH0wwRHazIfEy0RgpDJ
dQqZzXhjA4kYbjS0dceiyzY5Z5ng0utXFLbG9948+96bOJgcMyTtQQ8c6RCWeBZaY2d7ZUker6/d
DdzOLjx6RnXCxIcIXSErWlEpM6wpAomewiwfhftqc8QRXYZFoPqYNAz+4MJRDbKulhSBkuEo4wam
c4U0D44un6irrxiyW+1jnTMofawfbHAG6cZz2IHUn6QwuJ45BUG/4knE1oNXd/iGp9p3MVj0LzS9
tSqlP1BM5X2cg/NYrbg/uZsIsgIrj18MnZAv90i7DymEwn4IlKSrJQ8u67iWm2raAHBE9DYW2cXP
sRhPBhVnB5vzx9+ZOLS0qlKPZA1kxYFob/DEQAYBmVt2Mu7wgS6K/RRFq7Rv4oQd1q0CU5+Ei0Vy
CiCtpmkUXS3bh3+GYQMYtfKzQOKwCBvxyUrxXZvQusT1IwH6HQRLwrAa4pAtbn/4Qn372Uo5odLH
1eMScOBwJAUrvb08ZeSoc7VePFwoBCf5LDZxTPQ02pi7VcpdnTRV5hP6LLG9FlIHqSRnzYAxD5XU
PNqSIPRl0YCXo2jDQ6/Am2x7MuznwJf/m3vpTbOrTmn6QnTxwtSV/kbHuErCL/i7gYA67pFPVOy9
wO4cftM817wF1maiii/Ap9LuDy87bnkcjZ8Wfio3LdFLC8HjuMcK694wVdXalwMcdbfpRHodZJnB
tlw8J/q9vctQVrb2hr+zPg8FBSf9FbrElwyLoHe9npk+lt9bzu5hzztJ/0eptgL+cLV3lu1VUKqQ
uvy6mpZHQ477K5gAYiXmMf7bMAXrd5cE5Y1g/XBwW0Ly57LaWhuo1XYJbcOZrp7gnFo4XkEEIr7W
kr9QN13HbQ3FspQgGvquaqCLJONjMjGejVoqv/JYSfsdSm/wmDVM9BNg7f5AYjllVWpCW3zKY5qW
8Idcsyks9JnCn8uMna6lmGef9a11WsbfEZAASotta9X4hLQiRoRcgEHSx4wai6oBbMnr3dnC9baa
MZ7oLMisIkOrtE9n1Fza3oIHplP6hoSsFjPHm4y5FWoDntEmW4s0HuP+FPXmL4NhRfh+nQvrOaOc
ZZpsUFXWLOGCZ279tg9dU6+SzEARVHVY5ncjKm7DSWDMW+80Ef85OIE7/x5ligoSRNxcmlrof8QK
v1elwUdBC3L620MFs2dyAIOMGhgwGDOrI3HOvrl7ni07FbFgdrOr0i7+0QjACrDwv68A1t0aRfPO
ldaEDYc3cxVFhwB5QHWNEbN4th9TNwfT6O+XTLbMbdDvEdhcAG2j/etA/lzsUVpYQbnmHq6eROCd
Yb45DwbMHDmf4jrrUVVHY2L71iJbPIjVV2C4FQy/iLNqiv9IaU1d9Txoz6URvQBuHLNkgENZI839
uNlYsdK4Lhz5LwSyJsag/xYy5NlbI+VCZj0iRVl5NTqUESW+XnrYoqk0mQW384xh51ICjOEBy0pY
tjYnC6udhBNa4On65axej7YP6WxTkMPdyn/vTvVYi9sVtnts4Ztv/nKJvntGy4wGhwX3aLUj4OLW
/No2kzS25OPvIbvEt44U8T2vLlumcaj0POcuC72U7VsWpWAnCQiEa+FjrZVgCANHHeTGlu8MFezD
Kis7MXcn3Np+EFnB20q49bwn8KeZKErgtMnWxeH+dfGyWxPjaZ14Fo0ijM+t3A6s/e5lOMk8BnCH
h/9GPlOGH9LiF7i2SxWZFdabA8mbJYpv7lgRIjkX1Am+a3uFF8KAOCJpdFQyH/sgtee7fqPvZmx5
8NBmYD1r3GsgsiqGwmAjHq+ASYOIbtXo00VfpxDAQwVhwfWQMNJM+u+3sMmpEEMH4p+a6D7VcMOT
y/BGcLGSs5SN+OnJ8fF+SrydQpUzPGgn9a6uqsxmMM0yCrqMZNVznI9rxrm8LOyEihI3jS7PSZKs
Qytn8hERuAVJNcaKDuPmY8DjB8+RT19MMNUwSpRSTCwtnbl7HDsqqWs3Hj+RMuCfkw3jFgkxxB1v
zDQozbk0rHRhKovkpUPDjq3uywyoCYdgjSvdIjL80jQn1AVV5ORNaHsvC7/mSxgi5iQG4JD+6wjp
GG7hRA81+/xYOjvEn/ZXYi4IRbzCoIZWX9rVq4x95eh/EZcBSOvF+SUNdyOftm66CvDS93/HOWbO
CynG2Lm3Qar9opKF5HuasELpqG2WQcldclDUFxYHxNGqGA/pu3iTOpMEt3Bu4QC6y2vdbwElRFfy
iunytOywWUxGf5C7KGl2QdpOr5vjAfhAV5aC3s2eH0htjP2a+E7UCjJQOgP1o33/BmyzSgth6un9
Mwk8TQvgL7Z2IT7sLz3XuhQO6giuBPWb3GU9db2z+wlJT3BjNUQ/b3Z/jbKHiYF6yRdT3wQxj5Ls
jNfW+DSLBtJTTIyc1d92SnroCrHgVj/6SmtkStVumJu5vCNDGb2fcMgvg6P/YdtmJTZhs+pw9OQ+
+DjjZttp+SRxJiy/lAA03kSkex7/Tlg6q6nMezpBgAXt5SneMVfw8IgeCY6No8EbAlt6rm6BN5/+
+KFVa2Qms+iCWfBy8TbniTSgSgx7n4gO97a6pM/2Uh/NWmRTXgU3XJ99Tqig0DkQTRTyyUredWf4
4kpg0YuUEEqG8z1EAVJ2yG28pbONwaeGaHT/nFSB6MKqlxLX/Q2xgqoSYoiyvga6nQ9rcKjtZM2w
ndRRiIO4VH+Z4ZD3uaREDAu+e8CjH94cxr53BIaSuQ5HQyJyQV2tnOk+ZsEb4Ggy17pljcUrmDbk
79TpZyuX6ApmDgMN3k68jVwI1Dox4kW50iF2x6GPxLjP60ZG5b5NXUAHk60ZE4zJ59bwbl7qUlfX
H0Ydh1xP38KneaT9l323oFxyE8ao7FPJ/Dr02P4Et9crmC4j377/CCeh7R0o1dpEsghCHbIjJ27y
6IogkM5dQ/5MA6uu3tSgU1/S8NlTf+XOK3zheWBdYjl2TJt0cqrYD8jVdBAvNgL2EYKN5IfUXTux
NgyLyh5X4H6wVDdn7pW+P2TRMNN8OSKhMcEE7iapcbRvafKt8UcQ8zKilCDmsO+579NI202zp671
BnLTmi1g9szG1DimQvi+mdP5kCuK/He5z6DF+Wzb5nbce93UPUe5RoeysdaKVpzlH1jVK6dEHuBf
jHNijIhuCXJAjzK7FY2yvwOyLVyMqUN116UvcxGQi8tRIgQXw/QYsabcrO3yqKk/+mKTI8W2H0i9
vjCTnwrUT9jgTmoULWAP2SmykihG8wAO1/LxC8skeISqAtVIalWeFkQLJrBfeeDAf83YaJWrp9ph
UqDAd7QlBK4+xa77x7U97+cFl6y9CTSb4oG3Ym+ym5SpyXZZq13guH1Agzlt4MuZTOGN4H5VH2Dv
2JdFcsuK8n5n+WyKLT/usilw/Tuc+JRWuI+l5WZeWAzt0devgONn97CjL71Ykt7UPcitEKkKs/Zg
jBAaMnZw2bMeQ62gx1b4Qwt0Rabo0nxkiMlpGYzfMxedq5MGVwWMFfc5GBKQ4++1x2x8Q6mbqq6r
S+UBxB4UcJGHCetIBNvR2szu3ZSdLB+Wa+pwqKBywJKtc0uIHp6IVm5w8xDCU8ckpcJQcTpiyKAz
HAo2NpiM5OeCRqIWO7eH1pNuIJkPMXf3PpuV5ztAX80MAj3KOy4QyXzqcN1zNR7OPLr4yKO7d7Vw
k6WWjqAEvtpUF3z1uAzxF1M7nnJd4W7Ue0/avaGaKIIcSBpsbxTesr/4NEw+YffAmUbru2x9+uAk
BfMEB78JwWOGTZeme38doWmPxf69X/c1TLLbEHRkLsBCm1SsmfRi52URgIBijI+ZXX3WcE+29RQO
uPiHqLNNNYeVY/+u1IzPkWFdUCDaIeGWcovB8+9whilqHp8yfriuJO2QNznRYHff8onR1JP4smqY
qhkXTvO4SO+kp5PkjRgDFsCSiEbMPIz/0qI+j3+cNXxoy8yD9wtTrNQR0EgIN2q+Rl5cJuBnFY5c
p3HzA4xZszm6onNOsyn0SltqxgOIoZ9z/dKncSsnz8fcZYmIkdhG+tyjEC672B6cnSp6Z0Aj27YX
RgguOFmpYMDimAB4NOsKd6eY45esY4PzXYoJ3Mwxft1WtAR1QT625ci8CweV46TFV/KnF40p/1fB
OIBH+qIJV3nZbf63e8sCMd1R8JFnTFPau8GnQwOX3nFoX2+b0kgQidD5ODDNRhCIdlFcvccgKe6J
o7y4Rbp+L5yEtb/HMY3dK4KTPKbvp3+AehqAbKax1440JvvWHw4AKdFqV8kNMNU8H32YGDxruUy5
wIVESI3eqro/+7qXHEscFC3E9ouB70ZhFvDG79CpLd+g3iqagDSRbw3mZ29SetuPn522DE23/SJV
/7fzgRHkRVxx31ZjlPyK2fdISe2j//LcFjN7cWgfLl+NEsIK8ADP7ArIdzSAD+Csuom4OcltwS8E
sYb245DtbnicbWFdDyJ+egmLQGEc+vJWjfimEjn3bYapRKV13y6IZdyJxw6myHHyfb//UHrk0Xox
s1t81wEDnInIXMHviEy+/YvLIhdjgQNhLz3ZNdFPcvK4nUqvIhFU4A0W1aHC1KkA+K0CRsgVzZLt
9SMmkvoes5Tk5lKuDHycF2qj1Wlx3vEHt2QXLyOBnmyDjbyc6rv+ShtKQhewWb1OAwDeN9YK2eIQ
1M/pZVMWZg9xsTpzpLS615p/2FQEO+pSBXXFjG11T8dKbpMiqpL15fJ1MywEdJMBT4N7y7glnQpH
W2wo5oaicqbO1Hr53cSpFOKRqQSFxkhd522+hStnyJ7+wxp7y72drolWBHh1Lo2QmpOlf8LKXTdI
yn8quYILRzdZSud7kN2QYzNu24/0qmoL9PkqKyOZHrxzB+d2K0bZXSpho6LVqfa/kyOFm4cpU0Xb
wUdnoJvO46lraVtnhokGHn3kJDQ96p/X1N0OwmaWdjLHk6oWbz1UrNmWqtI/h1aXGqoYUof5rTAX
fNmB5053auECkWRjf60lA5qsSv+pO8U+Yc9VuhEWli1LNsS+k6/hCKuSX23WphUGWUHpOcWB9f5S
VokL9G0Kx9ovJqTtBBGdeBHADz5N7b04+3k404kuropM+S7KhTEk97L5neGpqhHayj5x3jjjhD+c
TEeG+Lmi3bkQXedwOZWi49Z/T8i5BufFCP/VL5YVYIhPWG1p6Ju/3H5GCOtw/5Rs0ZfS3GBXUEPU
unhpkgIm52YGdAxaHMxHfo7LG4GxOtM3M19oWRPS13XjtNM08sduNruiehR2dOl33n0N9NN7cCCF
Mubuj8DTB4EU3AeH2PWzQRhWqIS5vZYuuwuGInxNP2Ts4TujdIBENB/PomtgooAMCOwIFEosMZGV
flkHtNgkKokuDSECFaXzcLTZeqtW0AqQt3A+r1yQ+xp3v7qyRU2Zh3U4SEZIH1d+w0lzj2RSwVJh
u+YlZTFIN9YjlReNLTma68LH6zODr8OQ1m9KslBW3dFftzd9y++uL971Vgj4PkLvZ3FCQN1AGohF
KRa/ZbxmJAxQx4gXeDhAkKqBlFky0iUrkEe55lh2SLG6wOP/3u2sfEOsgbnIGQ/lT5ZUYifeW+Ui
MPAZSks2wgtprhgkinhKNLXDaR7VW7ZMvuAumffSyspRoCO66o/R9hsLtpHdL/ZEv/f4zkeT2vAw
eVed5cgOwRAWma3jgMsgzMIGlxZYoCShRTgDUnvHSQaozsbrUjHRDM7Uiv0lbh3bmiK5Q4sB2L8f
rgWUA8ajBmY9K02mBdcJgTGnFDxdJSQ16vTNSeE4xPrqk3zjSi36L7UlOGkCJtX+eY4ktOB2CXv6
Y0r/Du/dqkmiNld16AFjCJvq3NMo5KPImGdqr3qxnbzfDjDAjDzkFmqHkVSLKUxvXUG81OzS0fYw
O68I7VJWOOKljY5PzDq4nBgkqsL731g7zXwlDDa9tjWMX72L3cSZWW3A3o7o4mfJxB++dATztGHD
X5mALaPP3KBkkXf1KgssD76sa9QOo7BU791OTeFKWjcAK5VqCZ6kETQUuwhn+Eg2aON5HXAy33tK
1H9vzcl1A1kOUlafopj0AFv9Dsx8aSyGNu3FvGFtEF0y5VF30EymJ6p6fbEBQ3qfxFkPgFvGO1dx
Utvoh063/WhzluJ69SWv3jJI95z62VEqCRu854RWVjle/aYG8PTVNznQ+zCS13Bn9J2aOsATju7j
adjqzPXJhUtHw5R6nHWPjPH2x+FlPsoxcihmoqMux93m2T2uw+k1BQNr/zJyPudvt82j9GlwFVys
Fl+7jLCn8DYKrZTVVCS0wnFbjnUIATAyP8/xI61DTjCkzBy6SXMXlpww0RfXlSEQ9oGAHDAKmd1o
duIGWPbZGSjRnidr2b/VEX2QFORBoe1wNqCnGoWdWIyclang6yHBTWs9O2TYXYoc8PF7yeAZaE4Z
k1POZi0vVC54KyCqxo39XLcIYnyzxXcHViBbJ42ycRJP7lertShIL+PTsJIzhinCQU1l6IlMySSt
GNWe6Rvm21n5t+4gRHqf0Zz67pb8XUd3PGqJ0t2OhgL4AW/aE3e7zW7UHW8HQ6u9VfOc/yBUpq1n
BouqZW/N8Ji7F1KD8+flS0L2uk1/JuxnoyarDnb8PnPWmZkYF0zpPScg+ok1XP1PV0rFJdokfJ2m
VvZ/oYmGxxtqa4SR78CwMdnMm9IZgZkH8Lb7eupNFyWLN1qyfnzQDfsSJekyBL9AiTEKGWqjyJJP
5Zw0jt41QQ1yBBgbGPIDJEcPR3ZC+C6oltgvL73bxi32LpXASZQa1i0HEl1O0C8J4FiPoAK3PYsI
pRXi9kP3nCETBVlqAAW6TjKO/idFCVkkoHrNf6Z9wmQrPiA02N1Sy3I0biLItJsi5XeitaO1BEQL
kBduoV92PfALEm5tAOxWMGLdNV1KuVx/naGoWp+YaEoYhMDeqlitnbUueS89eVEQZsxNA2ll1sJC
FKGv9Ao4RgZW19wvN9jMuUTD9p9D0u7uIEs+Rv1Dao6ORNdZcqzN7uQBqKYzFRpGjy5LxJhRwedE
VVz3/YrKLYzXuWMEMB779QfAAtaqMjxlIRmwdFr4Zb1QERhkUDQ3+SuGYf1JrBbV31LiuYych15Z
pG0GZD3Q1JW+XRIBtVB9fjY4cbfj7kDZLlVGIUcW6tqAh/N0iFVP04CG1O4cPLkkvfg5ElMk3zmr
bpHaPzKC4adR/4sdJFKrq9BzOi50dlxqDDdxb10fWxSJEIbm3x7wW06s34473vSC933N1mG3GBpw
vHT69JzC7RWiVIWpD5O8mngibUMZ8Ecy+0KIFU0td/mBvQQBYoMRzWMrHDKoDytKgJJ6lWgM66OQ
F716i0yW303xFYTE7xojBCtpxJMHTUd2DzRM/CEzGcW5iJ7knyYVzUy/o63jEW0jn3/OhUjxC/9L
V+wY3HIIgqeuyiDRyJv6DVc6TrRFgYzFmZaqcudeXDYEybWtHz2+C4+L5j4/U9aC2D5ZSZSrUIqU
k4emt8NOkjhKYSaOzEB0zX48aZawgjYQUfDtVtV6Tr22IrfVAwI6sp1V2UZyvZKJw2YQsHMemRuk
QKC6zjbRp/LGi+u0np2lvflXQAQ+JMtzZ5BGBDzoBB7h+HxHXNcpSIflZ6U/CoMBxZwOa9NJg1Qi
xmbluUi/+HMdTrXObYypWjdZga2DP2KbCtvFrDc9B8Gi3VDZmM0wqbmXfi4oyo1eXbbzxywg5BVQ
A4+fb7k0CruGYZIx+NuYCl58NKx7kg04J9sHCRATTj0MlpKlcU8ZgMln6q1jqhsNlTSvYIeFcdlM
muhGzSEOdRiB56K4HV+C1RIAIAruMBZBtFF04E3u6kOBUb4lZ2lDZS8v8JV77Gb7exW7vDN3ZI4g
1IH/GdaCAYV3atr2SBJ7O2wNlmHZ/aq3JKyyTibeev1lLEgCXAoPX43EUM7yImzDEX/AfLTAKbOR
JLKjZqb/iEhEzJRcPHhSgmPcnmoUwOuHh6Rk4VHJNAbfquhY2BzaweNtBd6VC/qEY4OFFPbUpQG/
jVLPkEb6vFoxoK5K2AmxyBnX0+7Mf6u1Sl3olxcg5uS9iWPG3XYPYm+i9LuNAQMp7Ioze3gH2x12
KsDvcC/r3QtcRDvCe2iQoDlszUAzvulbxVJvJCyMQiWKERscKtF0tT5E8n5MjD2ccSci6Ck5P2+0
bI61UuMFTR6DLEjGAY5G19nhoVUXvm+1gbtC9GNYvySk+9OZljCeAZvkZ3TkSwYieypmYcOQ6KUa
7xyV08f9tVZMaQpcJ6PCQYquARCTc7x8T+YXlIvyGZdpTlilAnKb/MeJMHGJTp7ft9sBTDITLrzF
JekLImHZ00XIFmJ5Z87W2ryAlJj+86wnA9XbO818XOaZaAazkGowb/QyPDnT/KGvG3eg4V9LsEa0
Jq7m03YB5u2dorjm4OAcahayweDLgyQDN9UhAItMCQAD9vwhmrqb4ncnaFlCYnhVzwMvBAEgo01A
f7JJ3B/agngtNTLvGPuGgwaEQL5bAfuEwDhc5D9/k6mkNPcmeL8hLNneTQEFPG+Dia4IUOKeViC+
yMJRQI6JTJR2RYuEIhfZdi98pOdM742fqvH96uMJrsXGq+JrTKlKuwKP4NvwQIkiNJZynEbfKbFM
FGfZGrlYyAoCTmPF3SR+04sZKAQMqtRyylrN90+cdyPal45XrqVM+YdzX5Qs5GfEjnjWOeB1Zh03
dBF4K7jW28l8H0XduvsQ0BwY9n8JL/8q2oT5kZGu1xTPUYZhaKSUKb6peWBtFk+9M7+3BNgkNvKJ
pW6CrtTJLYkK5j2D4cWYVyXmXFsP4sDGyZjSdsC49nzXEVzZYIvAKiENKWwUzKO6UJOc9LbirgY6
zlJgwJKgxYBd/XzX/jTspb0oXzjcVkShQmyIQaBrHPY/80fhfl6lswcOEb79HB8ygDXmEr5LR7Ci
3wDapHD27CVeIVhDaJQANax1Rfeyg7T5tDq/alPFIiI9uyspllK7Nuz9Q4HTFgf2nKajF6laXZEQ
zA5MS3qbETKjglwN/FwToadEuoAJo2ScqxI9kgqTTUzHuu5+WTOtx5Mwt0hYSmZzikAwgqxEX8oy
GWBVBqmJ0iSSKSimm9BxtR60YDLNCa9exh3YveMxErfe64k6m0snd9M3Wsal4wfHy443bkJRiBMV
ib1RwUvO6NlOMrzOFGUzcPyKzkDZWrQi8+7sIwwKZxVRjMf6quEzRPxM0ja6EZ1k1AkieOS2xiaw
ai+xH22Yklox0IjcKg4mTM0UrVG546gHbKcYz4cbidyBkWAEALPjoAfjWfkPMEsFzv2YrOd18L1/
NtqJ0FQZHwKVBg/zmZygV8xIVtFRxPaRn4Zb1cLhI8xU580XFHKbnD2vSXHugxyBTQgY24Bv46if
Os5u5QdXkNiVSzicssh2wEcQuEv7nLic2p4/CZL1Nvs/dDHl7AsrUF3SJPmlx1xRomF3USNjQ3NH
SQ92/YaeImZrCAkSQiJ5RX7ZQ7p6Lx7L1SjJYtj3d/hzwivdOpjzpbM8K1pr8HP+OVgpsS6vj7my
1P4VonceHlv9Exyx2+xvVrmlPwJURKDkuusw6cxCyOfn8/KXXdJIIlktSbDtAeFK8hfFQ64KXnox
f96Xd+kXfOd1hWnzK1HGXubulCX8EqkHuGM4vrZpGzk5C5qpDFDLtHzoP2BmVv/2Y4G3J2MjXH84
xYKdn6jjJqhRYUsUtW4G40cKOmoH7x7OEJaiiGe9ZXlHcQD/Yq6uL9zuklya/5mZs+1Zk0oHPoNk
pzlL/9iCuJc0Gi3JiswHDWTyIZ1v0KMXwAUdJ2gr56LK46xqqxZV3keBEcDyQhDNRQ4BN4ktvwQj
ddAVrpZAyGw272GvBPyVXLW9ZCY3ZnaY9r3eS6BLXkBva1yPGc7yjl0/QBt0CyDL8mmnu50p6EZj
7WCEED++3utGnv8lpG79KzpfyGqdJ2XqrdTfP5YmtnPg8np7MPlgowYkajlY29LOC/1KjlRB7vqT
Sv9LBSQttEqPueA+viYP8sllX0pFsRfAPTQttSq/99+C7C7RgRmnP2qcOCKO8VWNxDxlPtsIBaEh
jzTBGqmCJVvusLpjluDYVPbZNb1v1x1dWjpAhGGaFO3D3b+XaLklwqeJz0o+8i2OrAnXiACFZ5aF
2U7+sx/IQbEct7D2h/K3azpCLp30HDbxP+fLO14g1wMbctNERwsCqKLBFbo5+0Eebmtgp7ZdAnVY
v4+6PKt/rwRZMmsCjU3CuWtSL9zFCVHIKQiij06+ZgrTvTJtucV/dTyT7I9j/0ETE9oxx12bUPYT
7KQG4/lrUe3cB1D1w8XGWAsI6CFfqeUWmDFzVmDr8Bu72F71CUPYjfTxK99PFv3HiLedAX+WOvEL
vgU93e9RlIpjIH/TcOfNMqWbjjzkwjqF8HTqWrX3LdhHv8uONcFcQlWhWal4Uc0eyAhwy3KgWdXq
lCX6Q7uKVzFsnhgDpGq7wEWpna0yX7yqWVnZHo1ZMwujjafrz4bh2SGypEGS7z7COsk9DPe6ihcc
otcuzzQjj3g/zredfbV/4wJjcyh1alGDNe4Pa96ykycWcrnM93oPcO51VLVwc5uDxQfFPsIoK09b
QoF+yHi9ORwveaEyS4I38ZDZSlLT/LWgjsvapOyexX2QkBhh/doM61rVFersh/cfrPvI6vx0gWyw
Bpt1QD7JwLqsIOC7NZ6fJh/P8yzxgGh7pXBPb/agsRVX6DO2WiXCTaiItDAGa4XoWwy3NBDDI22C
gEKZ8eqTAvXmX3rdI2DRrT7rrffyzTFNNxl5l+Q8JD5aAfs6Ww/aIgKU7IlYxV24yA66MyO72BrP
S6nYZxACf4VQND10x5rQ1WJosXrBD7H8NQvA7X6fAO9VSVvxTKIyfStIgLjNGVjE6+z3sPHov8vj
BVPbccIwX4UexSPDTLKzWWGrHdtGdJQNy+mC9rUFa3EJqXQcrU8/W0AV8cIZ3E+cU0cjHnR0WP6+
Azo3wyixMNW0l/ryDR1EdaedEAZ1eEUWFeyeXvT33d4pakwHWH/FUYHFVsRq5B0JcXYEZWxW4p4W
cmXcoVm5SY36MicWDMZqjJogze6AG9zw4JcPI8WW+ZJXJDKAKnVaRucrnsp5ZpqMCS84+GPxnkP9
XYQLb2/pkBw4iV0KcVpCxO3ES0BAaWcRph0SfBAnaMZuDfbXmXemPugvJ+VLVhmF/ciMsvCPlzHA
Nz5btIdmCXPFRqXj1t98or/ldl1xOYo7+I3CGM9uMfTZCkHrq1gsewyBy+Ykaj2p1LPmbnjR6TgY
Kv2WASJF76QKVgV1ZDn1cL0Ny6NlQ7KY6dWgmuIoqruqs5g5bik/Q1LEz7bveJhPMD7/drd0PMql
Zim/3WqIbUSvJytjkq+dYkSzYoNMlEXhevkSXZ6JkJC8WaqJO+YJTdd4qTpet38UATQIdvF/W+4o
yp3aPuH89HF8vnr2+i8iqiN9uILK3nG9OW4rB9qHn4pBRyLrafY0XnFfJPf7xYMJc7SeQEnrhKoP
fsfPZCV/uNhrqSurx/P67mvlM+ygT6nIU0Do9kHz/EgbzddPBQCuGYcBTdIQFCBdkZZKsuximi5I
x6EKe/wF4JLf/RGKowljKtZgpAgBRyU4sV0VRkMdG1Audfj1Cj2c0wnauKRV49QlsZOKdgMUqAhw
y+2jRLbK2aof3Frla5kBUWnTGAB5SrC87+OPmz1YB2s5o3vFIk0vCsDGvPEP6AUYLimGZCMY85kn
mrPbKyUoiLaCdmlh1UiO5xHftfTNmc//kqvqq3X+pWH+maVCSysJMn/Oa77c5ZTfliOZ+R5+fEk4
4fT0AI2e7yMglrpIj5qzL+3AWE6jQ4ha556OnP1gcDZeoEr1uyAhfnsgxXfRld7D4VXk8wPpLZ+F
WElibmknCmIeGUWxK+S9cdgeToDQGdnjFoFi75xs78xN108z8eRvh/ZMQfy7a9UGjJnZIyrHFoJa
jutDvjWXTugT5PTp4Y/EZSYnmyt43enRJwUkjfQZW8aLf4Y/SmJu6BvT0+Wx9AIzPbCc206j0f9c
T/eJJRK2bQGZ3v6Om+GeWvVtyqlPumEGxuwe/x4CZhPV4+kD2ZewbHbDR732uDQpxSTLvDHnyHiA
qUteWUWzcZEOGgD8UqQUGtJr1NOlWbjzDqOKCzYwuRFCUHQb4N2rA35znZCylbAXuGLupt4657fA
bKTn4Mmgmr9UIaA4z0/BDt6pk1hjqKEcmkuxRKboRmQQjML+WId7dgYEtwdwEE7AZOoa5n/l3Thk
uRWoHvtKJ0GZibXxtPcT/gH3G3SEpGtJQAS8yRiuajCPK+XXMWBN2Ie0FU0vIO0kxsegHZLEtGeh
fqelr+lZ+/CgOkctE0QKTMfCTEUycTXRP9amdPFB1QxqVUXxpOIFKJxSFaI500u7fVqv88cNrugy
1Yey5t/IyRcakYKpMaPo3uQx3yU32syFwn6UMZtLjaiz7nJ/X/TtP6dKZDYRfQs1uE5TdQY5VId1
dMC/16KcoatpES8BVfsZZqZffKZew9l3pwZH0gv7YzWkmKEQ6TuO+pW5CQX6EM2/bJOdtcTip7Yg
BCXxo7g9qTLQ+Svra1siUsrQ18kAGU7UbCbDRXOaqSbSspe0DKlqi7SvXGh/2jzq9RvY1kr4STo2
YGbZbgR6/7pV9c/IjnqNNkqnjhsgCLE8p0CRaLxkWWv8HbbwIZ26cXuO1v8DdTwIHDwo8qFrdNBt
PiQj7tVMLwFCHPnHKlri3OTWqKYWIRj4xgDvOa6K9olkrERb+Atk42eZOhtgX7LrmYUIIskfBdmO
UAFyimyUbntt2SADkAMcZZaxUs4I9rbT94YgrPK7YcBDz6MniYZ3640H19s1IxSMijBWkDoAjEbm
eapN0gICbIFB3ZOKN/lX5xtMAGZmU2zjNmT2puIJ6PLGz0fx4dMXqgs4i2h9Hl5XV9w1FS31y/0A
W6bQNZYxz2ytlcG2se9dMm/M3EzbXSfP7aJ0JdOvvWonsDTM6DlMQN9GkCRNJ5WguYXdzNYRDFVs
/VWSvZUvQbaLPg6zJM5WMzViQrxAKsMhbt8srfmBLfVqM457Qh404UMq18GfCp5QVU0D1RVtS4+j
NYBVH66Ze8Sc44puirwqw/VKGgBGoAUYNGUSpc2ay83nM83gbAbylMYTIIqoxaVnJoexmwn7PB2v
E8nmbEzgFZGeq9MlBCsU5CPLd211HHAgiE15jirBM+arptDTCqswjER+KniU7nPsJa9oiHAMXxzN
V8axWnvxS0ZWcg7T8udLf6lo6YM4vZwY6CU9HaS00PMlArvcKOCciGkuhJTqZ72lY3lsKBQNE5w2
nICEa+IOF9w+JH+tvoJzxCCbNlO9td6cG8I77/svSnHrtTyyNakG4T90mwAnZ37zIfwf5vKDDCY1
qwTdmo59mxrdGU7HOTojXF1E7yqyWVWhJ2DUZtzqSvDVJoB/imlVUOxU8PwMQdXKeo3cMrYylaMs
UqT2DYn1urFXSuupoyj6kaIGpsiHqPhzcPIntlEzaxtqPq2GEVbfh9TIXFIjk5/MbNvQaW/sZ0ZG
piRPh3GS48J8Hi6wW6/03UIUzM/JVzSMPoga4YCzH4K6haI68Yo6qUTAAgCNTF5hz6f6asyno3XT
kzrTz2njOnu/hnkNo4yczSNU8t9+6bD1QnIFuIRPtSKJ9rQgvr8wdDWsjuAFcDP/hWtNoEC2+M4W
IxUnZRSKQ79RD3aswTSeknY1ddlEAbKQHbmtCJzr5zGa7pt9OLL6dkR379swb+fdyMUuVGee0wIe
2ZnNqFTnpQ7a0O9Q2ApUmbJJiShpoGZmRGUjaVqVnsLBAG6MSYXZ/IOgm4B8iGh5m9aJCQ5x++ZL
q7xQcmxWnXMTVEO5Z4MHFcIcH/bd55gC0VBXFL6+Ls16Ib9sIBD4V3qFN6MWtah1m3dRdI94xmF3
KuBBaxtt07D/G3SbFNR307EFe/TdF4quZej/rXwbkQVNGteCtp6mvW51qy1tqMpQCBTrmMAXbH5A
aD9/lLENnIbA4Zj1OypYZpOoditHi7GvLAbbI6yVKrsA39W+kMas1ciuHbprZWEv149f7L09/FsD
PTbXFsPoSPqsEGBaY+RLBWC3l7LTFADMJ0DawaH2DWRnPk5BCrxGeBIL83Myiqm+KYdN8YmOeo4Y
d96pUv88WLnLRyrH67AEuqisLoZEf5flASZ26DlQ87Plew8/dhXoKhVrH7fxptgcMdPeQktox8Nr
hINvz2lvh4M0RRsDDY8q7nxEJ57T4gIpnQUEuhgV7JMoAWGa3NQKU/D5hpgH2jrH8npcMr9DY5/E
MNQKLhLsXbcAgzrWKqLEoBBJZidtJp8GcyaAx+CB/z6z5NDhWrfBVCdS9ELVd2wut1dyroHg8SN/
v298QOjdikvITCv356UWLsitB/iFjGJV4NCEFGiskOViHqcMTMoX6cXBI9ljbpw5uZwd5g7H1EdI
73527LEjpIosJDaZ86DJgu4CLZjclbX8usk/oRsMHT6bXEy+f9mRSopL27LncAeX1ZQGQB3YMCNs
fGJh7mXw7R+wj5+5CAF1WPi6wMisaEPKrQUhjWfG83blWpX5yYv0ZcdwsVgauoeSS8nm3kXt2vDb
waDuUkFViQrZeQl9dj1RJyxISR0iL3Kt1E8hqwDQxVBpI6aNDN8dQuBaxZ8j6MGijkFLmUb9l4Km
8PXVwB8u6E/T1QXBJpmcLa9WFacw6naWecPwSTA79bMrcpUc14nTxv6BOFq1ZUVFpKRr9kWgmn44
z7jyvOhyp1TxUJp/MYPW2uPnVDnFOnU7biBo4BI8narTtRMO55xfmRrpl6hzTrinVxeAA+Yb3kI7
BKBGPyw6/3/McC7joIqvioDe80Igi8+PMkQ9b2CzdCvx09+ABNIRUgM79XLAtZaTpHZ3Tj5fjz2x
iZd+BXx9Iw4IB/ZrQLfAw9vgcBk0cCIdCoFWc8E/8Un5cEIddNe4uIzFg8OsJ4qyOwN1/Sf2LtMx
JVZxOpztwFsTIZaA3B1HcCAUiYb4lqdjPJht2prJHALc+P1DVBn0RWCQmuDYES2iFD0Ikhicl8Ri
v+FyMrwsYWXAgI1QJKY6GbEzUavjpI/H+AhQlvY6LYVS0veOjtreWx5oLFzLRT/7566DDmPyS8CB
lvWQq2FYhFeHAJ5tPRGZQi3OOIegd9MHiVH+OJH90BvXJUckODoFoqRs2ZqAWvV8BPy2UCUa37iH
2yUC8h/EOqtyTPFT5wq1IUoJq++WuEfa8w34N1cN+8Rb6nP+eGFZp5PnWY7MiEv3bnLMS8RkwMuL
QXJhYXP4qSW+qQPM8SMkkYyWsjkMVmU7b23KrZ1UyxlOQGVcO4m3kPAm9rNpgf16OJnU/RVTYyaH
5PF4TtnXP+MrbRhY10qJvSAE4EFr79R2UE/VeWzIPNzwxnp/JTUnbDGPrFZVWdnAX49vB1FxFkf0
IVks13mEP4HhwB34+rkcV/EGCQm3drrydLvzN3voLx9RPtHcKX2P2JIsyziqk9j56p36cMxiV27j
eu8Nw+dizM8blKwOogVIgty+F+acCs9o8l30XAnqpQkGPHtO6Vn/R9e1BmJor4ONBX0FrRku5XVX
qo+7f0DeHrz295PcZHzH2ScnS7ax0RBHOW+dZW1KeEaX4/K7V0wq6RyWdF5mChrthXgRnWll+PdC
X619uhTpTdwe0JYC/pqT6ipTj7gMT14tJH1qaqjbA2Nk4bxACsv5mDgInhNrgEjR/hVhtIFyRH1h
jKDGX9/39pz8tozfU2l6tTkw4yrZ7BUHulnpiGIEe62N6cTyZIhrY0ULhqCcuol/jqn9pjejC/tB
zAXChCZacXzK8RR6Pp6snJoovrfbs3F2w35tF1UtYRusOX6gXSVQLJMeLsbsUSDs8t0e3cyXM9/Z
Wa2nNFsw41NYnYdk0pfKeYCb1fzLwUuBkS93FuYUtzqKLN3ppYFFyLU3jhYNr3cmPXr1sIur9Odi
ltD6HbFDYD2KYzdJSxUffQVOEau+5HcixccAw7mZ7FTJPA5pnawTYZPA2f+XZxevLrKrpEtE2HI7
y8wYqA9SSupa5cipG6GDCv8W9ac04qw3As3xFkTTm0srM45WSwDZ66RfZlPjweuDfNaY/B0vwzTW
mdGrdxWX7Pbz8bPzCXFrW4QBZ1HC/J7c8CRIoCkmGD7oV+unJeHHqcFmFsWK8oXyC6d+7BS25OnD
RH3jonNuc55rMCYcPRTSPauE9ptEVKHVsA0TrheKNQQ5PJ8YQkk42wEsc+Yh71WBI0UBttWiJC4T
gwrKVvHNdnqkqib+t8etA3rIEKrTzcAoW0O7K/1K+KSHYzSJWiLhfl7jwXrGvgl/onimZWZVSllP
1pf3eSTdVKewdR9xzczuOcLhsxYG03XhO3T/cgQKzfcTyyGFxoiB07i0BAiaP0WQHxEFmql14K2U
aOB8zTDLmivYMZX+9IC+7HGlxgpT/+gzF2u+pvXnlwX+Z93CjUOiccQg/ydrppQ7zCxhofqxEjAK
w7t+Tyj1ZUF27NepWWWuGLv4UlFDqi1BPGJ7jA7yGjKnXT+yeEZbKXpfJz3eOfTnp63hQT27qvMV
Ue76qH88EFWPQArVHOakk/58jYoTI3n5mLEUl6rSTyOQQgUMrIClLMJuWcultyGKKMUjuuXtgf1A
PwKS22CwVjeCUmKSPOQusakEKbJkqzNlqhiPGeJg9+o/2skx2qkwa0ZTtokbbe4ZLxmjbf2CxRyN
WyveIS7h7nTxUFEdmeKgLX24vSGUEZASwVfu/wLUl8jLFvuULD2SPckTys1SPEMOs/Qiz39ae2qp
tE+l0/ihNYgD3gG7SrwCORQWAgNPsWEduQzZblNLmB8luRsexUmgWlPUx0B+Ic9YC+T2vN965bHu
r4qXJ8099LCOiLT4ZGvaaVDVp92IZDl6YTheIBsrshkXmrt1Xh7ib2HQrzvz6d3ThzhFLFjy+0QN
5DfPVIznMrqtjCYyWqfXyMIhQ9W69vPTHzPaIH9NhRRbvbD+sL4uThV67PRoWxJZobscUlRzFVP+
XZJ5xOBZ357/MYBk6fCFcUayhQ6uWH/q9V/X7xMFL4M5+hGVpWZuVDobJ1RPBNtWZAsY6QeOIX3m
5oOcr4ktLlq4/S4lQt5QFG1witT3p6m/bdKxUJ7XLCBud32QbCFGi1JZT9L5BxMZuHEd6ovuVeZ+
7RMX42GWZ6YcZHnNRCRhM3FdtOa+kFdc/Ca4R+8wEUUX0wOcBVyrcuLjb04GAoo7Scg6zEP+8d7d
Be63A4uYA+GiA6zZ70RgQ+8o4ADdRFdTkhv+VIylZHrjFapZopLhSnvI9vVEriJ4VQ6E5BDKRV7V
Kp1VSHK4TGOo3kDIiMS+56DWyE8ZRJ7opu+4wZ4ZVjBnjQu/mcQ1DjhiwgPMRp4Fp//NTPUyKxnc
B9nBdK/QJOAw1ajYv9TJP1nBN5m21zp2XhhULqHnxJw2bLxyrlD0mfrJS22X9uiXjUDU3xM0DUt/
GcN8/0YhhWZSGbW2R904aLJ/fL1d+RajOZ2k+MsjSQUvcKvgJ7dkiL8itJWISpr7GR4c2GYsO5c9
cl9YX2uII3bBkV6cGuubOljHzuLzPLBjbZ4dqC6ernDBhjcgUER1fg4EmSAsx/oXB4jwkqDiVbA8
hd2rkbbezNbGwSx6ZdVcYV+DHXmp73toi1JZ2g+SBRHGQ4zuJdUWOcVxW04cXwk6iiMtr1zxlRFu
yFJQM1YEDqb7csSvu9FzY56ijRIB8jXkzNqUiR9ZS8fufRrOi56CEj/2n2RJA+AwZwEmYUXNWMqc
C+u6J/aAflk4k/7RRrlg9CMHW2EIFWge7CQhI8BgTVSxP6f5L6ppi9qbLEDZQrrdpeJbpFAfti4u
mJxVKI3fUQcF7cUbqH9b7Q/KdOeMjCzpjNMHKXkh6xhGcTO03WeSORy0JVqWTDjoMctTzSZWo7hJ
i6Rk/QxuFYRa615GNetrIh6DrOamjzqrhN2S/5G/3xZ8quB6cZP11wph38hg1pd/Wkx2iLoDf7iM
ftXvug7na0YbokP3O0yWMKYTCX27O0Oc6owYXOGCz03HExQG6SG0rz/Cz+OYfg7qTtvLzYwg9MtK
jeGdhKzmOIwP7jc4pD0N7OjkmWT9b+fJQheUj7/Mjw0kb/clStwJPI2ojJD4N2Ua1XROuJOvyF+1
+uBhIw2N4kYmaYHXxb+I6+qV66XAdBdlBfJSb72G4oMK8AvLqEPwnKgcNidv/3RTIQG7asTuywjS
T1adbI94uhrpCX4h5qsAeQL5oJ6T8HnLYnaTvtIYft0d9RBZYiXMPiv6n3P8mp6/CeaV9f/3Q3HQ
ovc+QJhstHQANPlCSWI8Hc6JFzXndhAbtBQ0iTCOxSnarW3l5XBZXQ5qkMtyl6eh9Vx+FLC2aKeC
DujV+xbPiPsQSzBVXhDjl+JdCWtqHBQwhi/jWsRIWa1zwLvMCHFM+k2AM3ym0uG6IjfCF9F4juhG
1ZcRGI/+25g8sS7kDuZnatXHC6gtHPsOJ8D//vOjkE4FPGLkfqorShYOY8xIDMnmAFniONFzqPcB
cakZmm/b+3irNGu4DEj5oyD+nQdotnMlmmYwwlOwSU/atbgWoH2D1sqTReNMXzb1bC96qQ8zzfKu
q/KGTkQJS+yF+/5/K4FihHkd8Ex/xBN3n6Tzzk8QTwnU896Iphhygx1YipHNmy2Zest53LLU5zrF
zYDWvY32yf2nB1ReO1CAA+dBtKdYBBPx1y7I1cFwfHvirsY18gsmMkFU6sa+dsgdq8HQqJaat+bs
aXfyx6g22vuQ1EXgncr7nAWc7rjsFNGhZ5bY7hyLDYqoZ4JjzZ+qEFgCVessIBbbfDzx6858DIHM
gLTAHdXqvzep2xR/Bm1ckaL/Y8qaLFa8VWu6+B1q1yoNNAOBLcAErx1BAXTaPFc02qSYMG0p/rZt
KqpbJdWQEm3nusy+DSIz/zDC17aEEyPn0YmJ1qyqFlZJ0gUydsgwGzLLM6g47z/il+V5UwDuCgJK
EiC0HTWR9XrfQ/L4hXnWZJ6t6fP3qQzBT9A8tb5Oco53Z3rkb7wSApWb6wNgjRyYEcz2FSNvEzBB
Eb4STlIzblCItLMTDiCdLeHl0XhaFF5HQfAxWfCARCgqlNU4N/YwG1pC0RH2DcpRisCA8ub3opAT
AF0hgivitUUcdq0NqDBixTe1KEKjh5oTjxle0K10pDCKZ63u7dFhfRUfR+z1wdyr1Yx86uu73OOJ
Aa60zmO7L0AoAXmHaExsRsq0cWLYQEOOeAbZTUi6Wol/AeuqredBk9bJhzWVuJWn8hSBZFKyrg17
Y75YNgp5+pweKfZPpxYjyLNex8mhhAY+rwBe+tfusoBJeNBTqDbp8ys23ocoiSfpltVqCvrgwGqv
+0ztnXqF+1rpZSVn0B8r0qUfRPYyvfpMYGXN3Vm7QlDN/V7REKSwwhaAS6D+WQsxyT/6Vyv7Z4ru
eoPu29aw1MD6cBNXnXCCQmmty9e9z/F0YEQ8KPfgFKBa3YqnO7cnPNd/DoAAanu42548FwpyU5do
HM7psVXdZ1jbpP4o4bpCjyrLYK15dnhqiH3KqvN19IUxdxu6OKtKe6STSG5DsOUBh8OK/3SjeCDT
WjeQlcqrB1IqiFMZkvlnWMYA1oBnrdveGqgkAcevIkgxX9MPItzlkEbsT4M3F3Qwr9d/JTA3gDxV
JDRXg/eift+wz+KUfn6NTNQfM4CeP3iqTDsfKBo/1OamsLtlEItkxcT2PBPMJerVAnVJ38mWylCe
+9Wuuw2qjDpZBL/t8z363Qx0pT1cevl+sAG7QhMP/RV+ce00zJOSu3opmg4OORf7992P9I+DkQjp
VDon1i8rYL7Pt1WhBKkrmBONi5pebuwFqtFOykxQeJTT14vkqspkZUGF9LS2RSiLgy+X7YDDWaLG
TaJOoLkyWbLM+HKxe64MIYti8dpA6uPmhIL8lb4NOpns1TAsz+pXgkv+SDBvgA7+qy2XjNdCf4ER
bq01Z1zTxFx5wAiWpVlU5LJBui+aWsT7fgmIAedssoj9qIhFwV5+x8eToPRTvrLtLNqkhGhmfcsI
VBa51oaclTpx0mU2pSzoDA12zDaGIMGlzvkvlvNv/zZHUzv5Ohm4ehRikN4AeI/VTvlLHu7Sy9aj
z5vhcpnc8f/viqPXAsPmPivxNMj9ETqlKPoECs8xArlo7QRIey+2HWkvQmr5he1FibZLwZx38O52
ofHqZfZf25vcL+eShvXZjC9F4bVzHrCF/1WVVV3AZZQmaDG4BzwiZ9XtghB0OIqig4cvUeoyWc9f
xDyntXXOlo6uakJzsselRz+OUstx5FPd7QyYdPB8G1vTbLp92mXAqxmEKZhhdhmjrcvKodObgFH9
QAoFrrAiNqMOwD3pHswSsfqeYw+LaD94saLAS3197+YOFmvE4t/qVYj+6dDpQBSTwf2VxTkQycD/
g9+I9T/MLv8Z4KbevzRCrB+xAL5AWV0TpuNmiDB80s91QK5d91dG+p4PW7Yq3SAd+U1ml0GYvisZ
5UxIpKjnAVkPA/+yqCb2up3AQ+BfudFvdQfwi9TTI223YtYLlFHbgiHlLvXYQLUYL8ysTYgnAP38
b0ataa3R6dyg8dLgkM/KJU7W5fSX/LeShY67FBiqzmtHUiXvisW08hRwOjkW3/iYGs3L/FOZ1ZKx
5iBegKlMCtSRkNdog8FzCB8AJ4vfIgDMIpN4J4seYVY6z2KFMjag9vijzkwQvH8mbMji/sxOR04n
cFUJ3vuoTSnC2tKihInJ6i2sT9msWVdUsBmYqgd+RU68v4uqion88SHdEhYA7an8QV1ofCo7sAoi
CDXDU6Nh/BY+UNe12/hOChu7DNMMuQ3fAkUoTP7CCIIcR0Wz//7fcIgwkum76GY1qRsXFERI9u8T
Hsld7lIxpro17jQgAqR+NkRvNq6UguFHe44M6itjzkwZlMVgrD3quxNpxwmXYnAl68ea/GScI2mK
riPInrO8Y6+ry+MGoiovZnQk+DKNQQDGg85h0jqE/+7brfTppA4um9pEWpPJeAM9//G1Cri95DWi
67nLsF9WhVrVkmg1rzw0PwLFga9hmeRe9CV015GmHiO/ZMxNLhUqBD+MzuurdGOxgV1PwuXB6mLN
epHo6Y+Nux7pNR996BtwqFs1sSLN7fZJ1cwqQroaj9GtbHxDx2zcG8KQf4LCOVRdwASMWI+ft09e
RzbCMYR2CzDnAK3+rTUdKTPQX918rvNr4bf3x92o3AaxNSSSjuKFL/zVBW9xHTHkF0g73bDBvmXa
BvL1rIvLLxep0jfuv4UpzuzfE1exqEoDUsQjG/Umo7qwIWLbGuXy8CmO5O7Jd1WyoKOqn5SKOIyV
IPz7/KBuZNnVVqre1I0O+ktFLTGI3P6xR+zlxH3FxAZTWixgO9Ms4hl4ffJ4KUwMgjL+66v2SpuV
OG01um7vucj70vJnNsKGKMVJL4Vn1hcQgimNYzDWQfhCJucHbWLZhjb9XJDxpqFfvgDsMN/j/hPv
PBSC7C37Pp2t6TZAjDb5KIwMxAVLgNWiwfHIssoygHYKkaJ5ISv7K14c/Q1G8ZwDWJ1Gme6cRNFN
LLF8y43PDaOfvGV94PKNEL6EK6EggaPWqoWXJvGzOS1TLqBV92EGqgZ4s5/Y3K3UcJoAAl+2FM2b
kWCtMVHdKhcVlvn33B/ftWWxgxKAtgsuXu37wgv62sxUhtKIeF9XXie6AT1ULagWSqDdX8kqIdmT
KG4czlGCqTbXIFEVlG4jQbvgdjWfxD68Yko6KRB59vzlJXeiv+GwppIa1QCXDeHRZ0qzZJMnPS5K
2vPkigQVw5ZMkeb/D2X+xjGEWPSuJemBhcrvpCCdkk66e5zzcFKXGWP0e9XWOtiGqywdlfb9AWkh
7HnCoZUL5UE0iIUD/3V7whqqX0r/hO+ayvD2tgH7wr5T5o7FA8auVPzjC/jCvqLOL5aYWsAT69Oo
MDcVZvU9xnM3FfIyHoL9ILk2St6qpFv7T2RyMI6oUwL3A91S08IhiGjEIX8L8Y8zwFCb+tZyKU/a
JWHexa5RUV9G7zKgml8p4RRWgrHXaquUUslmpbOXJ/8FuxHqmy4UwTtBTWkYuqIkMRHklhaMxSqh
tUruC3+kjbz/hPawBDHYDbOcBEfLGBpVaLxDVULDePm74ezALYFimnZYa+8iJ9wtoszkx4RMk6Ot
hldzIXwJfh7qkXdloJTv7couYvbdVxlAE6tdmWyzNU69RWEgRVUcxQkSeM+cQ4gXLeebvqv5aV4Q
/sDS7FT9ac5RC5geOMaSO6x0407EagoGr7AIKpmL3zqc+dbDWcbSV4Im3RTMIc1ZKpGoc91CsuRz
pWq0/I7l1vB6wBgxedQIKG/ilB02kcaG3IjidkUIgSCKtxIni27h3Q3I60y0pqkye7uu5sj+toql
Uqw56xF/dUWbZZBpU0wzlwCF4d1X0lRbilmrUpTbWoRyRcnHjzoMGXeHQgnm22SCd7dPkYAij8kn
YEnnQzbgF2sfnlyXlRfdavawYbqBX05lbGKaTcSDzJXdyeBkYYOX2bj8c4quffcfYKyzGeDz3XBs
g6900IjrzzF7oYqlQWfNnKXBAaI5ZlWWf4rANPZOG4e1A7hFcTJEAx/F8OwwxtEQSbBxBGZnrLbY
qebdJwTT56nFImGKbdGca7YQzjz2YsUzgaY4NWn10wMAbNe53JPzbbWimXgrCM6t/b6Jqr1rsCYP
ZimzR9zovbu1wLAe03tjr6PEcZbcqhUMEr6MBKCGBC20kK2BREZuIhLwMiEvkT5/OJzTuMzVgKeO
pCS0TZViButSiJx7ACWMqJQsUq0N5K236pCny+G7z+tLf3N+DrFeht//M1KNKBp/oxL9w44xkwSy
ZJxmk3TxXT0Tr8QYS6/KPaBj0s08GezC3vRMS4xrPrzCBXmTxQNPVyC60EZ7Nn0eQpUDirX8Smt7
l4b52aBDxPoITLae+FGhyAMW9vdZYjJToq8wkYiGIbj+LqN2qTZMhX1tvoonR+pZudGEksRPiL8t
t4r6UB4CvbpcJ0CbZCk8YBSpyRNbkrq2ZCVwqJzH6pb1Pd30S7cTBlTtYjB8+IQyHTVf4yVuDVvl
vKx7jo4gJz98bn6jSo40TbL3tQvOUOnbYYfmRhSWFyEFNJkxZruLPaLdUS5yX8ecDf6nOX0uj6H+
6iTyprAAnHWplKc6iOpNvq9IMccUu/Y+jhVVAkNBqwPAytIt2Ff1ghZiKlLN+rK90N+0OrIcEtGp
W2WNZtmmw6H+lsGfgieSxOBvtnazC9Zv4dGCAl5eltQWtdoWjz5EFNDPwJKjU7S3jJBtiOADE6c/
EPniZ8stKqFad0nY/qJWXf8J7uH1XpIE08tQrveU42yRwnpWlW1es7KC4i0pHjv3FAkoPWxuUbA6
nvmgbBGfg5+OKDivE5ZP3qW7o2Q2VoBSHUWqOZm0a5X1qcIWIWh207oS+3Ojsy2cf803nqJzLrG6
qJMB7tWAof67sKd78hWfCeiOu59pNyGdk6krRm50g1UZ+MV/BiWiyN3WlpVLnEKPlBeaElS+GDK8
Om5T0DFKx1xOR9MMQnksrFrDVlvqhdiqMEEbWeJ5zxLZ+/Lh/Qob657lMb0D0sovc7ChqZxyUzCs
pnZmTNYjYNzNn6Rbk26aTojiMhtLilePmIS10OM9QMlqI0JpiOb4ld7QOMLIf5zYRLxuxHAd/Uul
T8uAV3vf4aXK8BLBBOo4/PYPczz8B5smhTVyCWbYZezEfe151y2iL2P9szAai4+XWcRmdcMB75Kh
tnrRtN0IQcE2Nyxme0pbUah7l07veYITv9O+42e0F7Fdg/BefpCIhY68gRztwO1d8MiW2elG6jIx
Y4mLUk+PrdtdBTy4S78ewRrmeLiJK/ymPMT7aACQhstqFetlorCVB0D8PYtCBhrYgeLwi2dyErxz
K+PvFd2w54y4D8LoOdShIj6kN3avwweZORxCay3th6gOXE1n2W6mINGpafONy5CFCnJG97FfC6mL
wR+ykEmhzv+z42kutCTOldTk0Uo8CKCCQg0SjlITDbvP/Wg8bRI7iECzi18Oh27+6phl6sVEkqGB
c6DjJKgOlSWMSRlF5OArB4j11hTGDN+GtG0B2zLL8YTnAcT6lXDYGzEF8QtwiRiG1xi5rGc1a6n1
ysjGYfa7fd0ujsBju+9k5YvCOizQhJpH1uubpO6LriKyH9AZRsJdRkTF9/RZZ6sUhrHY+MTZOqjZ
cB0nbCDh5oCKH0UyivWEGFth4EWFAwDDIIkejoOJBmMisxw3/0Hw0ji4IYkVR+QL+OqTGh4xOXcF
6PLIUeZ4Th0BmMNcu7d6VpK2aHqJPyIex76IQ3t0z+5gdQHzMZcZQAPNg0B4iY06j6ZV6jMdrzUh
XLdvtQxXujhvAHLjQLnUt/SBk2ATxunBOGsurEa9niaIZ0WOLWcaeXJdI7iQUBBobbTN9eAWadYF
/ZoVD4M3wcIvi7qAECwnhHQ607QqrDaqgai1T5L4udV++D/lvmSgf+f7ZgJX/ECx7DfDQIBXpMHX
W+btnu03fEulfOi2N+tloEQBmvwh7n37Aj7ETlzGd5mWAVK3CW61MZk0aIc0oeEEelhsOiuYe8M9
/RkZwzLyBHQKZ0qpyO6+MZBV0PQTiS+Qt7M39J3nFtX/tJqb0a+wa/aVj0iJGDuCDcrXzPSD3A3w
9aTXRBKy390PrkdWGB3whNvR4ayyX3Ri35AqHnHPNS2Hqy+e8qfZYddFjy3dRKbijT6t9iYGMTRT
YR+kZ2SCyztLxUMw7ABoolHCaNmSb5o/zKvMab0CyQuzpLM5sc++xf7T9cPkAA7wxbgzm8aj+tUB
H38Er5Yu/6t/pH5JCPdlAiQJ/dSM/0NmDh/neNJDbLaPDbWNFDByJGzZ3235hBH5XtX2Cn0zfHTX
h2QwXyVzLR8xlspPYwh3IbsvEK095qs2luioMt1na4Sun3jxHPGti9YniN9TUWJUODHdeSCXxm80
dUKSTk6k7xSulNkzNqeM1Sk+qsQGI1JhuNEMmC0qBzm+24BilNhgY0f24rGCQZzWnbwXnG8pdfyC
81shXbKovpVxXxc1M0ns/75Svrb5fyDsqNqa0j4m0nlu7QhtEg9p7EDgTFBLS1J+HpUzQ5e0tKmh
aR+8lVBVxrbcDjwnBnyg64dfPeL59rSteq/ScXpLS0qIuMYid00S+mrGsbq+CjYrM6sfSIBg7u2t
0uAjYznMKEcjUWbD7lvjvEETH/mxroxr7etuyVYAwyvGmKLi2JGJhr5QxhWIAUcaIHRuRW+CC/wZ
TuX93huAizWrl5S814o42Gx8q2Uv6SpRMOctrsOriz4xyE7YomCbmLfOFfaGcdEuw1gZFXIkd1hn
lGwwDk+SZAn8ExZ0a4oxqu6UteKmjvzi87+GsdNTyp+HB7n7/u2QizvriC36y3HOZG6xfyt5wA1n
nvpP407aoSApk1+TKurEkcyl2991j4XDN1jDmiabneBfkvLy1Z8Iu9z0F7mg6iQOGkezkWNpvNfM
T643QHSTDJdXlc7rhUGDYtrR9/HLTesAcoOBgF2thy+7Q1iLrFQgfViVrtI+bocBXeaiUtnJgORE
UIb0UrUChJPb4m5AlTau5cRo87X8vvtQ2ZtgKhZuEV0b5JGufe59JzY8IpGxkfdNjD4YIFI818nb
AaydCcBlLUgN5dvkQmk/r+QPZ6qvfbxp/dotvKeaqlrSYg7v6lTYrdsLlYDuuGc9Ibj/C+DSc94K
NrsvumDFBBB0cV9aqo04LU5sw66ovo4upIWSvMAv48DZ+rBKcPHnquPqlKyZ60L0H1H109Pwp7xM
+fnfWZMHl6hiycf48EE3h7ASfjOAus4tj0kafoG3kcnnkV2LfgB4i6L6WJwhReUXUE0e4hsg89uM
Qk+I4dIzQVRpt83PLQdYHfpD9NO4hlLIaRzEYH0XcN3CsUlZ3iLPS5oh/Fcov4MZou4PrQYTgk49
Izywtl0EDBWFZtuRiT5BwTGrccN2qkgNlU2CojEyXMY5czEkWEA3GaxnfO2m+FIpwBjLEEHUNEdB
W8R1gAX/f5QRSM/LItvvbi3KaPKvK+8/m8mXMDQSGenQSRRK396Apv4Ha3kW1sGsWZTzofCggkgX
mBSSyaHPU+WT9naP3UxvBNyQD8tYMNR+VJtY3DBK4I7xm3p9LMl+zsWIYaLRs1f5daMZZ0XicoDN
RYvaZ6bAXWisZv4i25MOtZywwaS5LLQ9Zx1n0ixp90YHA1SPtFfMYVh/tS3msZxqS/Nq9QBMkbwa
Kwt1uTHe0XBAUbkRSQDPN03CNasc0IUNRlGuzOp/DaLjVyQn4RVZHGEBcnVfeE3MGY7W72t8H8gL
dP+hZNuvqB3/La21t6RI/MFI86XgATVIH4sloga+exY7m4eBvPT8f1irSiYxDhGV9vohLEucE54E
913hq3nTT2VYhO2TrZvK8eNm8m125Eq5Sayz+HMoqbsq/GYnDIxAO0QhP4FUDFYcGMUnc3wynSSh
jIxbCrcYANKKOqXpxh51K+0mJD8Vm9ZFbmz5ZCXvjo1N169eiN/r2HvOYmNZ2eVzmWX8cEYsbLV0
azDaHhp5xDlEcKNUbG+Jsxr5NgR45OpTkhZiRwo+ouTPPfXUZBIDjHhQBN6noXzFiKjon97R7YyT
+MovF6VUpl0FaaSujX3LnGEJjmekQttg39D5YmHEfbZhdc/Fs19aY+g4XX0MATQ52IqjX+xY+aWm
t6QtGsn8mVGqTn/lbjHz798FH6ddmxN/CgcAzIXASj0ra2twndHJCK7WmDpEzfklCwK//VPHuCa/
J66SGNYV/0z4RpeENyl4oSB55YivboAsvodRnlYXjt8LivriFjA4m0ynCXmzGtB5ux5qc4hyBz8n
kjeUMZUpuaCRiwKn/27nXhBh42LpQXeUfLw4RN60Zl8cfghPAx729t/kYIzKLnRrqOx09J9CXinp
SW6eMpJEk7l48g3mShMFK+kFvVEQROeGi/XypRVJAPsXFk030FeUDdsXb8+h9YWaCaVaquxetzWC
JuT5XEZZD05mDhRie1J68BSCgO/8YGEcOF/TuA67I7QWA/qh0Kd7XP1gxl6YcEl+gjDLWs6GZzQ2
bJakYjiGBfDREDxhhl7RgDyminfw0IUsDAI+AQnkaMA7j7W3kBcQcDut4WDZvzKm/OS9K/TPX+Xx
09Ypbr4jNlPksrvmDtFRFFjE2fnnQEt+hPWPoJslxHNn4ttVQnptzdKrEKebLN+zlBF7czk3l5Jd
mjDk3AF+kZ4VLS5KLiRgyjHAMKG0f8zMLHRTVcL5kn43je6qbTYQXp+TIObEq/Ff9XC4RMzXUQ9r
/rI/QyRFnw7FpbdvApysjLISrd2VUpA1vwA0Qc5OJIEKjmAkNtdYtP0HwR44UfnX9lH1tprOM++J
uOFTZOVEie758YZXuM3CjrIxnQScnq+fmvkn2EzEGpAE9A78CMaIg6MDGE+tyug7SzD5t5wWhTkp
xCfHGWKMFSGSakLeeMqV7CaCD7Gz47hcuydna91P5Ztk/SKvHOMLNeDIEaSU//G/TnZ6UJZevO4+
QKHpwWi3AGCbiv8tYDYQ14c3VyRuuMlPf1Dmz6ZffMPYp5rGEsx4bWB00whJm6UXKd9FRuKE38M0
0v6nWfQNA7wQSPq/6grzBojBaQG/UMNAGuveewOhesmBjayhup/aT4LMw6XHTgx53zE2icDCR0Mf
/FfwPxJRSXcvFwJGNsrfERtVEndjPsw4dlXlfpU3kar/rtfQLSJLrc5MKNikbtHx6s0SgX0IFPxz
cFrwcAmTRxFK3b6eGniEsNIBi4wLx4XijK2JZbnVTecK9Ycnz9Q/Q/xojumQkzI6SFTvunrfnptU
Qz5qeJdeTptxWMMiAQGqb08VcrHfY7tyhiNvADBvIH+Lv3s2dq28WEtqtr69qPKmc2BM/QQeGw30
vTO7LU9Ih5OdGpH1HWrU8ieS/2Md17xuBYn4AjZij1JEwcsSyzs2ZbLW2T+rBfyrcSitsug/8Sfb
YzGpzBN/Jw3LDi3f9Ng0KaZOeENg/4GCD6xsru9V43ENW/eC6WuKlEqgwDFggQ9LC67sxdCLsJsA
h7k5RkzBthqE7HWTirG46mUicPS+re/Ufd4Tf1C7ZpJUj9U5qJoyAnHCPlyuiIbBn8H75mcXezPv
elsVgishqQLH1RfFN7QywSl4AVlaJ4YpKDpQE/OQBRRObklaJYKXbu9y/hU2y9L5qkJnx6PujMJH
DoYCwpNiSZhzJHn7PaVGASMjbltHaSOjYRw7L7nK4ehhlE5qSm7XSdHl+sZxiNGMTzRnIHXAoaIw
d+nLYh4kZDVRFNxDPqeTJ7EY2ECMV4biaICxRl6wDhXhG+yISLl2filRlI8ZgvQ1+6RCtHqc1bBS
2osFu6CdztyGstgtLW7kZYjKQ4mniw1lFtwvPo9bjlolQQCU1Um52QvNKMF7uTubMomCypbG4rbw
JHflttyD+JcBQGL8V8zCctmjWTY7fpRi8URy7H/v9nZi/TSXz8cfQ6TgvbMIbpv/OAeTdThs6i0+
29d2QOlpWMhQFSjFYbUpV9qZCaEFSmkasDNirXSv250V6kQzuVHm0JPFVGJUcUGDfPdb45z90zWP
EF/2qgUNHX1DMz7zZIjdcudosLtP8PJ+O+rC83ncMySw8+aawtFRNd8zhQFAH3gIjlalGheKguJR
8FdHVQXHgZgSZ9m7H3hZFFXyhWcQQtGzU+b7SuN6n7XccF1y6h0TPe5ODhNyeMvlvscdHfyK+poR
+AMK1CL+AMHoDlovpT84mVRCz4sCHBMQoxBMTBYETqLBP6zC1OfA90+sImyNehShH0eKoo1YFNlK
/qlxWw6mzfC/B/CW2k8UYH8wa4jUNKPEWW29tSML1+NbUang+D8YdsBsBdlJxILE4MhjlSWr92NB
wt6XO9+GQ9RugANCJ4etVPUtkACOnkVAPK6YBu8QlQoT9AvIDif7eK5TC1gbj3wolDsvc31a8Wja
GCi+xlXR5MyMUVqWOflF+RqmvtLnxLCkOufdg7bZOmdi5Qh95q4GErkWM/rP1EMI2KsImgZrdHZg
joqHE0CfR7mMZ7mTR0OiuXKeLqKiQXn+hcQGkqdU1svN+UcNQhVYFqjW9zpck2tnt6nw4igScQ0r
nqBNdA0BFZqWF/5NxNOazN7LjmWTvxGXrHPiVr0AjbdWmubROky2w6ughGr1bGJy19RwSmDVbB8j
SISyMKjHMaSxob5N54iHt0MuR0vgE6SgIN5zBoFtm11j5XMXCOsqaJfKKQCisy1cyBkdYmH9Xnsv
UmEkmoZ/iEHn2zl2nDwn57Bo/ykmBJ7XGBAFHNjTSs1WaQOlm/aWM6wCScfHT1lx0vTZtIkl579v
QSHDVfHpfOYDeSzYESxRchCKIinDE0mcihBC9ia0g9HIGS/2aiuArfG4q8YCcMmaX5z6qei6IlwW
fOXpQsOleq/W8rDdG2zO+CXXh9gnsPbLvzYMvOoRzy+ZQkP9lIZnXyiwgWjOTSAVApQy9Xy3UIS0
au353kZY6/XoXBdlQr4xJ+kIY3fe83GRaLxhMsh1b0UN36+7crl6VyCndjsDkoh0VXRmlrwypZkr
3u96fi4vD258pVWKBhIaqI248O9lh7dUz9+JbZ/YtMQ+B5N3K+Emu+kBbWRt6+o3zALHBjSwFyaq
QyEQiqE0vvP+E7onDpgB4+/MgI0My0eT2WrN7enGRLsCBNDEOqJmv+kiRZg1n8WFVT2OV23Q4PLW
9qKO7d8I7bjUvsplHnZJulvAy9t6wD0T4YUHYzHCUU66CqKFcGVxhWmC7wgOidcZCD636tI+mZ9T
8g/WLxXO6c2l1zodqWyQAR3mQUbbhi3q8ap+/vX+6n694pMU8oF/7NHJl+a9XbIFhxtZh2iOZMSn
bRgPAjntwGbS8v4kvyltsuuscYe0TMYXyzgS40sGDqFQT1XEAL+7ie+6dHDUIrzEIQTOU5znpRhZ
SOvb8uRItF3zGKb4tgXol9ORKpisPcp3FkDudUtUvnkuCxYbr5Qh7be/KznvVFR3spRWmep9cp5S
lP/UXGG/IEJAO+u9mmg90+PpgSS1WL+k3rfy+Gf6RK54/1aSMI6PlzLigQ5f28Qm3QIYhR5S7yPY
JvaH/vZw7y+glKkOs5Mcq7+jYbA72aXuk+XW9EDxyzeOYIHMngQLmeK4DrIqVVRiV6MdKcUhFx1g
3ygzly6gioVm20Zuhj9pdpb7mj2Mt7wsVtsdvbvtDpST5GTjDTzabmRh3IJJImm5FVv9ENWntZC3
APRXX3QeIjSot34b5LNgKahJO1JAIvDZxg83b1CwI/X1K6AWgGbYVnunt4+eqFoFSEcAvGVETBdG
6vxvtp8O8FOW0OHAImW4N4Nm8kmTV4vuGipiDk1R1nKbdNkrDOdFTiiSa35nYcqYL+m8PGMKHY5o
AyykRrW5aqnHGQXU/ovUSMvRcxIhNfI7OzQ0h07S505hrnweNa7Lh0EP0MLpEMPgRlxtL9AiVsUM
W9SaOJ+rMWwwzu7kSANvIqVL2tbUqWKUOyVwt+oakQPtlJPWsJU2YrsmXDtVesRLgmoFiZLbBb9B
L4Xo3jHrESnhMStzItMtCdm+V5r8dQSpOX4qfHCqi/h/ChOi5+XKyhv0woP8b9ljP3PQ5T5KEYhS
ny+yvMjB1+KD2Q5shEIButdXmSFZsDXJ3NlZYzwA+KeYoyiNmCnnpDdNOIJydlNMs1886iu3f4ls
mjxDnEPPAlnQJZYnQwh+ANTKLX24w3mzCpWl96lrQUV++t7Zs8fyg9pg5RR96Daq2gpRv+YuFoPE
YU2OJNoJ4BcByrBmessypgLZEU3b+mubzd6CEqNrP+N6Az9TVWmfCZY2zs8HXgaXeKRkZxJ8Mofr
TV4nR/sTvty7Mh3JoZyC+Ft+R7/7XySxenk0ashrnjSGwcPFSH1OFVuBj1PV2U1fgd4T6ouMxWod
HJFOIxkfkKwYS3e/0u6vz30o/76VltBi+2LYdJ0KpjzzfBqcPKjNv67V+SxFItNct/ULsD0MAa48
UkDaEgAL1hoPQWFR/GEqVusQtQdtPQ9v9Y1zAhoJO+2B9MGETqMEwBULvv3RpxUNR5wY58rk8fO3
ocUwCN0cwARZcDqJ+8yVskLgFFRAcNplZWBc2X2KizHqL6nKqU51QR4F1MlaaO8KYx3ERDiPxFc1
wavwuxWBrkOtysESA1Yj+AtSAHgUM+M5TGek6CRaL5iI67bXV6EtTRHZQcCCjVCVMkxjenA/x1y0
oQTXhmAZca5vJn6YLpyCZs2dPa414E6UCfOfI8iQsGu4ILjTKGSAmM/koxgPVI/xMO93DHMKGE1g
7qhquwfNLda0fhxQUjk3z7HXrZc675Gfrgvv72AX9dJmTyC9Cv83xLxmwKC//Oyp/+M5wFWBmxYD
aqbGGyNk6+XKAW9QBRaklyQbloAAb9jxyrXHE5fKhkKwSZmnNgQ/RUC51VZsSQnV4y35cY/fDA1c
YIUmja8b8YrDECCRkGkjRT8Y5Eloj74NtyVyEQIJXCusv914Zua44zMkYurlVzHqzGIWZ6egNhG/
nmjOtKARvsunA4efX+ta3f9uxH/vN+xskf8FoXtfMXtLXxopxHrqQ1dV20l+vNt6IOM/AI3926hu
5ZHEPxGHCZFlTZ7KbOOjgz8E1C86XAm9Bl0pgQ0KxzmkPft8dCJbzRRRH768E75ygF2wDaemOFvM
qYEdQwBPWqyRq528rvKzEjw0z+68DBqd/8c4o8defKOq/0xy8ahF9fWe8BCOULN7ACpWdQVqXzTg
m1RosTxyNJLzrccfdGUPpKjnrAHheGwwKNLbQaUkNeOrZndaOQRxRAxM3+QMJXE9ygHHr3c8/ZYZ
jOVP5U+9CdEeiH+CHbfEsXC9mHZo8D+A1U144pgOvm4ENdDcocSfyQS2/ek3+hg3vhOxSMgA5hSL
P4QuxGzo5RRk2KfXVqHoDeOeecapfJSL5f9SexPOzvtmX0hsm+mWhpc+eyOyXNeZn5QNjeGobTn3
WZ4kGDXWI4dUN7ViwUcG76UNSUPAgwD/wflWTnDDl2W8ZpeiBywt3T6zB2o2P1Gbr7ZzmHeWZXPb
u71/i/YhMAK8Xr7J+AcdtkDg1qG3GwTQyIvAyNNTX59tMCCMeR1vvSNlfaQuWpm4nKIjKyOBx8zB
4SDGIzDOGHFc7GalxHkUrAqfm2bEVPe1JJnk3Qt0/F7MLjEUrTwNYFhwLW3rr0ZZS2g43hg/kAwG
WEF2fWxjdmfxSzHvVBfi8u3M2VM7rBFx2QLwMM0Vy0JDNJVQmoyK4AxmceWMeOZSxYF4GUjRql5p
CYAyA9SkUGDuoiuYyws7ELSBOO9cpUEd5/bQydUe/BuUnVYkC0a+dlKKqI5MIVMAxbpwQyQqjqxJ
WkJBarlArIhZRvWW47EjO3GbZQnz8Golz9Jq8T9fNcJeuHu8avb2JL23UcMYXA2PWr2ILtYNm5HM
sHzcCUbsxwVaGo44QPLvzNvy592kt3Fig1dbOMPVsQb2n71u/FcV1gBWxd3XbFXj6w3jOJ4TMQx7
VYBoocOG4nxqKTJaun/YWlKwFmbgDBeqVVyBXHTYcn/xDkz+UOZaHBr3QlgTx86TX/ZM+o5qs5Je
eTAeczy3WzbS8i8VC1s+BitX+LgZcDGB/eU3rtUSsiMeOaH9/hAJxDs8m13lyoxZSMNLIN47ehbP
0k6n/3PLMoa1jO1ZF57PqujN1K5Qhq61zc+0IdgcflLwzLeukU3TmiK0Wx7XCQZciERzsKBNP+me
LL5rWgCj1J9yhLZJKhVwju3jAiwjSg7lraAYXNdc/zOI2sQbPso13WXmXrfLHzUJxxPUalC4kA2U
/Izzer9xDBD4TGm+NReDlHsRYCggH3gyhUoBMKUDhJEEFhBwb2jRyzeLWDeaEAUSHUBRO1xeSp51
EwcgXf6zfU8bm7lDZSpvxr0Lsmf9GRp8O5Bf8TFS4oZALCjzwFz5OuOOoYGO6kKubh83+hDb6PPg
tMYmNX+5lWY78VlhvcgQqwQSFMFTGV6nyYMZY91Wce4zSmyXMnW2gvk7hvlLPo1cFj5aXiNv+xfk
dNuS9A5fXh4JjYlhz/aItoxdCtdA0QKf2DZCPmWDHDGTgAJr4dYLL4oY0kZnLRGgPP+bXQNEfoY6
ssqs34XC+L44GtdRs8ioljCY3dyhA02JRsL4ls9LmLaf4KYUqivanx4T2vWb61gxAjCxYMhZMMuH
QeJV9ByOFVlpfaPfvOPUosVnIitq8e4zXPWyFsRpHDWu1T+Z9GpzoK/G1ZKdMcbbmdVaZm1ptuYw
TL8k/cyuPd2RQx6ercjOHZ6A3FO128AWg7Po8m1oZ96bXX0+Q/IFq44WvKOsE0MwVVWN32KaWE6X
Ac5+HZE5jEfb/M5prcSYr1nlo44a3bbnp7z7Q/FgY36Uu+nXYsKse3KHd7PwBymG+0n7p1Okbg8V
uLec/Tuq60OugfKzkC+NhhcdWIeNEVBnQDQHhLEPSFjcLF1/Ruu7ZLyJ8gVJ5AoJh13s7/1LwWYs
4+Xc62psqgRh9pdGgNkWcJsaSdpAzuVZlOT0LH62vv7byzqKSA2JI8p+PB0y9dPxvYQQe8LTwEqa
dBgs3RsiKAzUAZeB62OG3Z6LCw5SzowwwRi3rBiehv+5zgw2k5MD/ErPrGfUUZuGkkQEnTv/I5Vt
vwIQAD2N1Q7Ow9STiJrqGHIxUtELar0qNFUHhD/lQydWOcqt3b0KL8Z7amylhOVcVz6v3EYzhXOH
bJJ3evmluG4VOwEzlXGU1cOpq+XxUDB/1AYIvCkI5Z/mgCx6OONeoVSio5IS6m68qElZcvL5QCo5
C19Vg74bZBZfoIyzOSEbyzhydxH5r9ezqxhaSwfxqB9jWPl9RKCnU+9v0GctHrL8nZ7PRaBMT4Rj
YMM3CyCVS71zRhyrP3cqZuKbdD7OFf9Dk8KdHx4S0p2u9FDkQCJJz0SqPSAqbX+fgeGwpPzIpIvP
K9S0vKkJeAbQeZHw6l9l8dGDd3K6hfDEFvSjqAXQ43W1V1/7haIQcOmMP+NJV8TJROiTE7yfCYwU
9b6HLBGjrFnHTFoNqxWLPn7xQIfNGVzbfizM95uoj6Yca+47kCKT1fYO5b16Qcd1tpd1NtQaSfEx
8GodMFI0uHGiLuWYVGhZ/+pUgyoZnmHEoYmIIQQY2a0eDoX64+LGjnD2s4Up+hdcWmIRFV0zgi2E
te2KZyMl1coxgkNmHjDuDPn+jhpVcGyuosABap32WbZ9lI+cxDV01GJAmFWrkAGesE6/DxYn80zP
/UQ2xbpgKDOskMQOb6O9SQ12xrsC+5WImIP/jWV+m1Kam9o6fZ0uR1BHTy6xcZZN8TgWvIYfry11
5q1XMEUqcJLL3j8y9np2Pnc/Oc9FQGaZNixIrJdL6rrGE8NC3wRvhEXciqPg5KLsKaF8UnOeBBis
4kGNnvvSlkpDAmHB0MNeimacg/uPvGm9+pDIMHW3Ueqp5SVjSaTO9+5c54flrA939E8lhE8Q5CE1
5pcvL9cQSGAnLxHDtTNxH/f0Lovad6rNyinqy9Ln3drFUuiYGphLw9CdXdWKEInsteTwqh5TNuPd
X7Vzqi6/jx5s3r8SMJ78aDPTRHve62DPXsSkSxGjyOefLvY2jhXAeDNj2FQXbcqFqzVWgvxWnM/X
p/U+zJG0WfDt6yPLJdTrMhuL++8JVvsxeYJs6PqEHSOf+e6PAdIeKtnkwA2BsJxscXA/gY5yxz3T
/7ae9tZ1hPJm4pb+tGqHYHOmt8Ut++QmtQfTGkOylQnbmtPHF1UTOK668auWXoPuOPxq246QTwx5
/rBO6ko8ogU8BerzYzETk7OOzmEAkIteV8DO/ZIH0gWxuPpUoWoCVVACr1TpF/LM2qgfC3Gjz8c2
VvpTm0XOvVfaH5B9VQnffoI0VUOtcwEQsxNPTh6xQwV/PfVDwkqvPO+Rkr+Mq66Ao955W8K0Feyq
6iPQ+zIhh8NOXGWSOzEL8u0kt2aL1ntR62l5wSH5kg/KczJmB2V53JfmDVzWo9X2QcfSEzv8Aj5Z
qbnQPPIDLe/o/wANnyRsJbSwW8JRIN4adWFa3tZuR0WA3u+vc4E6pmQeFfPKcxYA6lgEDHi9MuRO
VoCuS6Q4fePOZUpMvzBXJNfL+Cb6LljfBaiu/1jVYZAH7IZKjwDmTxMV1MwzF5Vq2S4P6vRQLUCf
z2WiW9hZPuJkeCrJ+AwsEKw/G2je+kIoRJLNiffaOA7/WOKr3sJib8TqQXxZ8XelZHGGxOJ7P8Ux
FIqOz0wYrwytuvE446NTlIzcy5AGrKxbU3Rox6zhzEOjdPS4zRl7oD1VUkTXeLeeEsXRRo31NfN4
JTq3tG2lKrANDt9ygVqpK2Lrvbym6rFXFXP4xj618bMwXUpY1WbuxlzHmHSDt3aH2cG3UEcMhgie
j5LCtWjemUzXm2BH7EsiVi3Sz9rQ5XzalaqRHImvNECjX08Js7WNIZNgLtohcY33I/j635k13SX2
RZGaS0v79DeTT6dJnQ+kGqXcwu5z/WPlMsxG6iM1BzvlbdFtGUMv7e9xuq0SQpuvEA3JIjwTjxrK
r7lVzMeb8fk3Zt4vlKK7G21KFHr8pHAvfY92UZDVSYppBECiBrCV8Q9295pX2/J3ei1+Xo/uFkCR
M42Lppx6MGJdVD+9tBEYQOIFUp6+9Gbpf2BLS91hFiGZvi18byoWxNY4lorayBOQXx2fwX7nAk8N
wxYIsHCK+C5dBK4npArPYf9idZHSiwiBaRzsO5lPPLphEkyQHjY+2LX8I60xuQSz91ia/7o8TGxA
lFJoUIGqdYFu9ZZJ1wwIxq6zEa5bM4DwDezU0T0CiMLIdSqIgnuPT5d/8I5e0/qSGuJekuy2c3Kj
N9gtVRctCN2A+wnA0Yl1KxNtm+qiz6feb/f1ZQCwJKofjxQReHEkSEA9yU4YH8gC5cspL90MEap4
jigjDoVJPEQcpGv1Y2exg3uqRwBeDhhilQC7ssitISKGZctM5CxSELvj6IIU44M9haeCxpN45vNv
2Pza8LDXeUeCJaWPIQ0dwblSUazChpQGAQ2SFjUcnaCq7Ocb+NXz6dF6PIB2ac93csXPL3qQ0kR/
FseReCX/YwMyhAnJDcTkK8RGcg1A+AZRDx8tbDiMQAMD/hl6P0Schto88KguNurUP6FLbYHnupED
QVb+HmK++Uv3iagvz7eoy3V9j14UtSnOz6sWYhM9UUXkwsSbITjKYSRVdL3FZTDJ35JJDo2OiwPM
i+uw0yFHMqcZsq5JF50QjSnDn9awiHWWt5rA+DPYeihjMYwZuqLaVjt5hrEPyLeMrvRjW+6Np0Jp
nivIs25NVJ5kNeQfdcQ0trp+ktRHyId506ehxms2L2sOnAAMT67vUT5SqQj8dRqJ3+1HWStLjfrm
UeNe22sMV1JWNCGdAiTR3181QRRCGbmh89AYY4J/vj0f9QnQcjVwDLjTIY2eUdgUqVNopNYXhYAd
7fLyw0PRpbUz1mfs63V5aW72MysXGOdYjGwVev6LOnXMsFiz+vcOQr+pjt1mbY++AjrxQAL7ZVgY
Ge0S2KmeGcr5JJvIFtqQ16a4uVmr6LmdyRWlhkdw4jlyOuBEaCusvqg91azJELz3chs50VLvLAsM
855jewMHXXqOWIhJc++50K5dFzbwgKv08dnL5AI+SMqc1rO1lHYvkxixB9OhXw4bHsz1O2pF6qzy
R6VTZ3ZobWx+wqb8DIp2UKBqs3m2HoJ+Tj/H0KnVnASH4UE8rtA4O8vKjoDRdsi8XU1B7zUYi4tw
YiJD7N9TGk1omJRYLqAhPA6gVs+BbDlKEDI9xddsXEQ8OXHWBgCy3VA+w8CPrl6QGwqOgL59m2+o
8eW283cDKUfL1VqBHiA7UDD7Tp9B3rpFEaWEjH5mfoCbUemyFDNExAovt+MNFH6fapL9Wfj3Az9N
ZGOAcX+hx5HSqVeXSoqj/Xi7xMDYOILdKWAY+YO+ZwACYQOqkLDCBmHtMF1ZA+vyinPcuJABr1FM
rE//wImk+nSSA5bnxGqSaY25sEP0QWsF80uR9lCngmB0x/Dw8cMcxl9Kd1CgVrYdfDaitFKKOOFe
5h4Fm8dwhTpZKXWCrCgfI+rUTlKTtoIEM4n4GK88edDZppFekF2xLqC6mJdIK1uRRJ8vyhXdiCEn
BY+54ocMcNRU7qw31hd5HITf4+KpTnA9Nr4ptB+ePBCpOhDs8qQdS1KCuCsBwi50EmYrOKtsKlEF
1cm99kHmYEnEGS8AA2pRf6O3hUrA6SdfC7FJnu//v8lwdZeAm58ZFB6mScTfUB+tI1rvucJ3CjNu
jeXG/15xOhNYvgfg9jzld1SUatyS6KaUBwqDEZ4E72bbGlE7992lCJSRRBVpaH64OgJWdK/h/pcR
InPmwf0dkhUBqQ3Ki1GW49PcJg6hPM1C9yuy9BYydlWCuUZBbqYfTgfhETJtVDTPaWJRrmk9w6qd
sYSbszXXg8oMgOlWpzB4Xwlm0YNMavKu1CKH46XPfgPrA6N+5JD2IdgJZ+H7KFEnoT9GG4zH9bn1
b20HbybFQiTVEdV0UFQTkYvj2RXya4IUSB/0Ph//U8ZQMjj6e1Iv8c/+FklLSYvNydHlZB1SIxaO
arhtV8rzgk+iUbjn4buzNZG/axo9TvjojeQ6X7pwcbasd9LgY/6o/Sr8FU036gqm6SasxnpwlCN0
IXbCSb38uEDM8iWISVJWYVmO+YPQj/l44aeF8VDbzE7QXyuDQ89aU0xc5B3wmFRsae4W3Cn4xPMn
pqWkPLCFVYE8yWTd3KR5fKXY3fobc9cHYelxbXupifCA/d236OuKWtIuKGoruTNK5+YMqgr+vbfO
Pc/h/mLJTQaUwLa3UvKxZCtjTJrhTGBcBUgDY7jmyokFaD8jM0V3y6Dz6jH+6soEWTe2wQgqOdFd
vWCESjkDN+LffxIm25JXzXVmBv5mOw3GdSWC/zUP2BOXFpp/vGXFthB2oSKmxJO2PHg+fgrolrYU
A4Ux+rjkXl3cmXTNTXUbwEtMNvX2fO/YUxPLkYLejBGrDTYS0/9tdPTFz0R5nxMZk7adzgHrbI/g
tC5eKVJ//JTJNVv9hwfvSnf66wMq8PCPDOBwC0wZOy5fmJ4nIxQahFnUZMdQ5/eueXC55QjatsZB
cbB8o2BBlQdttEiR8rooUXqljw8wJY1CU06KL7s2BaHoszLkYom0HBX2mQb216P5wnGQKeBaKLGX
1LWWPf7BR2UqZIW7InQ/9wwYA1yCb5pXSxC2t6VNyUYcaWuPTkutHc3Yws7pmHQeOqzJZyuyQ2UZ
c7XHakLdo+xftFU5u897GGGr0swgFRLIgBbrY8xEZKuAYZCnDwmhggnrYRzFUYfOzI4dec+L9kpK
/TFSOA7WG3mpqtJhoMPvNucRav+2RI8ExKutX8+/pp6bqQ2HIQOQNRTm8pn4VLqc3FEfcgdTspty
VenQ2wu4P1aDD9dXcCrlKdUKO1Lw2QUEL+ACqhuPG8Z0XuhR5T9ZBOBf9xxndvFc7clIGyjlERBL
NQfOtBiomKWITsni4cbwmDMCADrJ0UhQQZ+/ziduTP5ahFXbbrWhYLKl6oxhfSVlV1/Ybw0uZUAz
IXfvgZ/watdmPnMENtaXgtYKADB1H/+YXuEWx3Z7OG87Z65oS2/ofrcnokHJ3+sexCoE7CAEH0nQ
N1dyzHKUQxDoQZZGP8qn28Ed0xygZNOnQ8ok2OAuuRbyu28EROUMq458inSCiMuXwbUEEj7kPIEF
EB6AUqykWBlMqqBgek451RHDraSWsEqMf3Di0ibt1XU+qtf7OS8wwoyf1Mjg6SLSFujKd/OzRZkc
5J3uODWlmIBqLAXwc+RhO6Ws2fNK/k8c0gZykdYXIQgjQdKtokg977RUgo5Vx8ds06Xxzx//xeBF
Fd8Pc5wg6MH6zzJGhkn33gdiOIKdKQv0m1eR0knDo9qO+Hfnwrw1jlFZO7ZwZX49TMnnwolyYwmJ
m3/USK4tUH7ZKF5nnlH8Miyuk8E6f4vVTjv1SlDhxFHNc1JApRnsuCM5t+2qFJ08J0KkoA8uP4iL
5xM/LmQ34TckasjDCj/NboThqHAcJE6H5+2eg505bS27QQSh1Rbqm48U+V5wc30omwoGm9gJ9v1I
rTbunyqFolBqi4OhlDkMdU1QtR71f82fVEtWimGTX6D7OJDdnah0sOmRabNuiCGe9RWlavyVcUxB
66OgppVuQHFUNiylNd8mEqIEDESHAHUvKoJuj1sGtvojqU3IGUL2dZ8sHc8fLDgudRmixO4+ChRj
c9EwJ/EAZWN5khpXpHDGK2pnw3qgrGJIdHks6gefn3kKqeKvC4uJvpY6EGt79divCAozUIzyFrXa
mMrf01HIUwm/m71V3MgTP9V4HG8fyonkT7jb5XK7ymHSF/oxbJtduz98jtDT0VjjKbdwwB4HPKsF
0EU4xTwIrzAwb0h5upqYlO2fUHJD5mRA/YDruIDe+V/6qfDoKbWikuGuhs+c0KRaJ9YXJhnwuz88
kZLqNvdC7D58Ex3R9O2sdG/AVXpPSTLy9mUu/snAQfoRDYEpGT9Q+CCdcZKpcNOmugRHFx2FELYi
0JWnTXIukN0iA8BUkEa4Ey3lvxwm0/R8vx9oPjjQQHggWc8jenq0dVxtsb5bZZjXYkcgfM83Os5Y
RzzltoWt1rAkcQShtk4mKru7ZjqwoNnhvZ1GT5wGC4pQwLWGTbBfpmHA4iSC35+FCeAu9tHa1ldQ
3dZcKlPurl7TwHRNcpKPwTjnj9LkpNDcbFIaoYJUIIh6ws+lnE8Wa/UfjPa/nhBnfyuIezWtkTAL
Hr9UTuDq4skUs8PUv4g5muPN/kAX6Ek9A0Goed3bo05YNUkuafcLjTx8ikShrkdC0IVWkfclos2C
i6CCgQ9rKFOkwXgNTS5zjD0b8+qVAndBnsQGWbW5h6KjXMrApuCdz8SRPiQ+3hvKL77WCtRJwVAi
ge+wFfBzAfUsfPU1We3c9WoZ6aijV4skViYqDOtC/AYOaoESWfhhqsyR3QIK9OKr27uOoEgI4NS1
vUcijKRr3d9MfUIqaO4tQGgSjIWJil4xJYxQu6xPlTLlaqmx+ndyalktMLLO546DDUg6hpwwgbQD
SJWtsbxBuCvOp5qOI7T1mY8zoFXYxQm7RSMqRjj/5ggvIlHGw47H/Msz5pbOsAkwVi0nQQCEJg8a
J+8Jb5ta7PBzTymkF2jZKrkUTChmQukNgGq2v6X+Bd0ixnjjHjlB/9NmDrA2/4qDDfsMct1GbXrQ
EdJKmrJPZMMpDyBhm2SIcnM6dbDIgEOwxG2zyyHOEu73tgfF1Y4NIX682KcNHrScxIOzdEY9Snya
F7wfI7QjBb+vZWh/3cmzH2S8XlbjYRo4x7hp9aVHqQRvVOAyWMYY1n8xFM1l/SJej2aQJi71o2FP
pe7h/vX72C8Evu2zN9TdiculQ3Vesg8mT0P5o2O+vNSbfh9sgkl2VbM7/cfdJE7DFyes1CpCe6Jt
ha05N8Y6SR7ryRvQWs1KFyp57KZUYot0DFa3u4NPyhtQhi5WNN987c1guZvbRoIfrzr6bH8I2jmt
PPm5lI3iqbctsAXvwwm4SX90zb5G/pCT/mUHQcZ7mxdeFuGvcGUta+P5d1bswRTS6QDm4gMHYvaD
QAspOFbl0Vhv6Sy2X9sQewi9lxST0fdEZTg0mdeBBeJ4VFU9KzCBkD+CzMKQZLj8k3prOXviNJ2G
mb81Wkqlqz6fzpRGgSlBiNf/JxNcUrUaKNQLnWmik4aXg7EilHOXn8gjsAWatZ8zocK6IySWYsMA
jgRXumqB8hXcXQfcKtwO/UxQ6VlWCL4HBqQyyPwZXjr/V5VfsweAVNdOvqJj4QZuzHy1skVxgIhh
S8Q2y5r19tCiO9CXlazc7r0T40lBznm19Imr6DKsdKoV0ApdTgIhu5+NfDcsvHlkwTjjOwpBEGsW
jpblf0aVZHuGkZispW12S1OEk6MeH0X9GP+YNpm8vuLJepPIXgjyLUbmkXVspX/bJuSKy/8vwdEU
77EUCH8PhvNgqydV2txlCPDuTjBXVNCwsL1i5Q4ELMdRQWdEUxEbBQGm3wlpHJnjDCfdCchka854
kXvr3WC/R6fPwApFO7xcZbhzvTIKe7uYqENqGqjdORpo8BHnOERXQ5NQyLMNYyaXmV47NKDWIFYL
efSxO75Jbo1NrL8DeTacMXtfhtw9FyiGS25k1kb2UzFunI0vfg1obr+5CfnHsDiIHxQjIrZa+3Nw
6OXP/yEc/6PBq4BnW7NMBNkK0svajjmu923+UsfIF9eTFU6FkMmVr9ybzO4rSQI2RdV9OxXFBtfF
AJsWXcUiuQQgr4ROhfACiFgV7dnwCwDDaOqKJXWEO0dIIYTFPUD38uB2YNYFdQwzn1Sp05E/LrBH
9QimpcHrx2UCoXNB/7TqZGr5sP2OgfXluJ4JA7Rp/rPkdSHbS29JlQjGymuXd5JYlU6gEl709ryw
BswVXCObW97lHa3PjV9AoB4CuJafAc4PziDQ78GEfAhYGKmot9Ge3XXfOXkLfW7Pb/H4Up1rVFYy
MGLdSRy+iZYw0RitNUMF3Nro3GG5KQCXneP93/0QKxh6t3OxS8yW1mcL7P0NoQ5nRPJ7bYUf51LY
SxYfwZFHZKyDougCC3+5CDwVHgO5FYEx0lN4QlnGSzjey+XaJZlgLLt0f02GZnuUMVnYwd8A5COa
vP7ck6aTJAISVLFHMzfFbt5mzyqctcyoSsXn9sFvJTuObuIImwSHeGjKb6/gKQxef/TiIsK7QA5u
2a+UqqFzqqPURsO7DxysU4gKnMkcQPmFPSwupu+hvYXeWc2+lNo1cKNI/C3nSDrlcAh3ynTots83
SEO96rV895/PzV7Jsz+64N4yNhBc6LNF2qe/asLf8tEeHd5MLg7V0yg+pRO1Altqk1bZKAF1T85X
NKKsRTzChAKqVzcZ7Ph/a7JO7IFmFBwqi8AzxOT/fUn7nVDYOTMLRqnFpBh2u5q3e7Tq6hagRy4I
UlliU2PqlVNfTt8ZrEtWA4/Tn+9X+EmksEFoOzASSeM7O6pAWbbM8K0yV2MLI5rCI1TQ9T1xlP49
EhfJNAMa+sNzdSZqLPvBXqXz/oNucTTWwF5wZtJ8MNnTB8ZqnDgOFIE5+hdqTbXJ2vyt8fSQbiNQ
oog1VFqYT13/LwAa/Ar+6lGXRvyQOqWBM5tnxRK/Ash0pToja55f6+4jjHzwxxagGBTwGef8okv6
R16CbV304dvSe1LuGyA59zvFmSgZ0an+FIUWImmm8KPVdA2Wjgbp1LkTmP52Ho3+8bap4G/wsVXk
FVDPhmLgUUF3lLFWQ+hYlsWTtOWBWmPsWg76V+2JZLBVDz4iA9F14BtdC+G6KN/95L1GWvi4mtgc
dqZZ9Hylqd+202a82OmbFWZ9s9eujeyBQFSI64fnFIzHzJssTCHb4El9I5+v0c3PswNN9dXK1gzs
rWFYKxebgiFmNu86P+2Sx2NyYXxKKCPmle4XIYVSLBD6O34iN6pRSU0BeSzARbO23JaEQLKFd8jv
M7qOTrgU0uzmphSI13dhTohe8aRxySfdFu7jGi9LRYAQzMwVFmNGkHFgplCdQZ61DB5yle3bDa3S
A34z6MIJNmgIjHQS7MQBVtHQVsErcBkBaYQjzs/Zt6uvukfZLucVKDgapFff9SjmEldEMhgMrHcL
HIEsBr5+thWWJQbrhyBk+yVxuFhmOt0rGU2SWtirHljd4JhWRBCvxOx73G4aH+V5tuRCytKBJnUO
DlPy1zjahf97hYd0B9tNlnFIX8vVHrJ1FST6xhxiORIUzMqNNAO9Lcp/reQP3pOiZK8fGLfMWFQa
Jt7GvJGaeavqHKnM0KlGZs8DbGuUS9t+bgum9/P1hii+q3Yfj07FfRrsCvfCN5m4U1HUvaPQPMeA
OWxWcYcYMGw02C+HNBFGC7LrV+UZ6PTa+CRwUp+/bjygtD0oCivtnr5HQrpHu/OxCcKt+OhRIpcz
s8VZGSoX+ARG0IHqHp4yzG7e7ZCzlA+CKcP3XWZkq/EGdksCf+l6NC2k5j9zO+0KjVuNABjZi0Fs
ExlHRqoECe/aFzh3oroAJBYRiRj4AP3G2WAX7XTNFu4H8kXT9U5C9Mp2NNKuUM4dZaP34MKRW7Pz
dkelpEbeaWbRqsLMmWGid091vC190oW2r0wtEicKWjeSJ4okD3Dlk6JrKNz2YAJBEFeGsePo8hvR
TPslhT1PmKGw5y+shKt9AtrjIg1sU5pH9o4cgxF2igWhMT2M9toor+54hLfJJ52NjPva96L6go/5
+lYn0lVRgk+f/mriQNjwUkFNB+j+OR1hsRoZ9hy9KspbdKfZKZ0HJgtpqrPmzUWNYlLqwF2CSJEN
p1bMH1ogY7doc6s16rgJiJW5iagsQxV61HSaYLe60SbnIDq107MYHDE/oVMiuGFM+7PeqEHbpQV3
jgMEQObhScHNzx0gx2qMtv2cJMcytKKyeAMeZlvmthmp09lL9tYaaf3nHffNn380bzpe7Zk6O+r3
LQsFJf48SZbPkwN0DdnSZvmEC8Fmg7S8MI4lvmH6xid/nClwOBlAQHcU6aGyhauyxrGZb5Vc+rMb
Tqbmh2QUNf4/Ia3mq1eCH6WgOMijh/ZcQBeFB0InhozAGEuzo8Td5uzjY0DRrcYnS5ey4AZ98Gyx
gmpeWLX9PqzAOuT7WFDBqTD1AVjCWNzpA+7Ju+wx5Y8Os+lqNqNTwp7lpCuvqZJ6sowxXbHFgOiX
YBc1UNJ62T2A6zqL9Ve5WshLPllPQ9mNDjpTURHdWxithKoTr4KAZRm3dktt5y4WGOY2VjFLe3Am
0NYjQi9SqY9LbSZ8AoET3Z5naKdQzLmtAlGRy9tP7YIUnByZNHMGHTB661H7/+slAcKaChadRfuE
E1bH0JknEj+pU5CIerh1P87d80ZQQtW+JfzED8qvG7+u8iHSWJnj+8qRzsCI0Qo9i0GzwqaSzfEu
eMOYYSiTf9IrKvmF4Y7foZK9JVlcDCSOONfCWwB0Ws1eW8jypHEd1FRBprA6EGa50ZIi/3ymSp6Q
vbx+CEOjt+Sf+ESMM4YSjCk6Pgs6gtUiGE9+TyPSqRe2XW/TKX510z1ysmBszK5EmDIP7qrdMUF7
sPCdsMLXtOWUKypOjLPCk1UNAqy/lUus2CoK0ElcNAbSRwECTr1/yV3+bkxW51vxMlPcFl7MFoGl
sxgoQ9ZCJTBup2NxyaiHbAJtpQJlEWe3vilarv7CkUlkk7EbWztLho7Odzj6OEII++ap+oIpa8rb
c4b+/UPzG1+tuBoX1FWMVi/zI/HdKjI1nW8ZL6m9JEsmCjCUvojT5Hprs3z+YVcZHbyxNaD6X85w
b4c+lsgEu36pCnAaesjgGxj0nEohq6x7hgqVaMjS2acqKitCEbYN9r1q5ef1LrBdOgcUHzdgh9TC
0dr4v3WwviNZV4llG3EJtiUhy/vlN6N6acWchL/caNMgwApfD3QEs71YzGLvZlukIPtnA51S0cez
tfyEMZt7IqkiRJo7212XcsGLw3IZkJZjMsTTrRDIA2DaHxN2VfkThnuQnoW6qtPcxHrNBL07tAKa
FbyIbEkp42XJnR9GZ4vVu6gSMmN0VWAugc4hYicEEE24QPN8AubOOQSSa83rO5hgoTzAphMYR36k
6L0MQ8s58POUz4MJitU7gPYnQyPxHY5aLaTFKJ4tH3ult/bDcq1W074IvpAlDFEz83gaLRf7XeEG
We9OsY1lkr3oBrXBvQ8q8QNIKN6RxRSOaeWoHUs461ivbYOA9YhVIYrkzlUkZKsKsurF53IvGG0X
U11r4LXlfABsK2Zm797PqLwqk49KSVilSEmOTfZ3NL/jcVFlkQV86CzX+A++cd3WijtYH0HjQlBS
tvFF3epkoCXQiD3MakZmkYNE3r+/QzpPKQkoigb98LB+kkp/4vlkP21lPFesp9jnthswkXGyLEYg
KxGCJeUU72NDCEZraGjseQeUR5OcEDNXYfHowrlLLvewMckPbdG179dAAoCWeZAfSEk1wAgJ9Wrk
UZff0paFfNZrRb/IXG0T6puHn6gLFmAvCQH9KU/pjtPEiFFbMr4I9IPvwGQDOJUxHRl0Jgyz2ieY
ILrCOf1IAXsDvFaAulgarUfVRDw8wuD6lF45jgEgsFAJZ1iOYe900GBcAtwix9iEVGMtV5IzcE9n
n4mixmk2XqElapChLFkxuQzQBk86/a387owjjaVBCae7uOlXDpPz4YR1GQ3ksAE6xqbdjG6Z8Oue
vOrH9oI5x3g1R92axbf30bIaIShpK4Qs9S178AtmTF1iKehWWMSYITBgmpoyL9aRRMvzQE/m2a+F
ddxyAb9BE1yZ4FnZsgeqD2fY4TTsLxIEJ7gKCn8MkxO4sG6V8xSvGIubB5fV8eMlHiSNWTyoJTpf
vuah9DfqYOpRSAafBoIVvO0QpNZnlXpxfLrFD+S0JsZecOyrUIaN6QiDKTvkBvAvqIbWkACjKXfr
sIQIitsWO5iyhu/q215BqQ3tV3ggO3Elcg+tZG8CwB4H0ZtPdSTfu1E71z4YlT+AkoYdkEtxGV1W
Qa2yzJYw/nUaXVn9XJLl/ssjEFNHmMsglcSLripeT+Gdeu375Wm/K2bSIg+MVl0Y3iHt0YfBkDF3
Mncf49k7IgzdPHj3W4PR+GYYbqwo/6JVOl6r12ztg/WR8R0ia+lobum8Qzw1sUWpI7GCkYlHMaz3
lnNYFyS57zNXgk2NNWUAVYDs06F7P8LOkcxrx5shiS2zEGSCdlLGgEK4XAtlKnPujm/M6gOH9cSc
B4nopSXvuwaj3fGAfcbpBwflBXauM0Iv/qGLZj12gTj5mPqoyR3nlEbiWRtcn9UbQI4H1IhVBY7j
uKpWBbGKytrrPoaAxHeaosMuFJEqXE2Emj8rBU0w5aZk/jgXQw3n6J8ASKyKL8maEBxu7DitW8qC
JpNffdcP4TBT6OOAcOE3xs8EtCu7h53zoBbAc40EcH+iuI1mmgGUhhhBJYUMMq2MMQz7ZdLNEYLj
fOCGOSWR6ROnUND3EzsqOmYDthoU2carQvv0rHRLzUZZT58ej0sUBberEOcCUuA7zlGmg6kI7XpK
G7WeN1GkFbJSTe+8aTNmQ4UHW3DSZ3U+Hc4+T4bze/ShAu0HB8qLp61UZ9xKestk2zAlJYAsKJ7E
38SS+EedhJPVnBwNc0uX0PL52X0dzT2W/V+DE+NmmONFo7lJAcxoVUtbP+25v4wwqZctTnDhXSeo
G6cp3CHFKqgz+iFzE3CRuIkQdaftGXMu0tiZ1juX9nGSAKeHqX4X6CEb2TQKQ56MdO/Xp9I3zZDk
EWyfZPPwms1K9QS634VRP6yL9/UD1OwluIBZWKYDOz16eW8/KADiedEmYSp8OBEc79Gvo/eZVCMr
bPypPvRRX8fn7BoBsf9hyzCaOfZqN8rGCbMOnsOtbuLJWlvX71N3lyq3jeJLMxHTrnU3LH9I0pm5
eHCdKuJLbzOqtLY30+mwjjpLK3wMdJNRXH2/Q74QjkROxhJKrXD2DdHpTpbdeK+QK5lpe5y0Mh9C
kMLUYHG98A7Gfgb/voO8FQ86Hmx/51sSkIHtNYU3XM7lYelA1iNNZqgshQgbu5qzgDziQmMGXmUu
cegG/DYwFmyUHhJkpLH1Atno/mI4u03zla+ESvmNnwo/tbziTysWc03HQ0oaDGMA2DIJSolBTlIC
VDHxhWDoDoYeIJ+iyQaLg4iDsRT32dDELSJVYS7JgmefRxcztO8at6gzknYGxtX/E4F43rssovIT
S7WVTJeBHYJpeB8QfHd0FyGRf4sYaPW7WwHT1RBK4YQqIlfpPlFO5A1sw439KFOTeO/RhA85TC3x
0GfNAGVrU8rV3+mLwvwdVOlsIGLWYaqV5Yr7z7Yn1T3QgCiXwMh0lFP4f7F9U6cq5MdcD5juyMQr
MlGD+7lKfg6/fHxvWO0vLhaGCriDgZPg/n0KIR+8bOex8gLsiwtqsUOwrZjo0K8sTKiqGWqznNQG
fTBHCxzZbdXvR/8CFpap2XeOQWNPnl9ZYozAPF/aBecGiPN4oTMPvHpExMTA+iLucEBalUKMaub6
NC3tJto08yTSrySpLoM4I2plJhfokflj6hC/hghi4N4aMz/6DQntDj8LuiKTcQ8HtZMRxCgToXAn
TJJ3EIVLwAxx30JTe9kXsFf61xNsTpGL8zzLpd+czdcMP6iYmE4jv0l77WahTuZqMTR2Q3sJ8F9K
merXW4SZnftqcXEPZGpMYLHkxiDG93IeXW0FKkeSEekWDGq4EVGzLnaioMlZTFdKM5ifTGR98LRG
EexJn7oGF9EMPPvDjuUPKF/GOgrAmeNlWwPxh9QsYnDpsRPbl6TI/XkOefl3ONk42luiuBl+rjwP
oZNDGON3n0kkJ+eHzVa/VRILvOjsZoyP9ufOurkW8o1hZp4oXmzNhmKLASbeuE0dnuMb23rCAHdV
Nc4Z0MUyzMgfM4VjP+es+A/ngR1Qdm1FiF2VEP0b6JnmIrS9RVfJqpMiWkN0Lrym3xRYuekhDBKa
CfJnqvzgo/MG4AZWT/MR7BvwPObujU9pjLJ9hRYRQpbAgj7et+yRq1nEKMsJKrjPQhnrdGGF9nlc
l80hSQPtX6UN7a0E4E2WIyZYng73p0q13hfjqW4uQVpcbIBR699S+oPzrDSZlPQHRj7rfmu2o2ix
ehUrQh4b3gCKAM4T9czxGHBsk2XsBcRU6XaVin5PCPy30TYC6mdecwOx6GB0SBot8gnwulwvS+vb
H7AQ+mQ+wUeq362KcJQjJ2jqr03ukGyYac2cvJPqhxolnA9lrqod3B49rTfSnrigFI6uw+elhibN
CVMGtdicPj2cPnaTSVA7Hv3X9lnVdDVfiJKq/NnLLRv07pnZgJKlULf6XgkFqZWbd8M7/MoCQqed
ynpyZWWx0g1ha3JPFDca/r0hHEC1gVOm079VKyVPuA9FjoVT63ybUrOv31iv6LZfChlcRZITh6SU
dfXMulvr2BGbdxqNjVRO2HVzi391Rz+v9AwHJSeWWBEroYeXtOiKMi6tRjOTQcDZTKXmjYC0XwTg
H7V52yW4Q14DfSOj9HU+fdAPifl4eDH/4l6Cl8/dauyA4MzYMpYEakQlRQ4CxgbDApX0ZdWxEIdG
9gAJCoGEAoLoZ+3hkgUNz2lSGeRaCwgpehPtkxBPHpXpZS41ZUw5ayh85vdIRUrLoUpnyDW9vo5A
wL8HorlyL0PCEwmeVUaHymiuaRViENcMbyuUtITkGb/tnx4tr3/q0WkaBZt5CUMfTGfIrtb/SQCB
D+g/mHFaXFgzTpBdIjqiZMpR+3y5sTfEwp/OrA2HXgoFEu9Yt3/XcWJ1mzIraY2rcKrWQNnvY+Pu
9M7KBrm5/oo/ljHtRAOFt1lSTIcWY/+lfQjEXuTBhmzpsM7a4tkl2qOlrl7lyYadBUwUcW2h8/jK
yqREOvUaOucDCj6jZUvVSlJfehYqdDuG+zZgM+zVKn//Y0LsIP1ot+M89xoJgkFoh+zvQxGPDMpl
AF1FnsXUt0vG94BajzbbXrtky+el8nKfTz2ESC9eAXOKiEOiZTdSxcqQbKlW0KnAgQ/pBV1GwvwA
ePd1EHhoJbZZc4ABhlE42oawFXAUO9hjkJnC6ei8GcmTUNAC3uz2w0A1/BmnbY++R8N5Rq1+6JWc
W5Mr2BRe25lZZ8X2gxQxDfH9T8B5xa8iFSqcLYr2JJ/vnLc0GvO2ighZmj9hvqmRhsxGf1lXe73E
Cwbm5cuIEUh69g87rLqdX82+9WCzbY7TAlrVPfGvgar3Lc3tUB3W7IGzcllPIMU20AMv6IQrGSb3
8UYsObRHQy7SLj5mhOBVxqYGC9qab1CZ7FOOUN+oeSnAtj9awuGwCtO9WZmPlnJ4SRE0xDAXWq7D
Ron51Q+KThuLOCYJNkCXjC8WQ4i4mABoP6oilACACr+Sk1z8MhY+R9oR6yq6joWcbpEZAkA+uyjN
4xsO9mPn/dx6U2QBCvGKgvCMzjyzNUgf3vB79Qy4herSoOT3kcPHXtBCpmp6Jy5DfQ0bQW9DOTZx
EPiiyzgWDR1Zrrmj/I6WEKarCzf/xNROYGIW1mZ0W4PXeM0tuBGFCVEsvUma7NRGqFmLNCAdAePE
hK9wSOMxMBE1GFOkEN00B4ztNgZojxoLowZJz70eXfvhNAf9KQSA7HfnRskgmaEuq2Q6w1/oTGBQ
czoyCCSkklnICt8EnXxPC+lzHMl1M8EjVRQxxFeZMtP2B8KpfpE3qp//69fgBF/flcze+YAeS2rp
ky/2LoGwbHfy1FBstWSmEwhcSW201akikqNBBfygYsV8Xx7ZyA2LLNv5AA3h94PO127c4muiwHUc
7tfF8io5v8p7aRzBMotin5psmgMMOhUI4DC/iM3Ytxyi/JWSHdWH5R+ERLeyygSJ93rYlSyatO3U
LTZg64K9NScWltYmUNQ7V28ucqDkmn10BgO80jr35AvU4rXXcDmVD+uSoe5925ctINc14+zUR6mf
N+NjIdy0tc1FCEhldFcz+cHi51IxJSQxKJKQ5/D+to9M+REjy35PzlEfy00DqWhQMwUVqVtK7fPu
vaEAFATM/7t0O+bc7Gg5qCU22S2NhHF9odHig8tUne3iN8TLDJCMYK0zaF3ckKPLBklYhzNXE9e8
RbeJUm2524sQzeidpRjKccwgP0krPRnlY3X6+cVk/qaE4g8J79ujsckvmz5QRskKD9tzeK7qB1ML
xEmFQbbyABxnrXbELqXBrBi51Metj3yNlv7c0obwo2F2w4UGTIiJftEHv/DZWBXw2zzm6D9U0efZ
UWoGlQdeVhnDBwvSDAzoJ79yHN1HAy2lDMG5qn9xDxY1cQsaG9qsgSpWjBOEuYwTs9OPEn1QuBXI
qdP3rIsh2KWIC5mt56S8DP6oY5WMqTDsuQmrDFWhkz0Z1hPQWuqz2gCccRL1BEw80ZSTktRKVvy4
aEHwbI5LVcQUbpL9NHfBBVaN3HuvOfUR9MFX3/525CApK0+1t3CZBXKouFyz78xiHZfqzSdHXXf5
bILVdBFmhPeQdAVBjvtrEzTMvvNk+DEjfT2PjqNFR2mGWEP28rXFZ0FK7O0l3MlRzBjlxiqsOxN8
uBHzzajarX/wAexF2QOKhZjDx4T2CesRUFewX8dP9C2MtSiWfoxdMTnRHEJ3fEFb0XoMjJww0qkM
6/kP1D5Nd+JGZQ9/SoNk1rL/DpOIqFWv9yhtKwMMsgm+wJF3EnOz2hE5fHXRjl8ISwbHhDBr73s/
NBkOPWw8lL8JVTyZbT6Z2xUFsZfl+5kAmeTtRUbF4OxLyvVQTc6yunb19UmVUKJwDGc444NMxCZr
X1wq9Jx+bdjUjBeyZXgKWmUzbzl8Z3oBt1zt+t8sEB6uvN9VcgxAiaqO4dwWBQhzSFvfYxGE9sST
Rk0w9xZfOBOXCCKX8bdsRkLZl6nZhABM3Lc2KlOsBA0JlAMI4s9HAZQsinqngkCSq2FHLb9GhssX
GgcwPDU0yOzF02yoAoWs+6au7JOu/lrGbAVIKH/hZPUZY28DWoMZoRpGo9HZQ8XfhHqv48iWTfyg
d2FzOf1wo346PPZDDZ+lXTC7EB7sLQMr6EPPOL5lUV1AwnmW1YiQL4hvq8EnTUuaUmIb0PddTENt
1dGIF9pNmuEjpo9eDcILtS5rZUPNUv8M5xXHl7my8hPnYxsvhLodC1t0krUnQGDDPUZieqlKQxNC
mCQArFWSvRY/lMf1yEEQbBq1eXI7OFZDcH30HQrc9GT8zj3MWyp14Ue+1t7TQDIoXdqw5EfT18A7
upp87CfCNrD9hiZwgjsXOrvXkezUVXFydYIhDNWEqofO1j0UTBQhZHkNEee7fhO/J7iH8kh7TimC
W6hMmvtBRvM1Ltvcma9HEQW9OUk5bl8Mt8LTdI4r0cCk0gGexe9JzRrAQ6NZz7T0wLp7a0UOsAIM
AzIH1++nEXxSYw0KFI04QIaMyWb84Gwp5+tWzK1+6xKz7MDmP+8CFyc7///lKMdlINuwbeVns5tW
ovYrPs3GdrGZz0wRxSRerkcUr2Q1+TJvd9ALCDkdeWCCumB6A9Re95py6Tpfb8QeCuT4TOEDTKAO
qpON0++7WlN4b44VbKj5aCJ5dN7AecCRptIWLGGEbwlSp8RpP0MjLnkIq4m510dxgipABpJ4nnfj
rUKil7dSjxe1eq+NVaw3kOG/3CLUDwMVZvMVPOsjYrgTrQzYPScNifb9SLrnJ8c4zuaAkNdPsIe5
YML9EeCC9b6SU6VNbp2t0DXL5Jas6rOFIgmS8/pjeXfkClcEBWbrUI1pMsayuCDnD/8h5m/qINFH
2qDiMRPsYGQACfqR8ueo1G3ocwiDmHMuHJ1bv9fkYr6Zp42GbJWuthVWZxqdFoRWSOtv8jVIwBS5
iXdicR+rFNHQyvwDn75grcYO6cSUsxCEoNYGP9gZRMZdY7thZOt3utqJTPot1khTsxvbwrg3jCb6
omBPWaSO96sTrLr38lxidcKLsQzELCDM6c7e5yyM65XMfYNVwmGPNjKXp0YGi4AKB+LkcVwDNPUB
Ll3lpuh9RBMQnuUXNNTcdmYCe/4tH4aLetux5D5oaz2iPhA2t0G6TwJE0GfjtQs/hBtBkRBYzmca
+sUIdpgh1tcCNjzVF2MOlj/r41CeYJD0s5C6VdT4m9UZ7THZLkE2aVqXULzXQnEM1UtgJLySOSTM
nLw2QOlIF6Xa0V+RwsV+rl2XKz7hx0T54oceTuHTNE1dPAc+QkhtfpzXaWL5yNFjtaFHqTd6Q1d7
ih/QSV2V+/w1Oe5Hiv2VWJwRKDHos5OrRxCYSASw0ISWY25JuuokA0i8tYYvl2l9iGN/2+VGnH3G
dPkXW8qXR+7dSuaY2Aa9D8WYFGZhBZLi1Kiez+NTf4QklIrgJ0LKR+O4oGcYpFi+8sgl7MLQePHd
ygy442Wu6bFcV+/8V+WdzosVMT5mtGHT9+cb8Dw/QKWq/f6WmIlIGb8X73NRhLxdBr1Wfin0ZqXI
eCpWjEQabXCG4eX36KdgGkzhmvFTeo/PJIkfEYEBNwDNaUpo5F1avrLXJfxbOV9JvvPcr7RBUKy8
QhABJc2s7+OOQ4nqedRRibBrSvPuXp16lhjmFDlAgHPxKvArwximA9F+fkbOwOK/NFsHQNBtBKMU
I3Z7K0284DS4xcChGDkGQtZc4sWup1NIq9VFHEgVjon4XgBab/MDo4oQyKW3td6ytf0D9OAXh/UN
ciCjO72J5KA8UH7nAYjNveN5c5sVuS7NvMx7kGyQoj7bclxhY5RmsspbmVx6THZZ7un16YbX13lp
pov0MJ5EolDhqqPp59tQsuVBJe81noLAneOy2uyujb3JGtWV94UOLkRd1xdKMH2kJacLSL/VqiKH
IEMr8EAy6QcRAPHwDICl/FYG9RQW4qQm0vcGWkMDYEMUoiRNlrfyOF45Oa8bbkSCTC+KYPge7UBS
nvSTNeUyIVqR2yfI41wtcyV8l7m9HFE2zE2NvZYsY57S9l1Lg6tS74vsiUClzIYwVVwXMS6ZTKxK
SyAKlOMJci8mmXEkwysvOBT990sggaq/CCbpXAFN2FhEYfv3uDOQ3ImrBsyy1HsPxHsW9WmmkHYA
tCsrmkHAUm4VV+hslh0pW8xPOgJWizbnULcxmE7fZ5f6Gp1Pxx5iIKEvJ+hMDKPNgGUaebIDcZOF
JhCi4Vm9Pvuw7+VpnjGhtMt0aMa2mCH0FvfuAwy1BuCjj0SdvYcz/Zsg2j1Y965GHwfryb4XUU7z
HUv33e5aF2yxFFbMfWXbyNrCfUWNK/PEZ5bYlsEXoB6ZOHLy/O0tDvxf9uzbayjTRtR23Py3OQaI
KxVMvdR482HFasbbUQQ6aroNtWmI6LY8PGrmFqldI+uIs8FPAG/l3rTZAQzRnroRgWA/TOCzGuuq
OY2AWAe0M4f/m1R8L50lVoY4fcGp1gysn5S8b52G+pqecfCtqn8v0Zpc/GlThDf1n37MpJV/q7GV
9z/T0bcVzlgI6mLZi4rJq3RQyG6+VzN+pOUfQuWyHpKEzIApAnAjrzLUZSYFXUAbp3Ga3hIRtRoI
wD6O8BX92jXJzub6OM8kJBJiGCRWxlMpG4u2t+sp/D2zgt6GZSGFHEm5pkCuLqEqGtGsZP0QFxHb
e1TFMdVSvYJ22WeJpxjogVHqk+0zvn7lOWmaAHfjb2QgqijRT1wLBqc6zS9+FdU2a1cyZ+eoqF25
ycgiq702udHheomoYaHRrjmaxfEL2g38i0X/lwiKQXGdHAl5AE2rMYuiVlWbPnLQAktYL0HwtSwR
CtUA1S1Nx4qYof1ieCx+VrIWXi89PQamNqtHCMVQUrIe91lclHI50SiWgNxsZgcBG6BQhnAz59BD
2fMQl844rPvxFfi23LZJaylVOw2/ER+oTgDV5z/tYCwfv6TDozJrEsSMGiA6UfreZ2gqH2mKrUad
gXbDOm2lEswTQa9fqD2jKcQClHE7MsV0OYoVEwpqrSL5jrZTx7ffY/8xu6RPBqcprRIPdYoWq5NM
0mm9VA2CWLGMH5g1u6s49X58a2y4Uc9yhgS8fHlP7ZB3Z9P5dJZcMybJv6UlWYlVFXWjB1+zFQL2
tvQw6h0Rf8aq0PFT1V8wKdRw3XXJgNOWRoD8rIcSEFM60/veGtPVy9l+BfhKvIVgmU4tSX09eYXu
I5NyU7TC1+BMop4T4ySB1cWraijK8VvZuIDpBy35XGI+IYBLb/ledXG83d5H8g+v0ZT0OwIzd5w2
mM5Y9TAWV5hBIzYYu3I5vv2q2Tv08j/gCBEawbXBt0+D6Z5GAv26Q+cXvoKixQUklmqLB4jT2vG5
5zC5Gj1pbzYNgJIqouYM4vpCAKnCO4+lVTZr8PGfB6zK7POsTJpxtH3oqrri1tbSIxBPhdxla/nG
W7xPCu9ZQNXeXmdS42ZD2ztX6e9+S7N0c4eTB5YEY3j2xz7qhcpELDGMNwRxCxrGzTsSXKVHawW7
ZOQHkLIQdMh6X8O5/LT8KX6nhpw6QpuNec6WTIx0L6ZCy2Qu7IFehLg4fup+pqw5aP4VioPVdkIG
yuQXOZ//o5wMUjB3jDy4mtyN7EGNoGMU1KBpAhprGV/KzaTwZseKFscUyXEnKQjqtY35j2yUX/5N
3Y3klEc6clAxVSLqv1E2pJ+1mjDidJidfpF3XBuI2wkyVQtC82eWvIdI0gzrlzbvYKpEqpidiY0D
etDg8PqmN8ZP6Z8q18pl10Z/hxuzRczrpiRl1abcDdgXZVUWYdqPc0oiybjX0KDsr8rn5brKYDOc
bnEtWgJuAa2i0RiQqRAHsANrvGaTNPmP8qRi7rj5hh9zGbE7C2UozZlW1jpzjn1VzU9+8Ktv/PP+
3D/grCsvfDoRiomhjlqx9rAjIPRFGPg2/lJ5yw8kHLfoBpp+5nnVb339MsQJgp1TaWvFA+ecac7u
FiaaikVsw/CfWTvocJ8C/6NZZjdCyRsVr74+ZH2ttwOSo122BNQmTEvvxIGyRSac1FZb95Uj/QmS
jSK1HBhPmpq474GpRmVzsE+hQKt5Ce2F/N5pFdGgju5C7cofBeNPlPFN9dqlz+haYC4qFKe/jl/Y
l0YcKc/YW+sXEyzfuRYusCp/S4sy4uM5fjOoxU6i/6FucOS8aDN72JRsGH6oilv3iRr0cD823UE0
pHJBurlEyHBgp5bGqMGY9FEqKLaG00RzA6kk6zvXd2pvbjbTYznoMjErR+O4+LW8MIS5YYTN13Dd
Qjh82MGFFJ0cRcj7ZpCDj9oYnm30/xylrq7GuNGHFSUBpr5UQZOZ+ol4AFkiYqol+qxYxWvid+6n
skgsdSFBR3lUxr+SZ/AbjF5HKfdz5/Opqm9uP8xZ2bUnzBhxDizwBoZ3BT0FVMO6unjsaj9qVakJ
/rtsKlUVnYD3e+/EICOInxT5asWJqOsaTZ2iUldlwhpd5GgiLB4Nm9c1jYKEFaUkLHUBp9Ni0dZ2
aFDOpMBDSWS1m0KgjuInasVwnNA7yssoyookYMF3h5xmZqA76UTI6yGwcSIGZjRl7WsotHSnpI9u
4u2mPElVhX42iRAR/Nu+3x86nG4OCNqc/cxtjyOhnbAhvIviXeHa6wB5xqhIwLAXWsW8Hw1yLGyL
+IOaWt+KYglpApIDlnjVIKqubq/SiaU02p7+Iza153ekYHAHScZTSxzrBJRq75Amirz74PViR1KA
PJ96NtnoSc+fepbRNWeZCgHeCk/Dr0FYH1LwtVvjsewSgxH/vESOsL6V4GChFyCVegNva5mmW9mk
G8cX6Oo8K+kdE9ih3UnI+/OtqRBNgUsntYjQprkowS/ybottSmmH/g3q/Hxnw7VddWNmno2kdIdc
TonAzmoSnE9UObsh0dk286ep6a6jiixfIg1mk1hQxCVo3Y6le2AK/nJDch8b+1CQFfsy7KNc2pZU
P10V/m950LghOTSZ2WWB6lmw9CGmkjFRiCS5fWYUdSbH3veBNec8nG3DF1rX/EEO8n1EA7BMDzXw
e7MYcNp0U5qaLnwHlXc6wDPXB6NHMPcKvzg9Z8uQkMrrC/PdREdWKf5yWbL5B23+jL/L5QkVKIAo
zv/hAN8EkHGcPdUYzzswLosNVVYlzlrdqJTkfok29d1ol8iyB4hW2qqlEK70lOvmPIO9IIzBDIWT
YYdH/TsOj6BKPwdxPX3l9zwAoO0h/+VYWXEM1aQbl6vHpK7Dx3n4NglBqkeHk4tradm0Oeg6U0Q2
epPmZusZQqfkZcCvvVAh1tyEh7wFfkgh6Y/B/5i0afXaV1/hTi79Lwg7M178I0I/bJm0o9us2EvR
pFeGvVcue7mXfSq7ngleZ3uhhoxfqh4rSuBbhBiBiTeveaaFzi7O1j0CsONQGSfGqVYZoxR+x2zU
pisigbjp/HXckpZ5itleJq3tvPx67OCqXLyWJfvUHwreScr3BdwwR9PZMNDHs3ylgTe1sG8qY53B
BWULVdR9ehGQkvvZgcuRbB0r3uQV/xjDS0+aAfL30hug9rBwfhy6qPvSshOaPOFneQbMJjqzvG1K
+2q+sBEC/XCLVjxDR9Jfx6tJ3y8ZZW1pyBmwY4ki0XaGUXCJZ9yksK5dIX04EWmGhMnR8xKoJD/o
hQsgC/XKPp4Iv54MaS/G1HQMpLEmoqgXFvDC5rsUC4gPlsOyR1FFC7vEW+y4tbsoEMYr8pUrjYfI
lV4K1wy2h1vbyt2jitD6hdHWN1bKZmtSaRuuoIylqB4twwmGtfi4kpufaCK/9JBi2FW7PUemFVPe
5SeEtquI7wc/sMbpxY5vxliYp4MzgF0DWP+XsaddXjJvzXRxzYbdQyrbH6u+578mOFAEib97lLuY
4U2PfWOfWgcVfK6WA+I25EnZU4M3j7cJKyEhg6aDyfmYCPI00Jc7eVQS4GQHnJ22PIIZHne49Ii0
V8wXyKomGaufwERp5+jmc7WEsg8HnOJq2Gj04Yzo/h+Ys/E5SSrHx9IJ09Tr3Wv69MjQhX+xEQam
ELepp6rddLNEnmuV0V5lkZLYoI9Cx2B2SgM+0/xE35o9rJR8gsQDNqvlJkR2Br61NDY+uVv7Velu
BRSi6BKJESaQeIWTCBB3KbTAn79c2dcv3MyPsTxItToSbCEe3eGWDeQjFgg+fkamIywRfbx76E8A
RVel38ztvzR/CPbO0DX6MOrE53NbtG5kF/Bl1oT8xwUpwzYDot4/MDnaN4t7LVGyIBNyeMaW7wlb
qV099b4kg8q37oCuDTVwC6Ye37vyiQAOtTVBfwvXM9xuQzZq47SSk9DjeacsuLmATjCtMuzJseJb
PxWhcQVUab/aJdrnioEgrmghFk830AmQauMEz6tv/rwmiEhSVEWukkxKvdJmeLVEJS66qPDopgbr
vtkHw8WrsFzkRttvJpcGF3USqrf1JsQ3zzCq/DdjOvJ04R5e1K9hhKVBXfQ2i2EVNJUSMH4yq9kR
74q49zrp567h1maSn0Frha7k/73iWqCDbaAp1DPo8GNzR+1cLqyGWnrnEV3zNHEbyUZoJBF66/LW
27U2vTUvRcbDJfpyzyhWL6O6SWG0agNW5lS+zEAtpxtl8NmNBqHgEZnlHnT78/VzKQurOfL7ynFe
PWJ3iBuCdZUFNSAUyp55UGxQsxMTSadFS/e917jn1GvtBvBwq/AzhICVBw6kCl1GEcaaeFKqTsHm
UetY0ufIaktZbkpbp7W5On6lGEaYkJreTzyfk/w8OKWy6ZqmHBGgtRBiQiQa2txOVzSRadZwpMQZ
sG2D0tUz8TSJm7DLH5v4r+y4Z88ysVgX4CsEJzIXUymzQMQRPOFAsQ684nNuNowoSvaLgts4N3H3
+vFp70MLU8Y4DEQJOCDfq3/yn4GPRveDG8rxeRjQ4IRCYVygF0sDpflT3CyV+8hKnNDpwCqh0G7+
0Lwe+W9gMsDXB/J1tBOES30zJAbRdkxqP1wfr2oQ5pdhsmgsT1d8AKuZdU52mex4M8jdBLNX10o/
JzUfJIibgJ8NE68fplmOAT7rvaXhqI/88cu6WcYRIR+fLP0SPuZCg7g2JHt0b2a16u+z5wgcijci
3HdGyOGxefIDYs9zba96sk2UqcfoZLCRSqzLSrtrODd7jAdLwHmcWBQ0f6dot/rn+Zb/SvolKSNf
2dys6/0MxKAPS5NrzFJAdo4jrxsTeuNlWWsfCtU3omrEHuyik6i/KTS3lNOLtcNDt2pjTbpnFjFu
+VqN1aYtrU+RwGwXh7piwOGEsAqcg8V2jOtIceo93WtJXKnsNHP+Ca5gZ5Gu4/BJq/nTpWwZIXrI
RAX16Vx/tW7+PRd01weXHzHQpUA2H35AOGqi8piUTgZZ3iuP/DeX6KH6wzyl8OReHCkxY4X9cGxD
3iC2aU6n+et+Hdshws8uhPLgvbHBIkitPqOv/nKqxAFocfmnLtHPDZST9UV9XJls4zfCnY+ua6GV
FMKzT4hStpvl5n72+OhhEuel5gc3T3KdSvUmq8KaqbwhIOi+zvwfzJYoxdxMyjRFLDYpdMEtmwvP
FMvRcBF0af6akz1VzJD3lw4ns3r2wlBKsZ/5qLKM3Wh4BJRSmz4WlpKNo2yLk7/g56S1w2f/Mrs1
P/6V5U8AjcbVnv3ybENlmqMloUA11azjW9vRo1XFbWX6mDfgU8UGkS7l8JEkfadh1VLTopnSZeRy
4vN2J4wWyyhftVEq82v+dmkhm31nx8PiSG0f0eU4sNFEZtmGD0Dj2Cm1YGvDoXwOkYW36haBmd1Z
FPlj65v394CUL+7QnXDr1lWQrLHovtts2X678ULVTSONTL8wAAmlcFnIFWpN4gtJGPulEfZAc1eJ
arLXQ87+vc/22lZYO/ug6j+eoGih5yjzKLv2fxSw4Feg5LM2+uHTcHwK6N7DnrdSiQjY5n4t6VO5
Z3XYpWJpHeZYXwJdB1/wM7WrQNwLrXaLCOp8DklMSsA53LIKapDfN7mhoNJ8cHVhmmGDLigzhB+A
IVHk1Ne4gMZww3i3PdXp0sANPiNiKAIsOoseU3DkKctCWhbxujIzzbIdKNgsiLa9FAgAPFA6nIdl
UmDmtokFiDot2xoJxUrpOuaRnljMNcbWZO5/4XdcVircBvlIzmLLMfWixFiJBmyNtqN78pyXqZ2S
clFtnQ+NfT16Rlw6TKg27F9zP++fzW0PuBFNH9PkqefE0NQkbfjEQzKC5+/ZjAeCFNYERiYdmry7
58D2y1+aNIjzWepCGRKldfgM9fDgabYCFn24NuYYPOlsQ/ggZhuhE8sA5lLScBH/BJ14mb+4gb9Y
tTFTbgdW0VRPCrrdOm+1RHML1es+qXuD05v64Jfb1o3cq+RXjfdM19IrpTdO71Re3bkp9SBfmLK3
epT7eb35qPKtlKUhgmC1qw9H6Y6Gmnxpw66B8mDJMfEclmxPQupjpstSVcnaPsApzw6zR5ejeLHE
AZZ+DL+2hN2iohUTD2p+v0rIU/Zg/2R3dDEhc8H6C4vHausGXj0XjMIO6WwrIG5CGPYfyNCkqUza
a9CbO6tY5grufIfGdCTzCMKieY3P2UmqL4Cq5TqbPNZBbga7tinkPobhRU05hHFhJufEn8FDba2I
lHARKULUXdMsIyjiZ63/ex+jp5Q005H68GblDAFhX1opXTcZBafLuP5UOUBWFthfRz/YYXj5yDAr
z9ZCN5FvCiLrTyzvHfcX2WfmCYm8CiIhGFihuuSe1ME3voZPeYZHKrvMS3eRMueordVJxhlVSZOE
qU5Y9bJaD9F6g9LXWwbNjKNikT5B/f0EnNSbPfaVfYTlxhC+sMKkm1EyerUtSw57Ui9id1PV1nEY
dSeJFwoGDmttVPQfupSq+og9QwoGs0xw91lqbBQXSjPZQbS070O1XhOHyd7g29UdeINL/f4U5Kyg
mj7rAQNhLmhGSN+K9YYc3fbjNGRAnyqYZd3aSQ5rXXkfI7a1N71qNtu87+r352EzdGqk9B2h1hFW
rUoeR5KBfty7wMduUPeynbpKlRUGnTnjz+xL+YJ0RUgxn+lfYtwswXZ6WFydNnt/QNlPwYhdZmso
syde0gi9DbvefIWUzepIRx5610GQzs13um5pHKhQIRWeSjl0zDcFlm98GDxUbim0BbHprByWEGOv
rz8dkZ7yfzI9cgmbsiXRROsUKcu5x/oWQiM+61SCY0OlgvfVU5xlwCzH4keVoVosMYb6qfqqmjSO
/XT3LoFmi/itKmchG8t5WLurOmrpSCJVlFk0odEz60RyM231yID0gdI9t6peJcEzVPrWHkR3/ogS
zgbwIQV63LuN0v+7WSTV09cABd/hE+AIZjzmOyY8Izn6SIO5mQbzXaD+qMnLU/ZfcWKP9ju1Wkww
Vrs9gSERF+g+GHs6/nxwYq+t0h/CBu1L9AaIVUZFh86DodgksE1JQOA5obqT+S7djphwLFsNHzud
p/nJGMhR9lS/eZ9NGgbhXhLS4dYuMXKCNGS022OdTFhjPWrRBS8rAGw+/B34YsIwCJXidwJXYWbm
8m8Vs7SHthLcR3iUOLH8v4aqdpwli+eOhFQi/VAqVq87pxAsw9WvcSqcMFN+l5XB7s9pcblYEghr
CY1PizrOofHkmYKlx6A6sEuYOBOQH0fJEVgUIObtvmCm7kkSLFlC4Ej9wXPxL9tyYSalKsYg0Lrr
372/6gVjhRI7zd0rpHfGa5tj0RGHvCI87eLnXpGSve7GVcSqpdtg5xH5SO7pVdbWM2IV7cpq1kov
wPAC4z/LNGPgCcU1N2C3JCOfcXYC471MHdhzlpC5U/9bcW5XTT2fADdAsWTu4aqiYhpfCtRKVKCE
343WOuk4ppiHIRptTZNshmld1slthevtzkBFIQd4pwN/WraC+b0yJQM1TnoUx2QOiMkvshawPjib
YmPOx8wUqcIkBSM1RYTgIHKmewuhowCBKkHsbnW49bJ7Fbxcl+EmUVVSvfRl+fLoLpuzqQCEm9UF
QyCMlUbxj6rjK+xp4lPo9QNSlJ2J93NLwAUMA1h9IrV8xC0bTRCfJWJ8EMsyu+hmDiKI6z9fXmYU
/3KTbpg/ZxGGVWVbo4KS1gjuNKVH7YiwM39PTYyeHmqbPB07KhyT9ECqnaM8oNUPW4s6CntD8A/g
5x4Zw0mKz6HW/ixPzHyWdFyoUnKZUCu0V6hsWZXScurdjr1Sjn7sQr1LHUccFaQx3dGeMqliVdzh
p94qw6BZF0zH5zFnWcp4Hy6iR5II1vBg4Zgf7LrXWnRucOlo7w0NtB1FTjcpyK2AeWprUQtQjGfU
XwOTIXhH2a6DsJNva2V/OZJhDT/sT/uDHQP/nrKtoHAaaq2vgCss/LAshlZisqQZILa2pnB9GhNy
6c5vjExuaE+Qn/PkEVo/r7q5zAwe04pqvz7XcgST9hTr3i9bSwYFcsnaHx5V8FHNYzV5QxuV1+7Y
LbbkoDpNUGnxnTsOmzDhXSOpL+yFSZgf2zmGoa7BCXA/gf1WT6WczGn/q8EuIRN3lkeWfNPmYOuU
RRTFLQxVS26PcirtoTjKRo8G1zOcANZdGjRamI9vz8weGkGFRkCyN68GTUoxIetJGNyJyDvCAQ3R
wUztDCkBtDwHsJ7PWF/Rhp1scGEu68AiwNoBirFCFNrG2xASmyfL08S4I1SD1wyIGD7euIjZz2m2
61cmmS8q7SvBbzgmjjCTWqpZjwXeVsRl8cmf1vGgCxIMSsxgFexs0tQlLBPY+lXmySCXADVwUJzA
cIw6HquaKial/c7IiNSVsMoRbj1ZVBh1Oe86TpkLyRl/chJSJgFBMijFsvoVLtFBic2ja9UucYDH
SwuL6Rh4akwq0GzNr3daRCy9cNd5uLLb+rAgeOS10fd+Bi1oJSmUAo5givSy9FZAKlMSyRD5RJZy
FiqPlVnyKfV4fyLTnYs0ip6TNik5i/I7rm1dy1kNtv/KMFArt4vRpBnOQnUvtUnUyS8sH1jfP0A2
8QQiJs+QIGmFItiu+e+Vb+4oEbyIuQEBeWUjPFlUeHHR/TaVw3niAd5NwqkBMbflVVOvCq3LuCI0
WpyUXbV0Obajg78aGdW9yp9a0CukxPIfSTptgTF/y+KPSOIBRBLsGBk+RFm4PVnIyy6qWVKlVIBS
olbnHJbrRDotGBimWtxW0GWoJIxeNYGfVA7/OAJwL7lAcOpc7mNHWxyo0+tSvpoa+OH8WTRBYcgw
2F/Fe08MNH4Y0GcCQ97wRqs8ZH45ipJylu4vYwe0mF50/RvUMZEvgyoCFBfDsyq1ANHxntBCeX7I
JcgGaGVAO6+og5o8WLelTHoz8UaTwIxS+LxXRXgt8O6Pk14tIIQ9gc2znUndpV//5LKoGXUh3E+G
c6bb9khGakuMOrxoTU7Cqi8nMUEVc2aAmmL/im4yyNUpPnPMurKINwqOMlDWaIDJvCR71Q6eSJc+
pJi9GHGyiPuXKVDxYiNQh/DYkFmKUDa6GjIsUVU4DcjDC89RpfiMbTzvjIFpK2sD7YphgjWH2Msw
QIaZUt/LUyY/iT97QhEmxhccRzrQ8CNWW8y7KjgMvZw1m1PDnkOBQ8hPTrCk97l18tIhjMdzhQ9H
+8FlqVe+RgoPBfrb+y2Hty0MlBE/k8TBYSpAQ74ZNQpTklCWcu4yisPTUQXOftknaNMO8WD3cYNb
nXafxPo7i6IbBFYLDI1DjjrQ204yPeMXfPmIY18lFTQzahtNx0Y4LTirBoDuRd5oBEmWZurLLTeE
5yy4uWh39PaQGZuJlVoF/ZDhCosl9ZvA6thQ09JWxG+6EUYktak0wkj8CfvrBTtLqx7iavT4V5jR
jQq2wz0qGbRAKUnwXEkHW3eYb9Vqm985VvBrcAI1eXg+RZzj9zsVDz0vObSF3k8ZV0ro6Veqdpv4
0hukpKcN6K0N0FEBnVN6AHKIOh0zneRHgQc4VN7r/5vInNmeEo8X7Gnyp09JXdjfI0ZdeDjeUh40
DLJ+PrB0lwv+qH3IAXc0lpoRyzTOTYEzVk67HSlsjUeihIGxGKnH1IP4LoBJ3pI96JY3/27ODUPJ
FTKMiE/YUazEwdzpwwVYAxNjffzKxFLV0660iS4yLyMWgaE9FW4d2cMjWMqAcV/ebMoZBQSy2dTQ
PpD2HrZ0glPyGD7rDd7AooncNsaS3eClb6DvQ/KTLDhpA3YBYwushBqgAx0rfZWgA8bSKTTvHqFd
Mg94iEdDo1rtWObP6V8H1zxJpTRbvJqfVZPZzvzsUxhgei1sAfwXWrigeRuhGChXNtKJEs+wMumA
SJUuJhRlZFpsDCEBAZw+sXH8H6hUty4fIRJxsf0sFK6PbpTIU/bGySmn8vSgsNrIHRk2Hv9Vhdnx
gMCI2XXtFdn5GwIREMDnRm5giuIAtLH3ElmqWWVUk7toAfwWTubC8DAmPDG29bruuxW6ed/IOlnw
OC3Lypho5OwD2A9GFJ8Tsuxu4drrEsITvNQveYhIegVMBJepyJ0p/siTf5TmxwF3rT6EY6gc+Sg7
UCaA5NrIv0n3kKd+bZcMhHVLfknW8jvVxH6YeEKvoQ1pJyt7tEhm5lD3ePLo+3UWSeBnppGCWvNn
sWBPF75wCu61DA8dqusIvxcvQrzTumu5lu7XqaN0ME5R89s1aCC3pyswk7v1TrqOSpWfj7cH4xVF
bFoyUb0QTN1xOl8UEVNm0N5eDDH2nFveqj6960Knt5X5qofjviKOFlCTMisRMmg4EDnMdQPTPO6n
2Pzorh4M1Txjovd1eEJ+HzWpZmUqR0UbUOs7AIfxqU5hbPi2hpfiymPKZ05x9Vk2BPAahr2+rG63
sNfCQigEyXUzwFxO/0ujV5n8u1CB2Ft8LfLJYhrr31GGULhiLhgAGX1VGSV/69qs0EGxmDmmkGt8
tjVNzk6rkWSLzLIyfzMI4B6r6qGRjmcjTYqNwSiUt2EXXCinhr8sxr9S6QIabl/O6NdqBaYUHzcW
3xHEIbPsDHKgYvyeGZ8XRKHM/CKLftSfer4LdMoHslylbaX8OQhD2XxBDBXzAVHQRRuUs/s8ZZUf
8pljLsEcE9H+TQ+gS5U5qNjiAFs6ZrqqzpWwRVJWWjsGnARGAhuV1nxbXdyKqHWtsU6vZuNNQ95M
nTR98GUrsW+M9HKwukQWWPzNjt1NHijYrD6hySTO3DKPxS3CApeVa8HuqYYXZXv5aNE9X2Qp6F0T
AZ2/htOHK9FkMPFQPZ3dx8h4+XCFIsCJ3/FXV2YLg5T+ubOOvgP+Ylo/hSKHJPoxnQTEBLPhPETO
obZ9JGcmHoiquoEt6aUwAUnwZcnPMt8get63Zt1FhNMLlloQtrtMarWGvYSF5w9//XpdrBF/BHp0
+wkksE+TWWI//DbK6yIK4TGQiwgv7oWRle/Mv6Nkj1lSARjQYxPBweD92KLbXG2PG41zE4yvUS7h
0RLbSNzq77Eb9P9rFgK3oZh9RDc7aEYrAyqVT4jVf068xzytzWiV9czTq/dPRjOZZ0eBNBaOzxm7
fJwo/ufF0sR8FSKWlCV3e6mNSQ08J3tOJ+z8F7aj5NkCmzMfC7w6tabEu3S5fUjFWtoC70LzqWVg
cmXr8H9NYqd57bTlzWyYUHhwZe8eD7Z1OGTFC0CjshXR2f36zQEh8Qp08CjaEwqiQV3uwjkqw1Lu
oAFaGWWQSlPLy4dAD7iWchMB87eNOMgsAD8GRYKYHgFGVGAyeXeonzu8WAn/Ewg+PrChRCXFIkAh
pK3ECzrKGgYviNj3DMrgM0Y+RijD+eIq8csszBgWrRc++BZuU5oU5EukMw3J+ANi+vGiD6GfF23l
fX1VkCLegHflwlRwFSMwGNfA2AQ+uwCQc3/kLH35c0O7FQC2BWfEnsDG7hBN9ziUy1N5koB8zj1B
8p6OknB+a7wkBur5okApZliOpelSOmtBo8mh/LDOcF5VW8cmAkebAhw7oDHdIMaWjnR7adeZtwyx
TOZL2Y3MO/MxcNrFTgLtrbtRLUtHMW8gDzDy8kqpCDGZtxU6i2h7F6aS6EvJ2dQwNAn6cJmScazt
07g/xh0ZQVL7y3BrSq/D1uXiZDLRiXHzwTOP3T77ypn+xi0uMQ0z1t78fWmkw2WP+BeV3q/EFT6Z
DyEiqKBXbEnstyrLEfZdMs+Ix6+UbMaLgyYdy8mHEJLABaXofEmrJUc5alYFUhF+3Jg0OgLdO7jB
jhAf1nxKGPNmFOOigWSug2Aof+M6MceEsi+0QOiGpkuEJHCZj7J2x4rf4bNRI9PlfNETYYM95AnR
OLJ45RmnqUP5b4MPavZyaxXPkQjjhCoKBTmjN0lKeujpBb8rHRYmjdcRb7M2trYFW/BEbykI+wRG
k0jZhbry0AxHIWA44BEeiuSyibdM/sLCP51o07TiBHKF0mPngPRx11O5cyd8RmFx+XRouDDTybFT
s5l6kiX7LB9dHK12EYdVMZHCjzlAo8LaD9wwxXyeL7CB3Xl2yS/GXlqgJOwWPdge2cuy20JfAtES
610RpI6Tc7yuQkO2KzdZsB55n/ioofbRXxPQmIMH4bRKeV1jbc4SneGF9k6cNf7DX96yKrFcHZQ6
rbiXtujYZgglhkrGw3r3Z/Q5U7NgSd4dkDFNmcAwA+iDc+W1yBkOB/gd0Mrn/7hyTU5MdhJdhTb3
ix2FThOKjtZ82SontJfaQExogq2qUulotMPuHQ3v6IfmZzwKUscYCH3niJIY96DXE+oWD4a4j358
BUvr13Ipv3YKRlNa1wXCwuBMtb77+IRX8unrZ9RiR9Iv+a732ElIc7xfxub4sIMsaj1RytjIqmwt
xhzJy9QCSyn+SX7N9+UXjictUqgvSK+kluh2pvKLPtxLX+PqBUjzi+FxJZI4qQK5UYGGgBGB2efT
kDmtbKoBpai8QQJgy2ig7d5uD+ylcY96lxSgx84aHLjp/ABUQCBMSwyByVi83u1oZT9Tqmmgbdva
af/DPtlU81KQ9f28UgIpR7bXVsGdC1fn6DCvZ6PxE0sgw0PzaLKCEnv7h2h3tBdMuzDWf+dilmsQ
R9cDwYxOOUCOHieXp3zsifojaoeZrrE+plD+ezSUNc/EdamvltsQJy+Sv7ZczfSRePHGyFmusfOT
rTMGMScsDZ3q9gWz+U8DND1aBXh6QQGfm5lp3WAkrakM7NN8TGi9b+aXK4u9kQN2vBExDNKIIBbX
SARiG/fpVy2JsWGfdfCO+JRTkU/R2dB0EFKWmBcvMUUc0yuAdcadJE/VGK+ZTRlZFz9jROol5JGT
sUO/hm8dRKDXzDe5EvniWneXY06gMl8gRJ1bOuSl2GXt2fodVu54qw26s9JawVs6tQ1DHV96R8BU
FIczLe5QCJMOwny6eKh4/cPXHGrkk8n66ZEujN2xvswaatY9LvM1vKixFUqKhXm4pD2NsvQXM/GP
9A0NzDTVFqGvGPdC/YoJPZM7/RrITXaqYofn1HLUkaxpA05NFYYKP+BOEiLvUlWAloiasv4nFB+W
l3spv+T5CLdGO9Sy5cDsMYDPsrfnkVP+Et1cqc9QR8caNDmkR5HciKDu+4KnrTEhI4wiqjBitOSu
j8sA+BPrRwt/QE/NwHES+ls9FsA1udYtRk6gn7xgrWFuWFRmOrJeD7CR1UNF3yNbDdbolWR4PV+1
w+J/xOgAyhScE5TEdK7U3DtlXbHNMg+Oq2MKpXWsKW1hhBBpAaJIK73p2XrsoCPOCcODMHzfV/vw
aXUITNwj/bh4TrchahlTFiOg8HNNLe5HLPqrzhnioeynUJ2y03qn/P2oJQ/nf30+4FhGnsRb6VWI
BFYcxxOaxILJWNJPltU9eVtPWhjQkyq6bs2PkcAjZ4nBsORcFbOOs1ZHV9wkqwc/G5A5ez9ETZQ4
yyZrGrMRuN2LxOwhbOz3MDEZGEGsD+bkIQB7ZoFNsLJ3M7jNljaARjuXoZRCPfhxD7fR51meFc5M
Ze/T/XLYfcQyBHIURRGGsx4LTinPWxAPy9oJ4tnKkluBL+/urH3IvDP4lTM6JpOY9UgCY6CB7fef
eGMqe2F1V+cXla0pbYkF58u/dVU2PloMYkxCmcIFw8tO2khEReFWuTkn1VVPHKpmebmJkIFBrqcc
5dnHx6ECELEECfSERyro17ukiygZbdq5asIF7YBMYUr1MtbF7B+eaG4QfMN2/GV4Hmn7uzvg0xkI
ZIVKdqb1nRv+8BWtKFwqg1qpgjVRFWjyQpWegsLL6V/yJ2+69lcZFiRn3eUW2Le6t6op2MhbP9Hj
85/yfxWE6zUeHFkjKKnF9T5Oks9BrHR+CBjbUKAnnFT9d6v/+5qdO+4g+HH85UpWqHghN9jbvuYj
KOCrTDV3LfjQdgBAlEahavpVNg/phPjYYw8EEFaxc8UDzqVgUX6xSo/bhLgZ9igvlg4ETNyzXzfA
E8Q89FX7e/EK7lDDSRr+Xkz1A8JdyhMFmsVcVMzhGA3rU7YnHeXzSmBFcvIE3we9D64r65IqCIhd
tSveQzZ6b0DqVTIlu/AK4GokfOMmxGhijtHEpsRiKpAHjfM23KwCsf19DURd7Yf2yWRMgvv0zVkx
sVSfEJgMuZdL0mDr2y2wV+EsTL+Vkk3zIfhtxBWAMVp7ih6+K2SwKATk4v4XXD2+Es0LwF5kZnsq
//rulWmt5Vxa1L1oaRcn1PuM1timFtUIY5J8xd8fncSKO46bHrPcPO9njUgdOq8NMBu7KFLq39gm
MqM4PkcAco9RR0LjWS+PPSaDVRWr01kSpTqr/F42QVlXEGRB+zaUSGGt6Q1cAGwm7XR6KrprCesx
4QwHeVnGcNNMEJc9JBk+a97K3A2Np/FM4pON57lbDolF6MqBstPM38b00JfQawaFUD5/SJ4j89g1
uxJt6XwIO2twHHzpXuXwKUVdB0Ds5ddGWbQe7i+orUXqvQBB/IIZh+pE4aom5noM2KaM8SadVoQ8
TchVTBj+EdGwmtJ+4Qv08f5suqJ5YgJFso+1X0TQsFtiMilk+0XrM5PihOYEB13CTUjPTNPS+Kom
BYUU5064WMQJxv8DadWf9FWrC5hYBZdmKJGTn9IWkYOTH2DgcKy3Fb9vBhdINpBlcbOsdo+OyNDL
pM2NoB45ZXQ/N3+kExVbYRfWt4SsIGbP+k6aa6ikljwLSjxH85B8z4IROLJAuJW20hwdFVRixCh5
arRAuFUhdlOa4C4dfJnygU6ape74KRKjvg0c1HsiceAZGDAaGbA8E8bMskYCZKvzouCm23emdWz2
zAO43SH5RVIP4ZEGZP8n3V90JEbcz/CtlwRxvgaTqtsJzfZ+nZ+16lL4ze1KYP5ojUPgSUl+Uu/M
pJpcLKfGZsBlVXwQH24J1tlHUHt45at54zplx9HS+e9MUzGl2U1rY+c9ACRLrG3FWLSrbiwSqF8B
DipL/PHFf6CA9C0cCS1hQwR7oHtdzVAFvM5dx6fP1/+UZQvVD6cN8zwIr2VDkeqFWE6nLQtBhEsg
Pb9c3agHjlInf8uQaGUrfLJoxwHkOsGvw+0HnXkC3EgNFodm/7aP0SzlNrSbTUEPf+0BC2oxQRe2
Zi7hWh4q4pKEwHDa6htJ2gzeFJryz7+q1X4a5hyroGaTbSObWpADO3xmDifN77fWAXGjXRncbJJQ
nL7zQOA5LkAT6mBjMKJ15JLQBLuBZP0IP6mplcHgK3j4+04cflXMZRRs3UayePyoZ71uyyFv0Rcw
vr/KBwi6q7cO/s7NMiyRhsSID1GrSvh+TncFzTIuwn01tQDafRVHIpBxxaH6j3QVxvaE/DKAZO9l
1+PU1IwflQHTj+Lu+/4ozoO0P/IT/znMOqtYo2i6sOpuD2RXubUdaYNMJTJohpuZOeD/23Kj4pH7
FCQiExIegDZSJms5jqobPU/4uRv0V7nv415gTd5mLVyj4kjUqFjkyi7m+JSVQMmpK/SGCdI7Hbbh
H8WY9n3C/6z5DyHgxc8mRoeg68gjUGokvQR58qUXOXHDF7XfC8qNxMPK2ckb6zgS9tmsNmC61pOf
XfNRON06CGq2Rp37aiVaaUTqDU+n214bRdrL5TCfE1OpIyk/zoo7GE9nJO7CNNIPUBeWnw3jFr9h
5ildx6bqA5V5OurkpajBt9c1yuJCCwg0CIqRNVv2FFRTyro820goMGjQ/KZNbK4T+uhCl933Arma
R1yqv7IeK3fyd+lnkb6BzT2wAIJ68zbZ/OWrcv27kL140eHqV5PgjoGJ3AXa4x9+Jt2/NcsSF/K0
kzyWtoClxqTiDB/d6fxgSvkNz+Q7P7iPY4OFJ+FoM7qjeeTgl4n45uWH7wcxjeSgwDFBIEOml2iT
WeoRfLzG8h5l5/A4RbmbkwHEU6ysMop4/DVxhNEeEYv/Cg4ohn2bS6zYb3mhqaWRn5BQQWITWa6s
jSellAcMWjL3Dfu/fGwRz7NZWUfcJXl57TgJiOX0bYbFMqaH8rJXQ3H1l/zWXFlgdKwkeiceh55X
3YCJLhsYrKVMVEq26JK1233SM55rUHnXIIRMEPa0/4MKNgdqGOQp5zb1uMt3SmkigyT1BPjtGP/0
DcgspXg8lENlf7Q+WvIwTCOEOL7oqvg7fHYqfPuQGTmLw1Yv7KB4xObJZjc/yqgk/5E0y/6JO3OE
3pb5c3o/98P/wkSUwDzCEGmcGP0nvUONtWzmhBWZbnh+mu0w24kCpEKxULvLJM9JkpV2MDeD1Wew
Y52iax9kEy4TLI0phjcW84EA/YeAW7kQpbWN2gYvziz8miMuT6ED4gjSiNq/SjOwp2wwJWHaYql1
vw5K0MnHzrsAqW9VdYwjYtrp8lUqeI5L3VjnkmeSx9Oi4ht71ws1eiUx5G1hz07L8qEY3wdWhKSw
0YMylKDVa0JgDYW99fZlh+gV0uTvjVd4xrbclszftjrQJgo7wLW6tRdVbbEFO2YrqHEw40H5Lfr5
HjjxFlgBsit6RIg6MP9Vnsab1P5oNW64K1BxMijznvVBXZwK/6eJvSH6d3a+5owKOWGkbgMcEpOI
L/0smo4tq3F8VaYoozt9asXUL9XB3sH+nNt1JTY803kYVwjx03inib+DstZsjSidEMTnGhhQj55a
RxqsUKHkJdADH3mhLYFZ7U72qx7ji08WpLsQ7EUDgg4mEWhN7pLFeye1PVLcK9XmBhUsK7fm8Me2
1Pt3yu6an9Sveb/R/TKYpjGz68VsjQ4fTro4m552d6v8xbUKME9LJE+PMoapE+6G0009buJppk56
NGEmSWkwWq/ANRGAnZn50/6NjY4KfjWj2IZPy2PKba8m3/TcJobtcUoILfSsNFWQ7AA9EgXy58gH
5wrmKVrQwOk6r39Ckrqs231t9v6c7Iido6ArCqHJultUu93gUO9IKFuDtbwbu86Il69FCIu16uBq
k7WP3vuRX04jaDGKVMF9kOJ3bLUbUzYg8oQo894vq+31SMOn8FrzzfmnvwQp5WsrUop1wHgFGL9a
tzcLqhsHPFj7KdYPOiwOF/8ieVIlls7pKY4g6QKt55DKo8/tUdDWkplfSKiwr6J5Zm1Qne4uP6os
MDxLF/4Kj9OY3t8aOwM+Aw5pDa+6Fa3HGnrOaIQgELSH7Gp6rktSRAy6igZ+7DnJJc4LZgSyIF4c
UaNN7oIO83uYegFVS0P3gM8jJYqsFC1pno7jCtk3YiHkP0/9Uxbuy9XUt23rgnefbMaC6EJlrnt3
J5obGQqKCxmL2Zr08NMAu5dXHtE+k+AjUtT9uiSU+9alKuoupGHsdiDYpjNBwbdXTjtlYLcEtcEU
RCXxAGzcSIj5qxIRp6dHX0t8CWmWjIQ3RP6wL9YcxRu65PJ5lxlZBG7POOhs4DdBrDf1qxkY5tJD
e5UYtdHlDljXa6MpXE9U/Z1S/Zzwd7tq2TrnskzlN8gAxJnwjOxIRWYhoimEVe43X8nSNTrWobFS
BedUOIvK4IGKbPMt54VaRCoMSbG3dFlavBT6MVbUy57bKeNItoCKHS78DyZ/P9YIuuoIiTY4Zs/E
jV10+XNkfftH4JLF8MLj8iabEvYaDsYFKHcEf+gTwLaQpvEpZLwt/5ynGzBw7knPxyqehJC3giVi
jOX5XGuUVyYCS/31XSZ775jlJHRX83yX3Gi+I4Nv2oLrfNQUMb5tUOHe2Fh5lAQMEXJ/8hLhD1W1
FG5vmnDInjAVlqEZBWS01GT8CoU19n1jDqQg2PKfA6D+HPD2NONA+Aau9TIAeWdW5AELsMDnb4m5
Za+Obhi3IsiyzOMWxHtRcUrHEBS5gkH5rWlZ7d776SOcuS8rvrPYqmY0VAy3R0BfcOj8zyFkCGiA
7tSmyh5yKWbQmLqQf2Fx7UBHISK8JLq7v6YV2lMAONvb3Y+Tn4UmDEZFIoXdg89+C/GFEgzCpIGR
3A4eKSpJD7/7FOPubmCM82EtwhEu3we4e5eX7EUgNh3HnJugzcBO1a/z5U+iKGIyRQ3edIEavfC+
WSopbuRsMrHj4QFZTy3k6kf69GAGbrUx066c3M2yr6ViTVRGHJFWNEpyk7XZwJEhhHNFPbv2osSi
wAu6ov40To2IQUlDmmv6axOjEBCc9PbanPaUZn7v+9zpfqS9FuBPaoKE5m7d91rDtOUVpX5UTVFk
E+UFn7N2D/Rs6u7mxiHXx1D0RrBPFYfCrp3YttkT1Kj4JqmpIKcCCdm3xaVfkR4GvFwnTf/uqlnM
gzCTal5hA1SoZHxfcEl9cPrtfg3mUiNddIOxQc8m3Fh2eSHg8cd8gr/zxfOJZaTRBlVnASDswRnX
PBr4812w3n5MwaEs75SW16i7iSsPvel9SsgZySWL6scSu0JT5ZLOpLdbPpskOVKjjknEfFl1AANq
Rbu9yKnC1hv9+XdaqR/Th+84BGTt0wDJdxj1TrGL+GFdAF2eiWeciEFkWNdUGeG3BkhZy5/DSvnS
I2kk6YTWeYeSuPl2IhunXXmTv+8+BcZMIKAobObwQBGJtNoBrZw6SYiSzwUFjEleFcWebegvJEx5
9+lCZlj1D2BU7WYO5YJr3BhR9ZvPiU0jlmGp+MErMYYaRhlGWCbw4b0JXEhVV7NxttppEn6ipB4x
mhJVj9EsZ4TwzDd9Dm18M53YRcz3l3+HBzkh0hTY19UIJRvKrnDvM8liW4IU3tFRhnqeEgH0m2Vj
byHRmBNmu5m29nqUU9Zz30TH40lbD9wGxtoHNVOU2Bk/PVFHkQGX1xTh/7V/uOl4nQHEURrdVC8e
uYuCvp41RtRFSQoXyqckeGn3zy9Q4LepsrGothceaNRtirDxxrJbQYTQpA0YdRUiq407O/+lmzQd
m2S1r7zarljyO8eiOlDt7VmGG9zQP+ItBwQfQebijnfgCUKT47BipgnmAB3F0wwtblBN85sO/bwl
uBhAxM9s7I6K3Q8+1i3H5N3C9OgPyFbHySNoO/Hmr0lGr73YB4PgSNRUuGNbACBoXXYB8EgJar1O
Pg4DUiAugTXwALSQadvkHdfBWEF4PO0gT40HUpRKhpa3jxO64qLZJRGnyabWo+moubCZDa+dcdtE
7egufOnisW03vi17l8OogTqsH5tVdyGLOeqCABcr5DZKfFYv/SovizQ5uROoSDCSBCNN3Do9TQkf
m3wauEVITKTDUIWsHSjIIawXf+GsKM73aoHV22Fct0R2yZhbddJ/XyUUk3nbU3sFByuNqv9wDGam
ZplA//JkO0sx+YqsEe8y7DSduEMfD2ZAIuaNMW/dJGcRMqOFLjCenVyxolfZL2dawB9KFC4V8kot
KCcHxORWGqMtofwg9juLX5Mfj8HvWPRaIIMl6Yad18ke4SzZKDKhI9nEh1tvS/nap8KqWqyKE0hk
9tZATNxUDlw3Laf4RRU05/89e/ueHWsdZJhYZwBLdPuBcKmSbloGMVHorEe+DkbCV4fud9G++0Cv
1yInbqXX8ZB0JfF4/rMGPLbRHnVLcNNYKoy3al+BZ+LgkAocKkaE9zqsmaL4TiM6R+dgfT9jvqrC
KGhEPw9wE/K+9mF8NoNJR9uc0i5LboW5/eer7pLBTAX+WCdcVZLRcIqjkMjeBjKvC/PP0/QjIfvQ
kwgFKPKtahRfI8cDLyftpBkXR2umMR1PR3XjuKr8VgN1wwe+vdOEcrIkWcvi4+TbfzO2Z7/W7pjP
eIsfzkTKn+k7HwVhux5accxje1BqClatMEA0mFtxVSnHIH6HX+qnRgmM9rwGKyWwwRHGUQ7VfVSq
s6RMClSeNIeMKN6j4U6dqr/Uhnvc6gErJQu80QgdB+1DyUUXdDDik1P64s8pLRKVlSzQzzfz1APt
BokWsYXh8Ts386yrhgJ7lMjiQtVot5nB2yi9TJ1CZEwEnCFsgeluSQXaugYzmaOHFRFYlDSwAD5c
P2XECis1i5iVWCRjjG/1nq10uiMasRxlz136Rsp8sK697x1Z4yNgNomW4+5sHQDE7ZzetuvXuH0F
XAyacVmEwimJ5wSWo2WNh0c5o+4w8dOHL/mvE/qKLgISqpTGhIKrzyKJ2KKAnNoKrgL4LI86v64E
pRQuOykihflSVs1FYLtg0g7JcVTIJlhkfs8ql/sRZ9ghuBJ0f8Ms8RG0xCIrbWl4EZ1ZGlymfTwJ
+/Gc6Bi/aowZ6K40Qyhy4ngoI5+JZviweI3eV2h6JV6ySehj+wbTV2pnxpW0y3KhwC+piKjoFD24
cof4T7Z8wutfQP0y7nvBg/3szJKiBvrj+xDTswZmD9VzhRdw89/hCVxsWCuUayuzBf7wZCrTHrRD
WY5XGcEi3afZ5WNObPDE3AT0rSTrift9yfoTC5h21LhKIso7Du2GJqv2BMoV04JjQO4rBI+yASOA
d0HoomTDBhBSJrHXPN05gYIsLU3/HywY7cmdYb5YVNHCelVolSUSIT2dNRGRx3NsX8Aj4KeUUom/
yXGhiBVX5I3Wf5hFhZJaEix/LTQPRRGIFbUn+SYx58ONd4bsqGYNG7/bLreBLQWPYAsaaFHuuvfB
A1DaNkhN7gS70nQe1Kp9ZI7yqdYPWEYPbxVNS/LmjvX9joTUwJsMqKRE9+8FyIcm32/lvwqDnY1Z
rfwu+kePFba3BUU+7M1UjqFirhW29Sorabb5tLKS1tBY8jg53qEnhbsBkTTTh3DovCdtbOW9589C
AYoHtpaAbtq2bAEwakK6Ka3W55kYaTNCZ8zTv9IKNk8ZIxYYtuucBhPdR5vs+ZVTqfJ6oWpH5f5h
PhgoCYRuDxH+FuYytGGyOvS2xh+Q/s6i0rNIeI37a8UdUsIWBzfJ0q+g3prIvQX4Fh/J/d3mK+ah
KQFufygJlZBY1ZDNipMmqxegX5WVGKeSjcqVgLtZcl0DkJ06P4292PL8kywnOdhzf0bAZMv/0dK/
MKc/DX5mEwyo67Uhcc1A8rYb3GpcNjql5R9VXIyOMU7K6XF56R9Yg00z5SklMBtbx4YcOftF7+42
YASfiBXnegiJxJfQACNsBbXnQmlVwuWMjgivrZWnsSqZHlWAABZtFxMr+pn/gj0wHaLI6qZyO0oM
eehmlszkvQQIu/LUfCixO5sgbQMkD0z2ZvjEXkPXfdT+Qz8etXzeBYPy6lQ8ClpFaLF/XWczPop5
IX0Uqrmho7R0ZWtyNv1seQL3CJW9XgT2hL22G2eNWV0R1etgtvN4lfjKFQuv4IA1jg0ptX0jo5EY
vZtPjW0thKjguguYg2XNotfWKu/J0WaVQ+x7XXEeAG2GOhMqHI3EDZSqRusRUZ77oRdxBoCJ6H1+
lg/WwAT3gIXOPn1o/awZi5y82IYFLIPSLBAje+9m+Uc3H6a4h/gqdBQpK3pYD3C7UHIhgv2S3RCJ
GvNMbb67LQklNb6fUNf6nU0ioCqd5xQAa98GHt0+MnBhDnnYKBKKms1XjNPaHHeR/lkw0ZtxpJmY
h+tnufwmkQFmMAgDmCDorTNv3OVDNF0Tz69pETp/i/6sOgJ7ItSORN/pPoEAZGk83o5gbipU9Nnx
rAPhk1QAKIDgA7JvR7pLA70OMkt3CUcsSd7F26t9+Q1IQcLmyW0yP48dehw8x1QqFocmqUgJjD3t
dwjft6SaTZ1pOxwl021YyEOKqMtKu9+lahse8kmkOYzxOYWm2XLsbvIeyB4Swt45DPs685yJyLGp
Vgiirt1+aNAUOyGfAIcORH0CKVZftUlycYKkOV4apsgWWVTVyfLZAK3Mjp/9t8CBkc/f3p64rnAn
th9lQ1OjYL/bR3EeVgkrSTaWjisXHuJ8QF8KpTNCrO21B3+tcDhom7K38x82K3oA607eIcIEBBXr
i2Ml6DL/W3HRW9DgaSzl0cZCgSB9AXmdBMZagIYTcxyPoZwYIrGQgVwVLBNIYQVGZovZa/AXYZFi
Hw4yxO6ZtDrEclOgFw2cUihCwF4JnJQqTWiOOTq3L0hV/9ry0GUCYLI6DP9h1rM/1+vgWaCyPtCh
/LVaed+e+dHxztvGdJpT9hbnVyVO3kycx5DDtKmy+WT9Eu9/Jpeg2mUPS9lHhIL6M3xgcFGcMUnk
JaZVA+q+2pQa5lHg34zv/FRJJVvfdlSI4bYL7JbjLntXrtpexR3hH9zslbZaYzGhYwzvhK5eCIh2
j/XzqPu9GA+gIbpWQhA6X7/qOPzYbsm5b9CZbqRA2U20J8FSRKU+QrmNaeVmthnhf2fGoYPUMcTP
Ob1uFhnNe8mGSBpuPJalNUR0Ath7XZDwI3saaO3ePdK51ZzPi+deCrKMER++DJ+8cPlGz8O+V/vX
9Yz7H9+EM8lHf9zvt8kKqEpJctwVXr+FyxRD+5dRwyeeWZarp4LYOCnm1f3KnxPxXxQeM89URz5V
qQiRqq4MpzmKgDApwFSjWJ3Hs7WqP8N0aEtBDTeM1h33zmnx7anfenK22A3gSPXjUqLfgnCDnJ6g
I82JuwRJ9aOfUf1ycsL2FuV7sjqfYCBhEIXEeMSFuWPpnyjBpwh8ADGb6/UleE5HPziiz/bQO2fe
NMhvADBeT14EC8ZqGbzfhI/EZxpPpacSIYgd4omyHEkm/qF6OGcnMUiyz1jwf8ZHVea/xel4Ej/R
+NLCS/po6zhEaDyKkXuwFoz+GI3Zljkvj8Ler1roDl0M0wk/j7x6T5Re0tljubVQ9+KnxclxrKev
1frgiznbypMIkg0iexCFy8o+7bS0dRTewSpwiX7tIjio2Cc2RGBgQPjwZ5YAM4k80QO2ukyeKkU8
1EKIVKTExfoZ5EULJZIIm7HyNdFfnQANrjHOfwJmPtSWpE9s5BAyntWwc1UFnI/cHvVTYMb7UZsw
R6TuzX+bJzif+Qb33QIgoECaH1C0lx7Cm/EhZT7aWBPIgQ2X9Y739N0QmhWA0xkRYZpz9MjVu3aa
Ti8H5UEM74PpbV94qHDwl1WxYhwDRILWVmxgqKz6TpzLc3wuRVSbWvoX7+w1VFWa7tbIyHqy79KK
DAOSnGcf+5sxkwHPQFA7abtopt6dO5wtBIO+dISZApCRRegHIuKsCXVtsi6Vlyb5IY8q7GC1xyn7
qsh3V6VHTfZfdQjvsVgqi8cfXDUT/+utZoRf121R7ifOwqs30F6iJwQ5WRQ0QMXZOdwDT1aLH9QK
qaETAgDTOC7PLdn/g+sVLxaA3SNMJzFj7stlpxx2CrkyYPFZYFbPU9KSOeeZ8oJHmiQkYg0i2lMf
bVqtdrI57dngZzh1e2UOekhvHIk3KWDeIv7NFXhDVaHpZ3MhCYX5rkYmWz3/KDiRjigivDqPgc8m
qUrRJVssQuF0TpuuZ2hkIlhN/Fn+SUhZOzU7fj0dCNcrYodbesJwgn1j1OPXktOHMa1vKcV/m8Hx
S99Dc5kTnPqglyte6RgavIxh/wQs9PkKgnxuWVWmVxWv6rULwFlr20N2ngj/hIISIIauE+PYN5Qz
r+C6QMtA/rxYT/9QkC9RDEeESqSRY5DLFxmFtUqMbY3Srt67lgPDyfRmvcdgq4HHv1807NahQ2Q0
JLfbEAm+Mya3w7Uqpt9afKTrRdPbTnrP7N7rP6P1D5Mc+i4KBTnHwLL+K5Gxj7e1PW/pkEfac3OJ
/0lgLpLCcHNSSO2WzvVCzY7M6qKQxWQUgS9ya5/FOpMR9X+c5r0vVkd2m/0DERgqs0XmZlQ61CAX
scvscnXjfsjTFm9aC991bDYoAbwKpceBxj6QRiXbB2oTEsTmLGSiO+5VeqQWeR5HSQVeM2498TP1
SybXG3q2cMDeuCmqy+v1Ic996UD5aLzOQrxqjWvqKobT3YpyGpXy1ADdJJMEWbutNGqB3OayD18C
ADpyF8v+saxgQnph+vs+nhkk4XP6oA0bER8jXCTlK2slR9Ff5Cyk/Wbz88/e/6mCOgIDMma/CoLI
GRe3AonXEAXyODDrEv3Cak924on5sumqmM1v8wU9e9akCqfGmYNbMo60qWOGkcLqzA6BV6IaZ+RH
h8Ik3k6O6VuRIvaIycenRUhOmpWZzBipRKdU+oZRQBA0MrTM1/uG+ZbQOG5sciwYX1KMCKblwBGa
o1b5nPVYaW6cEv9SzCsHplrgzzc+67cWzoFvBFYsGFG0IKQjgyF1jEWp2LTQ5pnd87QeywL2sD5T
dTeFmnXyWt/kgfQI2iFRsbKCbqy32vqWEoMdzhJVLc8/uKAv9pzNjpXsAU/4dvWsvC2/Hjghpvb+
RTP8ZRb0JdhYTjc8ScIsWVeBv2pj3SDDYzW8Wp8In5EnSj8ARX7nxYGdJmC1Vc6RP+nRTjGBs3I9
eALMZPJGwoxdjfaRVNszAkC/ws8y+IrSrBisu739TI1tECZEhRuDcyuvF56pI1CSS4oWq0dcO2Ii
OS46hEEmIGtRAt/MDO8nqE6PEE4slClsIZ2wgW+MQLTkOjqdHUKuI/Clf4bcPdNiEAz9AnzWHZUC
JW8nPNBdCC82v6tzvulfDaPT1f8aap3wMtp3OTc1aoiCpQsw5qeMxk+JZQpwrXx94DtoObOYmouc
7HszG5++kHpznPeExzJBVPXvV2OoFM0QZRT8VKmX194WpVKzhXDWrD9e0qwbYQWqJS7n0od/zE5K
m6MkzWNYLPeLF1mCgDF7U7UErh09z44FFveqPumbL9YNBxq50JMIR0e87QhLIFcTV7Oyox8y/QeX
DxN3T1T7SYst7kyEZPNzmU8kD7y/A6BsMGz22Xrtzr3f7heq3/RRpmOJLFhZNTn+EzGpuPTFN+8v
iu61eIpqc9GFNo9a06I+v395eM+BpxqAK6/uu+yqpLyqbvON+SdTk2VnxvCh3qoQXRLOSrEgsfqa
JoN4KwFATdGfYBjTZ5obYdkr088+xd2hCyCGAZIZPQQ3+jN0trac3L5ozTj9qI9jfvhx+xGApr1o
AjkTRqS6megac9Zd8vwEHWgWYP7LktYpGK/Hf7AMPJiyxbo47LE1oAT5GkAa21bOYLXL8O5pYBxf
UcNvoHmpM6Y0+3q1dmV9U3JLoaYpH90dU7Y5G2JijyIZ1ZNkrSzIR702BbpLy7N4/reJ2FWL8cGK
AUP6ChSZMrf5bqwqp+QzrQkdbar7CHTQSKds4XI8V0rrVcLK7ghdViG+yam2JcXnCXeIChtqcsER
8tS6SbNJqOI9BQ2W1CuWoSEV1nkFOHe1e6wK1SB2womO2uc+vYuPCt4vlgeJSaDZZHJqi9OvvNcx
FV4mfIDyFVgmgwc6r35qGCc6Pbv1EgOqKJUsq3ktHzLU6cAkz9l3NZfGDXpvJby1QnkSCNjQeQ+L
CoQJ5U1roJE6J+PjA+51rOUlEpfXW945VAQmR9r/zDhhudCrX+PQRkRVR+X/l6/SKMFTr/M0a+Gu
5kL05Os+TEevBl7Ct6lDm1EBwDLnN+HlsvfNP6MFl07ptEhG+cfZFYkrYpCj+looYyTt0yqJ6drz
5YaxS8ClLr42cQa0gMasCAZRHEBSILIT2VgHcVPi2Xl0Rav/xUsSf4fJZYgh0qkTUj9f09rd5e1t
0mi7dqs4ziXGBe30Yyxgwee/fhHiyN/wB4dxAUwq+aoiC5BHg84F3XA8xBGUcpCBV76j2gGlF9W7
QQBc8HqEEY3kneG/pggTBKrknL+SXy3o7iGMFUeq8KbZRVKs6YxOgIcpoWkmbVTMsxBbAHMPuxvT
M+dCr5sYvRNj786STBCv58QnYyTdwgUc8AlAvJM8xziaeBuKHe8DQK9tN7FOAFX5TA6tQU7vAdSE
v3JVqHtBjqtaOzq7pNZTAJG3KmD4yijx7r0rtuF8brC1ykYGdP9UnVM4xSOlwIadUKwzuBwWwo8D
YzS6ymg/zukD9Rz8HyKsq/i74gRCxog57KIbc86XgxwfjdUwbQ5XrFfn29DciKTcyVJM1lyog5YB
xpZ4FTAchcEgPiirt2IJwpXs41Wlq1Dw0hsnYmzOM63KcEgsHWGuVwk4nNaX7XbYm/ez7t3ywWFL
1IQPRA0nVMhscr+kXnUEQcSJ6rTy4m37pJqJwEI5hQ4usdeUEg/fsaemMsRxxb8KBRvfsgt+6olv
0HXCKsXZm5XRgYz66pbgasYWrlqeJ4zZbhWQY6Lb8Q2G/+tezhF5jsk55QeYimKXvU3/6MYQQtJk
LcjQMymZ5uQ+VtFtxAqGym+4MLcNRSJrK1WaOsDWXpe/Iz5U7G6g5VbaFWZT8L2OKHpphh0NToLh
5U5Z8cb7OOijD1x3ckE8b7eZE1+Z5aXCbtIczOETdpUNbsES2xxUrmHwcZ7s2NKlMYkrETh9sCeF
mbqkrN2Eiavg3qX0TG1wfUnq2TB2zk4KH7BalgnPOTy4GXdDFFBNNxZo6NFKEofKGMRsGPq0rIOF
6uBXAFwIadThc1y0fbHvlyd5IqINOLoeqATNUkyEzJpUCZk9Birr2YPixO/cSkUrgtsPuFxcAvj1
Dap4icCrDLcGj00h+crhQy/22iZNtwmLQRKHa70iPASZ8SWDD+x050XazAES8//xx3kpBTJRpFtj
LTsXbqcHrDZLuPw9T5m56riD1HqXxZ7vQJ2UlK4UY5T05nmdCPcTfpmb+/vkVP2U0L+iWscHajV4
dxdA16jmIJtymjrskPKdLkrctOsbA/B+SxqbBTQVrCE0+ZJ4bSkSqPm7vRZ9pEukpHD38L5IzDCc
zICz5jcNr6ALMedogu8QFP4STc6YAhY7FQUf1bsbkJObgFu6CqmONwB8SFkvYPiumbeM63kKlcZp
folQg9+y/VakQm/3LdmN9nwMVruS9lgxxuMfAxl3cbwKjMVJSGUZPPDPpaZO5Q1ijJSArGlCMynE
/aJyLegQDxytE6pbzzLLwyQQ9lpsYgVeJ40iND5WdbYnLbBAPsk7J8CmaspNkBQUsdJMdUQpBPyk
iNfPOWev1W2G1LkoYwPQMXN73WvL2Z++jDphENIeqVZ+zDZvJWLJrWa6r5Gy+BLCXO9lkHFXqt8c
1r/OcT7byFa+a66sIjrTmH+zXeakXallOqptb8oFwf85WYB0Ae3zhZlZBbC56VU+qS1qDzUhx+Yv
TwxHlnoKP7E/4yFCSW63wPTpRL9ESJlqr9lFVpao+c5AxxE8LbCzMrcAmkPfXFH7a4fS91mAD87Z
cajdbn3x8MpmvItFqu0/Xmqwjyf8FYgpPjdIcHQ1u9NHpPdxxR3kHtuEatAGGXKYnYCkUYcaLEyC
jSqKBxgXh+yfk/08j/WOSEOylDUlQ9S3EDNnv5AV8byggHjOlhiRQDzlpkAFvgYHiwyLHxDWHg5i
X3ux64+1O8KZgr61HCwxAz3ODHUKFAncbG1EA4G5UcI5+xH1HCpn2oI36CSm364n7RHaiBSw/NLn
uS42mlNSGji7VfOjFO8/QayoclRu6PS6oAUd6+IcFyTCDGKFYEYvS77SSogdKRiZDVdBxcE4YQI0
rgoYTvZ0fSRqia2KOVedXkvApm3JJPdWvziLJ+JLFTa5hmVSIlpaRuKgUpxidvrqO+TtXPBzpdCx
IyUgyz5F7wtWYTUaPcyICsiORmVZ/265p589Far5N6qvtKOv/8lxAvjHy0JPDevACslubDTqLUTa
JdZeyCge9B9j+qXi+vJ674rbcuoLpBWfVXfmvMyAerv3dcqQxO7C2fQV1W9T4LK8XRsHf8RaSD5x
pD3VDwlYGUILfRoIIWER5f015Bd0uwD8CFg6I4xfUobP+8LThM2xU5QHydzwbAc00Kb+n26fqT2s
ShKGR1ZCHnITyxyKM6NsmQcWZvibO5uHhpp+ajCAaAQzNik0E+hRCqaXHM3CxG4Q5br+ozryoF/s
U4c3mqcRJQkjs2ha8VyCzXUyAMZlQ/TB2f5lw8ztOuqJNeyj8fpsgSgaU4BbI6OqvkbuFQUIdqxV
OoAQljsanCPEJhqlVrPd978z4/tWYLMiClXIfJD52y/xr4Mz9czsqaItHlEi8oRrFVX+7vgZEBu4
1Yrlw5f2NdoUaCLzJRJTsAsTlwJp6KpaiWKXptQlLsu8ebPdAYLwFvB26AUG2TaFJ76LMfEZ1MCv
Q00Xf6MOOPT2N0+3E53pTz81OOc34ocdU9aiwfl2QehzkIe/CQ+DpRrRKOzgaTdZ05gWQFwu33pc
f3sa3NSwlHo5yjBxPW0JHx0yjn+Hpy8HNE+yuavPCNMp6zYTK7w1RlqEdONl2HQvDOFMmRWTE4O9
e+UJMEknb7CSm54Xs330+Gx+3pdJDOFH7UuT45GRybK0U5Jj9wmDANiH8tVfWW9iNejgait29ZvN
SIKFOm1sy59aXZCGFJD7PpBWHUmMJC6iBqHO1+1E2FFf2H+ZW8qT9yeAedlY5NXjQLGI+VhAeEvN
1Ir8RXBDj2dN1ZOg+gr+eknv+bYfeI31vKKd51H4h6EREv4CNX0dMzAi8bPivSMm5MlYrMERWIOU
+j3qKMGtHZSxneu/v3l82pxpVRK1+FKs7Em1EhOp8sUcu+k1WSetNg5FH4HuOrGw2Ph6GOMZqLhx
PiwTJ8sv6TXc49VJLm0Ln/wL721poQXPR3n26r32SxKawTntzk5bwj/8dSzGgVQTAz2ncEPGDhg6
RmvC5YX8fy99OCKHFoC/hd+3E1HmeAySfbDyTQWd2PxtaiW1g0lKoXAMRkoZuo2wUBu+F2D++Okh
WjfHeeEQeTjBXA9uhZtGOr447BtqXss2I8p7SgHNsPnn8ZW9Au4JG8IpUgXL1mf+doNxfTNWIsW/
GXftRUDV4RQAXoegUQ+pRGLP9iNwNCOjb0ZZshpertWZqtDKaYzUTe/gNTtGjWPL7926W6w3XjvI
AzhfYjER0jthfGM0ynFjmqtjj+zECWkJlaaYwgbOeJV3MtrI1WU8ce0WTDnG5eGLpGDa3d3i7Toh
KGbVgh/6xebooDwlrMenP7AhXCJHEL/s3gmDd4Sj+MP5ilZ4w04jQ/gUOy/w70XdX7CHjE3dwff6
NLQsNBn4I0XmS+Km/lxtI3Vrsh189IrNgPkY2C/YFVVZOopNKDw86jHXS4ItwlA/6B9e6IPUNY1C
/VUabB+/dOPF1sVqTojjpjymRVy5Gj8dPpcv6A3CW6DbMgoEXFigWwI7NPliePOY+GDqlOetKTZU
2r+MFcqrMA3ao5D8tlr/FLLk+vl7qITXLarLVplQ5QOWVMm85pFt+TqiJEij8WHpxbsVbizz2820
wnjbGn/5O+HlESMmpA1T3Z1xuOEeQ5ZTPsucfveSmRlPlzVFlVw1AVlkjODByNLt3STct0Ucckd2
bBh2mTmBMpovo/rw3+Lwl6Cz0j1zy9p8IPjtLWjJHW0JGMddHQ8ktcOVtn1E0Qv4fsS9P7nYeew5
uygUcxGNkXyGJ6Kyuopd4PlzWmRDacutdVM9Plu4RBF1gJmudsf5/77Lff4hRrXV1NhsHe7oOPSX
6agmEqh8ZxDKq7F2iv6ji9ciEZMbzzNjiav5xnUN1zE/C4sBYHcm9LogU6F27NZJ/z6sPzNr94b0
0ErejxDH93jR8lLkGVBazM7JIiFWcgJGsgYqXA3qgJmaOBLQTEN2Y69cuw+TvSC/+mReKVKCUdN6
L1vlUJf0f7JqcXHzcRqsibbFrGNxUYV+CtMy8r83guYzTXzlPcJvv/asI5j2L7mtE9a1410nYQma
+AbZv+LAh8u3iSknOgqmjlpUKotzYnUhcsOgxQxvtp90WSHqNKb0N8UWOXnwpJk0BgCry/ul164c
PjhLlO7ImUGAdPoQNnU2jwrQ9JD/9UOO73JKDGApmCY/ecPR+Q1y561ZkHxJGQToQ3cItBCGDWlj
sLlNuKxtSUsrPrYHP3AbM7r2/2+3lO+VS9K2BYeJjvyGucrXeyWz/qWkGzHYCSqfwWvis9HP76Bp
NRDkXB/qI1SDzNekQJWA/qB6AeZDhUYJo/O3G5PIMDtYXGk/jiMM0kCQ2eGuinsdGQMFD85J+aKc
fX+rbvRi4tVSHZY8msyxE52igTcjX4KqFDnGU9+bR5uz8zGDXT00ARHJj6yaWUVgWx5Q+3PmDx17
uVn37ue7f81KqOgy1c6fTl2OGeITrT7lOy1Z0fTxqynC0vqD1VkUUDykCeLbJrte4lzFP5EgMSB+
QKQruz8iW366LUt6rb2HWA3SjInCNjIjycNwqsDuTomd3K2tBDvhud2X4XoIURUf3MYMsiGajR0H
PbCnHyIiT6sxiy6Z+u3CATL/r7kS4Y1lSl4zj23WNxoSOTT8W4kL6LZkmyHiERZxQbX2LWSuPBAB
k37I/CXCe36gEJVksbBafRecOHBf26uOLn64XcT/PP0kqOCe333TiLPF4orXHVi/Q8QiJ7SAiYEV
CpX6qbAn3SHhoMolQQOVvfkJMvnYLRS5yEJoARpEoOlUUSNE8Dc8tKfeKS2Vz78WuPJ14CDaX68C
zGsEallOnJG5DqxSElJrRy7X0gQ1hmNBhcJKrp6M+z71LBKSUv/OYGIC6FEvqxNUClQva1pjKibc
o8T+opQug12g8JEAx2Yy9rCUhsk38tz1H4d9ZNOcPPMOacTpMG5wPgsrBD15Wedp+8lSH8zSCdUt
0Wb8NFcAG07AL1aAriM8nnVqj0h9smjcClAUFEGjzADy91VZVlKxRuz6OV+hPAmczXGaJ8S4v3Al
IhQu2FiLCybu/f3bOnwdfOqJzaep3WTt4C9W0kszoTDOd/akwIN8kFEZ+bYOZ49YLAsHUJIk1gBo
yAcpPSLpEmDpZzO15W77Cw7i27cQJJoB73QftwXoKo3kizRQYA8b97cQsIrbqDVWrMsYvAkT2QeZ
BEvPyKjpLw19ctxH8BbuIRFCKEa4MORmypzFbWQfr/tLTgpDwRzyZrRwkOQN1ZdAmp20ATIkj0Vu
k02kFFVFy8geTgTCki/QlycXDq9ayXLrk8AB9pqqPrdKHwi9cph83km7duv3SI1OYDZFsxI7rpxS
Hpl4PNEVTuCZ2G2b7RyE7mAqZLcuVAAcd9kSlqhQDqWcIilNPckr3CZivTywNqZZJnZ5pob/xx4/
YwLGSQ70t4DnfLSwNXy820sILObzslJGpvKLyxgBFp69KRuI89irG4v0Bakc9BNfmHkncXIkhVuT
gSYpKu7cktgbdCzyMTtPDQgj5j9td8ZVHpwrN6TGCRyoFJ/S6slqc7bWusr4BX/b7t/kKcBwBrfj
83L4yqW1yoWGSxep9+Nnz7bg9xaSG6a/y9fEJYbZ5zHhNCvBGjdFNGLDv5JNqh4I+dnopqtdVYUA
r8GADKr1YVuxEwuC7J7rAcCFBnTCCVgIycZVChZJ1M626HgcO3EVLq9QiTmPupcUUeXU6nYDp/a0
3JFUO7HVxlGtirmEheR68OjKNrsN8kfViVsfZ2pwKa6ZHhLqzaGpyylFeG+TppDug5ILdEDirG3s
+fFTQvCoc57z+YY6GYV1HTvMNQBksJRHubQv90vWTUeyz4IDZRKNs6nB4p32yA0+jHOp/cxaEg/g
1A5YeMzc+so2xzl9piGnVI2MnMqKLNqc+6yooCzR9ev+WKmy9VPMI+dgAKrASo/T4x58WRjhoYwn
ZzKkBCcQCNTsPrQh1wR++SDMY96g9fs/xxzJTFjuhGARPSqTY9fjpB7j9/3bp5QwrEd+xJckEt/N
Lg/v1jLYq7lw+f6o+1mXrwCUthTx10Zd5ov2OPT00GBqo/U8kO8Iff8kCIteH/G4/hblAabCKGkM
7tHDWhuvtKGPfresPtUjpLi54PWR+Ap9ntVPbPV5sug+8uDguQPdBFCnLih/gX3qvcQe1+v6SrKc
r4rJmSg9ZVlbkOjPMxT3glW0SW3/Vr9wW03vd1Epc3Am5QJbcXOrq1lgxp9xrGv2XTYYTEw0MfYo
HbrQYlJ6lMdMjtlndKTqBe0LfeS/Lk1lbP7IDQkb473KJneFUGhyBPvpIswDwinEOdiB94UUKi6N
h2wqu6/KLr3t4zIROuyIl49dPSwwH82b1+H+W9klWskWWF6iJQj//KTzP+35ZpQE0Myi+7+jfB3v
PRa4lFiZuXKThFRRcB1pGbkltehxKgZT23V6/VaJxL15ZImXDKV4vGl47l1AY0gG9tDsKYYLgrZj
DxPcVI89fFzRmJZW903NRkBhQIVz0iG+WREu/UMd86aetDMILSGIqp82hSD3BpG5GJqjGSEB1LH1
y6yqonp34BBjRvZxJlHSymMg1PlxnzwPNM50gy5TuScT3AWw51duvPLynlQUicW/Yk1eBnBVH2vD
NT5R5FhEBXzeYQMfHb0JCOUJjram0IM7YqgUPJo28oXqWLLXMLtkR5jvOaODcA9pzks+WRFDMHU4
2igH+iCku6ShjJJYcm+uiDNVctRHC6C97mRH26r+V5iVdr9bIbIXa8X5/4k4L6CF3TF3zN5GnLyF
qjouKQ8rBsleuvn5l375l29b0DDlykpaoyC1MU5Za2ymw6BnPMhaIyLc1FYx+DZ5QLdDliwyb1tF
htdfjYpjSJ5MDMC3KvvsgiSsWZhZNhPRs6c2D3oMM0xWsxZ2so0Zk6ys2H019GeS2h2OM4hHHYFM
+q1xdiY/yKAV4cpo+tjW6oKp1sy6egl37u146y/tZORlPbikf0DFnp8WOLkQcU4DC3hT7uPUh0Ag
NQQDsfTOAvuTQNCYomy79Nk9tw7MnRjEJ43qDuQd9M3ywnN1J89HY8Uq/QYk7ItlITDHOBpPrRd7
6E4f/8/s1yEHS8GJ3xWIu+UW3u+//tZvk042MGyshvjx/T9xeZUi5DUF4V8Zt30lZxUTrblr5Kq1
v7zjbMLa6RU9oi0uH8ySCBJPjERnrlA1EhHEG4VFdLCR+Hwfn+xDquczPIEHHPmeONP3aGQ9LW/3
eth+VkF4hNWb64+eD3cnfk6H3YVfnKPc4SG+jGZTX95zsYs9T7PmpRRpZt+LhFEoRGkvyb2i6v7n
8nayOmDcFk/cBEueZo0dOwif4ksGNJ54j+pTiIZr6ofUHA7VfRJfF/10cLS7hSmRpccTm6ubsajK
BESEBqGA7MXdjfvH5hlqxVNR3x6OeWDrND+FGLe22XRc6h1bzzlt9VI1gl08Zy4qENuUYqIB6jug
zeoRK2qYTjlqhAHey1Y7Gra7g/CGlraVQEqc4myingPNBz9yRwdOq4fGQdNUIyyCaCYgnfv7hQXV
R0cg2qIRcHEo+dt55wzRxODpqII5opWJ92WahN2+PHjhM2C93jxjdHTv4CsKtTYe7imtX4rwpeHl
XI8+CV44OoqsBmpupVv8tcyPOMPyHQOp+81//DqA55tGG7RMWbf6IVasyrSQWUMzKwhG83L9mCPn
yUNFTUmwc3wZ3XXENrl0JJvL5bYjgwVZ3iZ6NubVzxczt4I6ID8YLImiFV+q3q11QN/v0FRnpqHl
FIvvlURNjxSill7ctEjSTLdiCRDdVnuzy1yV9VRNnw4vUItFAj+pfcpisev68/o5MHbe15/uO4gr
BTZwwnU4XkpUyG9VhFZ+wseg0GDjyZqcxnr8UoDGPWULo+cYVoF7EJipGiEU80/Np1jjFxZeRSsa
zAHbcESyBGKGKuC5uRrxrV+hGlM+k4ebVksiuGsAm14AB3QFehNzXT3GqnHPpuKz9XjgNen2z6ZB
hUoQhHRGKYcSLQZ2qdxB1QYYc2U/9JrG4bos6aDpY1zrkYpAMhxwqQNWROp+zciku2QCjX/P1HZG
BIJEoXjxS6qjEOdPQvbGJQ4m6El2yjq/4W1GXx9mq8fwwYgd7PbYerViDnghlLxlS2qvRsFCx9yU
tJ2r0U5n88WpuWL/zInBvBrwRjpfGqgkz/o+sKJuxZot/4PTvGAxZsjbB8ZF0YrOsxPFFHwVwjA4
L4Jv/YZ9dEEu1DV2msWy8+ABwOTmzP/4sIfn23CkDfM1heodKzNMhzn1vUMPoXsAP8rIMhpxySNN
ksyQ96GmUuBsJnNVnmk1jxFGt33lY9HRVUSUZhhhd1q+NsEXcbWcq/joFEUdTkBa5tpRqOqv2nGL
WSft4rkIcw08I65I1Zy76J7G53NGH2/AFhjZDRXPsfSplqCzj/Fi2L93tY+aBPHQkOjxVa8tJ7/g
dSwt0zfL3FOeza5CYpq4LZMfXA5zmw9y3pk321MsN65sn3qcT/9WwhiA5jGZUBAZuwxrHfLngj5V
zJWxoTZnpuU1pvn3HY1pi+Ij7LBB736yBC+jH7Y8CYIUmaEM2FKN+WAWfeJpfNUpgVbQDRPMiFed
iovWRsZkqupIu707FbHxkgrpWe4JAnZQEp80jjF7gMK9hmIsJHAh0b1BAqidmpvns85ve7G+p9An
UqHpo7l+hUpe82Y9YgIO2JKbgTJObBuPaqeIqRO69VZ/JQwqrxy1OPoDIQEii3BTzwCi/yTqB9QO
5YU20rNbTg2ijIhYe9fkgiRZTrtZ8wB+75D8KXbuRBl0rTRmhSt0+hBVVJDlMMzqlvV4Y9esCGoK
Gzi7S2QvVKMGCj8Bugj3LbYTCYr+CcfwfP/TYisC+9DqtZVevt2TreU86l4PbTaArEtVfaaWerZZ
aiHtka85IxKvvwidTAq2poFAzRbCGZNhyIaKYX+TksBCpn9ej6ZSduyOE3dHVgbirzUIdLHn+24d
bjllPiFFVQyp6FbquuIrUoTxVH5fLKjO3hhyuWqJXv4wGCzo1ssKqAfQsQukJDFrgk78BR4DyQZm
n05dRQ9msazWqg91PHEMXUo4agT/+/ptaa0QvXf3z8vH/lwnd4kl6cXr7BbkFsVG71Bo+vu3WxII
D8gMHxSe4JgKDegTPgMht6y8jRRV7nad9Sqd2rajFOXTptMJpXAGyDBrxjO76O3zIe4bmp5CkS78
Eybo7m6gK5qGn5iofwVGRQ1e+AkGK/e4J3Vq8hktTDjtaWOIqYeHuYWrnAidlTcH/Ne6zMo/VENT
a9fpuiK2wvsV7DyqSf2RilFGJqjhAGjEEB1OH8Snz2n0HMd0gV0qw2JCW421JXJDfBgpeyYVwaYM
aHBfwvDdjIiNftJGO7yMEF7kv9Tb8yJNYJj/sstxc5FijryKYeDZ3OwOSb1iSIeBvK5IGPm67MXv
v48IF8EcPCD3szlVMRFHkVodvM7cuPgPKZMN9WsNXxroWMBhflU7JMOtWk+LQd3NltxIe36dSYNf
DGjdBCPRDZFOR+AlI7JmZvHuousE445p5XWgz/nPWde6CVwJbtnygzvuPksDW++ad9AgbCBWTO7y
tEdgRLLay3DnWq9IJMvOx1iD3lqKg/9msxE2OzBOeaWJqfhrnRCWYcQJfngTMkTJphIv1HAYsdbA
BZmr8/6cTI8/93AwNl6rtiNHwwG7Sthf1Dz5c3CpwgnscV35++kx7WOjjOKLZPolHIJ8DwFqnuhz
dZEZk5F1h4q8k/2hhRw5Aq56oaKZvaCn66KceLwA7HMjH4lAN3bzMXBaSJAICHIaUSW0NDBrdOvk
j3J2ilRYQadfrA/3gy4I7iOxIY2hYuFR7soX/qp/C82YdrYBw3XH/RxvTuG4Tf0N0F2mJfg53/CR
xtuF1rAfb+BRyqrDluhkZOCQ2Wan8XoqnRuvSY5cgwBYelJnePgWtBPMZ9GdJW09BKAK4KqHUAn5
1bZys4D6nPr1e3ikt2AtdT75eo8OlRLQEV+LUxMmN0HrfQM9WhK2Ud8yh1VeiDWr1JpqdOrwuD95
X0jWy8P7mVP4ZEPI6ADLyBqF9UFiDsMdwJDCa4NYRSkgZr8cliS/MZFQuPO28q1pVF53JPIv7jvN
4eiRHg5eCqa5upkaHMXaTP0wk4FfsdMHo6LmhoPPcuC4JuSl7isVtV6aFDodEd7nhL98gynVCUgl
W3SBxeWGnZ30spDbT9MQHcIuGH+fJ59AGxVRHhL5pH5Nyfw5HOYcIoP6Sqhn27VwrL19RmMpiXhC
N5P9WYFTY61rHuIjJ7GowK2XA0apdXHlbpUgXGKNB/fCzCtWXZOum9Mg7uu0h1P13Fyyt0B88CTg
KCHE3BP8B+D2QpQHr8MkO0+W7seCVx1f1JHerO3aNmSaWM1kQPenBc1IRzHPTjtVic3WW6Pqf4kc
/9p3frv82F7cpoRA9BvELSokZyB3M5Yu/liDno18OWLKOlBdrsCBB/QbIYalZHLHFsaAGESLnf7W
1/ZiVaaLiFFxQGHa6KENdRrwUk/eEI90ri1HJ6t/Osc4KPQLI5zz+Ey/Yq9+tNqyf/uTlgQq237J
oTkpJfdoNwc16GITjUkT2OanTOSbZZeOfp0VAPLUxECDql9V/H2e0UlOSjpv72nydT++FFajy2XH
QyIYKnh5nUFZ+eXw/sq83pZxaWPD+UwuVfWqvncWn4T+YdLFg45hZvKCaZUGM2Fe308JX3/fSO1n
ghAT0zQUJrHA2zvkce4J3r8ICQI7Dxnra1C8Dmrq7haVEg6BDCeAy416JONtI+aTbwoaibx5r9oI
bFeSo/Akxdgi96aH9Bc+bf76d98u772X0HDDekOPh65G8be8oAknx+UB0IOm6KmtC0bnNOTCoopf
FTNeQu+pIW/LNAo2yLPd/FPOhR2D8FRvATPsswrRewmBvogRIxDZn136KZYtBkXJtavNTItWu1cp
LI6gdoUp1UQX3BBoO+23R9zF+TwL5D7zVZhIDdne2uHjnUj3gNVwMHYaqR4UCB1G/NWKRxGyYqeh
1TUNZNt9UQPr7VRwmmY7W5itCu0SBBNi/brQHRTaV6qrDCxJkOqvVfKjPVokJXS6oHpEejcfKceA
I3ZRxhGAPWTze8L6zlBzZ2B//35CY6mLmbjorbTeyNMqZlepFWZe3gqBGn6xENj6Svp0Qvrwkyz5
hK88zvxTNChl/Aee009PYyAU9FtQT93uR29m2s0XB19svrMdML/sh6FuEOWLg0ueq/zt1MUA4Bmw
2PFJh+qGu+cbqw4udq47vMlPBHW4tKCR4/NnedAEz2Gtf7hj23As7PjFm3MnG4LgKJkwQchXoC77
d1+d3WC8yimfnqa2Hv7fRxS219KWmx+p1cw4DsxJgvYVswY23eLuahZ7nK6VudKovsZ5lKkAz4yn
Nu9+fx2ocAz5O+czqBsoVvaYQWMs/g4KxtYa1itK1MjG9fHoKjqF4OM7wdLioeVClCJU/7ihzLcE
wMzkD+5HgXpfvs5QUslZ/6qwjCvENCwXLFT57M5TFuSRspzvLY1vaiMA/mMxY/YYi/b7aNWwfYq6
EccMNn01K3zxSsBp7FOgMloe4XQq4Rea6s42fhuZKzl45T76sTSNDcWL3pYZUOD5r98hSjHJ5EzG
9r7df9/LWopWLhTSHCkgUx8ZkILyr2X73nsB2D/cWygjng9ssCI9tOhhermlGw8KO9E88qTtVAkw
/XQyb2AQjwVE04UoKUrfP5G7Q9qaFLRvNdsQsAXQSrM7FbzAYaLtPmL9HvL3ejUpJl2Gz7a1g02m
KVxBzyKVE7AloD+VKGDZjjnKeV3w2XxOev5ZVUX7cAzGON2bovVBqUoKmPNW7FcU89WEHfoXOZHb
+q2yYkUPqDFdmt9H9AgdBeDJojJGhXeL5sV+6ge0nAGScESVciDiU+pYTUTn6RN76xviOLuDvXbo
LjbXngK4U9Eb6b9fxy9NEqfDEYZe7sPQ2+OjcakBPFz+SpZI63mE4AdwFyOK3n2aVeH8TcQE8H/l
t3C8+nGDqsaSRA0qjy37Drsfd7Os4VCjnMIjAIhN6w5u0L+WnrEiQLJ4Ht0QSevSn2FcfIkvKu9r
aIu3g+CiewhbBk+MI6sUU1KdrnE14Eu/sYdCzarDU44vm7xocCeN/qMptH3sGV2/4LWKYieVXRGr
wF/a3C2ZeNhVVRPfs8XT7aE0T7XvDjogYoMHjd2xn7AHuRuaikSr6+2e9C2QTS0JgACD1TX9haQ+
JrvbfJUpFfgmGKTQx2g6fwHCCEIrgmjAXCdXsZz+dcKxFYZPgtQAL6pLi644SOqySE3L8PPI0D4+
KDTWled1Iod3r0C1KFiEZPGbcrW6s672mIaKwXOXqZ/NmrB+qCdFsMrbWGvzSxDtLampx3qacQM7
XFSKYURf/g+GwpFVVk2FpdGo1ilqACB1+AG1FHouIx3vMi+Nes6eXHedTHjw9AmJe97BgB5+9UVM
3Onwp6hEp/uWqKDGM6VFA6EcmaC52RAmoslBO887EHF6HENlAobmUT2X0c6wVzkID8DxVlE9/Pce
x4/uZ1hNRFqIZjp5BxtfB4f0BD0TkFnksY1KKb1rpeH5+JPnuzCHdnJjEdF1vrZbzBEG3zAWPQI0
q+5KJ+EVRJrFNiSbKBniuzwpxm/NoWHUHI4UBqHXziQEfa+RzZbE+g1WLdTAIE4eV3WEbjGUA1aJ
yyikEHwvIFyperm0rjYYAJIpYnPFAA/YrwsVoM3BeWzh987oGp0RlgwDcbl7ovKCwlgStXcJFXr9
FkjkIuvzi2r5dMNq/ckQpVP8YAG6+hs92RKllQ07p8+1nC+AzdPohSwaNNEpwhZRlZ4Vannh8RH0
04+Yx5hJok7mCQL0zyQNDDBUInXClHx6BVyaC5WkxfJ2Yn3FL7AnoFiHVCkzkT8UmuKTFkA0kyaR
3jfMIv7M0u5hrWXhHV/NUJd2bN6X/5FRlg564Wejzt2wKIaeYOg9WZgFhaVfnvENW1Jr5M7c8vwY
2RXSBz5/YZC8CvCa2qVV3X1LTUw6xOH7n65uXcx+xiWSdZx4goJQMu8o2g+s8TizTW8fpWAcxs28
6Aimto+cHRrRTG5xLJSc5xR0H7uOUqytlDySeJ1qIOUqHVjGn741aXKP4wI/W8YAibXk/h4x8rSk
6fqkoIr2iUxKY39Zs6O/o0OAIBUHum3IqIAso5dzw+0YBPODWygA63RUhOMAA3ZIhYjOe99ewsjg
MtSFULU+Hqm0EuUOee9gGlMKmcQb9ou4PBaeAU6v9tf0M4IZ4RLwuKv8xBfdBEo7WmNDaWX7xNn8
nrxIXfRD/dXFd3au4s5KonO8WU+EilU+s/N+Ffr6GMiTEFaHJq1wXJVwsDCpZRHyot//gzq+e6Tj
EkDXw1fg0q+4jCEx2++B0kQAQWQqiimtHiqUDEjfp1lNV0o3irul0CfIZPtq19uxeV1E/3tmMet1
DiF7iIPL+0oKv9wfkaU5BUWGYdPchdbC5riTFqpEKAhnzS0S0cdoN5m356BT1zFE0Bllk1GirnW7
xGqHD27EGf7SQn8e2KbDzdL6LRLlODItC4kYc51eq7ZM5V9dJqDMK4NEkeurobPmdtdbk676U8/l
2ZjMaFji4prGkL0IA5Rn7SyrAKgrWFSkntIbYMe4zgMhp90oF5ATP4zOiFDGrCQzVgaRPAyRGGYR
WJiQB32BhIAnD5nLoyV0Bw2IkMftX+UCehR5MGrg2EWW2yvDbnEB0XmfgJdEzQpybultvbo9D+HQ
d0N3Q5FCX1egEBCO9fL4pobzR48pP1O5HoalKDAynZsDxIkd6irO1jRPekZMxxqEQCkpAA8LN1tQ
nartDrZHHV9s3SUHKwYYeR3Yjm4OSiy+Fx69DWw37vmlvT1/LnJ4DCcxJOurCrAQlQY9+QYDJe1t
rwsRjKqu9adzWZAwFrn+oDfFMTnLP71MlpJfP8pL6ntyJ12LAG/PBvTaxkLPTiiPn/HMkaLe2rrM
Z6CwYD8T8/r9elWG2gujXWf0s3GQ5hT9Ln0LlHuSeV4nl9NZu5uJ1KImyoWkXevR/McosUn8pBwx
JVenS4n4QE3CPoD6QRpnM+8L4wH53jDgbEufTxWPTH+yHvCpQQMANx9Eqc0FxVxqU8c9YfYG/Fpy
0ITMSuJjFKR4VUlZ7Rdgxr3lbgI6p2yr8PrJjorkrDffHzS/KINfOImRk9pxlzvh3F1TwHwiPLUI
MBFB35ddW6XJEoLE/9qVPsGoyYRdjCvhijeF77vZAJeN1z1zcwePG0JI9w+d/TMeCn+3zNFwtLau
BHvI9c7J3lkFsJSjg9luXsA1Vl5ivzqqEUXCwIIj0Vb1UyvbjzphaLclF0l6rE2qHDtqhC7fZiCh
kyP7e4H2BleEF9pcvCbds2w/R1WnihR1/oFcJ7UkNYNQ39PBJeHVBqypkQMKelz1ufAIw8mdg4Oy
2rlgke/rr/ky/KLJMY3tT9zuugwnYfMywgmGHMSAJ7FYYg0N63K63sL+av/R/cfUvPlR1sHO4vg5
gqVOrq++nfFqEKdwyb/kju1iJmhFgqMtoY863bajhvbvpMozdt2JFzlJ3NWjaWTxUwoiEnRvKhBQ
QTJh59cOnfzJpWXZTflkPcBNAbO1RC1qqfb6z7fspANtU+HzR6hNIR6b4UDWVBhcqs9SICzjHavH
+bbJZWRLS+AEUesIY5B/0q0mJoEWfkTLKdvvkA1VEynR1q892KkHXUR4gvRmB40TTRk9MTHTd23y
rtoGPi2n4tCtaqWw2kTcgShJjRdSnfmoedGnphu3Akw/IR6qEzhNCNFHDG4+JkoLNHHVMJfUU+5/
4a8E2Edcv3Ayl1STUMZj/27jNn062vJ9YJFQ/M/UF6Y+N9LH9x3RP65H1KIfknc0v4gZpPJeYfU5
nT0A4vvMQxac6JfGehsQQs4YNOGq2MkH10yDvZWT9K93dnVVpSBEJ6kIcKBbf3UivAIoRylCd9fn
iweG3Sq6QUQKEBhlArHzPFGyKC1bVOkxXLe9GQs7/NpI+aMwJw9vPtQlHpXS/VkUL8DLzFPDSvpS
rwiK5akaDk2kGVVmgNyCP8J9ZOKVDVh0tJSvFxdKAlRP8wQty7lkfovS+rUvn9n31UoIjwgsG6pw
KhpZTBSFpJ4xOsAqkoGFh01a1DutO0AegXVfQ6AOtsKYspdkVk7a/4MFRHPIB2m9jcv6CpCE1kAa
RVRjHBIKNhOiPDZ42yjoKlu7wR2NkmNBzvoSlszGHXqJopLElqeF+ZwVwT7XrM4gCDy2r8/htwmQ
DJuSJVPK2WCFxQ1wM8+fJ/ADo4qx9yaRmKUrEXwI+Pf627dF8ZRna1Gly4LOlf2I/eYdWRFlMZEW
Ki/EWLNX1zwqz99zLYCna4SShi+WLTrJWdZZWUhc43YZ8otlgeEIAOwcIh43ArZkf5rCPXr1DTn7
YIPFVnngSb2VzPvTliauUOBmiPoaR55fx+DQ/BjBvCjb0lL3aO9Z83JdRKH3enS3SyBCUIcwJDEx
HxDfnc7q21uS1y6IonWXIe4I8KQNUEcmxDJF5RmFLc9/yovVAtdl/Iqzpmg4g/EuDGn1nE55h/IJ
2TQhwohVmI3ninVnzL0bTscSoxf0tDsh6epsStwnBwH9aECcCPF4YxuCe/eP7FktMEG3BcXq45Yu
EodfAxGsqMicUXe1aPzuP6BmwoxAnR6c2N+aaZuYcdWK7ciWQZNElUVMOuRHwhvDaJlK54d1S9Kj
5ks5Rbk8NheOC3Nwe3q65h5OSA9UFX4IUG5ZsS4QWtpYmeLe1GI3QMiWYgeDFaDmpl2Ifm/SHHXY
kSPHgHJ1A/UmwX5UkwZgpuDpfs7VB8E5BwPv28IIaokh9GuZ5IHBJ6uTW1RewCRb759bmqwfGQ1l
vxJpuVXL7BWLMWEm5Qa6JlYPpey7vcfKMyMIw4VA2nE0/Ctxfm7UsyCknXf7dqj7S1WW5+FUrJGi
ShcCQi1I58a/v1ozm5wujsCRtTf1cgfqpQtu63183KKPjpH3d7bOdEUIs5Fvc00aB9NXYE9i7kEk
fzzm24urTNMFbP8HY8b/4+zMsgGzIDjLe179SPs8s0If1tdkVuNSoBs/zbUwMSKjgk/Gn/ZBEk5C
MWHkDlF0ojLz0KIeOhjmEpmVCz1XFRnOBqjzt5Uw9PT7XvSamPTnuHrRRDBWaaZ+M99EoFo7oPlq
zo9JHkesrzCTaJM5NgLFkAoBISXBM1l7q8h7nBsYPHQlJBSki9ebtbyXPsv9/gqBJzkX0cLmJMdE
o8XcpHvhtuErmmq8mJfABoFjs0nArEZvDZjsP612nk8IUrwQ+8vPi/nHlnLZx+VsnNQucqPMhlvo
sY/zYSLikimpF9+O9GXzm8B7/rEECiXjaEaEVvGn4lyRwV6IpQphYM/PANFDPD5uyf2Ti1UEIRW/
Uu8IyT0VfgPHkLFXE6CGVyE9rZ6p7ztN9vO5YV71U5Y8NPUmK9+0uAoHVAzbVs4SbtbDGrMSg5Ta
w79RufAG028vxo9wjW9DztdmdduN5kIUEYs1KjZYw+KWHz1JzUFSyCgvODKHF9Ejojq9PiS1GE1X
Wf0lyw5DQwKcMvT5LIOnvdkj8few9p7jJJyFMf4sL4k2RESSC/N0tzfvFV/d+tN7Wb3PE88qNGi0
dfGTbOHRUAPHbM8Fj+B2fZafJHVQZJjzp80r/1aBA3T5aBuMpCxXw92N/XSu+CyjGLZJVskqsloW
hWS+rUnQrEQIQOxcWREpZIQPgwvbXzJaLVihgCO9q5L3ZWWJf38zMWiu7w5Ou/CG9a3Ls9tGBrbv
OZiLqMldU2rBKCQ9aD/J5KgdVNfiONUvwip/rVNzoiGuQ/7UHpC+Q7X4YwQ/4rM1m3ezEVtJKLxA
QNQxkGMxdCwhp04M1I9+JLeLiQSlM/q4P/wPbihc/yScQimobdu6b9D9owiURiRHgHdJPzxK+Jzl
BzCyylzzcdSGydQrP4gZlyNaKz+hbWxi0rr8gUNp0ZjOV+og7GZ1zqJiigoTMfDnNcrL2EpT1wDp
cQXV8xSfNRFnbnku+0J/v+q97w8DvOf+mhKsE3v/9j4ErWGKAf+hQZ5KG9pdttR1CvEtA2pp0/oI
PYJ3y+UejO9D/44kE9aJLFB2po9WuJRCz45quB9o3qVpoW/WQw79Syj4VWueQ1lT2jUticCfOjw5
xGdvRURiwcEcvnk+vkDIlL+KXTVMzwVHZXvb7dSbfCMeNhTrQEWHhKKyLyvqqWBm9GdTCK5Bo15M
ShRXBS3KKQptJfqXCAvFEgFrdb2sXf1oVZRMeHwuA0jFYV8aLZw7D6p7sAauLGjD9D0B4XQEucpS
yD+gzbxI51iqd9RmCJNPFpSPAgsRM8wJ6JEwSKQs2FimN5nB3zAeg+1D460snjd3otMC43GblXQj
YBlBoNljKXtT/f09l86b+9rUNVgTwlQlOWOaL27mQA/539WYeAGyXDt04bJDelt+PnB86RHtsgwb
YdnhGTzjSFy+yEwciX399Uoaq9dBLTG4RvR7hnfy7XlXK2a31x4lSdX508kujOEL9sMbL/ZsV9YL
H9LacH07J0mfKx2+S4IXZPEpGeCyt3iNlUtv1rZTCFB6mYLizG8CuxQAoloe5W7RwIORdiLidbfA
30bedsRQ0qlVvph3dNpUkb3T+sp+eKUm0oK36UnvFIeIMzRYGRuOgzqQ10OZazxohvMVFOLp6spC
DHLEnKKZ95t+cqbmx0h7WjPayxdKZkVLvbC9XnvEVF5ZULZ8erFavIlEOLyGYO7Q/fPr+o9hFV+w
3N67QgPxtyEhMKNb0YE66z24jubcgPCGOb4Sv3LYpxVuZNSzgFSo84Z3jaR9qrbUqFhLdfnje99u
147XVZZptUWLnHYsQSbNNBGmDvQnQm//LDYtePNKg3eANv43xNrQc02Xz9bizZ86Yvjey6kTDlDI
2y6BmJ5YXOVzuSfyrL0/sSygakDKfRXhK3WC5zwgzdjYlgQJEm3s79xStU1SLWiI+xdvolxfKhaJ
ZA0NzaPowE8HY7te/rab4QPhhTybRC4WJhwFPUjzT60/8g87z5fHdS7v3F4Ty0pi5lLRZQu/+xiB
RmT6fPuBsWO44s+FkwAuPex19wljVb0ooQ+FBKJUtO5V0QBsMj60p4kgWX9CCXUQDxyJLxmzyXzb
YdYNR7JBcWRwFArga0/ThBYyMDWReH1mPr+8RjDHwAU87hRDBx5MUBIKU+7g7+qdjjtpSSGngHYq
4F6bEGWkWhBYbX/NE3LUAizEBQ4NwrezNgvEHxLdEwhkOQwDb0D4rT0W0GgsaaT74WbFggovIbRd
6YPYaezVrT0hQ+fLGHWVk+s8BqQmNtPu9N2bnDqXXX0+HLCdLiNi6QPX+VNMDCfNb5FB4nqtO9H6
+4aMJwY9lJjneZVgc06rASkTPcxYVJ/4CKWS6pNOwteNL6RjqHmt9ryt9guyb4rCSdjLObh1WOv1
rxIY12OeHYNa2EeB1pNbQ7wOJ9Jx3ZTKqVtevtTRrDsvnF1KC3LZu+5aepxkXGUfJU6qRKB6TeRX
w8m90foUuKXicym+RkfHJYDaVD2RsO5gVumtHEPo/12bo/19+f8G72vI8/c/W0btf8+A94R1UKpM
PObYKDnUqlozLii/GRU08WIWE1EurmkLqN0Zz/nMcjeZk0s2UjE6FDgkqAESsIwgKRr2s1D9FZmr
pFmzZzDlcExiL6OWbLYQ8bcRgeYD5cj/vDaOK+45vODnJfSTymtEUudtDN2js6QEsevQP0j2r+1v
cnH62rdnnWHPReQi7ADrUIOoRMSJfAWb/k4bmkYTzDqgTgi7VvSdQ3l/Ga9NKbsIORk1mPcUlWAl
pk1SPl6V+vskjHPlDny91jBY7MTEGRCYb5+HDBwlfT+WqlkUchC5qjPQNgv6YG+TCFaIhpywg+wR
rpsYubarmFFnx6qvpXf/qgZ20CTWO5n+BQLeU28meuHsbXFJ5Ko/a3HCMzwFyWKXVB0sNVzDT8Wy
XJpsH3wN/RpJi19CdqBjpm8Ijh/8bUeN7YcY6/XLSYP7RrrwvJUw4KXo+hj1X9SXNeTekEBlxDki
Zy6i+kTLdH8NdajbJhWPTOazTHCK0RraXPDmsLs5PoqvR3klRjhiHBqp1IUbDrvDDpPAKv8E4JiE
IBg9YJgOg015ByYZkH5hESNYDuTnVWITHLK8VS1ao0It9qLBDL0b40pgBUjH2EboPtkMJ0i2BC4k
GiuWE4w8AenhZkewl+MWm5LRDibNnpeB11h9zumwwGn1Wm54Y3vnnJ6dJUkaYOI32BRnnBNAi7Kk
oL48O+SBFKbRwxFjF9aN9mz9u40aK2KukWCCXrE/nUg3f923ETnOjFcel1N+zhshUS6eYPOu5Pqh
I9vp0ZKgKcmtu7bT4WL4eHY0fZcNgRE9RXgTORyrokO4V+GZzmDXQUZnMxnmLJQb+D5zhtbRymMZ
7g+bJYQjShwrH/oXDrZmkvkOyGZEswkbIlBavr+0RSghLMtocsFvbBjUv9/Z9Rzf6M1u+vISF2gG
UYtlUsvQflvXrFptyQT7TEjUbydEN6Eu1ncqgyk2gt1dHhLz6aTXDwvbEQNtGksS/5LRvkmhobU6
2EbofxPHe2QUjp94eG+/91a2EOXZ6+dInWukgLh5kQKGwI0oUcCIdFiLyeih8YCvg07hhDQ+Dazw
JMzoumnh9Zh3Z6pMu3VQNpW/z04BS4W0MfLSPDC0PoNsJE+JfSd/itASn55YsQipkkhJ7YHgadSM
gkPrTj4QXxEl+oJj+N7L+PSa5nyK2PHOkq6fUZ5AVo89XRWdJ1Fn3jT7Zneh0j39Sxvfsvt6PP6Z
ZtgeKx9rZ1NANzvNP5j73wgapCXhnagVdXEBueZG4CW1PJBk4unm25G3Fm+qGtiIzm2X97PAqRpl
Pg5C0ONFhjy5z6Q6oZrh3cw7Plp/DJ8mVhHTFmramxox/o45Ip6SxUnzoGYiTcgvjZZmHQktXgLy
ifKIrqrXbvWSkLaJFQGNnCeVq0Zu5GELEG6AQOtxhWp84/VzVzYIUky4/H961PvtjnY/0HxVrLi0
8iL72kGhaEZBEOHe5DjJgNad5dFWy9UPPjthJn9K8K/fijSQ+qWzGDPbyYonuQQayMcaEe+dw07Q
cuE4NK0EKkgA/osOxyzWfUkbX/zi36Pw0MDnDGcKEO7yjjyf/nrWgzIBmPtl59lBn4Do0NNxI7wi
/EXENQQkPXlkCc+/B6+yPo/xtIYyr3/Vxsq+h65GIfS5eTceIIrZYjQBMEWf2ljoSIYM6KX17kny
KMl+ANppBDNCpojF+DyaVKPEwcUBaxtOeivw9NBKZXSdUwRIUocQc+sbKagXJ1fi/TevJUwbm6wa
R2vhSomSm6FeImDc7N5EiIOvuHSHsr4qwHbvFx9lUOwYKz7euM6Cdtp3FABnC06ELSKmJ2RvHcOe
EsOgOl3IU8QRRG4qLMyqA3IQcy5Ldh3CYr+vaCMwRS3skZrsYm3VOczxS5UOilvkuDl4TKlx4WTd
LXRllCs9UC3vGdMtCEPeW4QcTST5zyZVi1pulsQBipjfn/roY01UeoeenrMK9U2AoRnY8okSYSAx
z+hWprRiP39PUMaaC945AJTuf2cN3xatZ66kZGzhQInS316j+Ma6glr48l9heRbFBy6YR9ZgsPnj
YorSGUYMCogHyxj5twvxRrZiFK1jDxd5wXbtW27nHQVHp36wv9PnBVq/101WIFeq4Tiwkz5Xqvhi
leUP5AmJKVsHGjswKxaJdBqY+sNA1YINWDn0FlXzBAd1qb1onkFojH41zIYyhzlV5GJt4IcluL6f
XB7dD+5+Ar2q+XOxKpeC3LFu12Zw+AU3zzC6/Fuv10vAIO3jrZnnbK5hhXTVnuMEkV3fkiNTg/ls
Bi57WL53CIMijbC4MDcEMMyZf7toglvw/HgcwvLfUxRZi9fvu7LgRcK+QJsqcUFIt9gXuXLsWioF
Kne739YjOIjJtEtAiHnpwG/RiEFbpLzWtOz2dDy1EkHvDJb7Dcv3EyKyw3HNqwrRE96Smi54+1HP
NJyI4+LsrzI9fmZaz+c3PQjtfIj/ZdXRezXJ8bQ5R4OJDgOTgtHc7ixNc8cDiMy23C/dCbnggtFZ
PQRVTA3QGpx1FLg2milXhNxk6dsLH4DAMfZd+OjirMCxPm+a9pwxyLrkDwoFhtddn2gwdHcKDgrS
t6ATLxn3QAd0XJLtK3kT7gE3p9gafwpGgzuOiG0mlToM13EJBkK3S79mFTsP/+GQ9fFK3kcDGx40
/hDQNKYKfUh1ooFbG0e5yz0XYMpo1ZYdXw54sXuBNeox9XoqPW8DLMTTRa2wq/1GmpxJ6FRXqWab
fibE/OOJ1kBQ2txLV/0zCHmb1rMD2YqANtZmi/Kmp7573mTBHoW8hOvwc6bXkMpTgayTEjuGHbM1
g8Hyg4ZJx71/6SR0DiNl4GoHrn4kRw/g8cy5IKgXNhJQrjm00KTT2wBaMV6KozhK4P+P6AYcBZtA
YAL/ybCXcxXPYcmmcr4L6rCJpV1IwHrz1Ko6/g/98S/7rU6U1OqhaMJz2/UoPXf8H97Q/Qhf4XQy
UfPoklHpDJgG5WYF/P57BvSPc4okYkho4iRSiLBXWhR7VBO6P+BcW0BmEzOB4w5TGy1dzq+DS+GH
kn2UqGPbSRkQyzwncU2OHN4vlUSOdJzrnXCgyyzW4EMDfjcD7g5ZSCqTKR3p917H8pFJNQ97wvue
w5ew6A6A7LBmm8nFnvn/52j9RlpgtXCcFUWI51SLW7gaqNeguoc1AGc9pPhm68Ryjx3zGf4PHxaB
wvBmv29mac/5EFW0FWGYOCW9J+SX1Lr+DyALIXnhTHluVZwefYt0goBN3tBJvxwuPGQX0sm5OnXC
WDAh5Ie3DwIpVnkJj09E44sZvVlX3EkUNZnsNQ6Kzqg2AeGG7L6Wl6xBL21IGbApko5b8hQXLQnw
lKLK51hWiyC1xJZN+jw3B9Le9jOl8s7ezfDWawy+wCSdfst71BwBwuREld9KkpguUI2dRS6W6R9V
xrbdG7rPywNiAsgeHsAlSk5mbD47y56YzcI5NcIre8k+KllaBuyEa0EJZ+ymx1HPxZQ8xv9HZlPg
GWx253gYjbhCW8H5oJByiK1tsK8TVd0bSOIa8c9twED+GllSPbWGvSdB6q2T9Ge6ZjwDvfi0hmFU
1E9VU+IcbaqDenPpduJOUm7v3gArEl1bmDWT2Lqkql+S7yKuD/SWfOWat3YtSLSwKdw2V42DjGWC
J561LHNnbzQ2oK1IJqXynXfVxJqDltsCU2hDjF8pJlnKOoMqMrB8bD7e5+4/sUe846lB1GREIqCG
77KDzK61GSKuS7kXQAjNblQa0ksAQ569/Do2Gtj+N7x3T3VzmuzeFCAm2jbEJdE2qkLpIJT1I9nv
BDGbnVlQNMA7N3VKOJUVwNyAJ6wuQQ32D1pwnVsVr5OemI6GXq8zB6oz/FNmSP8AJPmaov/D+nB6
e6mj8dMGAY7+a6uPl5IODAgB9QgxnRSQdbUtmNFQcA/1zckGfbQcC1x63gF+AwthmCblKACuZm9b
Wyb+Xa6meuNa0f02F9LRGivTaCDgFu8UnBfPqaL8EAyvR0TfwLnFWK7i5TM8tR6+PQBEn1jCMTP4
O9gOpCXgqbqFhaAphA4VG7zAlqj+vxvIuwWMmILwVRGEC5Uka6EBG5gERFbWgUbHa6sivk//BrLi
4ZkVLaDFU7Jj02jYHRjUMTNllURFn3KLs0X2Ii+r99HSH0OFLG3qaTFEKnnPBV3mIqldTshULIbd
ijV/MRep6vmwN631RnbFOX2Ioj5se5t2/BjicF2TBXatZ5ncBWdmeoOl2+T1vwFaChY81bzDcS9A
cSyUcpUs9Shn0OuMbUOa4y7w7PPdyL9FY2UJGSTnt4UrABIO4mR8EMPOK58prXc72UyQtCYvpUUC
cu6EKRL8mosiVNeSPzJap12r+XsrznnLyOq++n/I7nWFo71LaPNoFHXWKSjCdPp7bmodzKZUnRM1
H9v7EC08MofREN193/n0ZUWBEFE2q9C8uhTjzA6/GJ5z1T4rPgEMYWE5BB48wn5PuhZbyjgboSDH
Otqj1+Qk5jXZewgmtBmJQ8Eml5SuAwkx6bpbZx+jWi5zNhAqpboKGKLH9IxseBLvfZz8i5/5Vjw2
7wqfbRCR0tWSEJoZcsGUQ+Ov8dwIhHuS+im1xTRTYJHwgbcJvPWrhNe9LKRCoAO6EwGFYKZ+8+jj
8HE8l42/CW2pmcGm4+kcbyeS5KJgHebxKYhr5Xe6HDBk746spSjJKAkUEZPc7K3x2RvqwAcnH6kp
zzsLc7z1QbxznVPLm9noMBXOXvb7FwvCnhnRJdfGV0hSkpvoFLD6PBQUu7wMpqIk7Rxx7Eiji9U8
aNsB6/BohvXJHfodhS17k4pApIbIaB0WOyX0UrN23F3nrCT2enersB8iGPzHfX/sGDFdBZ9cy8qF
km0eNKIJ6ZAcOsZWBopTkhdcYyd3RkGHvDjsriHtczJ11Xx3vg7zGjLJavB4CSzFkuyFoD31S1SD
HHSd8KCq8XZx/+NkyY+1Nnw37wvSAQQf5xEzWQjUNhf+1ALXXbvXB1iZkPzxO5dqbMpHxlYS+WWE
/B8oXfzKIR3Zk7QCkMI9w5MgiDK4mGetOpdrkQ4sbdnfEXz91F6OkAppMra1+0TYW80OLc8USBHM
CtqZUPW/ZyTaro15IwUL3QfOMAJ9YQWJnUNG/j2v+Hj3ErW4N9X8rDUiQA4/F8mr2HlIaabYZYNm
fODGVFJMx6e92LNoWX6iWXeypbY+jZOeWKyQPs2bvx/j/bw8KF/laj+ERQ8bet9KEEjsaPtbDE4R
t2KCGMcCHT2b05J7coQzwNQndjSgpUJlAY0rsTfLNygowoiA/f8sMbzim2vpiwEc9PAb+9rUPgV4
OjK98CSKaH0ms8oPIWeezIzts9Xf9vnMe1fetmbBLbI/4l0tDhEU+WshbzMKTOucTonM+6Grmz73
hPnUwixSOia1gsjVB4d9+r2STKdZRjRxQiLalHAU00oCXWgQiZLrqlNio++rbgZXWYJkNyjnGqjU
Dx4dMamuAcbVUni7aU5BdhEEK6coxBhEmaTrNC//bj3K48uuZ7iL1VkXlNr5XFjNrXg37k+TesBX
1kd6xxMFb2HqEwWx4PNwWd7KrmMDSsMtMsfl8gH0zc/nSLznLLUDMQHGkQhZ8VQbwxEzXPzjvL8j
t9qxSwKTvRg7GlXDyQQyqbF8pA7hUyIi0wShSKmurZQSNMlJjCKkTh7C2Lr9Stf0Dr9eb+FZUIbU
dCymAh20VowNBUZNQjiPgv4BDQqN46P64wWT7uX/42KQsEcvk/UVG0BKEAaFIkdgLsJmUWoe51bK
ZI1j8LXC4EOI9Vs03Jm/4ysLURH87L+Kw8eaQ6O+1jMrqeY5MTgJYMxsl/ykQXK4b9yXH2SkMLR5
ln1+frdCPmqCFmx0L1xk4l9H9gIC6PdeK78gpAZRubZUJLMrMxVRinnT6IWadRFgDI/sTHy0C3jl
+R0uVos6Ix8tSQCts9l/9KNDY2mmXATNVmcFvY0y4IMeifMAmTwydYytBm1O7kjlWIAo1pFS3vDQ
P55mTVo10baBS/WRCrcFF1bxfv2mM7w1NdZKXCkl6ZKz8UPbnWEGS0cqPv5kw1sLKznHJF5stpnM
dM/z4pe3hOjb35MBWONxc9g5fP9VOz94Se+eQ1ERLK1y0Ag3dLjVFdo3HDVYT6nCddVPooR8EsNS
o6oJW/gr2l2OgRpmX3u4sE9UXg6TUUKOpiagVnqUJxGpMjYTpPJO00O1EOm9gmid6PcCJqiGhDk3
u/IMWlgvnLjCXd/bJDwegqllzivDtA7Nv0ygSDjuNEERbFSY7CcvjaBQX4c36R27Lb9ASD2GQVHs
Ft6xcLMhezPoU/ksWVEjZXt6HnpCXRloRSPn3tia984/jTKovWiSwmQm/Iq5USGbxc8dglCWEN2y
lw4wU5TWhkuafB0mPt3HXqhSZYh8NWcIQtSxxoQGdFYwg1qy6zaquRLW1lNJN8uiWmNDbSgHOzq1
uciggFcmDZLayLkZ3BT1cHjocXYE2HS+bYpNB3f8S1guq4jnnjsZsGWlCKB4Ey9cCybwCusBYM2k
PxA0WKGPU5amBae6BjLWq90K5yQKV/0QEeYqbQqU3hAE1G2MhyXQiNN4zEf8mJZTbZGpnLzO53pl
XjTGf6RSq5lSTzCFcAakiswBbPnF1r3Xb+Mi6ls0qXQyQzZjJrC0mN9bjfMxwSvTHBYicVMOMNf5
hBOIZPc3/R6qXjvRIgBKiAGuoINycH05p8qqPxSBwHdqXpQSZOthPzMDRTCylYvFOo+o43V5+TaV
YUtNg+EIeIihJUvZ/Y5dwj7ceeqVDB4AcyWdu6U76TK+6bzDm9ZsSiS3AWfaftFNyNIjV8A18tT/
4YSZW0apHQvhkV7hX4jeXZR2oBPPYYoafe6WejQhCpGJ3QEmp9DD/LVoE9b8S/abSX1e9oqt+OAN
kfa+/mDE/2hSBeqQhhVKCFZWb+MLCGvoerUlO1eDdrtYMghFEJ1tTd7KkE+EeY0ldXl3cWLLga89
YyNYxzuCXactupOOTDVvmjudK5pC9cDlldcgdTX76cY4Kn03DmrMy9O5G7pGWE1hES1AcCdHbmGd
xw5gFtKyiFhwjIAw5U35vNmbPFq9huhno2F+MiU5YuF6DebYIrj5uUWgWSehsD77yI2PtUPf+D4g
RQI0L0O0Iuq08ou73UkK4NSd02HVwzHjBcuxIevHp0Ba3V7F7EVDuFG1h4rawevfwv9tJE7/ExBU
HNbFUKHI16ZYif7ooq6/XmthLiRs/O4HYV9qv0O55hGs78M+GDbVoxUjp1PZ8H3+msRBPJdKdJXk
zrKYH23q3migA0QbHtDl4XvumgsOn4UN8+0gDwwBsmG75yVkt5NMlwQEkdUFF6ztxiuzP08w3Fvk
N/IDN14vrtbj6U1Jz6Lq+Qo/6r8utSxiXMMH1DsB16sMLxfyTtn+BeEiIdIT614RzdFK8cOW8ylK
6mzWp/JMEwLyjvCN1MAk8awCQd3CRLxFwbZo7pafmo35FCM6dJRnae//Cn6NijP59E67JadY0Z8X
TjjXO8AsLdGafztC4j5pTPVlO2BBObMFx5txC0YXxn6RpML0NbN4hPZRnzfvFTVjGsaNhwRUf08p
veI4V8JswJAahvYLAnCpdrtxl8imwBrIOu50QvY1UMdhn9bazofWSnDjJ9rWF+dsWG2q+eVqp7//
S2rKUb+MF6Czoj+zyL5+IwhQdNGv+XR6P/i+3MO3FQUoD7BY5HUe3C6temo50M27dFxy6FRWUscl
flN0UzkQveRD5HF0A1UpD5yQgFO4tKgOWyzKFv3KKlaLJTgwZDPETzX2HP2W/XCqdEZ8BHssKHX9
WrbaDFAckR/i0s1RAta+9ZT6l2WqyhRX7KkciW7l547QfmS4ZYupLP4ktVM0N8tJTXKv+PPmIHpJ
o/HYhK+HrTHI/PBV8La1N+9P/TmA/sA3tRbfYDB2O+gc1yftrW+9QjSr+IVxN+ZmX29RmQP8ymun
GFG+Y/KmKkrovzUJsyOCz01ULB84ZQeYbyeTR87zhHT3QzXPjccyj2ECNNb3eu1dEO4kDHJYG2vZ
q8CNBlNUh1gxDq6Efy19ICYsoFr7ZhUwHVBddrAiv0l/QCTZgpoYbAXmrbYGzOlfmtRU8YZv0wO5
A11NtqaqC9ZmGmu4aYlMA4ZX6Iii+BG3ojjQp3e2RffhYW9aPnyMjBDemlw2yTdjqQCkGhhYrEtd
JTMEaZChyIgVosHxTVaEottS54IpUMsVfmPMkmqYHh8GE4OZkglJUmevlWLQLpZLCoPcYZd+5SR9
am2pGUNKgRWGFYFqa8gcoP0JibgpHeTAZkDMnWxROR/ug32vSQqueiQtsshdY7U8mt2mVQtDDWkK
L/6MMMtr5ZYyygGRvsavxQ3/kSQDxMOtnDVBAAmKWEpydqmJrIzj7r0cphlyUDehZkF4u6iGlrCZ
9kGIy40UVI5vQue6YV7+1Sk4eFvSPrLh3SsI1saPVC9/wrSt4QMt/6bqLnSBAwGMzxqe6sU0GnRj
ATgJED7dys79AdAAIiiwsbn9UKVOGtmXxmEQ7xZuOufrYcH5X8OlgJf5+HVQ5wQ6x6uZd9qEQQ7n
jZY6+EJXymcuECxcB5gg4SkFjPdYbSN9alWUQ0+vTHugVUfrMU+sZd8UGw+5jdpQAhGMEhhWxlbE
9IprDxSILETU99SJyIvkOvyd2RJBVHKuVVsP5Qne4Xp6pgp34CKLVOq37IGea+gzp5YZoGUpilye
dV2TzRIxzBVc1MXB/539O9P2EWFoiZ3yhCezGiF3mmevkUk5eFFDGuFKqmSJm4+HMzO93Ow8auxq
IQA7OXlF2ovTO4a969YZ5AlED/3INb8We3jxC4xvUVf4HiHPQjy8vdtiGfcaFXUiaAOdk0Ih4eGd
3t1sccj7kEHqxkg3y4cz2mjcrBU5cXVc4FpfDh5wHV5hYcBaZkCGNr6Fj3enI+s8A8dkgY1Rog0N
1dX6/MH/YGfu61vC/EkWA4gIkscpkYI1QW4LWyUjD28juzRIs7trN0jK+9rfo4A3hMOmFwEYij8p
TLm6DinerlZkF0MK7cue9om6EaJKeiwF5ZW+NR/H/mEcKJzmRh81yu7psrlaOHqYnirK7bdagi83
IWpwHcNFOEpmIz2N4uoALZBxLTo/AL1OoGqY7LFISxf557TE5ha/JJH3vnpxATVkwG2gwqh42k52
o26acvUcObeGILpZcavXweY7uSTjpIL4mqddj5S7SqCZNk/6Abv/SMBPF/6pb5mt3uce7W/TpgH+
m1T12ATnkQGTACgDxVaEbo+ueWOqVY/twhB1dGsLBXvycn4nVGeO7znQBC5HYqpLs2R/6c+PLT3G
8APbMDVANJfHOzS6RuYlRtFoBIpefdCGFi5YNE96I7bzLOWIX1ke0qem4lWkBvuzRaWSMuR0yYo/
9vOncnofe1gVjOKWhLCJ/vObDO3ptqrLQ9VvM5IYUsmEWQ1PV6W/IxfpD9KlVI2fd/cu+ZEBX9O6
fMCy6anb0mWLQV/A6freTyKOLh63Tm1cGbiFLQMEl8JQRO69otPfgj0nyttfbWRbtzloPpnKK/w+
R8fGCZ6+vmzHPXmcPy4Ch/wyTILFGCgYxLTyRQN7E4fGaZOCVoNdH/jHG9jVjljd30d+xzhPsP8s
t0H6SVNVdHWzw/M5NxXWs1XC8Jl9ohvsWzZnHAkFG23tVXDCpLlpPnGNcIgTgneUWGl5p8rvUao+
1ovY/Mbqjh/0NlUGoKEsHMA7KzvGjU2TetbBqaqTBaRP9vOnlGSaem6WGz1Ya4XuooKbc5ejck/D
zy1/Ql+L3ohASxhfbHlm9C7q0HDlA7Cr3boFXxfI1NG22HSqL3Rs30d6PnJ5U6UtfzOkMbcEqPkW
NQjf9RDmt7aVyOIV0q/hDXxkv32iOUU8pgbw86LfkmGo66mr1ioDxQRb/79bPrs5yCzd4QB8eoTC
HE/P6JLNTS/1UJfM9ORPJqJ7LTVctEmu7rAgLdIyWZmmxHpMraEn9wo9hsUUFb4j+lBVerE7wGH8
Mxnhdgy5CKyhuoQP/2xV/ShrWPY1u4LNoWQtfWo+TT6/eX8PFXg8sDZXXzkVYIP98u8+6evqrxNl
GqpYF7zFElR0974zI6vSN3pGKz/PMkknsuJhtit1Uv9Jcl0BBAcBuw3imHw+Z7MeK+vzsOZUzO36
YVUdbGlB9ObqZQKlDpfwUQh9V7+H9p7UI71W4A7C14AMuyaUJMYSrrXHUcBdjW3/vlg+07TWMDyj
dqDDCByqed2bNC6aIDC+A+tIeqb0evaGQEBDlSD40hMn9aDWXwuw9k9p1O1cN5LC/nDsLtKzB1ex
IQ51jQTNkPv/sgPhgCZol5mvW3QWVKqhMon47eKavFKc93dLMGfwNwkZmq1W7l6OZDGKmgnPxgTY
QT5f8DOoh2GJoVmGhanvGgzX30y8MzSSQ2mFk50zpAdkdHbom2xvd7XmyxTvcALxTYlSGLGB1ylW
eyo4J8enFdzaAwmeGXa+oSU8LYsdx1yVFmeVza9TMQ64OStoJpFaLx1tIacI7MbrqR6nnI1zjrY1
II5EcQxMLPGvvdiIBl5Df9JYiuhQm33+V6u8pI02cq1n0KzmtcP7cn3IfJ/L33WvXEr46IynEXsS
CgaeZWM9W0QcT2w25GiFK98LMJ4HT2e3QQPw928g9CfacovFLA/GMlBFRi2fEODX1vz+aJ7MoiRm
HgxteBJPNacwQEDOuwVg4EkQwPcrWxWQvGE7dHlhcEA3gCM4YUMnX6auDoFQm81efh+2DL5vFfd8
v9ESsrzt+c6J+YujCqUQqZyapsqd2vtS7vxxVtDEBxJtLEaegOAgbiTfkIAjbpDvpRntSR7hwsi+
9QBKr9YW8Z6oKlsDCYAqfatH0V7wzqmGnK9C0DEfY4TR9I+f0oFvU9i8jLDZhPjQG1RiJB4AINDV
UbwBVzaS6BS4Tt5U1gR8tIUhi6Lamho4aK905eHlsju5AZvjslSoqqLl9q/+xTrwIGT+u1aLm1du
5TbYU/RkcVpnOwcfCZqxMTKcxU4+aU6+wtmi9R2KrPV4/8RUf430cdbyTMqermcp6xSmAmhCh3KI
yAYXmxHKdhp5iV5J4MQHPtGyQHIuoQOuPAmeg+3RuWUb5dMdmbGKbpEz73Ew1cnxTmDkslvf/Rq2
pvbayjhcCvVogpfkpxeYGDw06BIKkJXJ1nOCK7F+xN6DLmedb9ojJ7DqOjWKuV4Zkcl4Pq0AtDvZ
QQv76szlPrgT52vKM2VO0jPwKCtjKkMMrMh4C3jes0r6zXsOXa6gPRvFKUA/IXVsmx8YDOTlKJET
+IOdMNXNHoaALVJTTguD8koS8VwUyhsWHnUattUgaIGvaIHoVFLzUC1cxSmfVGrDS1ZanlGnAjPP
XVY1e/iM1yyMb93paeg3kznq5Vwl+qt75QnPNkQOZkq2XSLPq5nvoMPBHfwcCfJmjUWiTXcnutW9
8BfCLydQKn1iqaNSKh9I5CyPaI7WNYoVQq1jQ8kzvlAgc6nFH+s8LuVWRP3vgGJUYJYob6ZCeq7C
rNf3RjBc7bpJZ9zd6ARIfKBbCHgOyCLDF54S6T4CIV6A7PepadmF8mS6YUaTHDai2mnwShVvrbUF
0Adi/oKODowI969G6CC/30IR6ZR51/IW3LTtqnKO9+FdV39bsSEuNMKgD20gtT0gXnH03obfeH0m
+s1BAvosaxtyhr8Q8avbb5COCF0IHiBWytJl9CqqnxBEt3Ux7Cbi44OEaXy8y8FQu0tLdIx7GQCk
6h19tFkgcjZ++1tOh/WGDUew86691Hbi5wVzJUZ10uGjmPUcFntns7e+dd8Ub/fW4baLXVvNTejY
GLjY3ryR0GSP7LGBKjyfqfKrJNb6K9j1v+T430GCDfO6Uzy2Hl3o1viHQCWcuEhyjOYmA0L1WjpY
yEUCXNmR7dAy657qn2OrovhRwhZUCSVKaMP6POJnopJbDISztwlF6IdlqmwjxQgK8nD3CSaLB1y7
jtgUzQeyT13NAmA2FH711oWoiXmqQPrxuPZlh7vpp6yOIrR160DXjhvYxrtQsQwCcMD/+ae4L/0Z
FNTQVzOzM5NyN6Q3L8OIdwr8ucmRzS3j33oHPD82TapluWJXuj4gV5zBR0RiPfqqW/fz+x9uKgnm
Cjm9JcqZJYLeHNrO8SxW7JJiNoJSf6mztuXPb9XBIERUeKtePU4r1RYnK5XB9ODZV1bQbU0bsz0Q
A4wRlQQcgUArNTN3PJ5vYA9ypmfl/vW+9FwtIJZs81NxV39u6fzF1dCEn+g8fqpU6x6jZkMcFToL
QdCd7TIH9pwLyv7o6VSLMIsBn9WpMvv0U/+t67ywR6D4h/XZupq0eWb+dVWlWVQJcl3dhVH89gQp
Hbh5ZNu/INMnsQTqUwnhMC651XNCHQjrCbMuzrLxcTp3rsklsUzzUZZNxiDOZao0IhsQfVcjsEEA
7jeOdc5iRH38vDtQUEP/cRjFlH0LfC3kH5STlSQFwfW1icYMXwKpIquMMST36oWPQNLq1FEbQs3F
i/7+OD8zIPQHJ5HT9gioygtP+OwA+v0LkhxP9LG/fI0iq7FLPLcKXhQtmsb4UBQkG8tBqAB+HeIo
OWqHSZ0WQDfkM0qDAJjgYmux5BmMKDy6dHl+Eb/Dobp5eWaSIAGuv1toz6lUjIjG2retOFfjji4X
t0JKD4uttZdwJQShvexp4eNJ8RR7WlJDckkaGKTO7rTdNdMo5H+RN/FShsSrB3c3CXQHE+CxEBsk
WpDTazF/NoQq3oheIFCBiQ8QJKp6azplEuZ1KE65lKRGe4zBULnk3r+ymUjLN/Q6l60DDipGoVSn
Utm5KTNCxSVlwtym7byEohdh3bOZoghcq9qDy2ijOTwuBd17mvbu+9Vf3Ag0cuzIQiz10xRLXYYR
R4q1bXz+lINn5VwYMHmfNSUPJVVqQXwINX1/AuKcRTwzCNGkEteMZ7zgLhumMz7D1u7nLQyHvxjp
vpojo3ldZ9uKyyyFX84Z9mtrKGBJODGL2Rn/Pf2WYCBAv9O+LtL5H18tm9WvG5tsKYOhlrB4d7wb
/IZKgAPnAN0Pt7Rh98sBvwEsG0HWvb4GwOb2zC/1pQzCQtt4F3dQP32ydMW3GnSyPOeivl65T4za
IZxYh5ETUU8mtIWu4AnWWrJwM3n2MzVPAPXjwp+f0MTf9Krin22SObkoDM8/EBNadvPvwxPTX6US
lOCdQ8wnb/co08a8ByfcZGE8qNEk4HxmjeAB43t1kFoFZtfKWwpCXvnB9o655uhR/vWAJqu6t9jW
ZcmdGFuG5mXyNkQU7Uah/00ChwFk8jAdrEgUrL+coNtZZlRbpwl3wjfjmiECe+LuDsdfJUR4o8E/
X1CNDen22jlxd8GFzpuKtMF5zqZyXYNzuhNjmgfWBRN8h+hFcsvTqymoVAySA54ULyA8n8pVzdd8
1uDpWi+CDqCPkvj099T7b2K0CaM88mX96w5QhTe1ybQVqJuDop4BxeUP2S91VAss6xQCMFzzyeb1
37Io3Pocpqfq91lOC4NBTRzW8FoMcti7J5Rkl50VF4CJ+vXyoV2Yqh2VKFL6YYwDJG0CL/5KkRvV
q9ZDbZFRt8tRsXtJq2PgzU8mQMgtdJioQOktuq7I9DQB0XA0NjdqRo6g7UFkkqxwpwwH+Nwf8qhi
eVKjM6tCUO2QaTh8oDDw8SRC1yKrt4S5a++/9r83gWTGHFZXeGHNr8bCuZbWxVsWnlSPOUgT4jJq
BUG0NQ7WH2/mbnrYRN70njgth7Cs9uMbJJJ7p2/o1nR8Mq1TIZ97zSFUl/ulqpEzA/HskQFY0vBa
xc85omThcY3HGKajyrmcgsJ4LCdLAq/t3UCXMAH+9XrTgKvlFSzisypErdKJxQ79F6UmoQsiqCls
IdgtljWxsudxGWv5jYcoWemxy4jzaKFixYugBvt6eBFWArVGD03xnUxW//9dbDQD92KMKQdwgxt2
uEj6i0vrFwOCuWM7XFlouMi/SZpTeAzXjVlZmYWAcnNdNrqomryH9SBnmA8Fz7XWAcufZOlTbx1T
b5KRBE95nv5XHUjMne/ehYMZH4q2DsSsOV0MPVdCrBPLL5fLl750cVM9tyGeEun2HD7mdHItTGz0
Ljf+BKFxi1+RkWWDi6dqn/eatx5z3TwdPS+lFQRMGvJ9PDTq9HvrXTyF27XnK/zgDKvymdmWoOvX
GTWGpwcclFh93pG2e4F+Qv/ZUGfEyS5nODr9p+UpjsLoWGfsTaQnK0tknVa2xymDe7o53ZvSwp0N
b2M1jVqlhZrLu3cziv5Q63O8Gq/n0pHx6YKFIODvTjj66a4dTvHq43A+oJh4AmhgUt8ZZsEIx9by
ILCIpvSzYu+stMHHnocNN1qW7X0la8dj4hoDHksb6dwNhKjxKIJVbUZ3bkxBhtnhugBTRzns+kr3
5TPLgmveumTIhcNtdTZw1UVZ6Ds3nZSHA/GvpenVmcKvJoSQNf1LvKB4nYez7vidmIUGEMeasm5b
skgEXIBH7kiYAOGe8YcERl8MiJE8Ao+9IPV4zVt6+0ce9/MNIWFRKcPsZqJsN87pHxbZh0khTfd5
5CApm9ZJyRECYQgjcDKFPYlJ44eLthEush38OSA5wFFWPPq+3eTHsbqeKuWNPjX1+AgjkoC2Q673
RwOI+DWmhjOXZhIM+PS/xeQZqviYKCbJM74ck2kzI3UvIEwFRpGykm+/lp70vqKIubEUYIm1Dphv
Gv1SW7zqpYcj0mhoNg6at7iyPwquYVPlblZvR4wJtbcqoGTG0TLFaCmqpXEf9Pe5pdnrZgni66GA
On5YDxYYVdBqGUyjL4ZpWyCc2/99m4raV76dPdEK6DcKXEmfshA7Kjr6IrUfi6+YgLWx5BbrLf2B
7mn0cSgnzVRyD8IRMn7vq8BlajgW2SvqRVZ+t0rJgMZ6Md9myOcbuaDgI2ynt019vKBu3Dqn8uQD
zU0oOm/KYGqmYmTF3LX8Q5kFMACzBgG/apD5ehnDMJCJQ87Rnf3+wxVwpqsAVIwZQOKLL/KHS2Bs
1c5ULHE6S1Ud+Cs5QrSKNhefe4jXtGTsW2ANCsEFd27CIG7abv0eoW5Z8TSdXZWq63N5LFVo7rvL
QfAupWW4hvpOjeidcKZn4+qfpGvJPagvYOcofnmJwHE5lI8sw61JXCWaWzO12pZKQoYc3SSRpI6e
GxhIseVKX3jHxzt10IZBovXshjOc7kd68n6BbJu2iwx7bswZBOxw1qnkyuwAmUq1bSQZi+4HQBoj
TnMyaf53Bjloo/Y3TDabjIr8tIvkEEs7J/FcQ57wR/c3woKliQWSpf1oOBgIXg5lFlv+6ym7XANm
k6O0Cj/R/BKtdMuVtOHPxqFcB+9xpGX9w3gswJ2XlD/I0LypNCbq48SmizEJwBEhY2e3xQU/7dOr
MK80x+bIezdT+/nFJst79x5iJI+sTrevEayaHKv5PuQT5LMMJ1QpbfjPy5rcJFVZCv/mNMKkZmmw
dJoBJKQcLiVz6SsaOCqqAM4q5PssV5JpSCM50nQbrc4oVprL3L5b1tzTpiyBCa/ai8kGTPFxe002
xK8NN6M9A8+qN7WqcFoxr6ebjOP03XWVlSGgo7RdSqgFRJMSDP34u3K1MkLwVQP2pqAgH+C9UkAh
ms6pIUpXT3136g6jg+qQ5J5yGbLr/ExgeFKVp4kfCv0+7a7lGp9TE9sUPZ/86JkhYc37z/HbFuSf
BHhXw1qutjoPUVrtZ5B1Te1bw65or2K4dfjYoWhLI9Pi2Cu7ebPwczbBWfLCuDtO03oWh+w96JTY
Wi2z6ic8hykGEKfKWM0N5H6jq0YoF+5Sngf/MrYxqDuYz65+lWSqEEEbfRDtbpUK/tB8Jap2RWNf
4eg1If6PsEB48GLwHPHuZ2v+ReBBFmFln8hKjWbqPe18XY8wZ24To321eaYsjcp4XI49dmaKGIg1
uMrDUQM5vqbvN9GOsH87K2FadE4k0cH/5HnVJEG/wIfOEb07Ys34oqs7Hx124SAhvcnN8pwFYQIs
ASNkTlPxobAEzgRjDJ2aUib5vsu+pMTPEKZs0/2h+2wIKk1C/dnxIMqXd8EKC+QPSP8GF2vyLWJv
Q08zOhDocVBsk3tu1NJDC+TF4QrHNW9/2G8EkaOIhrVI/d1UOaJ+Whs4uD5aBxmK8dvQ4Cnl6sGS
rJqfcyNmZfOfzpiOF1/siEWtCfQp3ZnGLlkp0rNbdUWB2DcacoGi/mANsOEFHvIiPc94MGZlUWUu
bfaZvoX/Rh67EWBDdiH40BFLiO4UsGm1aGA0d0K0cmzF7rFhqFfm3FiopsU/9HEKfsDlAtMxMgEi
OEHVfiKMFIIrBG9fLlKOaL7SfwRLgHUhbZPvyOzz2fpWea2YNW4XLbbIHnESCRts3LkYnC9FopRB
Rk5LDIt90UFBkwuaQUQYdy/gaVaWNYyUyk59MUBL5QxlKdT9TGaCbsAAT3CjwvePFwOnGEdov60i
E1pMv6GS+qNjroVH8bS8R/QTS+ZiiedNOQMxn6FpJoOssyU6tpZzp7aJ5snRbKrEKD/XUh6GsmBu
RRa0YmsankbEIcDuKPNPR1OWuvXncoxUwoSqtg3/lfLb2zxA3NLUQjqeyy4zWpQaGwgUCO9ZL5xH
1VEYCK3T3rPqvPS2qDa2FczmVIOfN6pKpRy+rdNuDc4K2zKKiFUkk/gzdvBba5HwVCrILbYyNqD+
MAmRr/WJuzLFpGn9PJ1NkfklMO/US1csDaUJPcc7bKx4iFNrOUZzRTJLcbvTwY0YuYuGjkgm00+1
6R3q1rI45r4Sz9V7PbBJ1AB8RMs4Jd/n2zFmCadke/EwJy9koGfyAVTIidB+KoZz84E7M0JrE0lk
dL/5LeH6zHRxgmD2gNfabqQh5bs+eS8VbuN//g4xXr/DePls3/0ew1aubFCB5+G4OwWUI2TZEY5c
S79LphWJC2z4XsRYd4kJ8BgMwRnea4I+wx2HvrhfXG2/hJByMZn/yhiAw6yVRYU+6lcAYRGBTyrV
IbHTiS2I9lIPiqBpyUqzCZ1io7ux7LfRYS3/vntG8NY0rgh1eG0mUV8TSjqrfLTfnmhPJBlj5mg1
rAv+ZmjcEc+4zJW5TawuFmcoYNf208uyaaZLSIksv0ymhm2kJ8yhf3D7AdEMUwT9Wtc1E/eA0yDy
BA2LoRBxVUlSla2EdSnSIjDXTvj374QA5O0RbIOgWsHA3ExwRAXDDUXldWqrFVb5JiA5IhUt7PMP
NaVQgZDj0tfACiwlPnXbofvu8UarsG3G7/Vp3OPu8B3QaPtwYt8KyOPJKbWJ1vzxpM2yb6ymVQtB
RrcXMyeEvYbjdYKQE0f9Yz+B/W0XLvs5iLZmQ/3UwrB7849Np/r1jP0C4n/MrP0HrJx8BaVqJBg0
eyxejuZ8W0EQaCWID30o287upk59nXt+1u0uEgNdxx+CzVJsgF99re63MyKyOShlL33s8q/1e6Fe
zMWqnsTOsUIOVYfr1yFGJCLzWd30BtvmvMHWwtNzWlP7t0PxZsb9/sZU7gxY+AkTOzCiwdc7h8oi
gv2kcPmj/67mURcGWpa0yHz+BJ2hgrp1FbjxbkYFv4sKSANUTDWiEtTiyKyRa8daylW2UMWUGp/d
xm/zqiaECsQW5Z9h+RGnOxu0iGFe8AnDn9tqjmYzvcbsNTs44rUrkFkepRmjYEYOMHu0/+qes5Yk
TVUxHV6YLsL3c1TwiZ51CZBvcYo8fpNdowVP1D9KWyk0njZh3f8pXI1O9Yp3mE0JD4EM0tAwC8Ef
DoesNbkUphMyWRREIWqXidMfwONh3yzETUSqDWYZD/UwzUy205DfLAN+zmU2n4+R+SVDzDDNbbpP
lF4QGYCbwMPxG03dQUuGvQL+0jMKk7xsxur+mR8Rj+2bxJGC+8QnwVaprwug2KuiBl5vW4BUqYW9
55F4kiMt6ukSkmeBcS7//kJTbKGGkaZjfGmQMvDRLg9wJ1pS4igDYIDsi4RXzb/eBZq5o8g9hebl
VFixRRVo6KylR21C5fSGwLJFDwuFswkaxKymMozcG/s3YKb3uTTLlsR+WNFRLx2mFWmmXMkyUaYQ
hyHu15PcKolOFbEz/d31k+EgzetJVhTjzNh5LNo0dfPnXfcMKrmM+Ip6Z3tWpAafO1KG+4kCuBfa
fqd2UTd+3OFvtnIuxfv2jXjNJgtDW42wFVQrjNgPDKOsxHs8B9aqzz7BA72HYJQQg3Tx7kJzDXkh
4FT3FCHYz1yakyNAADrOMZBynLkDrGKrI60W94SetPJT1Dmz+eCXNC0YFaL0P2feHv/xLp1e+wFO
9xfoazGx0HwtxaMXshXy6hroiabzU7CLW8OOPLc4re70hwybUWxTLUZF9gGLXQIiHWgRwfHI3tOE
O4sgLua6xe3wsoqIrMm42aeiHWfyKnvSdDRD7PNwc/9OZnLg3mOzKT8bEf7XBJWJ4Nj60idup7kA
Wn63K8Vqs47XOykLxU30XWNegBpFBtZOA5tFSxYJm7vQyoYVXiYOM9AawuMIegmx3xf84H/7fKkt
9/t7//CQKTzq37mIUjHUe2TRXuhnW29a6eS15svWmlAmwFT9vpxZuxraZnG10lhJ4IXG5iEReX9z
J3+261Y01qQf+aByTb89ciYZZ+uTWDwa93esXlR2Z4ZWh00VOlBahQmKYnEPn1FuIoN/U45lWjzn
KhXtfPG5uCMDHNFJM9fe8q9gJz32Sit0lqP/zvrnY5I6zczpet18jr3eIGCaFMPdUkIaXqBntoE5
u4tlNHo/ypbl6dPYGpMm9esylcVpI7SveR47Otev2m+KGkiSnw5Pd+u/ar2Nj11HO3uMtNVZzv52
ZVjiNZ1QrkBcfcpn8y72HhMcnPHc4ekOigA36czAbWR1DshZ4jgb2FikkDOHrjMJoJKwBROYz9x/
3tnrMBxfsGtkrmmnVGs3Vx/Y2zLpXvaXiPv2WPQKGpkG7hrft5W4q6H2aU9axKRFtmm1hSBR3bii
836E6/pI+Kw7rZQcmQtOQShI+zMsfUjQN7AQlaBeobMMS+WRh1yPwCjxtxfzeRoJE7kuGRP+9/YZ
hh7bFcqQVrKH1+rL3vsHUSuF0JpvbeAIGwWAlMjfcsS79J492BpbR6H+ZQ9zyJ9R7tXAnV9cfR31
d91Biwv84xUrTjaL7qPqzkU+yNbeGwYFzcLa8DCnroF1k/NnQjKBJqpJkYHF5/ZG9JRAabKdWzgX
MYGpZHlSICFYcb3XSO9ZCmx/P+dvRSFJXsx6Ias1UR47I1x39QJcYtQNoiEUxfvw3wvslwzCStOx
OYzq3MkR+Sqz58w+35hYnIvjfEBbfuiLec978JJ8ps4AYBrXz2Ndq5qDemeurBqZMRjMribXO3Ze
ZGauOOhnhMmrDXV4NgOhOTsldpZVz+MbYuL0xp2sy9aLlHHgBmUbxca2pQY2/0VAeV+T4fb9d2WU
3zOY5DlhXQW95YFr+gsQeaSjf5Wqca8oGmvnJ1rWeuXFkKcUcRBNr6wngPF05GGIw3XyJNGPdzwT
uRIkboP5uvoR9d9S9amDkqPM1aKKOf8SSTCihCMQjuUJbIiz65Kf287ubOecKhiX+w+08c5YHjIl
ObsaVlA6+oSGlv39DywSTIuFkLsuCz/fKuiTzt59IKZJSZZBtyAjdwRds+EQsq+AQLynXKwNVLU1
pL/LzlFiKGzw1VQlKCV9s9EGwlNweuSCowjdDX/IfCCVJjfYuh5ycSRdaaQrP+hcJCvYTMAeEGPn
kjqo9n4uWCEL9/gfgAawpiLDLpQtNwDV/wzExLIht3J7Dss5PdDtHGrricr5WFaXlaelHrnBP/E3
YJrN8a6grqL5Flr1MF4XX7n0yKUsRF4H57ewtNs9hpbuNUPp5wQCglb/ZhvvoNpaz9X3kKKoNRwb
bW5u6bdsOviVpMLXMpUc41dJKiogcedkS1VwVf1iBbzZtSSmqAusEfuAQp1J009bwNJLCzRXB23s
rO1ElZ7JgRlis8Ap5E1/mC+5iuk7gIJ/BMJxyKP/RVOrq9aBUMwWRMRh4JEpihqKs2I2SsYMdSrV
lWqfE2mtDtxpOJcRTnrCOAXtZa62/x3tqqW4onNGZ4DzmGm3DzDsSbO2z96Xe4gOcrAfSQWzzLLk
FHlH1e7HY5AXDfaw6yDUJs5yqhyTMxNPjdDkGjNY8FiPGnQnllRBxTZQ6lpp4+6f06KpmtVjDBf9
rNR3+xGdj4WBegmcl0f6IWoJPUfsD71dfK9WGl1j2RXPJ6vMSm8PTqpvoFEh6AJqf7Bq5q496I4p
Jggvomp9OHgkDK71kq1pg9Z2/r0ffkqVVgbisbD69TjUQudl6l4cAlWggECYNfNBa3u6PD3rrB8K
TaVbYunHKoN5h54Ci2dA/cY11J4cII4h+7aFwhVrBZFTIPv4DvB/zE8+GXqSS0YicK11hJkl3Bl4
U3GfObrHzEffyqWB3DhGbQoRYspXXR1etSdojNYJKclm9VsUlZlZFhIdYlKCuZE/wThG8qq51jZP
opcE+qLXPclvW3Gw8DdbT4m5AAST7hvWzPcMUVDNSXPBxmd4pPbAbOovRTivymHlIJ75Ckd+EIgl
RKthkfGpgWtzjEVyg03YO0mcoFyJawIni9WAxHGoHZIV9Wg2Ksad0oO/hgBQT4qSnKHYLqWybVU4
i6Qz4mDXgAxKqSrqZ/yVe8ay9eIyxofS2b2HiWegf0kxLHRQHAsnOziaOC/IEXf4ZQawyx2gM9Jo
oJObKTPrv1B0dQJrQJOIq3oX22PU7P31SBQ4F3BOxZ05Ivf1ZPsPQvpk54Hio+bQz9KWnJ0yLPLh
ohmhGPKBXwrC3HpoSu1sjwM8DkZ4BXH0DRE5sSbfyT6bCAcC4L5n3827DqmLNc1VwUtBJQQKME4N
Gx9SlObJaHCx656pkAprAI9t5tWVvRvzZDQHpYuSvEbEC0TBkUbXxBcsMj91+NF5ikmigiyG9Goj
bDpPNUr59H/gz47qklbpCbfT46G/K+YydwXnSt1g+JOvXXPx+JaU3P2wzeLLUGwYMwYk5BYu8A2u
/+ixke8KrNkE8Gz5Xronu+624gIsOhy6DOvt4xtCX6DfB70YsGjdwPQgUd8zIR79NIPrd3Aph4AD
aPZnIEvGbR17qLZ5ZbPRSa9DwOqGmjCWPOSN6x8ZkHKY0/rDEYZmA6HBQ5Bej4kyC3hq2WzMr598
h8yFEIrSARpEnvlHjI6SAe+hQ//TjXxXvnJmb6ObOoDpfFZieOjdXpFxLpx9nIt4ztrLgGsw6wrL
E/GWzVJdjDTRLOL8ekO8mpxsgGfY38j4d8Gl4EoSIqUIQQP6h7aFUnApbpfBjZA9tFh6Tmmjt8eu
kfpCeV+56g7oymRz1WwH5RkwWBYyqtpwwXez3e2aOhygpT4YLTEI585jgG1pUEcX3uZkwGC022Hi
5TM7KTsg1INpv7wB24Zcl94Gp/cD1eOXaYRZs96BEPOO4jPCTfr4rUE7iZTZSH4n52FR087SDR2Y
lZUFgnh3bRpq5LcRZMuBmJYVEJXM5x3qBUL536Fv/FUWeOCBx5y5DZ2hocv7iY+uMGs6SP3ItepQ
2MGXxSZV/lM4HiwsjxcU0LRaWhbtEsKy8FaZrLoU9X+32WVRZWZSlrssU3qA5fUuSq2EUPZSU9tz
u/RRpho4031QrciBKyY4/xf5AtRbudi6HKW73Q/W4b/MZFGFStnFHK5LfvF69mQNq/AvXzy1c5mk
mvGZgSbX+1pRBQw7B33+2xyTZSCYF2G9soXzV+MAurzkYc6G4zRRq7A+dzkw5qjL4mdX8Wkeq/GV
HjGOa5gOjmqGxHpcDi2z94qAxyE8YvHr12ItcM6Yt2X5rTLzsH980hbuIDiEQQoAfZBoD6GCWfg4
qRFDTWZWdrhjtR+Vm92VOYzJPs/zdV9kv/OPs/At9r4nVw9QDdaQmbhU+RJZdP5u0IM/xCemMKaU
HN8SVo6t0qh45PUfVgPy+I2ywQDTpSAKIpManY3leCcofD8cFYwh8HkQ2LVZ60FgePpIyy9Jdxvv
VraYzxU2b3tVc+sXfWnTEo3PAoadxhGc5dBDH0iyon6dOOqec1N28Y8VVlJliQWQD0Yo1VWZXBOz
k+BSTllhJM74Alz2NOjUyFZc4fnPIJwyfDtyJKucHzVKUADcXAuTPQPKMVwvM3YHJZsDO3JdmiBu
Cc5yhd6pypodkTE3is+wlmMo3jO2MIcUQ5UWUu3hvVjoYsx9lXpX7OHOxvC2nMbjkD3iSD7oa4Z2
Jk9LAQ86EnK+LDQtltTZdhEwHlm4FM92vt87yuvUhvOygvzluG9CbROSDlflIxvEa/BJfy8fWdor
xAx0nPFYdOKqNJNK7Sbvin3+rmk/DXLyL0nbZKqlirUXYeJu4b/HU9gMbde6LV73y8PJD4ChULmE
hab8u1fpqMHW6G+EH1u6HLCpkB7qmiIJTAp1ZglclQcd/akD5odvbwT3xPHK4NE7fT+LFsQH0yAa
Z1z2ltuY96XWvyo/kAIenRpNx/pGWcE9QB5xlsg3t1kr84cfXr9EkJjDQkrXHa3c67K4Zr/LjJfw
22a7OiCHDs78QUsOtuGuIo4++23gf3Kt+zQALUs+yqs6K/WmPHo513ormqjkx1JgDJsb1P54XJK6
6S1NrWH6JrCpGM4W6iI0IygO67lXC5JAwoCM+1igVUVxmjnWkg6nbGGZQS5Om376JRjyBJ09AO2G
nMAJwPdlINP6qrXzEfh9TEmwp6He/LXKWVg83VS5atKIkUhJPWKA+6BP4bQLEAaQ7buTBICqepAF
KPiozYoA+0TMvkAMEOy40S/PiO9L/CZzfbGLVIZaSI9ygY7mAHsiC0Y0TSGgBROUESFtJEPLo3mx
Wd5Eb1PXb8/RP6tv/3S1VMRQlSbklam0SLUXIbvH4WT3LHi9T0ILkST9AxOZiRuyapen7OjWsT7w
JNljQQ9B9wtmoWHuYy8dGY2UBUyfKAWFpsLygmiBhAdb6o/0vjpQ7yB0Ze6Fqn2u/94RjOZjYczv
W8HEU82P1BVsoMU+MG/PqUZATMDLEmUNBdEA23mVz2XTXSZxxISSFcvy5FjvZO4XS5TWXOOR6Sj3
zvgOyRBh18+lPNUAFG1WD5kNnuSlZ8jVFm3WZ5z3Nk3PSk7cMDgxY6WaNph6mtGJ+JG0u3SpI57g
T7MSkWD5jMO3O4meFuTO+ORWw3Jz9hQuRIJjxY0byxFhDMUTKxBhspvY7sJ/pMsRkQItY5MkJW+1
iOFem2bTnNM2lInJ/AUXot/TqYJF2tmH4mhnCmiubIj0WjP1OkHhti+mfPLu1x8M+6GXaNgZnKTU
fa+u9zohDVxWimeyEj2iV2NU/v5d7t2Vtmzgg8rMuAzKw1bMzWTg+LBiwBt79SaaCzK431138wB3
O/Va4QjkaqoVgydlhIyqZ/7icpsoUi7xOLCcuWDeGIuCLgJUp3XZAQo72vffRekh4O01S2UvoefG
034zcc7czmSsjwZNaPeiMIyM1hsnqPpuYOfCZU70BF7yriZeXitPhYPdydZq+WOEGuCoqJJSwRuf
+bPAaPrNYOaysxxjkzr9L8CYuhBLXtuS9dDA4NzrmCmKYKJyPoQ40MkF8E7LrnC2skTmZvlAzKiS
486v/ZD1d2DSpVK4OFMARBoQ1EGaLnW2hRwL3Xq/1qu2GTdCCR5ccJCn6NYNL/LYBBnkAy50f2yH
3TUTuORz44rlg+FIO3hfG4CTQmid+/HMVctU6VF6l3cVT1V3nNBgCUNO1/H9EsjgUug1XduVoe0m
bIbUm3y40qqnWL8NoI8z7MKVUK4Z5eeAI5nWci8cy0eyIbyBVsvfdQMWWPIj8ZZyl4Dgwh4W/SNy
DzSuwl+aYEWwSZXaeIBm3PbAHGO+oBcwIUmIn39HnMaExYynRASd+U3atWGc/73X0tesPoiv6I3K
VhUttmwfepLD186A9Od3206h+93GJqCH9xP/M9rlBtHn9Y2+H8weMSZQ+mnQEntLAfWdB2oN//QY
/2BHAUhJUtGe0KXF3jQ3v2aHVK3COMp9f7wADsPpsLVLbOfHz0MWKW6YqIM1HznjGs083+kVrxSq
2C7gn0+sabT3+A8s8tQBSrVIMwugfYHEFV3R5/Jakg0iyIAkqXk8i0JipPIW2z/JzhHz3tCWTT6w
aHQzAc2Pz0LA/Vt8Bsl6wkdjc4RtOqOCQV7809DTDee4wFN03r+LrGxSX0BE6dSUtYXX/orEcYAS
bIIA00talPjksefjLwEjhjshfJq/W5UXmhXTAG7V8sqlirBnyiLABScCtqMleCilNQwjoWNatBHw
UW/dfA7Gutp3CyPdctfv9mBLnvj60YqfxzFSsw39ojvJqnwXGWAx+5KVxAyDQekkaThKIj27Us90
s9EXEOtBLnXVTaNObgTCN3Veeay/h6HJr20m4CkID2raUeP4XCnzppKn/ntBYt16Zc0E1XX6Q3vv
EQ5h6vJdnygDQqaZEkZVZG6PhMQ6R1u7iX4aYcEq3b3xax4lERPMBZ6gnbW/WTCt66wszZb1xeIG
08Qx2oFgdOBMDxcg6Z6erYw66UW5SYDVUHrI/OafKt30qCtlFGMBtJZvYVPMQOgWAKM+4cv2359F
x7NCWd4HsQWwW3K0bd85vh9wlYwuCzLUYQF2XWIydQ0/nGSGHioNkSvbKRc5CVBVEV70zNPLsUK5
r6v/gWv28S8qLVbEanvfCZnHwcQ/ZphCAGFEjQhrKVGh4Pu2h/XjWQBmw/EoxJtoWVeuINrxfEK6
bwKjiJl1vdpn8iRdxVaSHoPLhS1IltAsMg7Svel+4ckCmsQb4Z6PxatIDlTk8cQ4niDx/sWgGsjA
Hkjhq5Tf2bQ7kh1l7Eh58W1aLOOM8PhSJr76HQi/NipbDArNZv94iEFwUGYDmbWlF8XCYtpoNVBi
BRL0703d2P/bEUor5vUgC3lwAyoCVHUHi5gQBBsFOng2StuANLcPbJh0EX/C0aViBSXClEgeuMAg
lL0EkMZymLnuwlFz2v7lgcJ1Rn/mYaIo7mGlAuV9sHannAfBoED1SG8PDUW48UPxlgw0iC6bxXrA
U65+rTEMVfFxmzbZ9Spq52y/STYtMeGZBZg7QS1SoiwpYkwqZFtsC2LJN1Bz/6HkF0H+f0IEG/YZ
cuUD7oeRYMF6kyhqzxK8VfaoJZMIpHDgh9IxvEF5YcHSHpPukKjStApcbSYTq8fntP6rKdHL4DA/
dyrHlW3i3vQhCCXbEw593dLCAYW68FTz/ymjGUz8jILT2U9+Lpl2f07a1ogB/UmcU1lQPRGIvt4W
Rgjh5+HSwjRSTt8ucD+gs7XbubSWj8duuRPz8odEDqCrDb6zCdAo6c9Kla5VSNftISoCq8r4pv9r
qYSQQWxZ1isvS/6o3mH5V02vZBbakGbkgs24EwQl8CC3OkXWhEVBgBOMkxoh+DXjP1hiXLDpuZ+x
QhYnlINViqNby/pUzAPqGqjB5MwDyB6h7LaMHnD8ia/k/eEIgmTePtYB2DeYq4z4qmfiZwauF4kJ
uzl20li4FHFpYTB/lwygtl/SbtogoKFOzBS+KhHQKwMMY2yUxbq8Wb6T69u5QFRT/zssvYaaO1wU
hUokzZZU3/HZvfarcrLJF/+jhtysm22S+2oJyzUw2S9ChtnptU2u4tAyJ12/Ojso2rnuSR2UvHHk
eO4q0CBoQtDv3Q4hcTCRe/N8DZ/dviUZQoZNiNBA5DGHB4xbuy1sQZkPEUpbmFcQZKX5V0+NCsBK
SRJ7dY1D1T+WeO3Hv2jC8Fk9kkdGjQ7kEa/eMSvlmhQkikFTemERtk1Qtvp8/NIHQVjHDkVNozqb
1Wur1wB//Kj1frDu1Vfy3r+j/tEUAYP8nfgMaTeR65Kym9ZRxrARwozKdxLFMsTP7tbtq1H/LqMV
EWyF5W5oTzoCV1E+/ylGhnj3iz/Gq1ip4AkODHz2G09gU7N+mMJ8cbhPUysiMafUuLRDYYNqPigE
MOBxI2NqyEWLJ6wrUCGhmMK95dZRIR69QqZC8fSpavnaX0kIg2pEs6WSVUwFFcnzlVQMfVSjQ9Pu
uLtmYIDh6RpbvIqv14t94L7D7Z9rP95xvlMh0wh2KQYS2mLDuUjtX9RQ6WQTk3R5T8tTqu3qbJBW
WSrwiBUWtx0hbt6R5eq3zwxh4VfLLAZyqtMajqci4TXA57mdJ6L7ldJ3Ad3idnSJSrPjezGGvamm
5XboC7LYf2/HV34KbV9Mf4tMmRlRMgDO+9bYLtUlPBLme8Kwh5ziocQ0ZrHHoLUKR1ES//zkt9YI
q9DUvQzBSldzXGh8p5lf4J9oSMaTEJCD/l1FOnczjpv3V7RS7TesWViU0+G/4vRntqEUstuKZEIP
mEBgSr6vlC2uouBieKBXyFaSpt4DBJgZy6VNM3QwA/Jw4lDMcq5A/EbnbA7mXx9bzw+uoo5/36gw
e7i69D+GsDVnnsDenhNZD2zThVDCgj2A51zyvSZiRWcRKD0MG8D6MIvx/4kZ+385cHim5T6pXENV
O1E+h1hlruDyrBfI4Aw9OCDbr8ttHvhQ4BzOJMJYQ5LdtUB60VUbBqFlccq8dFmJ1XApANxB/11y
22paEJa7y7ioxHnFbQpw8r+EgjtYn1SA/f+y/DZikb4NalOI+B66aT+XZ9RmO/rRnX1/J5ipnXBR
sdPjTFjObIDhbiYe3pjVKNigDtqjac6xF9ybjD4hWKpau0MIGujAL2/K8GK5ZP2rQWxf20sQA392
nJ2XvXDseB5PxRJrDCZbgv/4KZAOkLEJftPVWmbUmYAX+tpRgXN8O6f5Bm/nUYtRi9dk2DfU60AU
C3dV2awNDKnQI+IvwyKDOAYqrkpQ3Fpw2V70re0mzsXG9EXsVyflWPNVQg8VVvCMY1cj0qm0SXJc
EbSBDJaKgDowZ0w4ivGJhEnfmykEijTKjDNMOtjve5IfxRkKhzPJcyf7eJ8pUsw90c/kpn16dnq4
rRVDk/7rx1hVxJgujmrKYOO+94197vxyeZfMPGq4G4hBhuAHpWPypT+OKom7y+aBjpjnvXeevo1V
MDCZY6kHehL2VAA49VLpKVBSOTnCkF+g7mpB0r5u7TBWh77HGAbD1HE4G1bkQmE+ZaPGOCGYHYYT
DA27G/6zPkVSu5/pLHJrZ+BGuDHfri4jdxCweS6+i6ZTpChOkLJZP0Ssp/gYFfNKc4plzfMTJx27
a0oeqCWTHcPvYpAtp+VmOCqbEFG07++QWG0QIZHY7Y3TxYQQjexVa9JoC4wKhzfE2Zcx7rrDU+y9
h2sDK7Ot2smksJ6apZll4fZ1liNCHhnXIsnVlfzwDZg7qgygdmByTV6ibS6ZGNzOA78wGNMX8xvc
cE1CNKnRB9w4JPPQ77JPc6jCg2EJQSnz6X93qWckxuWLNXLImbkW4Iihrb/d3yMamGMyE5gEZvqz
Alh6+E6So+OFF9rqaQQmLWLpQmdE0v94lc3X8C/iYesofLYBEPl8zTQTQhLSyID1xBtGdnU7ZMTP
t4h9Suk49BJmAzncdY7KZviEbvcKMYk7Dy3NY9QkCx7aZYomp4ZNwo+fbXERuffyA0pNCo9fA1h3
FO1s0u4yHEpn26XF9vFe+rhyb44GBZuBye2T/aM3jyywOHqJi3OqT5sUi+2Df0wOqVa2d5EiXccZ
5w0QC3Ggwx1lw6h27URISrX2AogNhPMp6RF9rXl1YTNWCXRYozMSIH8Rcv+oph0wZZok/lEcQaNR
8+so+n/TmyGBpl/Q4ONxHRZccDYcQzDjQHsQPR00I69cfmM2VM/iogr/dtzXXR9RdgbeNF6S4uWy
Vyu+XoR076l9S0qL1R75ASZoJFPWD5a+a8KOW5dSn2d/V7YRkWqTUTKYkDtdbDmiWCsrXwAuSjBK
+SJdpZgHfBzzMK+U7uXoZURVyBe21eoCt3YNOzt16+2d/vCX+Fo4vi/P/qJgAJndDOtvYYoynUSx
CfhKwmEAd5PKivsY/NZUbpSg9UEyerLwI3JCUObEXhPk54m1SCExN8W29s7LATVpjACJonndVNvo
bFYqrW/LC0EGZsVSkgERfJ/S8lHyn4oB8VjycexsmE19FuNHq9215/au7A8zY9aziplGeN+9NfEt
K0zp7YUm9L7HcAhlllLpj6lCJELAFs5/KVilWElVPJ6hz3ZFs8vFOGixthYV1IZgGSpyfN1oMCic
9yHD+1qffFgrGFZidmMODybTH8G+uOirWV00fxMAQ6KZxSRhX14cMt91mLvK+7CPnJrTSq9Vh3aJ
+pFfA8owQJXdjKjJwNVFTvpfuuOx0Aq78gctaYh7xz2SNw5GGEFIudh8dIrsZHMXFOBkaO9bE0pQ
mIXCkYrknGKTpT4iyt0nfE1bDlVuokOnZrDlKExQ3IjHzCZG9Vy4uJBY/BHRR9/9Wylz3iDuLWrg
fzsCHKQvFmNchr7tk/m7sFsaShV1FrJm9FZYXwoV3dpAPuLXjje2GbmKic/QvVl2Syo/KesoBX+y
gex7DWjZ7Z3sqvc6CsrK7CuNtul65iTXrJQZP27oeuFpOfl9YotcJCzBtd6cjCytPzjfM2i1zfGX
SWHZFhHXCidrRBpzY4HM7Bpbu3tMHxK/Zj/v7YaMsBG+rLRstQ+/xXfC4pRxXI37z8gxAM7xq7Ag
AmBLHg5ldh9FQy0tRMDbd1M/6GdBEU+LpIABewRu35Nqe/fbrMss9hTFq88XFmBM6n/rc7gkZX+W
QsY2bC4AYCVHZoUEDfCpoV7iQdepQTIGhZ/kCd80PKnD0RL7UDr0q71nHcglkCk8GU7BD6cAIr5Q
SNw+p0s73VuAH1n29nNbbBxPbHIizVntigDp2YEe2MTrtNHMyo8ZRZPP+ncFg4JVw3xQu5UyBl/f
5L78gjAvNSntbh0byJT5iJzPFyrsibA3Cvt2QsYMLjPbTV6X+kh3yKzYkj1ZTFEtfgypR2nOCGl7
RcYJeVrWE5KXmsCTRLO2lm0tQA+gOiazSD/PUmg24ck6mPwgPCANmKjw5Uo2yEq2A9ce4tjKsRyQ
Ak+n530NTt576ZpWJN2+EyohdNVbEnsKObio2kilYF8fAMoWmYgDq9LjEo55KarVhXXFqOcEtCqN
HeO2BrLktaoqKidk4Q9Ryp5D8AIfTj8QX17/nJ3EdGJDfdxJ/6Ukc0i61yIamIO6iH5kqyOa5fnf
K/+EiA9atAHz1bVMTlxHSNd2MQWhu4d/9Ubg+19pfHIT+nwN60BODCAeoocN2vkAmBJ9B5eyz2PP
odD9BFXGqi6DMObk3e8kSzU3NY8bNPNNXgEmPdT+s2Fki1tWAH0hnYLaf1B+dNdq1gCiLEO8sngb
AZTqXktJRtMnrcaSiQXRGnu1f8kJAQf9R9vWtVukFcyqx/5wioolaAal+Pste0afstWovTOjY4o0
lhgzI0F0zPGV1aHOfiB5IIrbQAF0zbdssR4v3uPpu8wGOVrLExT0cPDvtQCaN/FlEvgXDxzYeNLK
IQTsOAPmvGClgUGio9RfpXojBq0bYbGW3urra3B0FKmPQNjyFG/1UiUkAz89azpuKt5GcjaVeYs/
8qqsPcJXVQ9Vr7HRWcZBppK2c1N8g2eKj7qDGiUFjICbCqIkdOPZWXqeRfUdPeGmFn2WyyPP9k4t
Yj4SCIDDwDLxOV0g0CpNc1XnEkXCreCpR1evkijLyr1A2d/nih2j59wdGKQh+Nd2qbYmxHihrZA7
6GC0uP6DM2YWk1CKcV0Qx3ZrJuGxlOVY+01X0/rQpVUslb+r5Svct3Yi6AOsWu44ukXyI+WZrSPK
rhkaD3dIeDUxy3prnkzdhIYL0Hpd1BIrbZPwWBvFw/jz6+6HKacfiRICQLV7k4Eh5oN69AkNtrRA
8amUBDCx3is+fwrZ4cOJAO+QzcxGk8HfnUgBEZAul1iEatrcNKoy3gGme5ctKQsps8PiR7ahXeKc
RvxEPikNp2UHr6Fjf1uVoBvw/KJbTSm6eo21ILt1Z970aB6RscdjwsP5bkqSSy9A/P4ulpzaV2gp
86YGXHVWzwrl/2ROc9y2DyAwKMxRalAM8Ei6TYRPiVN6Myb/FFpapzo+YObxIs0jIHgG7PznY3Ao
yomYE4Xc0uBs+gI78OqZFX6zFGMoMeChn0I9QruKLOJlbAnl4URvtsL4xqoXnQJHXRsWh/zmjhBa
w5FhVeSkr6Sg+dljBxELKlDtFSgsrFJe4w8yEVXEr9kYOuNTIeYRUiuBmoN9sUdG+YnjHevbqtiW
zgLTt5RXM0FrDwcCZqm9w9A8ms5N6X6EIPBCit62goVo0OPjEYIoDRf8b3e8kxVDzT1nHEs4nrId
638zjkn+0jNwM0SN3nFEuj+Bs4Uzpd294mtKg4LGjtWKyjy4xQRFYJGkNfRPJ503O/aVX7J5wSMb
Q+caVv1zb6QnNI1L8WpaSJhlBhgIXJP1uo345CxZTZT55bMEBuqOlNaxtI5ZUFUIB1zKuDLsO67p
SIORRk0QlgOJIjdgVDNK5BNKGRmyg/lmh+hhX26yMTmVD0PLIKiq8rvIQ+++Al6bBJQL2IE+U0ab
yfoe340mBLASg0WD6gYmYiO144bQpPSJu+tr+su5RsoJ4OZ/rIBrYx/3aXppsSx1l4AI7+hYaj1D
Xdq1lHsJ6CmNL/hUTwlQXtCjeQJHy6S1hMSnniB+5IwD9WTBraGG/qWrYfd31HLV8Vvbdypm0qDH
WU6U3BQ7sRImvetdWMVUydBkyvth+CGS3UrxEUwnWMMCqsvyqm+/3Ovp1OlUtkznPpJc7wSF4cuo
DAsiVGHqrkIzAB3YS/SKSP0IiQds6WnvTXA9ga8FTTc8IQP5FpDxPGKhdMPVFRpf3e50MLcTqFqG
vzPhQqputmQZX8QuA9wA6kdtBFpeH+rRr79jUnw9DGfjO/0OhV/j/+CJ1o1Cwd+fwinLNChpg9hH
KUVr9ffEh7/OZ4xja7oxBnJbLVF+KLQH8n0adqsKHUuiuXWhegcTCcBewRzLNjUYMaNEMQlz0s6G
iya+8d66BTq9368tFJILXzx+pakJbM+jLS3ynSvs6TZ2sLVopqbAXPNWQpWCIXY0mLh+G10Dx8Hm
wnauw0CdX8MJ9HJgxkkFV2fomEkHr4mtenXHd4IgeO84r759P1i8o/RMRyo0t0+qQHaBT+827u1n
wkK6dEJhDbygeGEoUKiY8C6yfdDpzBqvgw6OVgylf3o8/KgVMgGfRwC2Bv8joPc4+J1Qw3+w7yOt
FYYyNrDXvO8V1GRXU1TNeNahlNF/tQ3rAsfWEEVn9Dq7IYfMYLGrJkIsKacTA3KCnNjVxRemM1Bz
MrFKdkyp//paN2AW7ldMkIx+9XXIWlbnrhyE2xjc/7Ht0dza+9VTLxBrMz4pc60mq3IP8DgBbMwp
vZYj64AvWsHie1GT4pkjTqN8wRt3q1zH5Bt9UksUFav8ZYWNiC4uWKsJw8UrfxaKtCS7mVAoP9YB
eI0Ipd9VUph0g84nrOEzDscnTr+RJEoxriD1QebkPrg8OTP8KAob3/j5zar3QADQUcRm1t1epHaO
uxDeOUc7Q9wCK9QehkrMUavMYWnE0BVCHcgZ7b5m1v/5MTMzUZzYX7iBwKbEs7zyOA8lTobpppVl
w9gI6IsJUjaQaDb4f/JiA5kGjW3eM7GyWD5L7X9OhSW+ES+9PMatfY1ZKvk105IInAcdNjxawR/A
mam/s2yreWpBtABkywm3CRxbNJ6GqwLrZBGQzH/cCFs2WDdaGwotSjeq3k1kprdlaLRd2N/fI0fP
4boDSgQgP9bCBz3J3RP1IBNtfRDiw05krDFQMvCtrju/P2NxI3EmeH278IxlEyFY5b2hwPWBwd+k
V2t3mO2mZqQw2OT+a+V4QVNuFz+NQ7DavDz5qybgRcPiR0OzJRZ+YLV/zNBNjUB8fhax2CruPDOg
8WLGMZunqJjyAYknHPqrSYPCOO9vwKv1nHMMgtknVJ0ZoMTmIzqw3+Oy51hSpWHVzYwyoMyC475v
jSvNhe7VshKc0FZPxfzkoaURO978ivTmDwllpC5H/0TheBpkXTpSJ5Z9aJs9QN1xw9H9l9UEZUIn
tjADl44tDUshsj9vU+ZoSaUmMo44R+9K769K9HT1fWS5skKo1kh1l/pX/OwCvfl0LL7Xi3V4+Rwc
RaE8D80Ui/+bHzgicQB8GDhnMHOBXK1kbDxUKkNN3aFRbrHV/O5JGKsmIhOGRrR2s+AHtU/d+6NO
KJ9gjOJdRs8lA0uGVMDRVOC2Qx3dQeOxI7F10OALOEfFxzPaA47MEMBr2TUmelxwH80GxN9pFJYs
5K0hbYrjbkD1A8y9SrEVe1409FWkZn6W6we+kf6xFI9mvVT/Tie40nJf2E+wM7ZPb1TQsVEdi0aZ
bLul1jP29WC4rzpEl2e2i95dpmJsIbAs3uLnDUMNoQdkfWjZo+5Q1kMlenp8OkKtW9mTdTgNQN85
92/d/L0SyXUvXAkdu18CRswpaqorN8OK6dEwz1THb6WcjdrFRjSXpZPZ2q2FhhB7qrnmJGQPaSqr
xV5wUFjoHZ6kw1k+r0O/DUWIofEmlTct8kgddn4iEHP43cfSGzKHVWfHVFnmcC96+oueS9vIgjEN
UmGS7FwxrcY9IQL2yLVxy5FyRJRYbMxzROu7RMNtF/FYhAcBk626DVwJjddcfA9+ZEpfvweiTjoa
15nK0CQ3jFo0x7HM+/HyV6+OVHzlaShjy8eTbpyzu7UD3Hey5t/b6v939hPyUcoOaeugU80P5ppT
BsMUC2L/RSNYZvVpLMMsUd0cVjLI11f3969150Eu0nK53Wv7VoUowcYXSbrRm0RxdnHa168EJfvK
5y55eR7H2ETYwO2LcfuPnCwvIEztgKu7aoJKbIEQmoZU3ovx6JGq06u3raZbNcwQDJv+CBLamivk
0ooGqZ03GWwIpTbT0OtiXeDh2K6xeqpm1UYfqGL/Jo+nuSaubXMj0/zUdo87ubuCzAeM4USKKpeI
mJM/4zVmBXr5v8Uw0FbuJR3TZ72xxQgLi/DAkBHK7xmsaTrlVq+FiFP1TD99y/zLeJKzkkwEDApq
0iii91XTXHO9syXzryyhTq2ywLAflHf7bVDhHPoZ1zV9Nu8xJl8W6AgB5i7X+s9y+tkn5JE9A76P
QDgx/216wtbTrvtfPvzlVXOGp7KObe9wVnXgoBeexqEkDWnwkBxaHP37SHGZlG5m8xd/Xx8nXv74
aY3JWkYHFACnJhettESCLUl2XbyzWi4hYy/z6ES0iAi5bBPjgSoi5ASIDpTTZrxtdZhaPdkOZkqa
xRVpb7wAezk2UG0CYiQ2ZhZuSDAy6xoBzZH1j0wkmOUDmYq3lPpOidafOFRJode7wTsHCLyPJN+V
FRHIHIF6nsTveG/43Ost1ZARuPpDjB5Vv2Rv8gFbDUoa2SwyqbDS7a9KYQMVT8JZqFNYhVnlYnfY
H3x3EM+vyoUI4Vb1JltIHSgg5pNKBNBwmVU7ZB1X2kewajsSJesKuQGurEY2mM6To+h6t5Acvgtx
bTO1a+sZNcdI9hGeSPpJUgAD6NyOnbZG3xGUd4eBBRmN8S722aKUf5no0C8SNiWdRPJpBO+C10ZQ
aG4Duz+1Nx095rYZtwONpiRfsvzVAN7Y8tnhYl7tzW0gnQX7tARa5zipIw7qj8hZ63WDS4GWNQ/T
u6jLjKY/JkBCwKZJYZuI7ukUMmUF5+CzbznDLxVQFHdmuZdByfdWNX+kEazlaCUPP14abXaVjMdU
lcFjd0bzqmCNdMgss5Hnt//5b9slGBZiCe+6wuGAdt8dp0iws4TWfffE3KC0EZ90XjdaWdRky0er
4r44wLGFInd1kCYNHyPtky0qK2J+yX/CK7/Xs6i3/tTPMpmA12Hiq/L7cyMge3we5E27BJzQ5JRB
ubh0jCMi4gJET3/U/oi1quTFPaMppQ23JFyI+4D1KlLxV7hgjLVFuo8voVzIe8n3XTg2Qdgq0HPg
gAbtIvEsHptyj9vtoiLvtVyck77wGOPcbwOHjBwAnxHGpalDiiElEym2jakfk1g8HMT3d8t+maTo
C3TaqEwIu7S28Qqpve5o+VPEsdrdZHUQQXTDZ0aBM03bHteg5mivJK/RsJaAGWe+kDf0ilhuDlqw
gATCd+1L3vTXeIIqvPagrSkgv0j5RPBhMeHK88QUVYIDwEXzfwp3MlbqFti7KZkWF/+L4VAQhKr3
5RQhQUGr60QI6DS684RGIp2WhhAqCx5UdC0sVNRiLhnyXmUco6eIrQ8gvriSZMUOAP5tzEP+G1vI
tOXhIfs+GKUjFYUrzm6F+LAKCCt8655pWvfFbfBuvLje/z0Ro7eKExz5jWfOcN7CZOjL+uhETHww
SS89h0mjN89unhcj0XvBAKdbj1t5x2EjnMpo/xajYjq/00U5iCVyiCehGz2UtOQKCyMHe0FR6xJE
SjNc1LhFo2EtWR8Dmyg3zzHmULZpmYPtJvL14PSoa0U9akUJUtctX/11eUmILWxY9cLanHrChaZ3
SpFw2xwuUzA8VsR67ULkIYHblPiISqz/7m3sUmo6qEp+Bmi++dw+rteChbQGAWUEMWbbw/QVmzlo
HnvfFgIztLQxKp36kwbIlr3+ejbBK6zizh17WvCf5aUvxFSPE8mhHuutofHcEy77LiDsaLNwx/XU
tYa05JGUdREjlTm2wD+RME0IdHkhNVL3Ssw2L6LN6dyOeUW57mFL5nr//dgwOyJsIpnokG3VlX/x
L9JDh27aG8g6f5NNIyMrWouPwyeqecr6SC9i7/69MRSKV8YCVkeOsAo2Q43NhqHacMk392a9yj84
gNc1mDO7mU2LAAUhHlpMy065lB9x9W+yv+c5VN3g3+cQ3BWW2Xh3kE7EeAclDfFY30AaVik5ULy5
tNYqPh06hpA5PeglvtuBd4Doiijg+J0tFGUUuuZhZsgfk6rFT0detaK3tAcwRGD5TtBvBt3wgX7e
gq9Sl9m4ndxkaR3hM1Onr3RH7dvg7EApMEgq8KCZZT56tjb75mGUpGnITpKUETTvqyqyQzxqsWCG
3J3cPrpid48iLmx+rydTRJInglM+CELzOmYpJHXL61FPlVejrTVMIkG6ZcTnEY+3EmJv2Pv7FMVV
mFKqCl9cTrNdx/InrUAApJTKAWLrb/jUh2MhY2EvE6fX37ZrVHmsXf4XGLeFqAA0uLyr+zrvstt1
ZkEa4M0MdoNkwDKwDluMJA0dVqaF/LQgsTBZQ1lr1VyscHUDMRS88mt0VnEG9OG/p5Evxl0SJGMo
S37IXRUL/f3INCX/U/XrKR/9rCeFDUVHU5ey7UVgtdDxcPBIl2Et6IgOso8+Qf4cjZcGMbSRpRZt
1z8RBk2l5gPCed4gq8DTp1BOG04BfOIRueQa/uOmDFmek40bDlqlSIeeOudbewxbFLhW56Sehdzb
d/j9HYYyHpesrFYJuiLjGpVdhTyiaNSGE2wd/WuCqmR/0WnTb09+F8JS4+X3dXWIzYXok/c7TTsJ
V0h9EMvtgekCfb9LnORTZn5T95Todnq3cz1gMrpe63kfa+bCc04gXOWEQJOjuhZq8a80IZOdh/A1
THh0KVzhILDFD2lwqJ1wne7Cwe2fNtZC5l/EgruXrPSc6EqGLD0iKrQcGM7+BRZ5z3kKnMK+7JIj
wH+SD0vgTIkhzJZ58yhaRWyVXUVB4ADLWUmGFVAgqwO5Jg6TNEvDy7UGWJ2lMadJtqKjA42rACcf
Kw/tsrfrfmqTY8ra7TRjHwav8fMv8zHebbZAD4rS6KhbSSqmfM07UJCWNf1XwzpjDxml0u6A2Iwr
oPhaKF2rSiw/eh485WD50IblAQs+J7ocfRifofjzi+dUb7w0DmLRZd+goRJXsYkbseknpiPFjCLY
jqfZuPaj5SLsl/AWObjcgdqLqMBpkXDCDPwBlPHSEFp5fCQR5+fvfEgemKt9Em/C0TQj3+RJr9tM
pxhg7GJOwSkZfIxV+FUu2cM3dsmojvUlhKwDhin+TuvYYUbA50pOtr5BbwMJxITgEj5DvW9XxjOL
sPOtlmp88rS3zcQcq0W7MZyMFgwREy+o4/LaOoMRGGqd/IdhbO9GluHrQDvm8S7gFuGRoOSPEAUf
ftd37v/FaCYqL0J91SfrohYuR5Wp4TCsJuT5ep8uRvwZFRRo/41v9IwI6yjHFRiRs/23X6EBx4jN
1dUO0CaUWrcILYUUX7AcR1l5G52lni3HcszUTB4ooUCam8CEmh+0OF/+v9b6T0GmT5ucj+52FQaE
F/+VBt1h1+vUORjnr3tuSwcWFck0XkFLaHYFirmnObIF5RJEy4G8RAqqupYGqlDkO9oOzXHzFKeU
gEJNJssEmzGaseFEw4OOl39sbxJx59BGAhgNK5IaRnNaofoVoMoyo2R2Zk1eKkiIbgngIeaNPexS
wus68c0W6jlP3CujNDB6vVxb+iSvp4mWOegO6VA/G2MtqZ8q1cjM6Zw/oTf/eSPF+1xa+DD5uuK/
p9sgHEpM4DXbXV3U6BGghu2I3h/xFvKiVPA50Kx5VGrlRTf8slD3gTW/9QXcRASCCCxY9N8hyjMK
o4B4mRpbaMFFOFNF2V60OLeKsF5o0uVlvwVKwWHTNPIogvgtsSztQYtcT2aDC1eQQgIUp3j9b6uP
0IJm/vNmSbU3t7fG6s634O4CEKqKTQ8bTatSWvFll0mf8hzqTxxe5+EqpfRugM45wKPxPvLdpJZh
XyH+PHXlDMu2wDr+qdMugwYzXV3gHViPw3iLXlKytnvVSPYZNk7wfZ/Pfu+y84L7r/TuFqFgXfnY
jRJRw5VNwAnFnK5TDVCWSZnBZ5cqCpVF3yUsRz5ziid/hYtq+8iKZC88M8jKeW2ZWfjmEa9Z/PRU
cbJRwOaeWDCmC7Hsw8UHwcv39cdeh+MdihrKJeX2SOHFtrMj9/sPgSmQxA9XPTT7w00FMZsC+ECe
pN37dgj7vtWi0Sw9HPMkcPckqDRNF/333IpP7JTLackR5Z6SSGPNeTPVRD+CrRNvDfZQ8nWF6L0b
59E3ktcClaiyhyuyhNQ8K0wZMadLlyhPufuyy719Pn3h9JbpaeWgHM7+Mrzy5fUsyn6q7s4uOdY1
+wilpiAmDDTuV1tzuk0OCsS5B55E8HmJR5UEZ3Lq+GA+BdskLP8SQnMvzSUwy9WP+lvSxCVkufVm
TnHZiTjs8Zc0LW5tDZrt7DZO9qqzRT+Rp+sU6vDGNv2vKpZV4ue7oacSRtiXKAulqt7DZKE3w274
iqmhcDUe8KZ70VCEpcaRjxRC7km2HexnBhSih9o8J7w+JfhECPKfagucWqfHLNoyCD7k2Dh9Rp+l
KwGgNby0BD0vLI/xCcgtiNe8bpPGnT0JV+1b0F7rTas0W9omV71ci3Nb1fGrCM5zB295tYZtiG5o
QZX0gBIBQYLHaJxPRBGjEoSa4LnMchH/kXN3+0ptTPsndPceO8AlEauHKd4cHXUhCLw9YnyM9WUH
uiVY3q7q7e1xIAx2qgliQNpS+Tq70+UYpH6dH/FXFjKYfwOTwNQ1WtX5EXyau0Iz1gtxUij6mOJv
0LTtJzMotFyA532N4HYZEr/pWrUDhUmh2N8DASdmHPud1DDP9EKnhLyxWJiQOpea7mSCF1gOIx73
mqiu2RHgnXLElTXTXe9zn5acDZBxXOPNfYgGkp3uBsxYB3vEjmRNc5Mqkgg8QjWws2paUXbNNEa0
3aovcaEcdMcsevJW+FVMuPZghciBXhCBqDFhB3mXcwTteILyU8VcVX2KuZPAUV9NbIpqjjdHthjS
XQVaZx8cGPJKWLF2fsw8R0s5iCMoEccjmahRHwRNm4vsZ8z/jXf5rmJ0U2FR89OxA0utmIJFuYw9
jZrVOMtReIgt7QVHJ9WfHsTyh3/awgPnBMOGMiEd5tV8aSbHhZHIr6dtlxdpsC0A5irH6EA7VVSW
I4GsKCuXmjfGUyPVS4S6i8kgA8K63Kl+rMBxdu61eZP/FP/3cHR5rpV2IRsimQBWGDFzbDo+ymLI
Js3R6JB0gJwuxuwAC4PghqfnVuR00ET9aoplxiSP7dfI1BWhF+WdYJ9UAtM4AHq7EDsCUOT58HVc
TjUl1qGqY6Q+QqL2p8g9/6G2lfXHWP/lZmq5D6m2jdCVq3xA/8tSw4bY1K2HhIElI4XizZjXW1tw
EaNVoX/r/vxjP1GecAS1WnLnw2UPnixRsAZavyYJkObeNkC/ZCNpP4CSQYCAOkE+tPaVa6ocROpd
7QN4ygKkd21zdHzxQDOs6Qfpj9WaCQ2yuF19K9yb61LlNj+5s1zl8rYftxV7KEKvBGiTI0RYNz+e
1WT1qvxUj8BvEH/tpUu2g1dBvkLyg6HCCvKuBstOTmfRdDl7vPRDEV5S9A5VwoYJDxsFdHgGjvM1
8LJIwT9sPQmsrsB7Gc3ujF3IfDks1r4fClOud4x3YtJgQMJx2dHfzW7rfBXHcN2GqTyRmQ2xWqfL
m+2h8G/w4k/nW2dHH32/k8I1RJEt+pxNjTVqNQvbIIn/vBPzJwVGSV0ouXgN32Hxjz5yxwrU7/6O
r8d8CvxU+XiaumL5D5PZ1HCdyjHaGMnE79OBmtW14zH+wCd1POuzbxQ2xkaoPSPGoTOj2UZKNS7X
p7IhKSnypG7zLHW7O+LNGgXnJMk/izFR9OEVb7RX5dMj6wuz8FFIPjrLQW0e4uTY/JkkAoRlSmXN
EECvnEgiOoqQeR8FLuXo8sLSvFrMehQMLVR6Akl9k0DSbcloA3zsRooo6g9WC95/kujn0NhvFDAm
Te9CinbJtWkl1oeaL/G3wwOPnq/EN+oiYu6qYhaL6w/P0WR76WCeCahgv7YYoh11tmEC5uz1Nk00
hnVbono9diaYc4m7URKPM+9OWTGcLjo/WtVDoxBDpWOZwLXUrFPfO3VHTH8F0XcRhWq0Cdp6hJ7l
54AWbKHcQjs41a8mnNl4AT5Pax4vX686k0FPhFt693apBaKl4FBUorerAw7CR6B5V4R5kn8WPuPX
LMPJdG5jNTxBAH0KAsW+pR2a3/zcsyHDwHvXrWPVnLwD8qc0oTdGuLZWlmrwdTmdqBTOJJjkpzfb
kce+AXftUs1Ika3sY/IYz+Raoh4aPL7yKAkmT+ggDMXgABe+dEZqjlo32JmtAgvnfL6mIJsQrCGO
hbu0nxbesgWgPuxaOK/U+nKe25XxFdp1FYUThTahLRVeRNwc3Pv3NLlfmVtjWFCp2SOBcX865pyP
galgLoxBjzPlWxYqRRY4LwBA1Q3dEtTN5CTVtTpkM7oeLdYjb4kwX2PtoJmijpLFx1J0uE2xr3I+
vMhELWO4dp8bXtigktpprCp/W7MPJsMa4FaxtNFpClHr3Q7bOGCBqa8yArSBx4y+f+G3T+4pqf6k
2RyHRA7IO4rkjjL9RDkmjZD8ZwDGB+GPNKvucREWhyjmS1CIJ6Dm7a9/GbWyDZvEEFb8e3inZJ+6
U7GzsuUftnzGhBeKLiIY1TsumWY2svTwkL1OlKPPVSK4ZTbVL5v75y7ZVLyRkwJDRObvybAa5vsf
/Mlk2oGa7+0Nzm9noG0zOgDpKyNFi7tZgy00y/dx6tChkkl9Bz1qna6Wc5bcKqfQI1XmsbYZL7Bg
m1pILbLBD47ZWSFK8+Bp70nJaeAXqhWkDZ/G+QNR4NUEgxRodZRZA//fYesGT3VG07tLnL/tA/a9
M49OrBjRN4fbT3XKxzgvThnFaHzdzT0icwaB657p6tl9cB+EIbyKt2W5hxrQ8D728G9wwUAm85Ht
SlbAVszivgEC/+vC5RbJrNH+8mPCaK6sujTYfhyfqjtus4AQA1ick/kTxreAz0FLMAUDC0seG8Z2
/lmuyWbkcV+lnLXwrDZKOD9NADTLuYlsPOnVTljMWNdqfzClfWpKebLkmS11lZb9Ss/1A94bl2xl
MlPcm+8fCr55AcIIBCRp92ct8ZTl2lkzEUUSWSFAk5L6R5pwUh8id6dtC7x1H1izhc/hCKJdB+tS
nCXAtS5p8zaF2RaaZ+8stUieBksGVe7R5L9inHPrMFbxsuiYuHLmZr52K4Skk6fYaoZz5ZhGxXfO
OC0fcFQ/M5TcmZn5CIjHyaLZ2UdTbCN5/CUVIn4ImBQLlbQ1rcW8zD2641ubAzqRWtAWVMwGnwGa
+Yas4EGxfLrfgpcDCcSLM7Osx0QaBJAzGCo0l+xZeqCZUt8xjs0djw3nvj5Wg5xb5jwdVj7bPq1V
jzfzXEbt06XEpV71q1F9gPIWBEP+hWOP1qIAr8UwfI/s2OL4fZpl4MQQc223o/MMit9x4tkuSaRX
1BRpEIYmXRyugpW2UsHOXEXStitLiV1UTnOtfeH3OpX3Cq04qP5EdVlxgvIkN/auRtZczbJM1FQJ
PMAIS680cRY1G880hdwwH9CevXFXCb6de0CkGcP1NIi61XV2+XLnSVOI+9LEzkQo+ytubRNP5+CQ
vtiSkQ9DHoYPRDHeu2rodSoNxsq5BqiOIV3elx7kysv2nj3oduFEd2hdllrLsEkoI6rpnjq+9wTI
Kd2VIPSuiSPgKK/0H3SlA3q/NJnCX1Yo3bNBdE2bweMdvaF9f6WTXpLbvDYEQfwH1xTJZzS1kAW0
vwTp/MxXA6eM5pszpmAAqLSgKVnf4RzDqsCG3xi7WM6pDcbFP+NYez7J/69FfL64OoFG+qCS36+h
Kg0OV+hKI9JvaOaFr+YQVA2w8yKFmduHU9/G9cP6FdE5+cUn9V/BtSfimuF5uIVrEDtFsR9A/zyy
wRdoDo5Yz+cXwhAF3P+FxI5tArutAi13HUc3WuF56f5k66C56fogDd4jD5WOD2qxRAO1n8XaJ3pP
uCnguVsc67gSGFVRegCdVEDmCTK4MvW7esJcplXbgVkQcQmF3lQJOeo0q1y3yASk865OdqTwhKO6
9xBdi7NUVY1Bd8j3MyDcDUWeslqEsuSA+VIbXjfwvIvYSA4RaPsnnc/6+2gMEj22RkIMmDPhVPPc
J2K0kqGA/oDiHWSMjEUJzY3cwS35MlPUoxthb/YCMJ6fzgUx1oBae7OgOWJPrHglt5AGXCwpKF6J
MoVCz2vmrNh8Il5bljwAqVLbShV+bKVPAxLGMLMbs+3SGcKj6E2SbEVI7pOUV5KqWbWDoXYwTRTf
HZPBwXKYMqz1P+urWGyx21mSJ+jNoRx3z2lE/IENyJVJGGA7oSSTWwb8lO6tGHV1G06hpmGjGJgL
wEjXUPKsP5GkQZ+/RLtcdc77/CrpiwarJqDijju3IjEL+ETtdKsPV/EIpjpy3xgcXjwyCzzTakve
7dL50sG2u4ZvtE97wvFaYI+Spm91iQigVmxmo+5WYbbXSG/oC9huKPcQ/PSc7MayyTEtfPKM0YSq
W7/4H4XDifgyU2GVzAUTiA8nze4aaQfkBs2/3ox3Hh6W7UjFuUbVEolfCxH+ufhPrrz1z3I2rVeG
Du8HVNHRvSi0PSwEw35vNrPXeZ1NUl7Nj1PXm5SbcUtbTMPJM1E5rz9zptKOatOkWtNrbtkHzbvr
fHvkm1SYdqG5dG72UFYktcVaasJoVDH/Phz0yUM5dHYFsf26WnsPtzVqKL+++f5O3KeBQkl/GCz+
R0fVsPT+OIVhl+nINyWTtOqO6T+S9XtEXi0R7PYnjrGN5pQu3Uj50Lomt9FGEF23hbEb0wrjorAy
sjmK34teoKyQgKUo2+0YEWj53V30weoHp4KJmTOxw2LvUu4Y8VSB6EctWcYwqxF2t93/Dty5XIfq
jaV0odVFSxDCJDvFS/19at+lw18r8EoGZbw96c4B6PaP8s07mN8QlRjglQ5lmiAtEZjTUVGJkT1S
TaQk9hF7C3gzPKEDXYa16QOyekqKPELUQ+bntphJ1dOStwF1xxS2hyzyTHcVwH6LyHmq5iH5vnqK
W4U4BcWamllHnPYpFd+I9C3/d6QD5NX6dHpvX/dYRMdbShRiArIRG3f0uTUQO4Lj0415iveP1zt8
TIMts9lt5pTwbtfXsCKJF0AAb2EtMig+HiTNY9y/YTmfdI9BrLcAAq+hBpb+h/nIRjtoOemnyAb7
w5hT0Fz41jcgVKMX8lzjZ9R2EznbN80KRdXAeu+u6l9LeHetCTtC+Fa3N7/5Bd93Z/zceWk5UqYf
6x4df4N/8aTklT8VsaXHeVhEJFpDDMXFer9MMR8bPxjcuFlEfl6/rUFu+wLzL88IyTXZ3GU86pld
dN1+Gsrm+vT5iUpU78TV6LXtxEcJcUgxYEdf9wZZBtYBjhBAZFoHQ7/ioYyWxrcKM5OFrfUlSpyk
yaeXK0hCSk8K5vRV5iddfmsA85t1SlUiAV1ETB2w9vQ9Jq0n4Qd/T/vcCv5ruoFwt7q0iqWiRMDP
Xkd+eaM+xswW9Z2EuMm2ZrrdtdKJrA1YTQ6siZfKc3aIcAJZRwtWJsRrq+80JOnClylUzx9nKA6v
VgLtEQNRVEhhdD7QU0Vs1A4NZNUUmgB+cUGa63a3t9L1gX4TvTI+QAct8gArW9wRH1+1PTOAeBvr
/XxeH4Q0a3YlJn7c0lWePF1To/TfM31p6c0DIgVwm3nKFa1jc3p8JUoWp4I6kEqowYG0YQD97KUF
qCv0wcCSDXhudX0HTJONSVGqBNvdjAEgd7mJIh5wcCGpUiuKLhHiXxyLmdS3lHrkYmWVliv8hZm5
1+43KbyaRtXwFBp68GEAyxvLJb+4aI54y/spOO8X6FvnGyc3CLLGAHzybmdQKOdfZKjcvuBOqfSD
pOlTohRLsgFFO/MEybYVxEF4+GvmyQDLCDquOdpqDiqY2VNPxhWay/SHvbHmMrUnS5USXhQEVUi1
Vty8fs5PnACk5NGzjvWxZhKxISZwDm/wcyki6ASM7EV7nQl5zG6shQtI0T583DcZcH+inehVUdI+
FJMX9eQZS6H77pyAibRwu9bsPaRkvU4n4Fjg2p/7E293g0+ujasm+qLd7BA8VL6TH161rgmW8nWb
NwI7TzxSVd18raW/Cpv5yZaLnj5reZOFGK3PiX/dhix8xszkuAicwPTiOCO3+8s263fZfYkfXmyY
miv+GNvcbJi6pPvT3cveRkuK6SvaSlbV45K2uoFwqAI7TEglwNfw12tTx3cMtHI6HvAS1eL6KMpq
PyLXfj3CABPATQNkWjKHY7GOekFy0oapC6Nwh5wK3V3aGm0hieMllisCLN5ky4+AYBdBftn8j/fX
5qTmcICdae8p42/GmLwZtN5KKyJNR4T5gsbaN1yuifO8Z13z0NTsvCLaJJVf7/BT3WyPaV6t1Yst
C7lcfJ+c5CCnZjqUo+g8scp6KwFnx3dsb7XH+Qhf1BdRV7TW2Rvd8YSIxV83e91ZzmnqBcBtC6sh
2Y4WbbifR8cX445LQACrLz8VTH8D+1XCiCs8RbUOFMGqxHvywgWy643Gz97nduqixDYjDn0h+hob
+SlZ0/3P6yZpF3Tf6I/HrO4p6eqD7a83i/4qcKQLn6/ZpDYO/cl0H7odMpOX5CC44Wn+AYPRZv3G
446kiM0uOcX0DVF+7X5rg0vZjCqRdgMPCG/DeCFT9L06unZ5qgC/MraBnpMZUBW7sF6lQ6aK7tvz
dK/i7fwUVmn09sZqkIVqG0Z3biJugeJxbur9tmzEowQLcQXU23dxZsm/HSIFawznZu9jP7DW9cYx
yBSwCnZ/Y2KRK0nry+1zcC6GJKDmgWvULOJXXcVbHCoKdgoos2BpY0xuNYt2PZnNALHtLXGzLTv/
WVy6U/x/U3FQGAGTA0stEdiH9coIjD9dbit3WA29wWjEEg5zyuw6Lf216EzcKEJ8M90R4U9gmO76
Hyw+uYl06ABDTtrz6nrW+0QBD9lw9iIHIP1G+P2kQaIy+zo/SRt2hOPYzuwCwn46mX0eDwTKotZT
iKXpDsoy+jKlmu53y8yO3LancQM1EjQQ89L3cy9viliN1JxdQKTyhwY6l9ULjeRyhf65nLvQbr/I
2AuLA23WEPSJpmvlON/Lakh4PhOLb0Shqpmizxj55llx8eN3ifua6xdxGs6tfoh6G7WNO9yQsc5i
lT8o3Sq4dbGvHonS0vFzgGAIMnRy3dXTm7AQH1N7OW53oGQjTSeD2cv1Tb6ZKztE2F87Ymk/SlGI
zoSqtofLKyDQ7Z68QeJtjtLwfFHuESpMtfK6R2bbzsuG16GAP03kReCmngkFf94+FJoLHpnBFR95
gHyWNmqOp/6dDVUKKw1Pn3enwnWDABckDTY1vo7Hjj36RNUyi3vUen5g4ZDqBMYnzsgb2s5rXiJ5
XSW/nA1CQQ3C+N/jPEqPGme8DkduzvqJtmIUq+CFt8IGSY4uxgL7lwoSWRa2+QfjhMNQAnqyMdPt
VpRsTHEyChPT9H/exgUr+YRJs+M6jwRb67R8CRfPoYEou7PbDHXyuet0RWItM9EPmfyTOrswEgxA
nbesS/f6XGR5Sf0mP0n0LpJ745uuP3L8rPb6dnnJmyxOPqJfzO1+9TtsiUDE77TCtVpfNQoVlp0t
/c3CJQcSEiU2vn9JdEvL8V+f9mlWQATKC//aF0+mr1HG4D70xAf0VxwwplCv6PudFgsWXmJapgXL
kWEcg9ynxcE3QvPb3LmlQUxP8eSkxF+FhoqQ/p5LkZZxIV2WstMtF/l6lTzw+3ZxM39q0JH+u0fS
Q51zxaVj4cBsFMWQkXCw2y5d+OWuYVhdh3LVQ+RsRb7hq/WeNNIZaiGf2AGq9gTsW5Bk8m8LccGU
YYscO8L890JuZZOWLOjKYIuD2zl1ODR7bempycA25OhXZb4ZnSv7LAfCsVjyglyaKslBC/0BqLwX
OBC3q/TRBbl4Wgkbb2cRbSRQyGEqlV/Jmxsqm81u6StHh1HUfSnivXDpAJ4ZelGRMkaNW/5XLcrZ
tRJbXvbE4TYbYtMKNxDJ6myrcrY1t9QsewTe1dHchwsaoU45MMYI6+8JqBq5tTZFzEnJQPP8u6wN
4dVcrWFlKLLan4qmQZyC844mCSREqt+X8Itz1Wbso/U38Iea69JVNv/j2yNp33ImF5wp064Pr1k5
dxXiVBWq0EaidXCo77tPHikXohnv1zE+M2h+ag9y8CtJo83VkvMaf6Tbsk9XSryxvbjFmwkiYw9r
CsTjlLXdtfWZfDAvHoFjd03+4DQQTFlMflAebAjred0KF4kdSQQqrZTCMnMSqyKFykqib4Vw9KGm
rtRxOH7ouuckrl+FMUI8zglvAtpUKLE/pBDG3OaHDnsuR37bQKkcERKogRJyEwdVHwO7hKul32Gj
B6ccNPqGapnZgGJJ9W2CHiVkjX+oB+k1jDKXwZ5uEASnJPdeWyVk9v9eVI2hZy+2f9Ocpx9XpdsJ
lmBaykvyeIqk3+G/3F66KjZs7GVHK2c2ms/cV+LQv0UGdHG0OWpd+P1m3yJLgkuo9mqSisouG7Py
Vn/O6qVOLsnxmk9WqyGARyq2Na3bk//+HF2GHbD+NDHmSdjP9+oZ9sNzLQ+H0atmQZNUmpm8xm3U
NdEuRizHiUtxgdUA/eD0oZauFjsmJL1MyKtVwT74eYfUjjXudTMJi1D5CP8HeFpfwgCbxzDVJaLa
DkaBspk6x194kiVTc93435enniRSvCHJy+kipMZOhtbwswEAuD9tW5Pi2PeCB+rs6smXQYZ9xNe1
SJruZF8MI8vLztNfwtFF9nC6gG2kyAr3mLjkaeO/QJy35vlxDAYAkybWNZKvzHt8LTW8ejb3DBNS
8Aw3X8+z6bPGgQIa431LHixtTU8H5fHiDojBkQepv4N7KjpgPa64t+IjUwLLPmK84agsMEgelML6
/pKDLQ3nC4NfGb/pRlE9DcTTebf5lEv3tgYp4OFrzXW/P177PjsD0P/iJAkQ69MFOmurlv7qkDT+
dwki7nJDD1CQ5dVtrci3ZQDjmIWIfOvaNZx4iodqyr1FUmABSKOq0nu7X4gk3j5fb37SZa7M5PO4
NfN08GyogcG6tMnIn3E+vK9jysraxkJ1w1Bn9dZ2/Mpyr183INlJp5UrTITirEnkg3KkAy9hR0Oe
B8DnN5xDNFEM9lSOwlY2ohRoIVpN2RGEySu+j+LWT6pahgTae3JL8BPYZ5hY+0CqYxSBYKC487pD
LdERYUwzPral2sGWIuZ3oRNvLeLOenyHGw9WycZ/TCxJImUftaTKxXKciafjEJow8ozbU5gqJDzk
wz/HdQe6ctyJ955OMBQ9f9SKSl5VxpS7lrfy1FmBpI1EzQMEcjN/DyV+FE5Veco2hvs+YrbyWoiP
cx4yTYH8/TG2fQhvO5fhHmN74tiXMGhKf32bZ/DOpF/DoEEqnwKBJgln1Lic6+gSE/Az+9GmrU0Z
sZPF1FXHFa6kROmHV7/a69mXRYACLIpMyaRDVHpnsYdOi4ySaxT3yshpV92dQg7BHiBiJ/4bc/sN
ZNT1tpIV5YZ2tEyKQu2AiqcNud3RMyO/eZ/i27L8Nznfnze4I4yfjlBBrNiIRpes40EOfQGAHz1k
mRWPQqD38sRk2Oyc8eR02nz9rmKlc3m/D35iqBZFhzTs2NVraQM983pupJOJOC+8sqLXCDzjK9/d
nDMx5rK+ue4vw+UWkdytShuqvj89paFZ+bT0G5b1fY7U0sg3KsFLp9tT+OdQu/Gzqd5oejFA5OT6
5LZhS1loNFcJNe5+FOu0sOaQbKz1No7LywijkDLrkvGpwmdHR3165Nd5GZihlJfsqc3d2ZJJ8cNv
NMdzWycjSuolGl1Z3Qg6f+8OQgmDwdJwyOJDVHhT6zdQKZ7TeiCmAQU8V1LI2Gq7fejALTY5SPiU
nzZoQ7EREAn/9ETGqak0XGJv7qUdcPQ0ykMzpYGBWKdKfVkhJ6cjJDO/vK5/r4wAiqi2/kENj1Ee
oq/FovXpi/I8l22KQxndc61QPkWVZalBuhRnGnRqpXssikR50kALX9P3HljA9k4czfv3xzNnfsaZ
QMkR2oUhhz0LW0YVJeiJaFscpam4s0f/2gTd+MQnUA2nW8AINEgo0KGwlDozJ1Zv9oJvucOzYVcG
Vt21qxT7Wwcgk6Wrcv/eR65bt/Xe07rjq+YIrrj+CzNYGjYM+PL67qUH9KIGQgN6gZMrl+w7V2yY
yBGiGQbbC1t93QMnx33QHwEIZeUiawnvcDwxhh7mpr5PkmyoX+EM0jVc9FVc6F0A5ff3YK1+8meR
+dHoK9CHVg4qiguoANW4up5sYQMOCJk7hozyBchXlNCzyS99tCSm7AhaRwGJTfO0B3Gb62r7W2KF
pwxFEha+cMT4IMseykgh3KKJn3TqNOmvx17rKruik4ewgG5y3Z9QPtzM7oruJmHlrJNo6jlHIqbq
bXgOCqXItgFrbHB9Ml/34R1HnaSjlFwnroLZKgLEn6M/7FgFyq3Qa+Rw77z/YKo62+d6DZmwh7El
qGYAYTxfvUxLV4hXtZWaw836uupy5be/9ENZdX/QGw8mdB9x36vi8kI+ztqdLlH5jbY+dWnOOh7k
4kfeFAaolovsBkp7YAPYM96a9wMy3ZKlobAqK8l8sMKdvqKu3qlpmTNnZtqxCUI3o6c4Deg4zfNP
jddsW9W7QtZOad3UbnkfSXBDHFaxQCwBSdSeqASUpHU+dBUzYHEnI+351O0OWJBfDmWNBpPP0tu0
bt+Z3UcORTaz/nJqExk6rD6adIhsO/NNROA5CjAB6LILbeAZJ4cZQgxJgJ98btgl6VkodddIodna
iEWvN6IRobXXbTvtWoRMexdo9HzmByDBq+4Skh2VncDrqoqWKTfEjYERGVu+GIRJotrvTVgKpYV3
sMwK3w/5BsCGo/2lyLGLFJ7aNyoO6LdDqKWrGufeuok3F2NNvExdBu+8pQD0nk7MSaKEi58VHZ1q
wJCwqntUxyny2XO2WkP6YxMgO8Gf7lV4moIk/zOfamggOVN/PdDK3awfG7SYOJP2GA5JBu0j78dz
/sMhx9+VfyXYi4pxlA4zt+pxBiX+LKoEHe/ilsBw4DQSHvOtYnGtRwUlB0qlniNzvyNjoeykkYxf
Sh3z46BrIK1IHhaCmy18dGncmlE27ccZsewIqUqjMd7vNPpSKrEqqUD+QAsau7/gqTyQnRDan8cF
g7IZpuIQaby90pyt0MF460QfjPL0VzOI8nuvFZKKBpFHH/+q7WOl134XU4zoTfvGzsz5iI3nI36E
HzW0TZ1M0hg+UAICWgBc743dA/ta3IDC9GU2OPxZ9TAEHfWUPAkp4DZLYNF17DG4uD4LZ351anER
Unu3PIiI0LEQHeZ5rFsGGT7Sn1Y9l2lX5Znldxs+OhCRsA6eQnoek7rTYnAXPMCXBO9fWN6Glwd1
xyeDrJfVfDQUT4Un7ImdUG2bU5N7w09nbXAC8Wd3adfqvtkizNkhAaTK6DKzCk2GrslonX060pmp
74zDfV/ojqotdPj2qGB6l7cO2uWv6Eom+P/JUjf58uWaQyMc78ZVKvJvnZkZwPYbpnPY0MYUsKBt
v2mAZ68Z1EulecVVlqAoZiReruzVxXcVATuqWEhe4xG/G3mYOv8pnLweJl87bVOR78XgMYEKlNHh
Rn24iRDmoU89X7u7eGywR0FUImN7r/OSJYJ1/Lurk6G/hhJv/+BfXeuXoFrUj2qID9JBfF0Xnyy5
wVcJwsWxP1mjF19vhSRDCPQTFVL4LIvFdF0wbFMLsTR3phWqyAfgsbbdYgJsB2Rh431EQhGggsbj
WynCqduiEZFPyuAKgTe6trHe4Z6sTsyXHALmWGpSB56/iBjcA+lyiE+gK5OzwUf97zq2G/XXAtwb
m4/zMFwc0KYwi62FFzw6a3e4BOWQYllaTarJXdMVpDN1VI+lEIDWq/cCfvVR5PDXtAOTXCs7HTN/
8brj/kHremCrHFfWx0Vm1SEI5dkSQbwCxZ6nrdypmF0i4PPU/cT5NvqkKps1sxWrZOcMGRKdKKTt
LzWJ8jaDZoPmU1gtKjV9LGyzK5o2lQtTgywm72UhqvtWz9se4su0RuXUrxqwkZHXyymlZMn7XTWq
Vc6/cuO7rum8Rcuz/PTZ6UAKyxYm+qxpGpdSmH8SLXvKYqr2hb8blcR/3pph5ZITFDCyoONBtTkc
FFYmePed5EicFYmyYQIS076CwjTdhkXk86u61yxPeCRxpR+v4oe3BRYOGYG1u+n9TGjPrPtVCRGZ
rp2QoIooADlOWLDajC5Nu5kWLLZDEHe7SPDBYrsUHCF23TB8gsI2I7mfk/WLATQ17yGCiZnI6gYM
sj6C1WplTujK0HZPeLAMbOfzLhP2Nz1LupevEO1WYLnmLberJqSZXgT8SnQJFdPgl6r9JivKQq3j
bJZJ+VSGbwl1gfJUqOSz/z1YGGvBtqPDncJccNdzPq+1OJJDfM/WSZbbj3NF3MTbXlnqtw3dOgd0
yND1v5FVpL+O6nJ4wj9Uh+000m1g4VA2Stb4jaKRSE0UXVffiSgWiJM77XlI0Z7mjgA3K3V/bMbV
zSUZ0t7mDf8J4eCYkdNDxlInBKfYorFoc6Y7alZa2HjD9zp0o8WYjIM3wuQEJ2Dxg/f54P5TXO3k
nQVytT7yQvemCpCijN90pwvTumoM8KIj5rXSVkEPBNY4c2r3+fgAWtPSAlP18HExshH6zYASyMUw
7OafLt8aq+JlwaX4bQMweuJCKNbgXOCw+WvNqzllc1LAcs+BNo7BMESli/T86AsWr2VqAp+TJpPr
NJ1eel3vCzXWBh0H67gms8rbxgjnYAHsSNHi5wq+9nFBWmRCOp5tg12pPtgP+NkmOdbx6yeGD/I1
8dsJoqPGM7cRxRyYqWN9NMh/fpP/76dS4C0DqWOAuino88d1jjZ+QkLZcMaplX8/emng5ft4PxAW
ixkUFhlfRdo77SjZzjYvkRwOVu7h9JBY/NlbDwZglXyijOUM+Xiu1D+aKVZa0ArXFmCvwC+aHJya
p0iBu9yIB9rjVBeUmypRAPVNdw2QycmiExegNuMZXMLlI96OYt8ivqiEvqEfr/WFigFPJy/duBD3
56R8ipxcgrzKgUS0L15P/0qsqPl3YreP1nf3k7XQ7W+UjlsQBCiSov5zhiK9hikrH+mT4t75zAJJ
ormEVB6BfJFQfKa/OgJ+q3g1v7y2Cfohw2JdNUCSo/ohI7mCdDk2WucojU/IdnkpRVquJ6QUsnU4
ZIS4pd8TdVTxGuXO+ikIVmlwogjK5d4Rq/EVYmnI8u95QckhlE7Motguf3Yka+0H2vQXUNY3CEAl
Zu+HLCVDvjkl4WYIlAjCsZ+/8694zCHQAIiPteF0vXECSYaTFC8icBltLY00ZKFjGgJrzIP+uRk5
XI7UphzCxkaHfVDPjTy0WUEkA8M9ND6Z3PjtqTo6oEHUJjntjRxztDWLY3LRHGtPnzeMv+3xJXZR
e8t+nCITVIe0ptmEJ2zxUnS1+KTr5qykKP6LdruK2IpVN1urzRGcu4/C0Dh2twjfayu0CWoDe9y/
G7f1u5KI1lljAGZymt9DoP5MMloL+f8B44o9/W7DroAMzX+BN7UgKK35dKF32QIav3QsvH2/ImU0
ayzW9ULY1WeZfgQjXXlG4DJgtixXvRQCZdqlPOEdM3yj6HLjxEO4VjIqJljMZ/oKleutKFCXrJnY
67h6yz4kKAQhChPmUja2cJfN5+f0Ezl0wMVgAMR1U44UHmP/7lfv61ORFeesaoZrizT3Bpi1FAB2
WnXlBV+eDiGVvsWqfG8exwwTsK1moirKQW10Hzg/1Oy436D8kdD5cuka1zv+DDgYEx+CXoCPQ1X5
Fq/miZHXFqLnnBRveUkdaaWDaOspHovx2xcnaRKVWNxNk4ffYig+gt9kDrQfXUDC1mDnMzYDkVC6
e6fLBg73xQGNyTcALAdmsBnnrUGLKxUMEFt5YIKSrEHU1Nutr8F9RKHphV1yDHeZbxdvTQJyb93c
I35/NQrcmduLF3cN57HODlyZkurJHJvIoJZPowHKTRmVtaHfwezU0q0uvdkanFgRBmDIHRGLYUq+
mviN6vo/LafK+hOSWB5qq8CTfo04eTu4W33hYTKRXuTVIHXbNX9Mq+PLr/1i6cwXg/oNvFJlvGen
f0Abt3PojCff+biVapTS9tYgoBn9typUwmWCMpJdkGdv6rpybii22XbWnU7a3ocRTJk3PgHO1n+u
/TrliNo8/uSp9qblxIy6k5ushtteigACgjlwHwLoWaynCvNLfKi8TKmZbdpBqOFCxQj9FNd+uUpt
wWA9MVCks2tVdX6+BKulni+KS/zzPGwy+ozJbr4mAFO9OjgyRw0ZpmbY7C+ojHKY7/7zu8hM5yV2
2vKTj6vxOrub0wfKkwbfDhSyCtb1shVN7NBsPIg1IxcuU9gI56hU4eUi8sLU/KChHGFfoSOqNx1j
lEGDMg5/zd+cOzb5IPjcj6P8yqr+7/+jLxzaKlS55MJAjTFydxhSvcdr1kKqi2n043gvW2r9zhkW
rEZXOqFCu6ivrHvyciqq0WN0zH2QBdtv7DMLnL4EG/WvIYAm8jbsjMC0zsbsLo+TSCnxZRZcJKmz
9SgdY5HDww1H29FTekVSF3pVc2Dus57nkw2XmUlx03yJT5nD9Wjoh37Ht1XzFD3CuxkFzzHGhK7A
4MoMFVC7wpK1FMqXusNW5e6qCJ3NTDXiaRA0s0SaW8B1S80A3BSuN+O4K6HWv1+mGCMi2b5TFFgC
mtwl9n9MKWo7/aLa/Mc/ry8SJFIUKidXkSv35C/N4eA9XwNRrv1CR6D0l9od1n/r5F5a1sCcxCCJ
c+GlFhqqjttdNoPcSl4WvO7rovpKHA9p1DmkhlYjmTxnDQLj+vkq7kH02gIOTfy2dR4d7+TVmI8/
ZTOr7vntvsuZJlr6CdX1ol1zY7WCX2CKXFi68oBucyQdp/SH4M7dsb3bYRKAplpXaALpiF/1/QGf
/lhMlLXawe4e87RKCp8OcT1VYgJPx4I8+SVDgz77V4h92B+0eosrydJXqVwcMhhaUszQkZpRRetY
W9PrgBHyFylFyObXBsXsvxFlDcx91Mfo8YyVRELmEv+CJSpN/e7hEJ83kl+5Me2tn+dPeKaLFFlB
Un8mLvxIu9xYQVw2o1YArCbLcn7+5TiKCEsSzevaM9Y/MIOT2D4ZgiWlqd96lTO5j7qad/TlIb24
ptfhGjYJJ4yXDAARxW9Tw43RyLaksDx2b7/7nq3L7OE8rjuYR/CbSgoPe7xNU3pwEObebBEucepf
hZYl7eiobfggp8Fqv2BPl5nPCBzfHHCt3bnX/fo5zvoOa939CCpJzwF+oEzSRTC40lnY7fr8N+LP
pusIbIu9EioIpT++rfJRJwq9k+9L2vUf7BZxwISKG9QAX8owyu6PFuieNdvFEONfc1mG2h+e6I35
C6bJCgx2I3BphY9OOn53/5g2bRU7/5LTWqsKjLHfnkg1CdpfyeMmxdbFz1dSSP7CTqsE+nzWXCIo
gUIAtDCmZzOVgVU8WAhW7/Cs5S5JZ+g7V1Xk3gVeesjVv99luKGQ0r9lIYV74RN/c7d9N6CLRT/x
4mSP+NhJd8dFK0YyS3Aw+RjXJ19ypfpTSNxnWx1D1bCB+imXw0pXYSPD0YmkemwoavYayWPGsdcs
6u5tH/TFtPiInCbihO3RjNaxX2RxVX5dAbMVMWcHiNutT6QyfRcfNfggf27uWacneVmV0yuru/aa
2HGQV7XkBwSENnNpzt26j42Aw3XMX3Uu6M2gcBjxhrpcsIl5uJI5zs0XrXNUeXZjKlDG/bhSXeJN
TCX+GojQvqdLRfl1M8tqFEEUSsWdaGYEZBM5aHycppNlZjsRLIhlu13EF6jrJyRHVIy6XgZ3drCZ
0jKMdenf5wtDJpAe2R5oKLkWa4Qq02l7oO7iWA4wmoXlNeo5MpCaNmLOJhoaGyG1JS9Vf0LtTs7G
UKEJ+coGWRnUxRkydxLizqfROjQEAS9Px5bHaQzZwanOBe86A7n5nIv4UzcqqUavnBsmKiYoHH4B
ruYaI6qJeGJ7O8iYXojgi0hk8lnp6hFL+dncVbl6vbmxmvrDCr7Vx3ZNQ+2mS/0L83/eRdFsL85Q
oQ9Ao3LJOZPC2JkJIh64FRuv4L7qSbUDU7LppaPyh9CNlrQNIYH9kUKyDBnjFYNvwYmZfFKUJeBT
Ec33c/zBuyF3mqrZvr4KiY/aoz7MEkzs8smQaWqKiGIV6xjfhcUEHhhLnw/JExLvkuXccC0k9X5T
zkCuVINXIzQDHyXYW5ZFSXTHei1Z7MA6PSCaiJHkVWq2l1u08WJPJM3jiasLa5nppQwKJ22h1zpE
NJNI2Ymq65vrlAQKNrLb5ybTjzyC+jwI5p/g973YDs9GZTjXDOC21HSJWEofvqsu7vroEC3wNJIK
4WyyghOE7LYVc8Omn2O1gx48sZiScO6+f+Z2ES8rU1dI9o5+rc+M+D5qZ9iI7q0ok8sSfKB9MXqV
xF/OciarijPBSJJPGD5vN/rQDIZHKbz1S1STzoGvo11ikrwGhP7S4dA8b+Hu8fudPCnL6JedVCWu
UayIZbNmWfJWGXPJga60eF0JRxx3UnuvSIsjcYwHje8B9u28roU6xt72NQmnkljuXMk/oEyqG2yB
YQeosN36r1JZkbwkUqddhjRj4724snjIL50HIBQ3Gz3K3fO5Tg+nrvmBs8Tim9wW/QltWLqAeH4z
f5rW4bgjHOfuYSHTLK4TZsSGIma97NPEo08a1UHOabrflU3RoPoubAkDFJsj4bcgFoC1rkg4D33m
rEM4BtRlpmVstwlI+aPRk77tATjf2Dx7oor2cC7O7g6PvmptqAg1G1gTFlTAO55UzMmkmhy67Cjm
f0aaq8Xt+igRlWaStJnga5glEBQJqEHw9PeTDA5Ex2dpVC0JMQFkKt5ujWtxyhpyTF9eq8+q120B
OdkEekJWogiiUrz/JdMJvaKBRMHjrbywSZvN08UvGa3hQnTpYwEKnhTNLZNrDiEoDPZavCsFBxjk
QitOWt8RZ/Iw4eVditgDFqv/aGQqxc+X77ikU+ivipP6eHh1epFnC17E4PXH4ZJD9hsHOQ8rAWIL
jlQ9Xpvji77JRM4g7ucIqGqQ36fXg5Rbr9UqSGJvx3SOiYrzBSeFWryIK3rfVCb+zqPVRixWYo/X
it0dj4RVc6Q+SVSY8irZqgdV9c2SWm3pfIRLIVcPOX7leq0BjRqvMtWzRe5Epdj4Q7xaBMeMHlTZ
PpRXwNG5LEu5Aq12uwwjMbKj1sS3vBA5W8dLYmNJmC6qE74xf5OCG0KiCna9Lxqce7JX2+9FXvBc
i/Nk5Y7HvkU6HcGn/uSsLWixPnFNC63qDOm3zWsj9AkYbsjtakY/65Yiw8ulncWOfks4BNd+NPzp
jV5jYBGniPMCxfO/VmOIw0oz/ikMpLeV3m/HfH881+Y1NVnTLHehaC80k6fA9+QDB2EidoHri3U/
sGf1iklaok2vACUvzfjSJauSXcbRQ/o8Mp7NsoYLUnze7sl1GHDn08Mu1PrFWwpnZYdkyr5hqLTc
y922LYyb/R79ZyiqwkFiJ/cWKNJmmh9+idMK+u7IVTLO/4ihvRk0zUGHOClhxGZfkdZKcSmBsZLD
XwgpCU9OMlAaK+nkWfnupBZPh0LMSn53QpwoY1FrqOgepZQWdcvDwfgcG9IV1QVA4VIwN0S69NUk
X9BCKCxGiM9JS0Pam3rA+aSmvkbmy+Igf4FZDjhH1UfiNUfrZM9WXgNS2rtFKzRj3okhlSqVVNVL
h8P1S5+1zJpijwYUIrjNvwpUxo1FHMmePiozGGaPkEvvYwiFfFyBEHJRhhM4BhzBc2cO1RMCaPwi
8pVQJX0oC5cMSAqq1B2NyoI9o42Icpctj48NpFY0AmLY3oXNoA4ul2F+aPqWVKw38mOksFagLEhY
AD9vevvbOJmZwgt5FrN9sjeQhgukdhNv4o1F561ybb688RGhmV96GjcGKza+PwtttfIidj1CE3LS
QKomgOSJ4u8QzJ4BqtRiBIsoku9PsChcGzDU2lJ2v86S11MAVOokEIv0QEpZoLx4AvmWm+MGsBIB
jELm1TJW4xMs4YHOEVWTbTb27DvaoJvRA/wOike/DjbO4T0HPkuuzMMTbQB/lt3seSd70UZyRUDy
z0EHKZ/PGOpxzDRwe0ru9lcmlnFsrdklZCWM0FGJSqapGNkxUUBec9/gO4Ks95Gv82t9jLbSiVrp
hoB/o0rQj8Fav1BhLJVCOMk+pc5taPYg2zHFLl9W6FK9lFO3LgG/jd7GB2wGWu203C+SoRuIqgek
tVDWPaN1ZhKLtAmOcelI8kGgxJleIlBD6urHf0j1PuILiEguh7h3bQyuCUxGlGI66kRoFYACWbG9
lv22UIrKhGMsjo+W2VLWeB8IH0+s9MAGVZ4oVzU1ixzoaI7jc1etJhfGRgPUoDpTJvXESmH/IuxB
WAZnoRjiHCfceMCK5jqyfiAg8nWdVm2qjJm6gTBndhtBQGlsziphr/76u08YO2bdd2Z+irMeF3sC
CdXH8c78pFQphDhFJ19NSc6a6Tt6jKn7vgVx9hfI8neDS0py36pOZ94u/pFeZrEXEgOZcp4IbtSy
kT1KCsrTzhds1Fu+bC3ePoO8rcuf/ICO5UmbaQDbgDX54c29zvU+65KURMArCFI26WQzQWGy0DKz
s+cwphLj9/uUoZGWkN7iJNhgl54V/Rs+hZh0rUyaFRHYtyNDKpwDATFr1z08B/XwRyN85ywkLDqC
4K5h1VKPurLVLJTOHGIXIpDoODY/JdVpy/FfHs9mMA3zoiQOoW+S8U5Zd4wRgXgfiLv9s5ZRdpUG
e1cABCvk4XWD9EGs9pJzSsfzLd4CJAjQCqD4WIuiLgw6vpeXKBIHn+n5H0m2umzDNBvVqJOX4gq4
02GBwG3oikD6fJZsOmb4JyoNvkoSF0NrC6m+l3/OZgHTjqo9HjxUiYypens+buf2zPEfhjb+j7tv
edfMHx/7luzAUc8X9EE9NV7Xsb0xPxiKK8SJkO6ZmF+nKw4nUKg0ub3+KIzUpcCDDHfLRTfySzmm
JMvDmTZ2gexDdPEWg8uxo6vT+vVPEItXa1GY8/JhKY1x41QQLjtCTIm4Hfz5l/i8ut3mEcy/SoCl
coKaUkQMjPdsByjS43Vy7yviKIhHZDPStsbT7CzRT6qjzeJfQMwOAF9WhSnC8c/MTsm6TinjfWc9
w5u881n7fkqSTjBCBGlkLU3nex1Greqj/NJNkmrWXnYjRzypVkIWg97leEO6XN4jjuLwC9gXXegI
ZR5S1uDE0ul9Y5zQpmZ7soFzdU3SmQd2fdutm3M6q2YPsGumWAzSo/4kDiI3fBNhHhPqjgHghxWd
OvXK61T8k1Iq+NGOQc2Nt/YJC4TenPL+gJUeOvB9YSu9fKHN7Eo1kopjaShtvT87KZpJbPR9LvPa
ws+CLH+ql9UyTtIC0arkjKKpFDAIshcj6O0uS4s6Ht5qvMsvRjsYAedVnBSmJ3YrAnG8zv4Dp7pj
QtY8T1VhzkooIUNXrDydez/JA6lQhXenwhpmrBKSgeeGKnbvqoXcpMfbqjSQ6/eG9djO2KI57oZQ
LrGtqPAxfUKMV5B/skgpyI300LVOhSc8gxos8HpAjQVnLEMj93i4yQ5fInUNt+UhlOyYr3ang/Pl
qDrxCO4GsZE5MwHa3i8sOqFtfvdWua3noHqgnbup8UZnHwq/Un4Oj96u6Na0f6yL2h1WjeTQXltX
x19emPOp4DYVWtaC25I7zgIjNAnmvn53nb9aftVxSIvee/Hz+brPfxq6vHkn5daeoNcqtUGclSN6
5U9X1OC5cf5phNvg1mBrvA92spC5i2EHkRqYLAhAjBBJZobLjyfqq3qSi2uDOwBRXY1xjpCefdOo
BVnl2I3j+mznMIi1LUcCdkSRZ2igquJERXozMGEbfGbr94YrDh8VgkYASDxSRSIrkDCq++W/sb2x
4mFj72nJp5kindvukJf+CY9I88ohln6NrPktja8s5c8E6BwetQZAWU0r7hotiF+Iodw9nYLImSjq
MBWe7lpR2AmZvK8CXbDky1jLs1IqjnJ8qYtAPvlFlzRFTF/ThCs8e0AS4t4Hb4uW2Ta553xgKOc2
vcYi2F1ndfhMDBR4lBgCZ3XIvHfAtgc69xLxmyZXd1jpfIhVj8MohILjyt5/ZhyxcHtgbyzdssT7
YJ38saiVLk97mNOAgtHaoICGjSeBuL6Jhf4YuTkrHGvV489rl47ai30ceWyOB09sGZDFk1RguLAo
/MFcoBU3PUukF6faEIOikQiA4mPqNMyS46uTMC8BLUxzVNuq7Tgp+G+zNui7Y13BD/EbJAgkPtjM
kmf8jB12Zj/SjzZUFZnmRkttng/6j9v/dbNoNcEHsx++EGXXYDl1Qeb8ZmEDUusQw0AAL+aWgs63
rN5A557sEHNLjztLE4LlbJF11tf+qnJatd/dbScophPMSkAdr3jLJuxQKVxwqPDP+fAehdh8ybwQ
Rx25ApIHuF7q+NEu1IsECTwmxDfi5xIdxzse+717zttrAfXEP2Ab7Yjr6m4+4/kighwYB6+RH2Ip
ivcT6uKsQKduX6fDPIZ0vFPvEbfZyUJY9xrU2PrcIoIcrMO4P4oKlemCZikki7zb1oksKHxm5jkj
BR9KriPswK2SM6pf/FFWEsBsi67coTSII3hP5+RkogV4Ea6Rx5TImjUEYrwbvUuvVsOFMHRZQ7a6
b5YXWoZewxxrbx0ELVvVRDl8PyD0BxkKi2D0l60g8DGvZRgkuRQeF7PUIARVp0vRLSLULJj4IxwD
rEAdEFWOzbrddUADrUr3q++l13K3Xzr9ntWdVId1GzYls/uFk49VC4IYHnaBTTPFYmuexKzx14/J
eekJn1elwA0mCrvyP7ARxPjvQyVQm/dybr3FZVU83aY9Teuv24LmxXWbh8E82/+M0K6fbZF6jKk4
orkIwSWUx8XhIuHlLNr4WDuWhSTTwVukwkKwi/ODX9eD7r8jTQ7k2TcrNaRgSVn2dmnvbiEQc1I5
xVlOJe6epDWEDVnkyTL3xGKTFygBL+xn2NsrWCaxCvUs8w6dHUHHhXfAIfXy//FvFKTrqKiAlo3O
1BSWtlvfEr5wO1EbMSdYhFG1Sgn+9UhApmxPiQoUoc/Rn1al1t5j/G+5XvJEQzJveUIqnqPTb8XR
7dsVgtXt4x8q75rBJkFhcijSOnG7Vs4m3tWNoiyU5Jsa69PWvZglRUW/VzrzVc43ckNRbWMlwdZS
bY2lH/3m+oy5GienmepCpbK6GGfEITh9IaemACNSbE7G1oqFO1l53MLmbMIgxLQVZhY7jqgzDswZ
9ON/Btd0yguFYjLM6C30nkI2IJ8fGr6wZTzX72xfcCGR1++vxoiFgrp4cWvL2F9I0uKso98GbpDv
Au6W/Tv0wR7gGl2NhS0vQc/kDQ4gZqc6iRmFAuz6xyL716WwOg6d7BtgStYtJOSMqRYgLbvPeudB
9Ff7QkT8iDa29iBTYL1/AJ/kQzOXZqXkVhZaQbqWZ9PagjpdQZhD2YZKa63M1wCuHw3tvc6Nf9Fk
RmNK7jMcCiSBshhhqSvf4VOV6/Bc1CKOkFDrDkvew1MyKmCGNO7ikb6vaGIeY1WEhkZSm3xDdLmZ
mehicypgOFdbz7FYnlJLIE6NpjynS7kHijUKL9+JIeY1zyWe+TgCKmIVu1y4PhYKQ2GNGKwpO2un
fxXWNs9fxLxyvoAvCJb53HNhfMT0xiOGy0TMN3XlqkdyRgoi65liOu+M3/uPiTJCMyUhwk/vIVfX
2LPFYma1hLTceflAaI8Z3PoVXD7kEEuXxW+MW2cZpAjsgEAomxLACkyJP8DzTJfBybVi5QVOaVEK
TK0wEaVtyyA+9vTbRykF8PCGpNwLkes9h//iF533rq5OfQXOat2yIcujm8rqwFzvl6rt/NdbSInw
Zf666dWEOX0l7GlxPbCWV7GAGMi1GDwuL6eR9LV2PayaCdjyME4hkXWJrmz5KFxcLb2cgDhvrY6a
iuZDo2P8pPSnFzs7IeNQld4NKwyoRZcRc5LnRrJobFA+JyxjeFmr10oLCLh7hzwNuM6APMzXmw57
STzRZ/uENwyHPE6yo63vxQUx77WM9lNm6fQKIDtr1Fa+M40xAUVK+fhNCiy4PL5n8DbXDnfSNx/U
kOxiaXex1+GHY0GMHnEz4d4yo8YxsyU9Krk8yRWEP/V2eLXCZhbILDcTr+v8u/e+hWdL5IDsCgJY
Ls+HjWjbnFthjYO0tDnbDvMzahMscCG95y0aW0JHCLwMeVOAoCUpKKGLVOUeW9RGv2h8QI2oG9lj
hgwWZJVmfmATUBrCUWsV0gtkHON78aepf+CajLoof0cFkwTe/+h+p/9gX4/DWNxmasWjFvj/Gf95
adWX7yDBTHUuy2oaIiP9kOg3HVxssOw8MIzERkKC6CHT4oGJjwUS3ATm3/WzgMFzw7VHs2fDJaRH
T04/iQPCPZO/Qic1hv7/a5r8y0kXWXRpyjCOOrRpYYhBUJ3Slhfw/B04BKpCFRLXuDl97GJXX79G
HBh2qZ2aA+mVSM5GT3yGs6L4yMQ5A6z9hWAHkq/IVfmmYUdwqMNrr2fXnDpO174DpIisFw8CZ/JA
uV3Ood423iTvUL9f0Qftkl59lu0wffqksleFNR1ESyCLco4DukkW8nYtboyx/ov8Ll0TptTHFWWF
UYaRUoV3eAQ85gnyLv6u4xCgcLjYNZvBsMCpRhINeiv64Uupjww2aBtRKmLjmxgfJcX8+pg7sX5W
9o81EynhSy6C4xVkic7V7BJrKTslRR7akNoCuLg6TiM57XlAIfcB7qdWrMDtbszRt7WU890PHYx+
en3U77Q4hD7EoxWGh+cKUaAgZw0xG9lgte7WcLdD7/9EdMI2sABNc0E67fXtQnDI58rq0BirUfIy
nVBbv0U5oKlhcgVRKvsf15oOjIMZMpnFexFPJXx4IapvyMAlvuwHSUKLRX5im5yvhUJXV3zHDeXM
S/eajx0f6ja2VHbv1vZmaO7sh9WeGg9MSm54Vh9jHSYAoPel/ruICfkGPEZEYe9hzP6T13JHnYrR
GkV+l6Bs2fxr1fx1GhK3WSjhK6Sk1yvQM62YeOIVN1m5CqtRrNLd0nN/8mG60bFlXIjszeTx830z
gQ8Pix9ab2W2HUqRs+pA9iD5162cSgm85hNWd8quP7ivdHqRthjpkXI3perqe+S2r472FxX+0TI/
1tKoEXTL37uVr094EajCwrmOItgWwUzWJWfoxhPtJmt2MJWK4IEUkhRTqlhb99/eCeWUmzSvyJ2w
bDWsUD7VJODSi2Y6hBz8N7Z9iwac217iTqw5j2pFiP142n+Iz0mqIIlj7SleaYhZ9NrWsYNNjG+O
khMhgJ5nJPSnrwpuDT6MsGt1NSYFBUCZ6lQHnrlKOTBsDq0usAsbKJoup8CIUtuckXgpfn01Uz9b
YsyVWVfpi9dw3MPTW25lwGNi2BPcSUCDRJktLELj2HhBvh8BUG4MgiTbb213V/0ThLpuKj6dBUGC
HxIhVVwQDPXFfeyoAwLPF4KBhg8mZHynAm+aSUH6NnPZQMwU11IwNtuX334bYgB787FLavq9V9Mo
UzFbAwVhcuFzTMFt5acIMT2DiBxIbFHAZYbdxuq57AtPfDos/xvXX2F7pO9coRkownKFF836Mdtr
lXb+jaKdqYJE7iqB+43AnejLhAM58LcWmeizftC1PO2NzDeqDHO7pIyg2SD1onSVWq4x5bjEyaW/
A4BE5fx5WNxOOYloXnNaRMh9dSUCc0sE99z9i6p1NG12Xfiy5r2gjEQymGX/VCkRSBCpm7Jv6osJ
vtK1gDnSdNFVdiWLLQsw6szXkkYRoW/DBeLiv6OvjGYt+xOIxt6eOto4wC9MPoz7ETSX+szafsDX
Njg7keomdbLOjzfLehcWWUcSwrpXF8czuzOcRwEx6APDVdI3WMpwVwC90P/01B9jTz77W7i9IfDI
ZgLXY6y+0Pj8ucF5/RN2+Q98UYLEzP8wLr0/JI+WCtFNSMDqItgWuw1KM/cgB5fnMt0iY+2E6WNc
QiJnkmuA8cLqNQBDFHjZhsMfnL/eScDiEcU6Zfq0fwAiWbXfh1r7O94WWDsNL0TK/k1GmGzeZa7+
cGOq9tkQcdsl+b9xjvEx9Cd8CwivODDQh0BzMSZJCeZzn0v2FCiVCBuWuo3xAQ9yCnJSAuEMS/J9
jQlLYwbz7LeQqomcJv5QbXA9D+llPmexLMAVbWl/BkqI0MWYsGlr0MYi9/VA1WIPHkDHfRXXeRzI
SIktEeKm3YEKWtAtcAQpjKe8J5QPavTQx0ThvqBgkxqcOQokAJPda0oxNXJkPQu1S2M2nJoZQR+C
ghLK9g7yBgZ8fagIMJU3cPPfq/wJghSGXjCG0tgUkG3WU8o2D3RaGdSc9VRrDWGt9A1Zb/3FE4Xs
0qSJgmgJ+3SpFspfA+K2TQLaoqfFq80aHlMNoGQrFER7UeIIAznsS1vUhrugSiz2dbZM69PCh7+B
V8nRfs6Q73is0yreFkITXhVN3mF/QC3hS3NUBJCHoL6WVlAPdjah71LKDq2Sb3SnAxFRUG6/H0Br
UYyKkwgpPU3PcX+VHJx6FvwcACIez95bAK3G1UxeCsRIRr4ldH8bb0gbxUVKv9IjzPBe/BATMzxq
BLhXw7wcLOrJLajNynvDSyIgdpcz26PzyUQt3yns1W1SgGHgHrxnsQvhlMtEU45NP6S+zY0+hNQp
4KrPRADar2/8/jKo81NvNwuIznHBsUFrsc82vB7Uk6QeHYs3wsdLi3tO1f6AkD16HAQfeV7FNRNv
R2skKz68Sa2T0jPR8UcZwStCnUjAreSW4IfRXMzUv54Oo5DRem7Wty6doF4YnK+wm3XG9c3RAMVi
1Hnc/0OA58kK7ylgWvvvo+vz8yjTEmpuoUjepL1w8E5sZwouSR8GWM9wsl5H30ATvyDFJ1Rl5v1M
iLvMO7QG4xdLxb52CVJeQW9CRAV0/KA2tlAKK6W82EQmswNH8cohXaSX36XQIiVp0yXQmhDzh2Oe
awA0UbIWAkujQKQBYeRaJs9iRpNdGLrb826qeBR0ujdoVPnDGiJJLAbbkwly31q636mpIxacZJBp
oDl0YJ8wWBZ70jM9GiRHFH0qqqZS9ytxRCEi96hymAw+d53F693aR6JtNjMqHzvfXOQD9rS//pmd
5wnB7DRNfUS2PJPVGM4ACXTnkGC8myJS4DCxwVguXXVjiI0mV+svT9O8rjHXxbsumzh2/cQqJogO
kK2qalcCtb1JcRwF5+e2UmitoDR+zB5zoafKVLD4PnUp0t/VnM3LyiRhLQEhvx97w/YJAfNzpGQo
bFpctXIghZhUE70zbU3LgqEFRwMS5Lkoew45KFIaoOmYWrU+7gMQqH1jbIO8lkxtQ6m70QngGkPP
knlWnyEhUV6e0XkNrGbWk9SWCbvThhB0Ao4iB7hzlHy5MrmT6Ov14CkEJ1q09sArYt+/iscMMtAr
85YwAy3Lv5wrbDPcQiW7M0vWsUkY3hywmFzluHZ18SuMRWVm86bAHGv/KcDUNFFqZ0o09CXdAn54
eXEWHvVO9t89QMhgr4G2Y9wiPL0UezTrc6MbSRO3D10xdTsKzbhDuAFejMlwb9sCWGJPK0Bdv156
Xjw4qEg0pyXYYIh0oVqXoDOZSLhsJlkfXP07IUGj7gUwUo7u8Zo7suB8PyMkTvMRdSzhYJ+PtwjA
T2FCGVB2H6rUnkNYGr/WEzUIPJa+wV1PtEtElEYeJiccK4tlsBGPYyH8pbe+zb/zKWHriMg2qEJj
gbY9KBJQgeSaHcZXlXvtrVKisB3hPJ6VyQzoZf+KKcbDYeDTPB9hz/0/ZlgW/80ioJRxFG/c2WLZ
/RWgvfzpLrwMBRKnrKB94QKX3d3zBdTLoOCJsizfHE9mPtBDQvqu8kiqsHOfZlsv+j5BZQUU74IP
nUfp9Pag2bqnKkAYQ3ckdqct+anQEF6lSLpAqkWOKMMcoF9Fn85nMjDDJcdHX6LJez5Nn88x2qBk
e1g31+G1hj4H/UxuQLHYRu6/rjFzaIO30N6WvhpjrNE0MRatyAtKN4wyGPQWea67JBQV1XD41wOW
3DAN5oPyIKKaHaEYF6Gx2Q7/rbCbdJqPtQBkYLPLaPqEZ2m4xkNYgSjYQVTJ8qjt9oYXldAct23K
RGGV5FonLcGtqTomFqnxz+BPEnd0331ueimS/jn+iLQxY33M/beOgOXZwtqtK9Ft5Ss3ZNNrwFvs
WdMH/UQvcewc0CZGeJCOTix52Z/p0Yk+Mj7hmzAgEcBvJOZlLbo7nIdNqKwPiP2NEhFDuMdUrVsb
uGBTazMz4CsbgdtCCa4Pjw+gEpaSzW3sNaSrjvlz54KKOgWCIP+MtELHFnNoZMxMiRzAYiW1/LPJ
1K2GA11YmpzziJ4L0pzLc/gYk/5BmjuHA1yLuDFS4a6LJysOl4JapjgQOcLrBaTrosS5frars6y/
Voopp9fASssjYfWVKmqa6xUf+3tsCb0bl3kSuoWui3yLismh+ZQtfRPEe9bCtLEN2iKya7YDxvhn
gWTvpcK6slmwJ8YVaGAbMNxPSHZo4kcUrCAGN//9dwuHUGGvjfGhILmamN7nZi2Qmnoe6LG1w38c
K0WVD41VJ9reaI93OABLbPzmit33WzxR7/rFrOkSdLf+AX4NrP2pdOqglraLF+ui1li8+9GFlsHQ
zfLIFmLXJUoBVSJPjfDF7upSo9FDPMZn8tKyoRwLM48ZxYR3EyaCeSh/FAHqzKafY59REnjK/OXj
DRrKSF3kZwcGiKHUyNUnyt5td3E5vFIRss3NukCU9JCN2kJzfjmFCQtKZy10d2IBwwX/ltEbpvGK
ZIU8kueH6em+1kFQ5R6siatoRxlZ6RDL+sO+Be9CX/vI1NvDDTbv0qFeestzTnfSrlwcJzZIhIfz
OvkcgMp7eBBxkSHwmvYPGi6wSe67BRQG2FlALfoumQl60tI6u99C9rscWclM6pP7IDxuKwSCBhsm
gvQGARupGInPFx3QUegfxTrcPF0QvG9gfyQIpbRVxWKzvv/kmt/3w+foHQk1B8Mh3yYjyeIT0gmK
e1TFMCvaFNXLtUG1hVqxlqINjXu+eESFfensKdFYV9apwnIVu0YVozWVJEJ8K2c/4LSelK5jjZ2M
sd3ZHEiPyzO7IedtgaUV6u3enNkJQr1lMpYYkzZ4LLCDSZ19qB8tBLEZSGzw4xu/zFgva+quxJBi
NU+mo4+Nhm5YksyWBrsUxbvYs+AQMDWk6qUS7zkFi5jyeJP13zJifAdMStKZBS9YDaaNbEyIPh+k
ZWkGy0w1GfiHuxwvsu0lc4i1rMSPsxjE6HM9Wo1ozL0N6lKQsLU/FEA28NBGhijUSnGsO2wr74ol
LSvboVAbqISBfrWLCxE1I3QMSBUFgS8nv/F3Btg36A2/GdPkObcEGsMDBMXN1dlGMM9MZwkrqoLN
pza7D2yrXo7G0Z+3hwRUjd2B1ulmDM2cuZO7aZZ5cyEtsxReKAamm19+HXnKS/3aK4S00M1o9PYI
Rmd4wi/IqTyQHuwqFujocD6gsRNl3qq2mJlJQaDqf/iztMcBWHHIDQM6Q3+zaAVYk88OtDBMypHu
1E7LoDUOoNh81JnTMJU1jc606JLRPL0XAr/hfDXcUk4wDNg5XqMGrJuhqJr62zUHLkunv3KVT2zc
v99RPRcipR7oDlv34RpSIKB+ZYQ+G9xyOfT/2Xzk9sMyevGsmUOyBRDJts9VyjIaDTKQPLv0NZlQ
D3OJU41BqAaEUtl6EYH5UpvMmLrnE+bNiB3bAYnEpTIwq2HbHXQECFccjEWquGvN8KNi0v6xUaOq
yse1hP/LzYrz74285FARjGhXBJO8sdhMbU/3SMEnvbaMl4dmPCh35IGV6uJjU3+gEALsroo6Aav1
uqHOZ1DHfrxfTTA9KMak4P8nmGETj9MKukodQaflaqpFPGWVhVDurCdjtZHxyKGGQ5N95aH9yRNw
q9NWpjDvnEMqVpn6+nGpupiJzzsHaMAcrLyYnmDcw3Ixg9IDgxVdEhtTv+pVR3yAf1Nx7Zt5s5c3
E50H6iA0sg+awQEeJzCA5zmMeMZfsgxXd4T2JOaD9SsB4I3kULF83vElA115YpLXNrW5pwFMT1Et
sM+gSXcA3r6OAGasNgZf1yBLyGmT8t4cpkcWlmAa7qgME9CJSrJC21rQx5nEtD3mxe6lvFNPrR6e
+vEpcioiA/13QOb5opVucgvKixBO5ObipYfN0EvheAQyDeHNQHpz0ELR0ekRKFy2rphqv3VktxlA
QlSOtlY494p0wl1rxJ6IDft75gSWA2wb+8xuxz4gk/X2V4mMgou4hcbtKm20Eo8AqyeX+d6/EylW
PZHyAZJbNCb+JrLAe8SoCj8LSUh6na1LmiCtp4iCbCNrv6iQhGDEmwS99fcydlF7E+xSGFUgSSgu
fI1QRsLj4mE4Q/LIDrxu9avgavViiBhnOqHvAmru/SRir56lOth96Z1eRY0WyexZeh5Y0NvDna2+
oi/XRnn9EHZnIx3nSSNQLNaXObnPkEvd0oeaKnOFE4MIhV6v49mHN03VhZ7D+E3QMMMWtDoTlh72
EFHMAa9J7SM9LOi+jJZCJqvAi7APAUCkNNO//iRIFDXSuP8oh0vsI52TotXZQKH7rT68kEaoXHxa
BiFpgzXQJ+CLGyHPcP9137gkK2/jrUKbxRdEPeCtQJPuesaDbvZHlb4Ze8Zl236sBh7Q2CkuIpbH
g8jhu/MnhgcXSUtnXnHzt+oLgLxH5eKEl3bxymt48Ay2j0dPkr/8ngZmr1GVEYnPVMQaDRbE7bI5
qSZmmUTaGm9aCFsmMnxdLYn9/j6q8Uph3FbXdR0w+x/sQCjKAPVmbu0t9DOZL0obfdPCLyjqnHuS
op20y/4auymDXSGGo94ERs2aH0opD96+d/NCwUPuMJAq9XfgKONAJHMb8awETGCZcQgrZ5MFUxWe
yFb6XEfwLmkLmRoIWmVjhQpVM4pb+W2hQUdzPAEQGlYvUq0azqSC9KHZtmpfNO1aPj6LXRqpCgh7
EQyf1BLM5eLUgPB0r15JfCGLNoo4l98fjIk3pIY07MqHmtKa2jFoiSL8rXYdeHzVVYSI4R1oMGJJ
MwBFKNWRaEg4GOrc2yPZhUkLDQlppuTOmAnjDd4a5VNGORlRLgKle0I4Z/kuoJJJ6yA+S57sKQoA
c1Us8zZRvAuy9qDicXJhKkM+IMUcJTiMW5fm1o+XX4TBXb+anbbxrf/zwcEX409mFXWWe5FRc7dk
9V5D+MMNs4oHlkRbi46fRy7T9+p9Jwexeh8mWYCc6TxglnGTCFxKr+8sz047OqqZM0hxoSKyOYEB
npS97OQk+/H0M0P8T75rm8NTi6RPCnyrBIjjQKhiGcUWJxK7TYWv3hC6mu9zd9dlQ3UFRAWgQqFc
1r1FDHq+O1eji0NWGJg/gO0z3md1yGy0N4BjJLBDsS0ydxW2Y5ei+yndpDwoWTd0xX6WwDT7sr4L
BY2Io2S9Mkow6Z8uFag9WXPZMPS0G4zicUPvUVZhQYFz5sLY6Nd3mEtJprWnrAzwO0QYTaex8q8S
S+3DXozZb45fX6Nb1MrVCjVXQJV2ffwQTwm6AxzGhPRusda5dX8gqoMo8BxvBof0Ay+uVTGpJleO
TeTQhhOIMW+W68plSowzzHD72D0O114MQ7Qpx5NQGuIynRNOI6X/bC0Dr0iAMdZ85qXhYpk4k8C7
pJqNjtFOVoRrXZEN+Zwi8PFHOoA9/fLvGUi1ctvWyzoAIQAWuQbbyg1xlZ5NIrBp9NDbxhK/6SQZ
dXg18JcK9catVNrfR+bl0kX/Zqmvywmi8edh3EqJBga9Q74bcRU+CiUr5hb44GvyqPz3F7u7cEYV
1rkoq176pwjPOREGmPMlnrJ0XwQnUGDjhpe05KLQ4HEMjPZRGAJpUbfwHrWuws25bKKjzWWt2Xjj
TsXMCjOp0MQ7Hftz9qWhiB/bGymEWHlTfrSpilDG4JGCIDYqr0w0VNdZDHPo05+tOUpgwA9xOejr
hJxgJUUFClm+XAMFyaoiNw1cXPlj8LqxY6VN8jADaCW4Xtx/hknzXXVf3dc9//qHW5itV0ElLEG5
FSaW77vLvce0fGWG9IWMSTDNivdtCI8kW1bXavwjRyqNbkMvbS/AmNiuiSvXu9mGI1AVRksfJXoK
cnNMqGjxVYaBxJJ8ZKxNk5gHsEDcoApjs6OyeB+lLAO7dp+O7v0nnEhS5mqFlCMl3jWsVKoqVq6T
6Fi6tP5UbWTI2mvUAGJprbE9DahfygaNXK51tqRUMMY6cyD7RnCF1HqkcU+1ZmhQsInZRlwjskCe
eb1PlOK9zbJK3pydMGxjH5PEVfUlLX/PeI1uzJuYXBf+0Yrw07kZEDNzCDbnuk2kaIaFiDBXwxL3
fdDhaDs2Oy3mQodwEY+C2tbN8Kk7CCjd5Bw6hfUcgWVEVwW9OyLBn5nmS2w0zzLncYLp/oj3wu/1
lUlPs6REmfIpDD6qviQT/GS/rSywocXx5WLbVbIiSjNIHQgLpMq0UfKOM6XXMHV3/bRwNtKK8pRe
P55bj8dOxZlaGTxwvHUqLzmDVgSAlA3LPobOzCQEtvb2dTt/y3gZFyZv9ZyXA6YJoSuzg7V1ndug
EvnOW3kODV47rQDqmTde/j22/4e1hW4Xg+lE4xRyrxqVl7kK3gOEkWHczzTetfSe/9CeJVZN/hsE
0j60Qr+QsiUyWQ2ti06vYNnZTrJ8NxxMaM9ZlBsHfD8pgQTbYXEIj4YgVfslNql/9Qba4w1bPjno
aFbEHvTky9f+CPZoTaMHLJQL+6gMj2djVt0rcwHLel95ckr9yVYbXXq9eblYJFfnDlSXxUk2+Ybc
vR3zjvPCsv/V8L6GY1S/WHRVRbVM4SEmb/qB9oKdphxW63ed4Bf1v9KpF+yjLrqDZ98ZZluwK1PK
hILUkXyhT9pKT/jQtjpb/0b+P91Tek7yFdl6/WL9fL3ktdiuO9NxefMSFT6w0bYTBzbFIgiiP9+K
PHlatnGyYWiNfCO7yEgpJS6JU76lCmZ8mULFb0u0jwYnRCdJNkhKjVJSBSxDKsRQ6c4DL7FXT9ZF
TBMHuPsDrcD/IYBNRIOINZx/sjWp7st++Gs+bdgZL4zVqAK3nIWazqbiOloZuAPtbUg5My5ugHq3
fXXzrRAP5ynQS/+FuUAJ4TItxeASSMTqVnU8MU1+Q/aDLB23O6WwPsTnAS8CQ8xjqbqId2L2dbi3
6AMs6DQbcuvxfXbPdwhyvZ0+9tMDFRq4NXK8IaJmw1Xs1AzeK5rhrJg3HQoOLT1OOkB0IYLtPTp7
KUK3uaxAC7+NnLINA+KtZKTaTOoq4FF3v0X4q4wzieFCbWMEo+wP302FV7PFE6W50p4cuDHoCvw9
oQXGPTzsG3srd8OHCKt+0KmbwhyeeIOX9fBc8RLQssOVqW4lyLPOxVpHQy1ly0WeLOoKzMaz8rJZ
fjotPNnwltBAtLOF2EbogQfBtl8yaA1ZWbQo0ocEs2vxAN+UHGaaflLVe7u2GgRuLSTcobMBjvfj
TL+wLkPGA83jKoYEsL+mUlJc9mvpiGvD++yeZOrNI72+XwNiGV14kqptxisuQzUjsQ6R7iWoDiOd
qodySliMRzwvrhoeq5IJuNOHhF9zgWn9fOHJaEqD78QU/g+/kDGpwhMfR81aQiXl3qteO8fSS3CY
QpD+6rtsFMiI49tLUSbufOASxHA3qeLXpbXPZz0+A5IPBeXVimH3HQ+pVG7E9dVjrJJVoOmuRuSg
gOdoIFFGeGjDdrNY/MnB1897+RoUMBPVA4MfQ008Pu3B0KsemDSC6MN8oFAPHk0kLnot6KsKvocR
JBWtlwjehMfb8lgT7bAZxmyLWVpquGR1I1ap/4gbHpMb+PuErLMyyE8zuNzmtiUnJebhotRYMKww
unIjmrjWkdTNSwHdi+Mu4u2SI0T65sY4DnsFlTDrH4W4RsTq4ed0eW8n1lkfHfFwVdefuS7kykrY
ahBmFFPe3wEeYuXvY3Op6c4AXjgDf3gQYN50+OkXm8i4s3YpOfY9Bj8KkYH4DkMMWtM7ntwtflaI
QCGcCz1WGmbdUJIREYvFPaTIZ/5zBWojg+gzxOx/EvGN64P9BhxFFn/w67SbbA5mlrZj2FLZPouI
tB3LnUVayZOpn4cLTNpxYsVIOQ6JwKI/uxuSQLB3VOAzK+Bg7BP5R4rudXmPSYsvaQ904Ec7NLvB
hvFO/D/8AtWtSDwvWm2Yt30upTruYEP3WJUyGRvvVdbuc0xuFiJUpjV6ZxkT+0NDxPkXum7wYyt5
RzSfqn4B5ez4Wq2XVCBNj9+j2AH5G2AmmLTsen1pnkALNGWRRaCwcS5RU+r5WKmsalJt7UaCelId
E5rgjwnHy3+bOU5IgUYM+hHQccfjWRfuQLB1afijIWRkf9SPLw8VyJJTexTK9s3PfN2UxWuO4nm2
ac/CeDTftjJP/M704QfdXpDnbKCKMH9xBFq/tNnFPmJCReVBVCaoWMyImfkOJH+9p0bfQOSE6YT5
wr/JdINOXWVv+B+Zp7L7Wy1g8cqb6s5/Izhl9PPLu7IJxwnw/9F6jK8FX/njvAXWoep4R7jdObcD
tai30QNWv70+hZAbQ8aaC946bZL2XllAF5JbVa66+ahi5HzhRQ/7y2UeUiMAVfc5Tsm8MORpDGyO
W4V30xRT5XYJso9FN8mW8WfKypYjv/u7K554TWe3gd5ZOgh0TLEDrZHjrOl3UTJb3JXhhDIJANFO
j9UKJEhPwIEQINz83IJi5dZj4NkZ49IDtsM6rcSWiQnZg4tmN4gJzrxzCnW9NK7B8E3LlhE89Nv8
UBGF1vGJgi8P2YXrfcQSOhrg3khGQMkeVPu2HPbSfMCpX56ZsaTFS1CXhVQjIWndkawqc/LlbePw
ZRyzqqyXhfs8G0p55v3W7Z+Z8RF4uHtuJuRyzxADX/XzBaAJQntwu/bUO7/GWfZ+p5g1qrCB3XHe
WnSHvCJ1VbkLfv8JOPaddubL2vtnPClLusD9adOW56mxxlaXbJF4kjCCVsxxVeXx4z3qu3FTEVtO
rwgVXqFEF9bmN4JMVskj1PbnrAI1SHqXSMfy2BZ3FU/ovzWiaZSXQLTZ6+F1NF73Tv3Bmd3Aa/UN
DSjWcFyIpQs/SsbptXhHEa3flkMqKPOZPJ04Kh6CTTO/TqvliylnWidaHEVAxVK/DGy9NS5NgLCL
vJ/SLRestzcFsrhcPfwk94Nen2Ye9ajOYmEpoV5ljO/CMJNGERhzKME4bvcggqB0eL5cZWvzcqjq
YeEOYfQduUXUIH4dOJJx7CnlFqDtuT9EBrs5EBZoN3ccE7GkgF2QW/usoz4y9YUH1d1XRKKaHLHx
ZX+P0nz1R2UGMARhHk9aHtK6sFi01QaSuszyOHn8mfxvSvEkeKyYA4aufnEOwb9KLTsdlePiUBUu
aJwjHEt6Rt1XhYpFQU/B0BGGXqGnhREyo0i2qKU5xO3N8lw+k9uDG4fA4kCaMqAcablf3pJTrrSs
d175Ktm1xCOJh8OqoOoaKMOI30K2C+utu55/4YgHDgwTpsj9LbI6wtW+W7Wl0DZqV9W86ZN/mV5j
fdKlDh6lbcEoRvyt6HjoCTsSsrrPGKhld2cHGf6p7muTZczamaPX7V6LPw6s7nbXJi0H/sMZGqBA
YeGZZ28t6NunfV2kNQoxRcslxQUc9OvE9kvpxoZL1CdVAzQd27cBTV5vAlM3AySOavdD/tWqCHU9
j2mwEOxwjFU19Xd9IuCsGJI/IYqbbnI90lcujrgDgfr7txXnDj26nkrtE2UkDhaRlSjy48v5c+R1
vxukmZM6GCanjleFru7M67iLxj+EfXpkj1z2+/UdAgpiqev7MqSjGrQBuDYkRqyAOJh1iTScWkT0
TACPIB2xTRP8bxdq1jtwCISNJ7A+nO829TmaAjSkphyH9UZyxP9w39KFCf70Sm4A47zR84ltzYJw
1VAm/m3GU25dWFDUZroHhZhLRYaEKahZIVQKM/A42f/sNSLh1CGWP7aMtTgq87kMupgYwOuU7ZdD
ygHvgYoAHOdHVbuMZhN9ZiWQjSJE0nknjhmzD+yXJqAZivreGFcW/i1Lr05crUPSMjZQtbJV4SND
wW0yrfxczbRwzxg/1PuKK7dP5E2pgoOTiVLlRuAAwuWvYZOUc4h9eZhBRTTeVLVSX8ZLAUfS5/Z5
MXe/4q9FtUrwLRpnuovFsKwk4tyquiAHtfKkbmNh1E5b4XsddTj2W+SY0Hw2Kkg9V81QA4sdLXgq
1XUiuMB7ga5G9uMRN+fNAzyzQ33yORS8pqshjpLAFCz2Rr0kIPsTXGk/0cJkWgosVvtbMik6W7FP
s2wff2kUzQpiq9luSowi7gEMeKZms2TPdAV90/jFoF/CJXYMhpaDmy/3nvgvMkanoEfujqhpq6dG
+idWXv7u0d8/HVorYStj5/KUhqr/N72726DKZbwyOQzt/jKYZhYbD2JkGBvRPC/6k5K1O8a6vEJq
WmYExGAEEI7k3ZVWt4FzuWAwyH1PB2APgtI8iUjzJGspJrLiIdaBeUMbb//Ovl491dv/JepGWBGZ
XpwOaGkZv7hZZWCFR7sWud4TP2wlWIQNz8vQP6v9kXgexEoQo7xFyJ4xyy80H1z104kbPBRyZATn
/2PdkEsc4RWftprpnJQeYTy5x0qsaHGsbaRuFPxy6MkYI4giiZeGE/g2dTJasUWNKMsFw0LhtJQM
ZftqGOjGct6Jd3gLlhOrZSDoNCGBd4oQRZXfbnOPtiEdoSsjrF8kJ7kegP/dIyOjpL1Eog8EBKu3
L0Ehu33qRdH92ACg8KRsEowRWLujQO0P4B/iPxQ8EE8Q/5Hnsc780kd4+w7J5kNknAp58lbgyHFH
aKUB77xrCiqndSEhtMfGon2PK/m7EmzWBqpHNAxBzzo2tcC0HxY0158kUXD8ILxY5cHEqjaNf+AP
MvuW8CenqonJsheCFjU7ghnfZ5PFNHK3skmSDU2MF3XabGlEUe2XsBA1dfuO44Ul4XMY61TT1YXQ
YKRRP/5+W9ZbhtY32iqa7CPLyKTsFTGg2wDhPpJEBd+fNOKlxjdbZtkSZ4c1VkQ/LV+kQQWKVIkd
ehyy8kYQKGe8H+m4XaGl+3L+MoucyAyvTpNJCpCItZrCWwQstgiCbZyZPf4HWFluhXD7U5XfzRw0
rZKPGgOHEi2ZvbqDkBwyogR9kG0kf64/FVZvPGExJq2sZ9BiuSoKN67VA2wn0jBaP/exgMaTNhZl
uuf9xfHbXOktM8zCfCl/MTeMPTEUvsQ73H3r5r4AVJ6xY3y8Pj6bBuG0tVWEagvCluPAsNUVoQfR
3DGdf7smlJo=
`protect end_protected

