

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pM5kbFKfO3wtGOXulGoIYDHxT/fNVMImb6qtomjOjHJTBKmaspVOVrLRvtERhMiVBq054LqIbCxm
omKrNl5YFg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U1nwoEVdavnV5XVUh1tYM89A8G7MJXy2rMRUKIK7FuJgaL4t5rCIdYkN1kpAUTpZsvG8VhYnoITf
gPx+ZnpNIDq89cJuuhnbNRexElQ35WHZNk3b6Ovt1Ac8FuCqk8LwCF1khosIaYp7BoOiCymgrmD+
jO8RHibk460SEDaEPgQ=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NeD7mL9dCdh6jQqPQe2Cm8mOVRJ7WUTNI60h+MOarPJlSGIW3YyeTFxAlCXG3Dbm5AZqyq/7D6Um
0dS3Sz44LEfv8kzilqYBNJj687fhrDd6nKWTLbhkImuyn5pqhBbzJ385okbxTHcuGgO/U2MuNghF
/4hyyRmJT69e8g8FPic=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q5RFAyJ3EnWo/Sxj9AJNS/u/nJ1a+topTW1E806I1FKJ5rh0sAqwjYvhfUB9DJ+MlgWSdovhM98k
M+7/SZuvkwd1k36lpXZY6i/uA1H8sfli1FI/2GH+4p4nE0BCNR4yF5NyLA4ni3SAAWDe+9UndYtb
WQ8eYNjF760IHQOpzF/U1O4FBcQr858C+AHKRTQB5MrLFEiZh0igcP08K0fyLcO6ksLh1OG/Tg5A
5LkjvMAndMWosRl1q7kbUtFhn9VB+3uHP/LaHYhxdIuz9zhl4DQszY2TxfAbm62SNrnuhtIHavzl
BZa0VmJLpxgeeo8oVCm7UnkA5ETNgVvzyvFgIA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CwwODyIxPJaOqhXk3C0LWzZuCnht+KQbdmaYIssVWSWWhiBF07SeDxq6+8BOr7/WUBLpmVlX3NtH
C00zRUWg3fv9+q551nW3Njbt7SBWFLR7OyHIoKABDgjBeBCamlQ9LGEF7UoB7iOBYKuSk8CJ5Udm
OlrI8xSrsS0TcuIGuxA48YK0xDfcZwjmgil2FD6Fy6tQ7WVikG8CrdbvV0lyfGl8jL2kEh7RtrHe
yqNYxXs2/yw4uWcKr/Sc2VNpCsKbLpxTGFpGsQo6x3y+Wjl/pOM5+YQ6Y7r73Tg8z1AUMiPNHjbu
BN9r3R4QnDeKCwqPV6cAMGb1yVk1rwQ2l9RTRQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bF3xMUaKQqhrxLNzJRa5Xkh+JjnAh7OKs1IKf7OJVEuWA+FAG7Pd9bdwjXk9SCFBt9wbhJwHypex
SmUI0F+QkOhBdUtcKiYRnLyHBON/t5sUzO4LgYA5oJSsAdgYJgwV52GzeJEq7PWjnv6o/r0kB3sZ
MFITpDKyLwateefaL3T4xlnTv+EJjBSdMAZDiSsaUwdBOF6F+v1TwQ/iFvvJtE727/b2gHvPCMWJ
SIvS/OTpuvIqDl5nL1w3hIWnI8CAMt+BNU6/+GH9mSyKZqAjRamfpR7JHsMaT/vDxA6WTG9+HvCO
klJ9KJ0Wm8Cjlce/XTiDMdmEqMYjADeB3kxoYA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
CC6X8LupWnYoZolqW1eIcaebN3FMF63v7nT8sB5JleBWNS1QXM2kY/HLvOdlU4ji8BANLufl4240
EEYBc/vV+Ux7j8GZkGuqRGRJqe7tBQ4W5tcYGpnzIevUIuTqfowNlCfaUC53iwwVdqpTEnbA+zoD
66OUKsgJk71ykSWcdm0RAkr7h4lgYNzuhuz5iiolSelP3YLNVqWRkkm+eMfQSJkx5w6bZDk/zrpH
9lLED7hxyD1ANsmbPd7m2ulBwbHJfk4PlweCRAIrpExcaPfywNLABbfOsZdwL1ClNEA/t4Rg+B+v
giV2mldQ7050M6lII7skqKW/YiPzxsMQU0nc9gyMs+y34MhvW8ZQwp6t+1W4ZN09X5ioJqavC5md
D9sMm8xz0pAKFZkW1hb+hnB5xnsPmKlAR5Zz371KUWzdlkityFAHq/mlJAF1CBnjCzRiyv3al/AU
Sp0c2Ep8bdee0m5NQ6xAv0oYnHeeWyNm1ShyYA876x9Xn7hfORW1Ez9fYy/zzURqeVt1MAC+pXkT
EU9NbC4XpgsRGwXu4Km+JsZVZzolQi1xbj1jXd82uKijYc4dgGIQ5hPARCJ5L2KLL2hKqDRGs9GK
8aV2mWEEfO9SnWMl6ZK6Vr7lD3Jnn0xT2Z6mX67Cyj6hSb6JqGR1/w70wARG1zBC5NRz43eNVXvL
AxnF94UYh9hZOLiczPBNqPkm458g0IAm0OHRncjR9QY4KVuG6aSm1opgTQlzznNEzl+Hn5mTAWIf
pGx6LFt8j/N6noYDKzO/rwVFJMY/5ia2v5uLjHhkUP+apfo9GuW6QIw88e37+gECkf3bZ7F/w8gQ
4cESm+rzus4o12Ar6lifhOdCuWKqg+78zOCuOLU0T3t+GTy5e9lnj5xZkbF8fWNf6qr34MrLumaF
6Go9b125sgTGDtfbkINCDwxyWf2dY0uEYSCqgL8BAR/QeVpxj3T9llb9GV6LRMZ7ym8UDCrbUHop
LIrgBN9lZw/ItlBXw33HAFYRFWrRaQHmT3jZ1QHHdVKgrY+W+4WQEjPbqto5S/IJftQLBAHMG83s
pYDRqYmJGbFea/dARz3TS1YGvaqJfBKIfTFsVbEjD+4TFUX/0WZJTzFTjbGSkc3bnqU1cmL2xpGF
pStzCoMwIQM5gwMmLOHk/i5EUv4ZCZD0tXpuOSykgHGg2i7IhF/wf6NrSM8vLdQXifpjGHnubhPG
eZxVWaeZoZrIZBcI0pDrCxon9517DCl5MrfYFmBLAe2FcaVfPfU2YoDmn8zFtSFkx023P3ggR9am
De3i4a8IAflIvgMziwlPqbYmPQzNNAE5KlNXL1uWIPu4NNxIkypDo1hFIXEV6JIOt0pNRVKdYLGn
DGh5427qrQFMczMoEP/D/4eRKrhoFKWWCyR3o03hj1h1C9QlmI9hO8410svoBnFWA11r9wEu705b
ORT6Gbn5Aa5xbLsRe0i/KG/xsgMWPInLJw5E1SMoNHrD7E8Jy6fmQe4fCRE3APLiU+D/KT5qIrC/
1BhF89KY8m32Edf0YQBd8jhgG0RMLWAknBHRRx7COIwJpqFPCv3yZuqLNJKZMjVwVLq/chgP01kc
bVHZ9QyZQxqruNnnTdhlkOxVjwaNr/sO17shIDI1w6P/Howu48OHBMGh9WpulKwJ9h6uRN12nnhY
7KwQrT9SMh4hLnnaa/aOCXvxKHAb/St41Es+a6cfkzbq0gcT+L18LRbf3BxiEp59AIAR8op0xH3H
tVR2YsffzjNaaGmKDBY2jHDfzFdBJLiBZ/zoefGvSfoWIwMeBQxdtYvyUNLXBavY4hrOPRneXvrm
91QPUtIIKS3MX4mvPKiARUrrN3ZlBl7tMv5AuZACBtxGrreZ/XIABiMzbibLvusR7LobWDhXvxbv
wXJk1EEx1Xo11CJr4v6BtNaGjaAlj7NTbpMAtEy+boTTz/cwDgetQwY/VmtsNzDAhEBMHwOU2BCw
BLJjkM8SV8/3fLWgn8bEKr4sCkamhOoJc7LPdu1FrhtTKzywPLrTDvRBq0r7zH3aEmzfAXSc0lwK
6IujFt4EpId8YLqnaUHqGLC+09+b4ji+mGaEYcOBWVKZx8lH7tF1MxlljrWTUBBP/WU1jCL4/4ka
vH2X7h4aVwCPxCVUOPxFOBoTqN/0tUHkhxQPV6TVjcMDUIsQqDqWRTuVlmWZcOGEDIweBo+8MWwU
Yy1RhzrNxujizOUKV6CieCAsDewrLjk//uCpsO4i7HZwOjdJUehTDC0UTjXvrES040/SF6Jt0HKz
lDmEq9cL8HaQcaLN314HzW9Fv2puHkHR06nlLPwMVfEtCYKCpodeHkfxE0M81R83fi+Og3/WmoMv
qQvt0YfZ84z9J8QT+xye88a3uYhhFVZkVRCxJ/fnQewBHbGsLtcFNHR9Z1POCW03WSC0UB8AGXnl
LsmSRIltxopskBpfAQdKbMKgoJFogU2cA8/KgZ4rpQ3an4xwX53waMuAVbfq2e2IjrhYgmGrBAcn
GZP2HeS8dUwCR9dSSgrrYqKTeG/gF+ELRk/D9ZgvLC4d1YOoOk8lEoB4cH11EKjlXeoqUAxEHM9T
yxHHSL+srKjzsaDyy40eMDCMqS59arrff+UkHxIXETeHJUNbfCy8+jD7uYhMfyVKuJVglRQgX+Jm
b+pRPh94ZPV0XZGsVXq1Pd7NHStgKF19akOXk0PfTS+84oN8Cq8FOv/O0Xy7FmWXi/FYvT0o9wdn
ScPmjLq7bFvKDTYCpHytCOKYu3QctKsjvTImLMDAB42rYCKAvmtj5Ru2nu+gYmM0/2jO/9dap8/u
Q2cN4Ce6AMnp7JO+6+1E3icYnxXbz78CsIdU4WqjspkUDRTbp2AcVZAVfA3UbmH4Yas3j1ul04q6
KeVDjBx4XZ2UlAKb6GL6ORibXxqc/3isZsjiKr+ZsSTY+Ml4G/qQCxDu3HgAimCEIJ5LgJgg/rq9
g2ujG4U0xKWbo4Iq/ogKFrTFczFPdhN/ICFiLdqQkhh7wEzx68n42TWMQIz4LjPq9aeLgCaIJlWb
1K7zSdU0KyrpbMj1vu4w5+j3pfvFVmrQLeK209x30FzcZih+guaiILPfDtX/vC8cFF2eOm+iYpDK
guensJAsQoBl5VJGlnYVsnqs5JNzd6ScKXrfypBqS7yaiKBmkYoBD5DorsLTqyXfOV7VmJ9+JZCU
EFtLG9DRTD0Rm0CebOH4XeFVXRgp/RJ+28Lrd0FdSyOjy/3Z8Hr3E8wk+3wGWBvfUCVmkGPu8eSv
cNVEyNXFoifibrbfdObbnQwgbTBWLaEeOhb9Z3In0uuY/mHMmk34I12axxR5UMiCwQuPxvMLlkGR
zyk2Z4QuZdkgrrZDDiwUIWtzG3v2l0e4uEfPgCAMVxza4uoLx/QJpyXhhYCwTcmp8c6OhY3fYeXm
hpBvryZpipXxfItu7ncTqoCEYynyDuTqhWhIZWSM8ZoWEmfvnNpow+DmXthfe6sTpZrPkg5K3qoG
WqCl4C2iIBWuyESG2sQetR2eVHlAyNdM7NiHDAOXw6cCzgzmq2TA957vNfw01yeIhjecPMBV0JWu
f6LxSWSO6VAsqlQYY5V6Jy71GNazXkxsEAnBUxMPt8U+IfGJEjBkdev2AB5voPWggKEmZWkfdVo/
vnhwG2eg6jHSXbobmqLJot72gaB0y1CWLuGhsQBjylXOC/iFYGxWziTkWhghNYUql4QAiNMumf8W
qPcZELLtDhQx7ZWBPsKkitUj6x3owM7iZf0Pdafk/7iMxkixkkL/JPfqd0Gnzp7rIepN8aOOQJxR
MO/vKYP0dPZT554daaPs2hM8+qgrZvaZMDx0N4wCVyw0Z/BX3TnzThCrPzDpRyLgAGScFaPvXTRC
au0ucmID4uk3dDeUmyMkukD/gA++hHPFG/RQ2d4oiqp56DnBpHC1ScFJ1omBwpOx4pNBRYbfCkBl
Rp5vcqUPq17uZZFc/71oGCRAXYzQyqZwfvwJ+XaEUJLuF3c/lcebP8NVUftSGo/JwF/Skp9exj6z
gIs2DHGYPMDjltxz2acdBE5ZGLTeVCMFayFNF0KkOYJ36/QnRyCG1k9LScGPU9xD+5LmUau0ZbVE
AbAxGecObkzmJlOd0wWfNPvdzTaTAfBss4KdKWSKhkAF/eOfhuJeXk+fXf11RRZdCgEQ/PLpEexo
Zcj36oy5dNAl/Dd7+7D80BPPovU5Qb5BSdqALyenE3EO2dYfZk04sUZbC+lAo/n2R4FqnguDs8ie
/9cw2dasOL9n1yjBnlTqmeiV67MjzJ71RZGfTglIpGpoVE67fSe1tCW1yflvZy+LHLwLvBYVjPDy
/a+vL7XXo+oZ2y2sTmBUR48RyRs+VRnyEiIfSWzKHjM1P9pL0DYLciJpbv0U++hjjO1OgcbHFobd
gPyNNZG91p9uXzMuLC+h9GdOjbH830bpCh9W1nP3fH5YdaFQd6ehBlYnsLajrnmPuPHLpx6UXqhd
ANeilKWu1YMh83YHOfZzQUJhrzTuHp4waHebfbUSNc3A62bt7tDpqpmES2BftEKy02Mwgx9dFZcJ
dOTOlY4qC6BHbpR9/UFlaH5m/txTmYxxtS4gODFSIjmCtRsEOOKBTJ2BDi49ZGVgiYhdugkIpD9N
8cMr2keOtZhHfJoU0VxYUQ81rnKaRJBflGLulRg3TWVLJbUexkBzo4eALW3yZq0/4CXDwp1EMDnK
Xusep6QJHrvAKX0EE44ZK8ZY60a4pOFh/y+mZM/so12YwlNvBQfakq9wGniSk6sShR+Pd7PkcXMF
pxncZTAn9pMw+oBEKvalYdoaojMcxXJIUvqIG90m6mmmtQFESvQ0jR6TeOCQqyQfFJKHzxFPf9tR
VqEHzK0VDqIeTsWJs7CjG6TK0QNhpuRgiBwJwESO45J535+4qbiCMd8qX016X8nTh2pqK0bHbeFC
xxIqvzFGuF5/UXPA9XlwhUGhueVeleGfVSjYweIGf1dkHAkgMpR0ITxYgp1dDLQwSSguUmE7ncfk
cSpOnppv+6Dw/9KyXtKr/ldgBQRqG17i4MW3FC+Ufs/VSqCULaL7VZ+rdQH85bBrex2lYwfvU1uC
TbQ7uF8DczMSNJdADmlTWNU2rT9FXfjquP7GuVCopCOPOC27ilbeocIDj3O1+w8WFJMMqykbwidQ
ScrEXqs+GaPdwHkZaQuS1U+LsehkWXjXEy+VDs1YFnaGoBWi1nv5qamVOg6QmnbGno8JlNVu36lx
Ns5Q0fKBEM+eP1K/L+8Be6sd95HtndU7nWbBDVwDgUs7dEfMK7bzwxNZLC9Cr2Y/JLpTgKq1iQe2
Vdrk9puMU+sf7kqiwkV0ae8r75IIIrTpQT4UzCqPwZghyLteq1VWjCRE4sAQgqY+MJhcnIQzjppT
eYNvykQ8D7t6YGihs/i73LWRUE3Yn5cXi6pGMbL58m7P53EgJaJLKga8Wf9HwM/7ekYyawYUuP2p
1ZRkZvFLGE+vxNxFO2LIqcv6lD1hEMyfM8tB9a2kwHABV/pjgosAziXPL+cabwWbNAuOlDGGjbsI
XYte6zM+Xu/vUCXIRmHM6R29YsUUubD7H4C5+ImhhapOI9Bc5t/m9CnmlpIKn07OK9kC3M4pbVUR
Cq4Fn4cyPnrTsIo+wYAr624S/Vv9kubl4FClypu3gwnnUW0c2DhFvXQoQcXFcLW/kvGJq84MuSee
YZb1CQFzHGuSRSJifZe6z/42ahFOI9XNEOL1h4wPY6BWJuVSED2F3hrSTmzRQ9ZLhV3GtVi6ubtb
VYOY71hYC2hq9FW6d3DdCWz9HjEvYoAvzlZETvqg27sI9IInVgj7XfMGIkEb3UvW7XQTEJI60azb
lf3BpLBn7ZUxCJCiBsPzDuRJhjb4qNQK/yP776K8f9QZX9FZVBSrBl/pT+L5CptcNVOupvUUSOKe
U68FoSosg/S4+NSPRd++Alw74Dh6YDmCocGQlTgmB+Xs9wZG5WT0p81G5ZmfJILxjW5zDbuLgp5C
LDGxkqGU6Fr9a2urstCqyZLM5Fdzlx+fwvCxfW4QxKn1lGgaxMrQFBEYpLSAxgPr2cuHYCuxvMbj
rjO/j8DjG/oLA3u9sRbtad9CpOhedSlFhWWdkbiQSVettvJzJ7Wxc6Dqe3wCqEpDOeo7qpGXPrvb
jFEwXgtvaTxUB0oBYhk7LYdhMd3VF9GmR+VfkH000G48y0q0DgYZuXRRMxLquXWnHCIi1SDsrBb3
2c7wAT/G1twke69N4//cWZ94BhI116ae3YTESvqxs4mrcpMdE235OYu4CFNVb68UEak8mQSs+puD
Htj6NTloI2oiIU4hv/+om24FnDXcMUWHEbtLphbJmxIa7n7xGy/neEIWY8wu6ZFGAhZYnu+QyeOz
KElPTJGDUi+VWe2o9At5db1bOl4FT1rEFLOW8NyY1pioIRLCnEkPiXyntfZE6TcKiSTUCvpsLyR0
DWmbslW6hwe1e9n+4ivkThynO+fVMXE6ciLtgutn52an1iqDEzW1J2r9gTfWI6ChOV35Rhch/II8
uv9lfuV987658uVq+VUvWebOJrKA6yNM1d9fl/3oXH0PEhuJyZ1ZCXXOgDW16sh/D8b8Llv+qyu3
zSllbxIwepILqlMRbvyd5prLRLhYssBMUjQmuB2b6l5x05JXM55TMwnqg38IBRbUTtDCRorDXDVC
4/WUKKxxENzkNLi4l0HwQ426R9A8OhopBmG4prkfx4NOV6tzMeLOdPghtlMNZ6bfkfgWNSUGdrJk
EUGIliGvVWYFz8mYOMbndw9hytfg3GdimC/p+CDndUYiD/TBlEVj70qeQJ/hlz9Hy47PNu7VTzsZ
IsVXxEOm07/z29NLjWnjGU5BJ53S5usuVYkcxdCkdX+3nUVYtr+VRGsYKOHosDPHkqLfGiAZWqVx
9nNTkCLdXAqLi1QUh6GZbN9RK69Gajx3HK3ZkIg5m3gxRle2xsPedt3dtuAtvPYkkJDWpYnfLQW9
bMsbqVOIw79eX66MjYz+GIPHisG2d3agbqgZnrAQp2dbo1Ii/8w3pgaTkDiU6r4fY7uSuwFFmn0o
t38340jmNmJ1xMOM1UbGpL06bTldo8MHln5z2qnkJwhDkYvRb6zvjhYixo8cgKys3hfZen9Y1H3+
XaOPpK8z6U0vU821U0iNw3c7Fzn+H71uIdB0Jgep8S4tA8//XjpidESZspD+uZznFj2VDXaBSxY2
glYqiIzI31fkImfD/jFCVSQ03Czt94MpiS24VM1DyD4Jjsb1bl8I7Mx/bEnpkEEKtXqPhyEAc3/p
VC1iZ9O9rrWXFPbxScS4cjPBqM6ChPbu/crLV2kHD/1aIl20ajJ0xRuQCUO2X07wQUy7pzXyDxwk
1lqLnFmF3RUfkoxK91/d1o5sRuKW7MBynOBOMOt9GL00D+2DQpHCI1ABSL6Xhned/6ldS34mNoNR
LJRjcGUfcns282hVfEHhRFv8g2Q8HZVVONn7vLl0PxirIKlsieWuQUimtz1Hplyjb/h+j61zMqua
JF53ybzhMLENA949apt22d/oy2QhDdcl9FXsPj+CWNCfCzkmjFvnW5tjZeLdflhTuzcFlm/CSqys
7FdkfONkCFjsWVv3H/7nkk+qey0eMA1C94JHwaeTWA5NbnDaH3g6toLq8A1NKLbvlRQ8m/zOhgDK
2dl4SkeVAz/uhaI2YS0BEnNgNd3rDubst6049LYYSoJcdiv+aYVQxP27UzW0tfWpAi93y9ncYLLC
YKfsVxiw4w4Yg8glBk0VcowEP5Vduk0syZa127ANnOBks7MzJpLPrvqRWveH9QsxhLOZhUP6STEm
rzoVwrqTVtD7jbXmTlOztfXu3EHdVLLRnzQJlbIEz9KmvedjqY2REoYXSITWcZ3vmqs45F8MISOo
DedeMo0fNZBzhONz+L/ZhTVdPuVl0n7LX2W+AYwzdlHTfE+BGBv7rp7LNaMdyVGi0gku/4TEDGY2
Jd5wReeo/C7M5uEncvEr5eB44eo8zD4NpFbpWqhgv1KIbSGsvKhPY4FbkkvoVYrqmm4wIjSopgo4
F6xZ5QOyKommLrnJJOz89ntN/4n6tGnNO9dZqdboGc1lWiN+39ceTa3953zOHWwMM66qSuP/dvSx
t89AxPfhFr4o2+gYxD7LxWv8MXJlRvvlg4luIPDxOCMTvqlXbH5KbA9vXmDtPLrztTRrrfnhJWj6
9CVx8L+Oc0s+dEriO5NV8HxviDNYy22Gm83BI280uCAV/aP39GnsKScG2uUhMyqZq0gBb3d/vxky
Ca+NramdHdcHEXU+I32X4FMgDuc7GYrAjnc+gI/ymwFcP1hkYctKlqf+3mt8MDxnX7eYezOaMtZR
HbmkhVUjDXodFiJLdeIFNK22Tf9boSD6PyA1AoOnzIxhNSik+8uNvcehpfXSowrIFsxqYJIyKhdv
+FlqqN7aATeYyC3UYebhRw9dhHCorcykc07K88bP7Aq68zxrKszP6Hdr2VYl3mxsC4QUh2WVXqGi
nfxaQLqW1U8r/ev+8eMX3a+5N3h+2SjfYQFfIBtmOatJ5dToVYO4NfWhLAruY0mxs/ag0J71r7s7
DAyeWOyyiEYs8BS4PYMU1wXlA/GcMhaBeRyLddR99eDOitI5DJjQ+2jlRn1Va8M6m5ZYd9Cps9gW
Rb8WhSQKODcgxl3UEym4PQikCA7TmiXd7gSruPBdrVZpIQyHH591Qw2+eWYt9PnwlQlZDcpG2Cs2
tG/lcDj+7JXm2xB37DESAw1jEqw2vzhh676FCrGOp7Q1rpUWMxEIhSgHX3ymw5jgZLq/JsfIeRP0
G0QVw3nqtTnonuKtISY7NrL+SMPQnx1jF4shG8l6Ot4s5nQjptIrBimXnNkGzlsObzLPC6FBoZh9
mG0rU7APwE1iT/PED6VkLNRu7ZTVoqkZiLLzlQcaauilrylrFs8AD2YPl+K7pfY+7RJtzS+Ck2fZ
Q+ScD0UqBeG74sPFyMx+LelIFznOrSJpDaX2wjSfqkJ4uOsRzWWgW6c2GKW9yERSj9yIHN0fHWsj
6WHjSOuhEZDl0Znle7tTm+0KxBfpO+VckqcYIUb//xHg53NpurYVrcomlORJoGr3eiRnL+L2r3DH
gKaKb0XCZcKChXy85B3845OZOQqlFA83+ybal9wXiU/goED0vAKi1wiG22x2E4HC8rra/0FrHSCU
MMmPmvrIjqV5eAU/Vnx8QJDcslVxkNijEqihsmgIAHBSVEP6gCCvvRh948rRZ/ETdpXOpF8OleVl
e+5bZqVDrP6B8T7ZxYwue1ZFhuFQvhQOPrz6sqldJureTOcXy9G15eKFCe+NyU0gCg/wdgOmvyj+
iXnsdxE5RQlVcPoNIU4p1a6WvOv1Q4tP2sRYe3ug2I91AlCOgukBJbatSFpBIuwg+xLmr4F3jNpx
5j61ulAOiGhYPOHrrA7kALxEVI47DBUlt20FN0CfqO/22wGaD6zyw1URzz2Ah4ZD/4rkcNrJ/3m6
m+VFj2ax/xxnXaVAGAgoRNbFKkFULH9j84P9g4D003TqeiJaIKROl8NKRSto6IRv4YZo5a9K6hj6
ZDFzqn36dajD0XwUdTtss4mny5wrK7jMwgdqSoYgvSEXvt4Twb/zZQXGpvR1vR9lzrUb2aApCBV8
vSM6DDra4gDLicXAExUv+qsTGw7zQ1DO1KI468FXjkyGL7JIeiyBUDsYfMAMwY1gZC2NryOuk1wP
MUfFjQrnTqyexbYjuzs/OQ8uSnw1Gu6xIMzwQRaNAeyR2x+8+W5bnZpSnHDhBiULQYJHgJOiKb59
h2scOTLzwPJF4YqZq0cVCBYE9VNnIPqZVmt6wXp59hUGP+87m5oDuWAyRqKIgNoFi80bUFfz2anr
cb9rNoOuT7HFT6tRgMgY8OX+agBjVnBlp2Bp7rfAcjoQnh+UWq3nBjFNh/KW/jI+O1JA+dJY1NX/
/dV2DEeSL1+S9QqJD4qABegJEwpzwDDD56BO9UP+8IDqAUzP89AfmuE5dMy4lkLnbqLU1GuX2CGZ
3/blCy6RQveCB63aD2Ik0UdfKuF8mKfQY6jxW7OeuwhsyjMv8gIRMobZYyZ+OJw7Mr0no9nwlRKT
XJVWbbW3thNnJED620ZpTAjfhbja7tfrw82t7F4k4y+JmRHlXOz3PQ4lHUo/tGMQJ1r0E008hr+/
KEjxl0gpglcVLYb1qfeGiEX8zfYszRp42Xchrsaopf9IYwK52Ge1ekjE48pZ7uRlsiuXO/ABX2+K
LJHcHqHL//5jHGdBwml6QSZNlF8/VK2Il0xvOpG9ow+7FOcV6WKsvXUvlvlmKeOLUMdEmIgDDxg2
XyMMEOwQF6a5UQqKJIoAgKmFKX4VJkdY74qU8LgP0nBX2FAYl47KQmRmwZ2rBj7NLqx3tYx1ou/O
C34EHe4VkrkXsaf/6NO8l9e+wd1yRomQzvNs/DZJlg3S9PQ72enZpDBzkWe18yEZ0YtKvOmhbqmR
HGBqdZsx9pKZVxZ6d/WiERP8f7AzJxAsONKTxBVY98aR6XDjfxRMSNLmoroCLKyGEj1BRtRzRb95
JD6DssPyhFGOXcd4TvKDPkV0WOx+fQf7PvAfsGdlt4xa6MkKuB+f3JBPFs1sup0ejGF38t5zK+GN
bVYRN4OteDblJqJoHXuwn/LLl4hnR+AzXqFlJI+V3gckUp3eNcMB347r0/zxgHehBpIbCfxkavYl
VrhJwJ3H8y6CxAANjmWkm4WJzObRrPTBYx09RKgjc4JSHEjFjNXWfD8yY9QQwczVzXXX+scacxUT
VKLNLjOsmUBZIrSE6Chbjg4SsAGbnXNSujCRJNw0Gxl9642io5L/2Zukd4/E2fP1U2MgHgHUBDo+
wBB/+CUHPO6uA/+SjjgojRwcd2vD00O3RzgfC+/wPMtzZLOxtuurkChmN8TMSah8Se8hLoVKY45a
YX6TktKlDDghlj7i5VfegMPF0rJL0XdvHLtfJmu5o1bqYtxIXG0eUOnB4UnFKw5lYCng1QQSlVVJ
wBjNj2XreBOPIKtEEBEVXyhlUQWOF6sADGz/T8eXBe+ae9R6/QapdDB0ixm2ABnDfiYQs2McLozW
swgXjcG6cxM8nvbjj7kliqE+jB7q7RbJBU7+VTwmzyEJKBmTIE2EbaQQemOPseQYk5dPIwAFLgSL
XXRwJ8/0KiyMGgdnpcgPKvxw229ImQ92cYOojrBLF4iqzdiltljJsPAzBz8gpjq6hLADJaft7Lrs
HUwhalwOp62nVQqF7uTmlR/VbL4dVWQnK7PkVpGulHyf/n8WmMXSO1sLu4kHjeDl65j54KDNI9oW
XKkdeoXHLEAo7JRLNekipKJpyeYLyI1vDGbfP8j4TXwOb7Y01gBq2IqBSlNZMBtd2AASyL62M1+b
HlrSecha1WACac2Fi+osevioymjH4uJo6IH88xesNPLLGDp6YvLn19koQX8ZJSS9OzNeERg4ltTC
RgOGtO1I0fqhz+6HIwD2kc1WIqo9XWjV2MGSOUEgMN+qay8sDP3K0IbCDQkipGHXgtr24Y13YJiq
KIAPMKhd2ktadHyJ5MsLdxnloQThXpp7qGqsUFJWiccRxY9dG245fh/VmjWXer+ae5uEAMOL6c2v
mV/3yI1ND3CmX7sddPWuzJy/0eS/mgzSI5xc90Vx92rAjwPClBuNzusmzBC6YU8YFCcMAUd01Qzw
ktjJ4KQiw02A7DdGdutnB3Fw2ph+tF886mbkPY+hOEFi5uodNO+ubAthuKk7626an8K3R7fbcz08
yw1Nqi25d/Q9AnSodbkt/48bGR2cB+GoHdqnx7zg8QuFWz2zfpu2pkhsHfY3aJ9NANB5g94euhmA
9mmGHoiJqGNHH+F9VAoAB6ZzPDGyj+gTqRQPhUtOU7WoAxRUvAjtU2TnBod0+lkIOFBH4HN+Y18g
X+y+0YUlGn0fmUwbzm0++k/hSF+0qqY8+wabyMcMRW1QUriF5J8z5kwaZzucQ54Js0vlcTV1nEvH
E/2dUDGaerJodXwJsacd8NVb3Fp/3+r11XF7NFUnH474gfwZ7WwBUpV+P9W8ScAMBiXY7Ur0+lWN
rsErnhRY7/I2cwrlOymJRnpiat6+3XMTNXf1biOg98OPjMaIKyRcMKOjos4pak0jry0aCp56Q5/Y
yFeOJNh+yUQn6n78GZyQVbBV1iatwF9EgY/vCJ4jR/jctlnQVKjgHNUQaR2oif4Kcw3CjufNH3Rt
3EvrQYtKR/6DezJU1mJ5nXtlMx051tM04gUajWquNIgXq7iFZTfwB2TrlQ9zzUH2gO8wxt89bu8A
8mD5d58nHMSzpVXWNUMYtiASIeDwqZKGHL0cxrBo599OY2A/b9WEi6rUER475P/PgYqiTfumFdZk
XvJjJlmuq2TVLXLZ4PKdsQeCqJqLrEM4UQyb/8oguvfItwdM1CrEwDwcOHSAX1d3sd2XaIQMclgU
Bv0d1X5z+/vU8HqIcetyWPUqmLCSmCAD/gzgjIy+f8tH0Hv70kHXdYLywMcDoHdsgedagwXX2T4q
y4eTO52N5I24MoYH+Yz9eTX/uuO7QXPU+pucXYM+sfTow5Rhb3DKz64803L6Wa95ylKFsntpnwyG
7NeBZIcrPuHOpMhkm09MJsXj5GTzwBX5mejxy0dSMySzyhuvOBZ/OCR1UkGVn0dcpmyXVNcTEUR2
Thj3mZAWBb3xXmIg9KOjyVm3moQgD9qfiLMsy6YdRp5aZyMOfm18ktsK4SdIHRUwcTv9s+x5sfVz
HC3EF3cCPux/9jOkK9Xmn+L/wqOw2eZVi6oQmLS4B5yL6p8TuRPzsx0IWUNXC/pwecmgpiVa36xW
5iaSP8AUbFs9vHOfBNIRHiulm8rbyDzuJqO21V6mjJ0FcvbBO8nBd+/4QxeljnUGoC/zJgEKW0Yy
aUuxYTYdnEp/6FoOduoPzto6xxFpFmfWli7gx3kjh0/rt18f8GOI+CsoC5mOuofkCGu4xiqpR6OT
EYa5sNcaZJ/E7zasYbv83Tj4wBT4gAVOhtepsjWgk6My6WbDlYD5S8Ko7VydX+gYcN8RrKK1qeHg
eRiA9NvlTzJdMd6WwfSGZoJeLraO3nmhkIyivm8yODoqIrVBeGGZsIC0ac+7xzgCc589IALi0l9l
UbMqOcwEirFlK43MKTCU8r3LitVqYkSzLYj/3dWTXRr6vxYpMsDTo27cPBPUAHM/epy8DXbY00CX
OqNfasM/jklzsoLahyNqYXcKWa+UPxr/nkWS+DBx4ihHyMtefjwEzxGDZ61/z1J7Dpv3bSV4C34X
FtxeRlXkiamy/0D3fUzhLe0kG0LpwQRSYz1Jbp+QV8qeSunJxZAkxVvZFL7SWPI32HZCfvQ6Y65g
SXMn7GQFV59oXYw3YZyYbIUSaETdi6WOW/1Hj6x0VJJBZe8U1OMr8qohm4Q7v68Nxr9qEl4JUJyB
tZXfsB8ICKRXBL7qL7foSU/2MW2gmewk9Qx7JTpESnA3aV/eAKXiF7QxtctvXsbh0J/SG6+SxgPi
wjudz73QcVvL8UIJMhT3Sl0SmWjuWBHTdep1nOmtdC71cR9Fiptpw8q6LOoQ8LHwVvtoamo2tg4k
z1ey+7suOJFcv4OZaPxXr3MPiPLVnj16xviLw635Rtjwo/6hPkeOtZNqqrTEP5wc18bycKefI0Ca
W1vRK34bT6+GO0uAxvEvQKMiw2MHhmP7SO/5eQIylbP9rfYlxQeC9khUPRcRf9Y1aD6c95MNNnPv
mgV3rv3v8sFF+FwOmkwcgAeJUVnUzKVh1xBVZONKFGMsX5LKU9qjR+sg3b+myUfRCNtv7kaG7WE/
yEu0pJDvJmJNW7iorZUfvOsMCmHkcWAep/CjgOSPXY56rZntcYcoBdl/ngWbFSTlhx3g4yc1lNlh
rxjG1J1CCoDtiLRdFIYK5YLe6G2FtRjuLit+A2+VQHjS37Drad4l+tvb4/K2c3zQvVfuUFCwF00y
YSc06G6KM5zTif2M/LGekq1Fi/pjT5F9ftDzfooQF7EnVckaofz3yhRAFSxdtShjmi2LG0mRssS7
s8AdlRfpBANTFtiUyCUtxT8ZsB0LPnPFoMCj8fR3l8sDGemogAlQvv8yv3hXwPKh6TeEYNL9aKdb
CxYFqZDDPlVeJOcdfIk3qZNgbs0Z0ncpnyaVQ12gNEsnn7988bArhHjgx9rbH6YO+VMyJeiO2R4U
UN+HOl2l6yGX++Pas0CzOA2VV5bdeU/RZs7j+eUoaTUBDS/bAzHWsK5opeoWIO//OIK3rO6uUn0V
VQnB7uGlb4/is+GPu0Apo3u1/sAiO6NkhMUQaDCuSHPecEbmELTYunLEJKRgIYKq/6jY/shdiHgb
zRWfBWenld5XkzBI+H6qNeoNSiRsrMR7fZQ1iSJZ4ntQB1ImTtJjr+YKOeRT4yszGMBxiYIDap9s
R3rR0be15hzs4pBch4Ae4ADwmGJtycmIarEUSTMgVrWGFRoda0D2IneHukbyMXZ1hquuqEP/JGr6
s7xuSjJvhya42E061AfAN+o/+bMOn3B+Y1wtGEjehGoXGLV60bvqpkd6ZGox16cqaUup2AagNsUQ
IuU3GIhcXOpqSY//1u/FlAm5nDWQmvKHHIj2wjWnh5/cZjOkMiGvibRk/ylB9z5OknCTKbC6lY2/
cVCDmB/KBRQDR1ltGTnFgBVGA7T8gRlBck6ik4scA6zhrmvMa9Jc39OzaXEfxlXyPH9VqYk7eHdu
3xcmBm59Vfm0S1qbYj2/SXKWRxIbPdnuDQQWA1qoohOF1pYpB6w5fE3U7UxFpv03dPrb1i+kqtz5
q1qLicd6HE/MmJsXOCgnmNqH6MPIMxPxx5Fjjue6T0Siys/bqn6is40JUwALWWDzfuUEaALjGOQ9
3/NsFbzTsYt+peRmwrwRBXKc6684wv/VqzyzCzO+L36y3HnDxG7PWmyl5hj1Z9iUKBLmvYtgDEG7
S3gmxsTkEKsR7lot6VAq5llDtXPVITU2Srr6n73nYnCpahl04MX8Kqwc0YsIewjbQrbglSOEtO6J
VCeWTvoWJ6yIwpCCn6MPtjiIb/C3qJZVJ+IUOjRh7w3EE7Rfg7hJ8rbBgt1Hb4q84DvuvmaW0kj7
/795iGgB7w4YuYOGEXu+s5/a9G+0Rjkfu7MncsROMk1B2xewqs2ZZkrUtP2sCYulgvL2ERFNsRM9
dCE5+IHQCQqHhVOehImDMvO/QSARaoiwOFfeHaK7sYpe3XP8oiqdgRgrT6IFXe/BCLnHLNzXtyrE
Gk0ImRNguIj29UxrDOGKOMVsK8nWEZ5IFmodWgR/D25myXxTKRcpaSN3Z8EGXZkPApK4Cp4tSmJ4
82z/vkTiAJowRtwyEQ+aip1A41uMPMTaeKPS14xM1oLMb5AiJgBy6mA4K+uDtetS+kVg8zvBLDpP
bljx8JtjBnXdK0o9RnejIFTOzqUHy6nvGa+vNQVZ2dtGvKBWDw6T3faNiPTkr8XIBmmIBS/lQULh
5TNHEl59l7x6Yu4B9sdS6x9+o8XHjlW6dx/5EXVGhdI7DBHlb28LViO1HJFryR7auEIqcF8W0fKB
vJu6GAvAy1wrQEKoN2STBvDrlwsnK9PD2SlXYcNN7aYSXm1UT8/ftfVBx0m8BG/cpkwZB+b+2Ksx
WJR0Ip5RL8qAFpGQnYU8du7N1rmxuhS2bjIh23x/y0Y5sMq6NTTA2X0Ry3hxwXWPXqUDlTQ+OxaG
Uy2RqFQfUQ7W2xedmlS12s2JugzsN4VrLJAF257oVZWZMNiBXLvNGxOslyrBBAKfVP4/aBNwnP3h
chdJcRSbw/XaErk53xeGBmUak9nx1F94pt4E6O7aypvlNoHBDXs3Y0Mt1wOZXXnMUStc3Jc5C91g
WPonEvi3vyuIZXAO4lIqqafVwQlRPuQwrei9QqcHEKS4EZJ3lXaxYDT4b2Be9m/dTGZnJHZoGku5
stVOamjSmDcLo1hEtTbRL99hfLLVNgLryv4+l5sDUbXDUdY4zDxaWa5Cf6fKcgoHiPK+cSCN0UmG
X1bvizGwGoFJ3Av0nH0z6wWPBZMYQLPg0c2Vq2q5eVZ36OQI59kH87JShsQJStbzpcUACLod/Nmi
EEBT8sOS9/3k2EPK/4an6+4ZzXOFzckqKk7QX9xMLRTlgO/Jjf57RrMDZxKXzEh/TYN+kTOBFrVo
Y1KgWWbCNyMGDwwXTR+TkoOCb8bwGi8V8b5OlItxQbG73ln2pWGdHnAPqa/BR30zZC2LpioHR8UH
oHssSL4/mJ002wCdF3vPpA9qbocMIbib0wvpOAcmfhmsvKf83QLi3p5wXcJ2CUTbP9jTOzQVw4Bd
hcCC1U+oMUdeonpQdi7eyySZQR/P8oeEGuZEqAcQz/BEjW7FaJ9X26Jh5dnClVMYoQQDew2tdxB/
IlrgOkCHKTN7PWJYURrpNqfE5nf1XN0QfbPR6Ab2/zeFw3X5pyTCfu/5ApSZgc7Kw3VvBRMY8Wbc
PxoWx/GKBkh4WtO2fqPBXXxByxI4WnQ10SQyjAJPkRhpQ+UlNoLhz+5OCuPNgn9YrDN4gDjmLJkN
GoKUHGwQ1AgvPA2C9///g3fV2BQCZ13PzfQR+R2C/5RXUNNvDtx+lpUvNtHPOOQ+gKqLLJZvUXKR
lqU4jPtJ1P3JeTu7IvDPMBe6jTltqot/46BiwhU/6fdr+yfossFSe7Wgzfxa58Wtk2R0s3wYLSRx
2ChjSNEScDv+gkPWXywzL0qbgaYFiLn9MwXKFXz++wYfSijXjjS0Mu8cixwq7cYCH1qYIaPyiS5t
HVamT95TicPHEUll06JX6pesSWqu9Zg/33jwnOaHZU3sjIEV88QNw8Q88Yjvx1QtuuZ4JjiP3tXx
bK/wuA4B0zhwaGERSeDYf5xn7ePCOBK7E0oXOUSH6LApPjyE8x19Z9bgwcJLioTYUE3l0yAtQoWE
daG18LievaxM40cPehaLLtVtAgGzpOpStYK5n3v+4ZXov+cEc9PtpNjfb21oTikgMDi09/3NAvBb
eQnmXXYtCzSjx/cEpenun8moiyz2wFddkF/fGV5o37q8rkfJnidyjBDP3BrTZw+bDxPDHkx64IkE
L0ep0NArZCASFxytp2saiHbA/HgTr5KKTehHNX62I2tYDh8U+uNplH9S6T6rP7CpgW3TW301GLKa
yJRDlNRyrgL/PQK6ygZW9mTEY5Lsr8UDRPkhC0EtO2GDaEMcFxb4Rsf431L9wPFyrTF+ACqYjDTq
DlYRlpiFXPeXYtc03qel4FGLa6rTYPxvO6dVyPs36do8U4G/VGZnQZsA1GnVjfrn0q2E9JZl2Qnz
VPjol9C/cLOJ9CXOLq6TIGf8scZaqIZLAyaW1HAH9oCsGVYXPaWVKwJT6A1p/QJf0kp7JD/O0Pkv
dLZPtBB0DZsZCZtuSZAqTxycvgiuFNuzQK11XAzwQrYsxn8lbc+IeJwe9zdTwzsm6k/Pkci2Jmt8
SrngAFvIgX4QgmItmA1xNe+7Ue1adaqWNw1v02i3p0veGhUAl5z/BtoK4MhILNpgr2oRLhSWDb2x
e+X5wrq0fKDTtPh18VitBDe5DWw6GWF9SgPP8NX+82gw5IdfP0Imw79daPL/hVHyk94sQpVe53Q1
ShP2epy//gKzGfORqKR621AZ1CEcBLxnY2w2KpnITz8PNlHEp6q1N745hhNq64n3zmQnwdw1IzfD
INqeLXhpv2XXVqIUuzXrfNnbDGtsh/xjI6WahITByOMePawKQ3jILzgIVvw1okLqsRsvUSh1pMJ4
kEFAA7gflwiZaYjBy0qRuXgvjKgVT/4dQ8eRwWrm43O62YkIGS4OR+iR7kGR09oOpXgnbhHvsLXP
tj0FN/ZMYHbjYK0b5Xi3k8TfsBhiHTHkzOYytE/FULZ55QzJkhSJ1g4VQcnPB0WrhplSx0jrzBzu
jKd5mXB7aXzy/HMngmrWtMvMVlIgHtq1v2QtLHqFTRJsIijJpnREoX13tuFup4aHV7gVr3Zyi3Hw
TgyQaGqRZrIHi9djwYd23Jv1HMreE3fgGrJydIZGxxY0zePVfEyTEEmvVuobu9MtyHbmAZ1IMX+T
EpBc/rrfoqAgPHCg00sqc4p1Pk4692FsWfy0+KBuAK5dnHk6jEJ9zuRiFf7hPokODznGjtYWVL2w
M3KNwqcXD2QAI6xnmIYIaPJ0PNm1lNMRaSrcr0xr/UUmXuRiFlxshYKvTwdKKS165/kf7QGRnOW9
dStLkOLRADvR8VKXFSoCty25ucIi2coRxKU3G8qwcZXm07MRhdCeOJzJUEIMIl10GfdqYIzYphOq
0fXEf5yVuFK7kA/jmUXIRbCPxgCeg8C+MuDxQZ0IfwLN2/DC4rgmuYhO8J7SytI1q3yZGATnOKHp
TztBj7SGnnXb2/suBwGT1KMFLnQm+9GmSgiguCW/jh274B0MTzVuQT7dPDZATGlkuEOMsAWvtIlG
cmDbei0UN8f7FNIDfYXbwSFPMMSj2QPoYEq2C46fM9/1XTHi9mIKkwxQFMZjGqrRdsd1X2BsUEVr
s69bDXo5jmHtosjFGM+5FQIXnEHbwu8CNF/krvSPWrDVj4/cN2fMNLuLPTrid1ud/6AyBMpy+G+W
9DhH3nO+nCrHgLdtDvwEoDgpvOaRbszu09ZvozzeczuwhN1hd2MBz16izz0tEfcYt4IUV6z8CI5V
62ByrgWt6EJlB2DVP0EbmT2BASVp/Ee3ry7umKy+YI7BjOGK4v32K1SuugRP0lwI2Dm4bsI6GM5s
rLMKAPfQxZuP8VsgZQoiskNxsw9UN2xCb/xZmdLagZeJE8n9u6gTU0Tj68l+wIZLNr6XP9nqxqAM
xaV5SEU4tH2Ht/wO7eSdoqyzggOIxozGyWvHmaDe2peUiWiAE5okdXTouUMvRF6HJKJgDbbtTjys
ZVlTZJzAA4x8i8btoG3ufdKWGF0hrbXeOb1JUFqpPdXGtDZWsPnr4oWxUq2qHUwzena1/IVD7682
pMMDxibzFPwdxnLdHkC4zRHJYrxedNWWORcvmLTO+an96xRyUVg3yUUgBznkXc4MqWWsnUxkkJ/E
OO73cMOQf5qmohpWleYxps83Ew+z+0uQ99s0/jCf8IFPHq7ETw1DbqVLKICd7atj5yTrFB6RK8R9
e37A/q48o++q6Kms2Y1BzerFlbLQd/ZXZIlJxhTJq1Zr2HzazYFg0mbgJglCaIMz8s+4D8gGpuh5
z8WBxwJjkduS9VIBWghs2wClauAbNLzc4HtQ2PzyK7JriK3PIXJ6mAR8vZ0BzSfqSNMQXw13GaCy
zgMZ46d0ppdIfeF3gP0uTYcCzn4mq5OU+7hRhKXK1fSNMcyOtekEgssAkfBb98KuXTLev272Qt/W
tVFNPHFvgVB76r1G19m++yJyLFICSK+0Cix5oQ9DdFKRsfDGL01LQATcSP+5ijl5AOhgpBtee3E/
3MuUR30ZFKlz4CTDx2RX4YHzTXPGfxSmgjmcjDrIhq8Hd++rLTBmsbxkoxyxdra00vgGjz0x4v9V
e6YZeo9fO63kzM/EnbJGkmglTLSv43VajlE1CXn2sBjhWgwtvLyG6+AXoI2GCvD49R+Cd0PRH+fe
0gy0yJLLKQGfWNm8irv6DsMYQVDg6AfT67Yzp46hLekyJqwu+8xTi4DtP2m4FvXz0eWwDQx1dfmd
iNZNGPBeuhad+MD8KvMiMZOuhNN640m8l1S2LLc+or0tE6PsUHEG+hZbxfWwV54GuF9tAMrjjfU2
kBj63M5tgSkjX16DYdSsniv4d+UqaLKok9wq2k3TlwMeEIqgReo+OUGmQd3ROz82v3AN2aPYfLmu
+BUTXwXpD8N1Q7DUGgZj/N4RjXtLG/7hPpuhIcF2EbTgCLw4bROys5pccs+Ui1n7+LSmQxV1+v8Z
7AcpwK/rye0fVrQZJDnzzMT7bplQc57BMt8p+f9uQ4PeQB5r5rXyqYc6vtaN2/mYPLsWqA3cDTmV
dL6U2OsPDoD4pkrT8hMMmAbooRLfsEdjWT0kygOJXfzS/HcW/p/u3NmXLqO/7nTQ8MvkPGKYEsvg
TaFCl2UftFt5U+byEWsjEVFudx71505St13Ll9IE/NkN49MESzM3d3L/SdJkI/OmQnP5VRFYQEAA
G93vvqYTwRL9P5Y6DtaENw6RzxG+bXTHpmkpMBs/6Py1/4LKT/EL0/1YOmcngJBb8CEqSGhjcDYP
w6TaGJgYfAnOCBmv6yvpuD8p1byKgANZ0hBCOI7XUC5STxzt016TlAaP5d8Ks9xv0Ty9YiHFuzO+
IX/MRO21uR8WooHe5Y/WlFE3tDzhIOu006EPhkXL255NoXdp7C7hRdVEzduXca4q3c4Ziq/yUDI9
friTPuRwzASUZj2nsBOqo9kPwJhjfOd0UEiXUB3bVfsFZ++BpxedoUyfLb7A65DpFmYFGTArq8iW
H3Zf8dJ0Mkb1s09WlvV3F1vKuPwJlhyhzq9tdMXjyzoUixS8wnYGk7eD0FMX5KrqsOujhQCT7AvS
8Gyl0zWLzMF3Qz1aLSYUTl8bOaghKralE9yonFxQQJsbIlkJJiW6S2qnPDskSQHBWHjDDQab0CQr
G1b0tWDeyT4ROU0W4Do1TqIa0V2llNj5G+lB0ozM0W2JpBASq3ZYIZVrZXfNi72B0RBQe5JAV6yk
/ldD7beE6C2EQSGmGGe2TsnKIcf51vt+XkVB7VrKeHrF+NGytGZsGP9umSWdoLnxu0elA3KZytzN
NFhVTugRo8nZNitQK6XjS0bruPbFt0h2kRT9w314/MoDhpcMRy8ovRvogA2/0As+N5HlkOKPMDEi
s5Lzp6HWt/JE0xAJSABK95l5QPdSTQkzczPEoC43kek8A8nZKJXnFmdVoyWEM9NnV8KJ9m3bgvMJ
tbyMjQvUOCQm/9hNqdvFgcjR7hiSc0EGt7ZIilBfge+It3VMkL1wa6jf4Ow/YRKkaNN64n9k5+6I
WvYtpDm0ZVo20O1Dh2aBJwWva8ykxpxJ8yJZjVTMPVtL4bOMSdSiHKjIGK+dhw79SQ7/fccZJHzL
thQd0KWOO2HBJfok8dIbx3S3z0+FER03io4iZSeJLedQSW8oRuT/1j7rFyfeJDN6HLADHV36XJQ0
Uq+zMiDiUayz2ur+hF7vUXuy2r5X4MaYXXN7Vjj+LehbCCUUtc5Rknuhxqqd7g4uyH4PmEqQIbhd
jpGFpL5WFTh2v7YFr0OClJ4vJboAmtEDCrWR6qYJQIDwY2s1TxMXnx6HmZe8sF05gCP5XuHJi5f4
+J+Pn2naxUsLskSdGz7zjEovBea8lE1ftq8VpGbwZZFkU9l8+0MT94+ai8l/nFFzCSKnikmq1xZ4
NI8FZoRaQ9+Q65u7tW4LirnvU3eJtFY/8LcnaCM4ZJxH6oJ72hUaTs9iMWoyMcZcjL5SEDETjnq+
qkrB5K8gJ1ixzD13u2kDD6AVcSiBsgsRJQKsyTsDlahcv8TrtfMcxGqZdOSuTC6zFTXwYILPsIVi
URgnI2qDeGJvtd2TERhVxvTNljFp2CBl06f5l4b0ceX/aTGfR4DsbeOIoSqhrKufb4NuDpWEk/bc
kl+wN6ZItgZm4Vb0fWnAQ32tqHe8HcM6PDfN3O77wOe7wJbrS2OrT9P6Y7tZ7xN/oWAqMcVleRsT
zjNI4zImLQwJJXgtFeAt6LvbRZGkl82bJkkEMjg7U9qho6uF/3Nhh4BFkdiMxuwwZov/WzDXPIbG
K0DTHk9ITgFm/r4dESxqzqMcDflmmYzGtCSElcY6jLHYYOgOSatSiKs0MtcJCZg+KR1vDbtuAByG
iszrgn99nPpBFFFxKJVY4tXFlnZcPTaZVir2YwKTwxoP2ZrSnWhko4/RS/RDG3sBOx2to+V/17S7
tpmi0UccdIICF3/C7oG66OwIQTPMKfTyDu0vICfA7oP3MGRuWxktNcF1oT4JoNP1dEPaMWY8djVJ
CqhszpnliCbSofaFIKTQX6bc4oiawJjS8sMZ0304Y1DBM8nSQBFWYiAwEd9eQB3dQWabF5PQV+Nx
waXPIIHKFRp+CsebpTD0ZsOfNG/atFSjew/p9yCxYvBrh0Up9Y2zNihmW5u/purQWgA63y0JGtns
z8vFwGFE96z/fFJTTyBVaVJ1x2STrq4ytm0JpJr63eeV/OSw2HUtzfTykPVFKUc6AmapDyzDFAc8
KXdWk7mWjrD+Xic+VdDS+/bp31G5is9mnFIRDcskMIH0NGnuotojlVryystO2y4e3XNa9WKN67F0
crRiSge5NjDoVgG/K71qRELIgyaO/PrAe5dxKVW/CkJAE2P0PS6BaGAbta1RuDqxiQbRJpOgkj+p
qJ/MbThmnvKR1ktqe1f9uJXQCVXUvp7h2T9NFf+Vw5i1d7EHiNFwtG2zfwlbUz0KQ1eWRefVnFgu
avV7W/pJbQbhzwSSGUCqHgCdto9QrsIOz6yNdh0rClhHUZaVqxES91eihGQ/QSHFHaOrz/eBC9bY
WxiyJOdqpZZeU0X94wd58on/bbiYo8r9B7ipgg06Q0JbOyYh3xMgRIfCVMf9TOmsIXqR9TaZS+SD
rukJYl09RYLwA/bxpfN4qiIpcGDOEiMAbeeVYo1GmRPIlfQ5gn9w/37sLLZyPfH4Z2dvZySxYmtM
IAqXEB4SLiqUJxtvXdimJdZJ+o2HOtRuvDlPLyw5mzb8ahyew3tfA/YdFV2TVN7HL1ewlfe3N97y
FlIJWLoLJqaRCm+ScUg2j3+V4KdHOnsYaFUCPtpn1YNOZgkPW/hiBjE5BS3rfxLdrO25HF6ZtPXr
tB1KoDU0EXWFlmDI46amlwDfto+ApsFZHFLRcy9wrhmcmzIvMvZLL5w4V20Ht9Poc31OC8AshWTv
7syHwfyezmGEVRfXOE9/K1QXfkKH823rOJpTikMEF2ZhwMi94z/INHQlP1GGrDjE+L7Z55A/MQ8r
7tMEOTQxZ0/4XoRP5IRE0aetdAOTAh3Y7LQ/aXPeGU9csrgmN07hrHpjEH71S6XiLn4LWSRcYVGQ
rICtOIwFPOy9MLoibglsD8vmA/bWPi9iYc6tAkZIXJ5kfGd/8le29w22SDMH5mgKL/xi1reX7bRX
REc6xepdz82/zyAklsigAqImgxohb9PDxuArjusEBkYZVxnrI99fgxmWexJMGYHc3zz/fQQ8tEKD
k+CjQFt2AeLUW+j1n4Vyh/hLbjmfNYjPS/b8RQjhEbtqdK78MjJm/m/3R9ZwgBMWH/DMacpgBS87
wk9onQnQLLDUdZG/lDlLU1YJ4OVAswJYfU/MEb4Aku7TJ10LWt3e1pQ1Q+JBV6XAy5hHvG6rbtQP
WiCAWt+9aPD3N6uLfW2OjkUD6gBI7Na14UhX2H23ZiUi8UqPTCpKt3+5wBwxzNarK00jD/tMBjHR
tPQAD6CmzEVS5uffQ2z7tfHfW+PQTKqtK4c2jTTL0gmAmlKzkO9qt/ipnau5yU9rcKtI2awSSJE4
JTMylKcRCBRP1vCHqSiazPtUEfTj4px73g9+CA7JTFj6haRkJptFcViJiLEXn/lBUYohh6h4PJmV
u2op1ElPQc5yNYe6iGi6k66Nu60FiYjDwdf/NQEUkS84zbRs5UHaf9JOJZqGaKndfQtwL7G8bD4d
PNWxGUO1Z1aDXGZ3Mh4pSbPZpuUPoESE18kddbtVthtDDGEm84xDIDZ7059MX0noY5u5mnLtd0Q8
afLN6ohHoB0j+bRRW6e82nndtE9yhn8rW0uDm8HxXzNMFDOekeUIm9eNVz/Bzf8qbmsX5gVQw6UB
KGoy+B/tOcmmvMSy4kH1ewABpplDab2lQ5oaOm9eEoRXIxctfFj77cLkWKZIarzQ5pe8ESKM0u0n
o0ByBkWQnzgMJa1zUeJUhkdru2+DNp8EKmi3AH6EyvlZgQ3fvgs2jcIWPGJn7Jhhljtl91OgMsUT
gSyCOCTGTwGpAciPwg4Lv00u28ZR/RKfxblL6zCBdXVgrHzfKlCPO2N+y93Wp6eSIhLCydwKha53
oFkkEvZE5hEGv2j+ghOdpzFx5VE0sXzT3/XqxfFEKmqoxINF3aCK6lJICl/OpAdgCYvKFnCzQUku
VGAG8WROkD/nLQhVusXH65TN2jqW9uYb1582kZdmDdylyM6Ae0AcZcZq5hBgJ1v21WLYiWYX309q
bZQmkN51j+ZzhAyoQRX0VrIEUK7tS8ePXhF3eSlWuaMDQAAgZg3Bvld/QL4chfcelDoRYXZsxzgA
5RUVhHNNrd/rDP0pR77xBRWWqWa/21Fk8pHR6Z8qfCeRoyvb+8dv1dQ/6SLMzqWo3YtBvRODoCVr
vikrmcUj/GG9KLkJy6Ld+wp7IKlPXbmg5oXiVDwywSc8d2IvbTboJdU+u6+YyoAKX/YnK/DHaKfI
L2dRmd0+DVNzq5GotCsQC2zDuvBrNw1/LabXGshKb0wDEWhjKQpArvqXzkH5gKnkwAcOWq90a5uC
kLp5cY8EiRlP0CMDEDa2+a1Yh+gAx6gmCCTGtVGHQNQEcvtECoxNvoC5ekv1wfHaF5aMOYjkAae0
EOXfSm2qHw+UKkjrFjR+1PeCcGCqpLXq2zpg2A4yU8hGSd78mHKU3W1p1evFO4cm6RLz5onJMBzN
zZflsGacw6qr52dX8QS3rmuG46cfcUtwmmWILEPNFLWMII2oIXbA5n+GwpH5hTl1ZPFUmLaOYJFz
Sdattfu5HbxnEz2CAWlFKa1xvYqYycRdBl5jaCmmmlwDAFSw5VohmWddWlzZVdP5qE4JbSMEtxBe
3VpVAv5V/HDNOWlezcULcT104XsP2AZbKmF1QHl65VTHCtd2jwmEfF8uDY5IZp2zBvBMnD+xrYnp
eA0T8oZNv12mzeBLUC2wnhwi9FkJf9GC+Aj6Ms7Pi4vEixkUfuSRucs2lq6VXB8UPRbFxNQHAd0s
4pgeMh3/fGufKZurpiBZBSEmcer9g7jH2IPmSsfPHcJOmsci3MpG7VIP21aI8l58zHghRzE6m3Xh
mprgaxmgwHFXTPzwKFUXrHT2czo00xhQuyTdyxcVIJNwBDMN0PKpu+H49ypFu8wH+2XP0sTBqZjM
CFDwNEg8XVZJwtDb+S+85m6WD5zQ40QY9H79nT1+vzav0UMICHwnJdg3MNZYLIWOjvjhWNSEevDQ
5ReosiC7Ou/0eYAW9Dfg0i7CWgUPtD9WaXEBALXA3V6YPL02t5jRM/1Epm7b5am01QQW42b/vPmf
8xYc1xGcaWXNAdRkV++gR28NIQVUFevxFN3B4yMfZNeNeKrH/8xxDt7NQdchejY6CWAfLJXSNvEv
xwEaia9c8VpIfT7vuJowQTn79ZFEiCd40SOayB8BGMbqNlGGgOZIAxlsSoZsFVw2wJV64V3FDNoq
obC/DzziaOHYDkwnQY2JsVubE4T0FnghLyvFuVXGzjof3phYHUCLXxIKZBvQbzP4/Oja26HB8zIO
akD1xKBmoZbJov6O2BaG8zUgw8t6Wg8S/NuXAzxNzLD8vBmfPMTxOoeXx5SQ8i6RcdoXbpITlQXq
4fRmSimL1gEK5cPVey23HY6Z4hze9h8GMfRH2ScBDXqY1Szy48Y9xPKzytgjFt/qn0wP3D+p1BID
sc4WGsTz7RCVOkM+VaINCtzMwQ++FuBu8egQQemY68+BaG/BPj/z+U8C0VZcf/09gFHvek3Xrr5m
XRK7sUcn7wHKhvDwddk0e7tHTYr9+zUVmSTud7kdaoOZCC8ZGAAd1e5OFHDRz3vnLU31Kiq490G+
lHTwKLyAiu36OHpXE2kNGcI9t0ULbAstke2mGmIesFoJ5wxGZJ8wbtWKFHumr+tw7VDqz2P6vVZJ
cSadCYMCQwTnXcfa3KfvcOvMXL/kmYVKkFjz/DsJLHLwu7GgGzZfEjLPxoq8x23Ld3kPaTA0GDtL
F7YsgOJ+HmaN/VgWM0zlPIx6m/4EjoUKUQ7vXlO+fJvwq8uKIZgwm3zrBBHqQtGlGM6OWQq3p4uk
AtJCH7cVX6u4W23GSSh8ufSqm9lrpQqH0w2M6YgHTjz+buxplnHDx6HyF1DVLeN8OhfLKylpuA1L
km9yArEpVz6w3auYBkW14ZRPBfdnum9s3agn0Su6WE95zo3qcg+GLusRRucDItApYIhEG5zNef6G
hZ5if1GRStal9f464bpoBayeOG2hEvEpTzSUA+LC9uRCmlWdRHLEfC7IB3S09mkiCQo0zovW7/5E
GzCzC8XZfqH8K2thXAaWCfcfu+/uV6am9j0MxnxHcjMIbbAQ0ycV4GYGalNlNgHMcqBUd0YJA5bg
TwgvnlsZuXxnvklZCWETxaunIXEX1fkLAdzUF93HuzvOuvJd965/FQchpk6cDK1n2zkARa51yh13
D0/+z+NwWr/Io+yEAFpUURGVaRjWMaTF4sciRwR0LPZRWGMB80iO918rrjaj4JXUgG16HyPvVlTL
NzClC3HdGxVkH8ozmEt3nnCyIloSFBSwbaBLZfF+B2xfKVxea4A8EyO5z5UlyDwo5HRcmhxwpR8G
QDVq9o8xOwI26oLjGu+rFEH7ZpVVbs8oopYnhDVRqFsW3V/zswKispRnxGG1Q+L8nKYvjXbhGU0f
nRFvhifViDebdgEbBX9jOmGpZ2oIW8tv8wg4UHINihZC36BAanWpSsGqbsZhwQmHQd5JYXI//FVW
QSSTkvfrJST2csE/xm1s3eTC58e40xmDzN2YeOnqTtD7iK5piMcYvpZGaRHRu5DOb4ASVK3vkenN
pAE1+wg1+19VQc5+GrH9Nj6U3/VBXrwYI8iDsrCnyL3SNYGMQUwh9BcF7Xkf8wNpI6lWLHTiN11P
ZLB4ZL1i6jMLrE/3HelM+VIBgE7q7z+YmKsHt0yUuhG2Ka/9DqkBBvVoP1aFoHzjyLpHFkOQIunG
03OhgOnAS5fMVy7EQcKPsdzNMl52grQZkhH39wb+a1xBUPYX7cVTuygZoAd3DUN2eNwqgjZctBRV
FK2xuW2UlIEDEwJOZXQT79GVHXTgQVPBTg4ZTV9xry+yLwswaeCru6VTB5WMdaVNEoZ7T4/T2niW
34hRM4N2cLlF52vnuC2jore//3s1rprT3JWepZTHv0FHQC3AoKfQ/PGNOfItJ3U7cMY+BGNoyPLw
4aqfwRxP9e32g5Z/ZHhRnZfENr6nqib7zra8PDsz9juztBFBo+o6t0SszwVHt96tk1yLERMknnT3
BbGsHUhorrVqOuzcA8/ICbG6NewFsEwNYeOqNzLoJ6giECBBfppMiX/XCHRcdZyawEKrMmc5UvrH
5opqkBg/gp2hwbozFUgCNxCXLvjeVTrXCgaXfu9A4WOsuHDdIh6UW4qQaJsIJxXA90VlEr1lSwma
uTgT80w40NBjOwJhy0qAhz7owDdDzUhLxHoP82WSxjBdB70TltFmHpG7g6YaWNNXEPmeV6pw4hTU
OQ9MlkxLMJ6HwXUldoMolZJOSt5Ogv9LA1P5L4L66UZnoN+cr+HSsvHICEm8l9LwGj+9qfuy91iA
fPZOD7gKctOFl/5HCdluu0qa86/bfS/RWFarUvRqKjWeW8nazGbm9ps0l2FldL/gt3V8skT1Pbv1
pDbAvh+BGRuvRZlMG3L+alCVVi3t6kS35/BLCqjg6ItCrmfGggXgb0hUZJZ6gTgy51VIJcL3USVu
BtU3+sUUTKZMFlMVMiXJzK4G2YSJgDM2uv9YKU6VB6FkBmON3CJOQ4okGccOSQll4QuGMnxylfvQ
721PTg2Wxc8CG1VqB+OexffJbqplb1x61jyw2plMIb2zhr7/sV2WdQvhjledUN2tW7RAnaT8mi5A
tcRq/kIcI+l+Lg6X7xnq498xl9SziJCDpGhfui1RY6k2nVGoY1oDI1fvQrsYyY9MAbCyhHDKCTjT
psqsOmUbqZ7gjDU+CfNsyA11DXa1qHZCTfgvOWi6rdzsmZ+/ZkwDqa6BDYJG8ReVQ3Am4CtHvIcv
ojwqWKSoGqlH/J/QXb/Ume00n2/YpTLdBlhZEMv5LCnqmNo2kKA7MEhgjCzvc/+xH1ke1bbBsC6/
QbQBjuI6f+wSSOxJndrFVx7IheHPOOcNBX8RgH4rJ3DM5+qsAhTS68q2u5jCe4n2finYtUKFPqqP
UMkmWbo7XDSWek0gYz5sXLZ6WceTowMfkvBHcaxOuAeyXZfbCalyYVUvOEh+f49K8AvUG9uK9xku
7DDJzoQQA3CRVxE0LwNctoXVeqStPKqcMMg7Lqble5+NkhnYlkC/jwztM6IcwEzRZKWP5Pf5rl/L
bRcAxyZNpcDXXV4c2LfHrxud6iTyA1OzoYKE2XNwiZqqtQEEfhvVl3nSTYIho3sIYFaa25r8dBPX
s2y1ZC2J2UspvjVIXRnhWTjmkZiLlXo19WS11htJfwadpPuAwXLNS1sH/FOU2D2WqeL8sLcmV3QU
71mq6Zh2Jcrd7IPk3uGHP+X9wOBne1R57hDruiWyybhYyM9sNJUcj0WbySC1wrHdfcIHAFDd5ssc
0yhQVx8MpEG8fad3kaAcQpBRjtZee2CIsZR4CSB1mssmjcxlfHOpi1U/Sx02EdT5P+mulNCRMrxU
gdDWi2X1txYtdeRgOEOCOtfVYUsDFuOjHuh6NDCow8H0hY3qrP4drqfXQv6MQovS8Mm4UdBmjFV2
OQj7Rr5DUfpN/Xi4ovLXdfLe3nU+JoOg9+rQmxRY3kP0CLpMNjAjvIBOaS7ChEI+AzpRTngYKh2H
t8xBtSER/eciiYPYujXGwawDCXASS36BMULGGhVh4XkogX9b5AXIVPwHsTJyJS3j6/5yD3yx0Dz3
N8cbiXQxV2lywApMfSJt5iZLTCTC3XXWhKnwvAyqvQZHjxvtkdAf/9ZvVvGh3Ua1Yjf4fNvrkf66
Lbiy1zLNjsgREXbW5AZND9aV0pQdytNCUPesYG2ecygBwGEET9bGjSeayQemUYq3TKqj1SarfpA2
iJCPbtLfuUvC3/QQZxhLT+MuraDhumAfCvtz3IVdy60TQj0ksqtQLQL2SJqmtvabwzO+9DBTH7wB
QqY7uqMs3nyMk7OSERC40pZMtJbeqvwo4stHTkTYP07fv/DurGcjuOig5hnRe2Xg79tvTCdAf3V0
A9NFRUdPWMFqVpRZVKCO9XmgRtStPXXX0lCjnA3ipsrJKWPXn+Q3Mipezgs7dt8/PGDZv1ePI5V8
CzHGZ+o8Zc+CJl/r/eUbTc18MsoKM4l8tdJQNr6mmtD6k9d46OPa41CwN1MUonkHYwUp6r/xWLt+
N4xla4G8Tjt56/PXI4XsSjfDgH77j+GW5iPyhO7wcIWDzvdS9TCGmn69CW9WU5D+T6mpzWWNTOWy
l3wQz64E7x+klTxeh2H4+Ch12khek0o6GO1ZJ9wN9pXWYFRpWxF1taYSQBoRDaKHFdvCU3Y0bpYI
0NvUxVDdoimWxDJeH0m5R90V7ufzXbDFR4lBg8gFrv5QBtturThvk3p0uvcVF/acAO/n4mV21jt+
r7CpsUr15dd77G27tBqO44GQuQCZR1reJrrf9hy3C/xCTjOwnCedBMa7T9I/1im7ihoM6SX/VUDR
xZUiRMw8T/UDL9Vbbo1CvEslvLy2e6+OvGczliLfrNXCxHwKKh5NDGs5dfmC+Ofdwb2pjJdZpgH/
wSf4BSkmthBomB6HkZddiK6JjhjUMNW8wlwzHDmPmh2x4IiNBWy0G+P5O6uQFWhQvLMFwBu+kpzH
XMWoT+7/YCmQRMf69kFRf1NosT6zO2lYTxkSD0qSbx3xh6TJQmXNiwVXn4r9yi+zJMxRV6nF9zxM
J9HRXZxgmCAwycBlADhPVqfJQSPxrczDp0mE5+dCoxRwrPLp+pNSjU2bYyLsQLfkE6R8yUBGDKG0
6Trh8Fp5rBKEkCBnL92N+alakpgGLRp2w7tZxdPurX/qSQRJpxmEjA5xHOaqca3agiNbpqdL4b9J
pXLjDdm6Ess/v6hmLFXZM3iv+FNT+yEcsFHDVqN7sfBTBtN7oEdhyF4vT030l5L7mKANbWby2zVE
3cv9XwYPAg9lUOtSCrw01k5CnOssVgJkGcJqZNkuEyPgxAjjfIZQVr6wXot8q5d9t35PTkT8FY0a
vex/G2DPuKffBB0KiYv9T1kNzP1PlKKeg/BwbuSyLScQZ0vEV79Q2E0TEY7k5qB2BwaEd0/jc2jf
RZX7ymX5JSgpwCNJakUI0KR1Qf/FrhoBCW7IFHL5eU8LUHJtaGXBjap3z9CU0yD6OaedZa7QENmP
mqUI81Ansam9AWZjES99bsr+UyiAQrKuJiSwThIOIE3UxTlgPoYpIbIR4iqpb2U1UXrZk0Ht6dMV
jlWsNgu9Yy3QCT6kdnJJ86ZQpb39CVLQBw/ZPfkzq/lgyWlx5fvuERimnl5PcKOfyzEZif+nvl6d
8l8u71dBgCQVw4QrQgKl0xzeY/8P9xm51YDbTLvgutWlrshFMO8/3YfRiv/2VBgvuW27A/qXWRYU
+z7bum/n1EsyUru8meoAQ/dBiVdFWZPzbgFAJYFGp0ZOcjGi90RUKfme+5IkwYK7yHbbQZv72tYl
a+Kv6OiiXm9oqyNUqXKPGAxUUJpWkryaBUie8e9T0YO3evZhNpdzr+XrUAZkoE2tm5y2OhslPLLw
1bhvSzQK3OQH11f2CIPEgPhLk21vgpejIH/rqIwbDvmTSBKXjE16ZeHfuSQ4F6hH1le3NN7FW4Fv
eTMgW0ntST4pUJntWj83P3KrP4kfKihRREFeGu5rwN36G/FlX53tFWG3KbYcdSXBCcaBlPO/IZ9+
R2TB3n9xq5BTdcpbmzbCND3aab4km5kdFZSWcgsKk7SetKDSuyn/ZAvp+X2ValKEX7dmTAOMQ2A9
ATotJtGkOZx2RtXN9f13rAFI0Y035S38XzUs90LJGEF5AmrBc6s1fVf57iQJZ/9LoqKERbA8cp83
B0EKULFPBElC46EhUSHaEOZwT3s+Vv+TgjhV/cpKgCNL3z7aF4/AVXApb/jCM8oe4LCKMBcXcGTg
4ldlmCgvTzlZsMMApWQPh2nsP96Lqdf7WGmroKJKK7/7QAMrLabQpqSAXED64pEnqoBvf5utGKJx
HrT3s3u6VqBybb1uNqfvmeluOyV5doZp/JOEg9oADMEy5DEBj9mhYm57nqh6LX8uyPP8s1icRbxF
Q6cey3kiiT9FNYPs7ZZ8tgdnGCYXboh9+tHFLykyMtE3PaVGheeGUQbWljg9FvPfzBhNeU7QimH+
2Pt02CBj3Z9KV1PmgKS1DiPUBNdDG3G6P38bXGHz7Fx0RlpFR1O61U8bSmIRifJ5BIP2xy+YMChd
nYWdZqfViJ5zd4LukxYIR2dGnHBZZYelNiiWoAwOrBkkTiAri3ejAXqrGXebU1T68Ist6vEYFcEa
9drUwCaUSNTQm7PeZoAfxB3jASNkMaabuE35dA1Fpk+AfPBoEYW/oHLjgMtFmxBuKeQIR3zBpnOj
fewQ/4WzIf3cLbPMdCdwRw0La8UgZQLHaPacSFwgK8oGJqy7r6LfdVkQDpe/Y70yJylUH2x28nmN
Fc8MVNZCdPoFJgYUeJaKNqDtk2tXAKLQUk+6qaLW3LfjSZ3N4RqiP8Doz9iU10R4/ulWM/yQArmq
97W7IpWhlDlnvS62/iErPLpdWPzIDbhT9y92EhxdmSU+u+TnxIwV6pkUIF5OxKeXM2P1fbXmMQ9K
Bo1nBieB4YT95gxhvV/TU9n0B6T+lRoIJaBHiyYLJwG4M2QpeppNIOt7kCC9UUXsVYd/46PPFgOO
58h989LcXqLYNE0Mh3GYWYFWJHac+Zaf296DHlGffI0t+LmXgSg80EBVnt7P9qDDsbHl85MfRnkw
+5TCJ+soQixiv+58EbZ2A3jw2ji+xCsOsxjjRbqZ35csPTm81UrVgswIy1hWvKj7eRQlKfILtXOu
vXTA+9DREW1/8gC5XESE3yB3T60OHyzS5eazVirQNsJeW2ku01pdEsLStcmeNl6oDbqOOK9MglWW
P/6x4TEU2chtGpAoEMTPJG3BBB1KcBvlvQ06da7yKa5Vpg7GthTi6+UADyhOBzEfZaJBnlnknjv+
MCoQLRNthO3m7eFO3w9GdaxFe3evt8emdJcZnvN+8+WfwHs1CkdUHQBPlYUXK6f7MsUvFVQA1VW6
k45bYvNd+i75jGB8nxHBpMp9jpK15l+Jx+trrcQHFnex9kEIcSdH9RvwqY3Em8RT3zQBHeUFd0Ck
uXsC8YkNL3oE0NEFMmd8ddTAnEZLbbIS3cfQJBQoZlke/9VraePo8sYeYwK0JbIw6NyNW4eFa4Cf
oNUJQVMIWwpN1hS+nbCkMDvekUAFY8iLdMvoMWUZTBanswxQ6XYXN/rbaBpfqqev81PwotCD5/PS
R82MZxWNFgE4hBAYX+RQUEIW/TYPFBEb1ygCMoCSIXN+QdltBfX9zOGAQJnFzWIiCcsWYUFAGvxO
YyXRaIkz6+8kz6xtrUvxRNxd+RiAj/ruw0mJiVk5V2vaq/s4f7S4DqKUX4DzdoMLibGe+avoQD65
DqFKrsqvQgPO1zK+D8I3jQ6EElrDsdeE1gSCb++rmMoZUDqD/rynEIR0qJHsZYPLMZqqk8BUmWXK
Kp5MDl3U+sbxUj1/jd4ZEmbILoVwyA+8JATz6gy1U3xLYZpb4ZD1uGRzy+qjQoRO8VAsSMEJzZps
4IoigUGXT2qep75HCwZVNRHjef2vZ7CPZO0uHIpFG9bM2HqDfv7a/cC6u4MB36KFJaXccChpxH5e
6zVuQ/gPbX9VfX+MOstt3cPM7E0P9fthnKR2PdVDNS9JMLPLTKrVJgB+rrgi+99OhWNZ0QdjjUOT
axvC0x2wkG39bSgLLD44mikyaovsZlgjuu+gT+pIE4Qo73SNZMNCGmsAGUUa5ywhohr62iYFY8LI
9/Y4H1ZjGIH2Q+hZ2wwRQAJ7xNVPgeT/J6Y2+4M5CzPqp9NtVDDg3JyzQuPpDS9xBtT4TitMINbm
iqQJ01dn4421dkrtGi6JdHbeA6FvTVyWLxoIQryOyKiuuSvOc3KEwU6Gl0jiwqr/c9KWCuz8clj9
vNOCKHP2bu3Q3m/R5+6AkfSqE2iTgakKdKukU4o5eSILjstFDzEzGU+SVwOJMswRLYvBlDz2rTpE
Vusfsap1Y6ikplLqbmyeq3yJpeCmKps28z6R0gVOt3sU/Ml0/EGJb5eQymr//m1ZUbmcTxo0hqVN
HBQmQYWFCs48Nj/vUbRCnxc9XMPc8c19sB0A3uMnSXAjwvXUhmXuKDiGM7X47jIOmvYevMVuoV4k
ez8qSwHxYL7VIPv92Org9OJNHMRcjcn0ursBxxEeiZXFqy2jpnGarX+Duo54187W6mTZve8meVGT
dDmuYezF7WV4D0eo98IUc+XLerWO6TcpQBlC3oxHzMqADoXakGdCrIehI5RIKAvZgZ7DChiRk6Kw
MV+/fVU7YqMxdVwytHvw9Rzw1rUoXndGz5wK5k5VMpAQG0PPaBnpuheJgcqAOdHpgSGDlnNu1ZWW
8BZ/VTqUeaxz4GxRgfA/7FzuVkq92vdzHpFSeGLk3v8YJw4JWYnCKE8ohZny45hltNCUE9e4Mdhb
MpAfsSB9vB2I7abor2ed3We7ZTSbbe0Wite7cK9YeyX9Pg4En21pI3BnGH6S8LnS4X4Q/UuvXI22
O4zZ55quCilFBGYc9tIyV74sybsubhhnaoW5PRc2YBfv7zOvn6fq5EqFRNBMPYd+p+Ze1LDniYsb
jkgACUZhXOe1tsVHZPYrLbFGXQdqO5HcBafFQXRM7YEYM7n5G2Rewtph+B/h0qSc0ukgU4IvtbxM
LRSiTFbFWB8Vdl8n3hibrl9rsOhq1ciJoTygUecSd7E+inPFPQDG5j+wblYq9KU1PeyJPFXJjDEy
k7O10Vpnio4tVK0k0m6mcP6lmvMqPcRwkWdqSYvThsvWgAJMgDoAL371GuGeAvpfd3qQhdCB+Awx
KEy2RtGTL9Y+UJE7ZGMkUBU7a/nvQ/fDpg0s1q6XB5GtWHrxUJkYJv1gmiT3C+JxkudZo9mZhJ3x
O2Ua6LamamfGV2siS/UIqwDBXROhZ/os7X/tZP3JvRTRX8505tI9sGZw28sWf4w/uz9pvseY1YQo
ilFl2oVUlGZ5umCWHyQpSJ+0gSBYjIaMIaKu/KVFIMSTLRqT5lERM/ZtlIzAfZTmqit2+/Ad+rUv
POaLsIlhzE3+95jYbqmAlfHCRFVIwLrS/dbWaWzO7e21giFTwQgZfur88YkAQbMljhX/McuwS8o8
4ePGeg+EeScE+vymNrNa/S1x4Z7gLtNOeEIJiwAiG48SRntsN6bLOwCsVN3dzS/UhGuDYe9z96BZ
7FyVEa0IjUw2glmdI2+qkoiXx9TXTsidKYL0PzAlXiY/cMUeiAWKfOrSG5jswKriP5eK5e8eOKRR
qJ4kZljC/3duQ8GsEiGvassr50vUX5aYc7SnpNMsfvVMaua8FquYullJnolb7L7pkbRHnSoHZxk2
cZRCTiAiyn3VMI6ru2eCi8NcUh/5XCfHwbXyZIp3cUin9XqmAV+Ag/LsynTpGGvntAAensUY1FR/
+ppA7UuGzFnU4J3qtoJjiUbhHxpwqVcv6KCKM3pzZiyg0R8sRmATYrk8l6xdxoqaJZ5quIuCJ/eJ
4542K/RKexavxp0TNz0fREriDFAtyAEnmAmPApOAuLtSqXTv0MW/G5MHOxIcjzoHNafg6EN6fFcc
Ov5fXxr1oR27DN0riRDH5yxZGgJAKuQ1nNWwE8FaU++NyDwLb96LU7Fgs8bK0InOZGWabDytn1Yq
Eo+qghvXs7z7oYoSY0Kd4BetQvMc6AHolDemRlnmxurCY95dCQ9lgJzTuZvWzl/dTwbTwl6Kg3Ye
sGsFPh7+/tXikb0tfMKQRAJjJY1mf22tD2E7ANgzsM3PtLDUDdw/QCVO7y5SmObqAKXE3m1QBe0z
7foE4U7+88r4HLgceR3MXg1ovSAXSC51D6OmGfTAWfiCPysvoKKJMt0JOf8WXl6pTBcE3cCdI5Ii
/lrxyz340rmxSWKDUP9Khx91gdFbQ5B4YjAYm42CKiTi1Z4yx6zkmOVjnxYVkBeDOl82KbsCbFN+
HFqF9kXgA6DJrlrkbEphsqJEhnjSvEIA5LqxhbY39mCeqsf8sjLqNdhsVnoqiDG6BaXKuG4U8cWa
piiDnhfEvyL/Z96Hc1z9Y7VgEL2fEGnRrBT0xvEaE3h91znbevd1NKOwj2rPQ7kmnIQ4y5tg4XEE
6hbP79KsFIJHZTWMDmTpazAQHdqgcDOnVlx9WsGVYzUwX6YrD2YzmBNLYB9yA+JfArSI/4YOlwa2
oi0Jh8fwsNMKVVgCNq9Ez9MmaZg87nyYqz05esP8Ign4CKQ7tU9yUC9XAfDchoN4FweKbXdHky6c
QzAIX/LBL5MgmB/9Wglg3xs2n4CyQAY/shWVk6SZ5CK/wz8bvkQxRh0sXsABqKJSaqCQWVdpi2io
xFrVP7d5DafS10vfRjODJ6Z7xvvuHhYEJyHi1J+xLwMGDflbFs0Hue4Kmg1wKxxDtEohWAh6DIXs
av7pHMQedXwWwOmqyqUgMU0Sv+mwGxTjG81UssGeYZodN5LZTDmgcsTJVho+ia3v7QlXD6w399G4
oaU9niKIQJR3hhsJNPJ35k27Z+CWywKa19AW2ym4XkkdJKJrKtbS5Gc3Ed0TLQuBRGe8O9jWoV8m
aTZJQIZ60CdvcwdzLnOp+LzjEkoSHEb/OyI8+r25GZRJi/XJJFBHS8Z21waO8aoiFTloXu4wQsWO
nc/vDCufv0S12961ObD60kbs/OtIBhsc8x0RKMfKmW/I3e1/j5xQJ1vFvEt9+43sFWf8dSKZBwg7
brdrTS5eAIaT6y1K/p50Wovhu3EcpyZVk467BjMwIEneVUzt/w4iI2NuL58/F5eCtl57t+tTPzdb
xG/zljkgDVPZehvG9j+r2G2aZv+bhC3vXTa446aa/YxkLN16JVzaXitNyM3wEMSlyAIHU29HSOWQ
cDkrkKgfqBDmEgoqCbC/O2cAA44UK7M1aTxYwQ0GVCDCu5Iu6AXO/uyoL6DiHbcwPrJzQsod9rGk
XaD3mFkNrmwdrsMhau+13javMtFR+hBrbiSuBozGVciWL/4GX13caDymWKA3996SmaH09mKbV6Bw
viImiVTTkCi3gyvD1jNIwKpKX4M03HMKai/yo++CuKshZUtUXBRY1aHOM2IPpdgXQ7s4TN2pFFEF
Su6AY5B9ntsNcX00LmfUcTawCCisuikoN4E3msZYzOCfrx6SphUuYfCCgRY8svCo5oIn5NJ6puRQ
Tvo1Mxltv84VQ4xZF/FeFqsTk9ARm61/8n5ktjgQxc+6DIGstrO0uN3eMFoNfL9LfbwTR+vg8SlX
KIjBfSbDS+s6aanENxuimmYLC1OUBSI5nOpSqQ8uTT2QW+J3gpMPgp23RSrC7vUwV2lwbV9aEtGC
YHuGHc9VzH8IRLEN22lunNlzczlv2KaSshL4x8Mt5d3tsfKvZz4iU/bCRSwzLWOeDDBt9lUQI3qO
8bot+fzVarPgNegGb/5nmtRZIuS2gwyCe4s1fN7TfQBwRu1lC2Y0RgSdFPZgZuRfcTvmfchtmccJ
KGXFQ7LW42DokujCphu2gfG/N4ZczjCWHvYYgmRMl62+v8MKRKQ63jDdmF6Xet6vZBYjyR3mcdIT
rD4CRRk5X6Tv40wNwe9TvzGLP3ZPeAQ/taNtefLORfgIq/cKgXs/PdKdnzzOiukV2jhqknA8EIXf
Duv1Hcl4Zj0Zpu1YtpjSKZWIKrsLYqABnLPKi7nviywkx4zz/BPOtnu4so1GFD63UvIysvF+Gn5U
62D33rZHwvG4binDR7NpIibgQ2VSJbPOPvvFRbFJN48UB1TlIIeU6JwltCXq92xU5yvsnvv7mwiJ
r8bWm4jIf0G4KCbOrmJGiHcMkkiDQntdlqqqzsu1BSm5dtFuxr17uy57fBb/W/H1R3u01ts9SqD1
6UwP+VeQe/0NuY0I1FznZjthFrfnNgzPwzRlgWGcChmFDqHo6Qk6YlsyejUQVQwFFw1um3hyL1yh
2O/Kfa1kSwTeyGvdJQWG6lYwAuc47CIi+pw9Qt5XSHCPhGPozvnso3ujRWLVTwI5kkYMd5EMqnTp
ChMyZHf9z6+MAzn6oyf1ZfYCaE8N4nSN0oyHPv99VOR1+QTUJJXUsVxmf4Wfq6GcU15X5yWsg3gq
K4LiI1gie4tpY4v+14sE4cAb1U5N1amkljCIeBymlJibmdUlnOT7RhKSrRacr5WcFvp3evlnLQZ8
01G2DLDKNQ70LYzN/1OdboxfwSg4hD4uJXgYc63r36Ou4R4GfE3v58ticDMOfvUof7yfzZehFp68
ifSpQHaPnBBR7NQFP5koH/KKTCDNAvcUqRhOtYOzM3SH17YWy1h3KkQcBC/4RC55LmivpcX/uUI7
NlR11S3BhbnCPoWPH5YWyjww4iKN+KvnRhfyQyR7PkvUDckzyvCcuxcnsPSGFvC9Cwu0UzFhIsH5
/1kddex9iEOFL6LeARQ6/8WHiqPrzpmfTjqwg7hazyRS8sBwjawAPn43cs6azv7QXsXFmrsnhVk1
EsFbQ0KnIP1gZIRM/4cZbNzidjkQKakAHYwkQnK3B0JyJ3ggaPDmnDA37rCPhHN9LfnpF3cbRXXx
bYaJUAkh2++j9plooRQN0/rEqFGJlm+Kjlv/dgGCocqPATiqy+eF4xlTS3V5hUKh1jS2gcVDYksO
BroNAaxNH1RtFxm31ZJg6rX1T+gu/F5Qf13uC9maYxNPRQvxL6Qidur3BJn6zzpC5Ivgzfs0tU+j
7zePKfxU827mRfpIYfeECs2qEz/T9jnTpXx/85V1PyCSqYBP82HkpXhAsf9OkLwP1fWhYvcBxF4m
kIe2HUQLMpv35i/69FBpc5zajowMp0+igd8pmGTMQipvxW/F8s0jbUyoSjYc13x9FQTxrclHOeZA
qJO5N/IZox7gwKHlpr46Es8sNMUVnZfc0GqD7WNfP0/kpLgo9Bs6O6dwPX5AWXgFHksZ/uuI8MYM
Byf3xWdPVKE4ESEJLL3eTWlitIezyCm4qlFOZ8wRWaVhYuIj37OzY/P66d1zyqtG86mfzkSyPaPy
SSIAIonwmDeo74DdivCLC/lV9cz8e2OpfMPyhDFOhXlO3iiR4Z7PQPuvPKHFZwqXK11XI0M2Mv1a
PaYZlFyptFZ3rhJcgYn8Sg/3rgkbCkxQXjZ5XJsaRU3tl/9/2KhGJm1DozXHxhjSFT/6RxQDajMu
sCuB7N0LZ3A2VzWTUEpyLohZuv0e0qjLDcwZfOZP9Mmvb66AdGIf/i3ndh/gkGgHpZzOUZDzeB/z
qMR4vs7MO0qpsvs2RmpKn13kVvXiTBihGbjpsXlJtJn/4dJupnEJfDKfWY8qkNo9kQDGRA82PFFM
wKLmsdfrm9ldgmYIg2ENLoUt/2trW6QBGtHe3SJrOKeZONqrROVdkmruMoaS2RFQwMZTPsheXWKe
hrNyu0supMUOMDRfrznCsdDD3l/QqZt02YsktwY1HbLgap7CrWyurJVfUIiNH/IGxcnKADPJXtXY
DpDyf5Fx3/N5EULjkEOJ8YuhTEwf7K6mnY/i0amjbYyet/nU16KmuLwxJ2bibJPAmaVRc//jDeFQ
yZRwVgUOEmN0lgQqByGiYlgxjU31ZkhWRC9K8eVDGClZA4NfQ3QjZic0YPX/7ILiHT4C2iObMq6a
ArS25U/+wYsTDtUR5F47wmNKYOVt2fAHvtlypxrpBJcixGbfRcmMqntfk7KxaX/bMZsZct0AvMDW
E6YnobVJSO+Uo3lAnZYoKAFIyCpXfeyqfuYnyGSbIKHOYKt/KSmXxMzj6BJfNft7iMuKEY/knRMy
w/uOtSi7Ec4SjQrSPnjd3F/FHsoCbYrZQbPBHxGnkcrK7SjQnjjbtjFmcOWHu6S8DbkV/YXkd7qY
JDXiRpTLQzDdKtr/+AoHVC5G+o6zKCbU/HLGqnm8+hX5yFBmZ8+F71cIjEf9wr9xXw0fCGU0DVD6
H1xAmVLgTaIZks9nsLFa90GPuOKYYr5Ih902R4TWqMTH+C82HAltu9OofVtqKlDpFjUJw2mbDnOI
dfER0PYBCcgWEV6Rk+c01POuqANVqGAxIdhWNf/fneyf1MdHrKFbGNEgZf+Fsd6lKGU4+eMPeVCO
YgI9YmecqQPLI3b4ZRDuTkxcs2INKhCwhHLFglcZTPio0ljAQnhckd6MmXUky+vJiQlOngWDZyd7
4UXSbO0dFNg3DQ4vr31g0BoPcOzfgO64ww/yhsl6jen2vNn12p4mw+X95FcuIPXWO1f0Qx9CFcLc
yls6oUBzkNHef+WA8yedzoZikA+U7LCKZOgMLE4cxFNXU7M6jb4zcMbWCu6wjR+OH1cng3Gngm9y
+Jd37OOId6BKuG9FZ63hefQFegj39AnZu9qnJQ0oNlzMhR9RmzaAZBbCBb6Ji8g9PqX5AHuXgJfA
b/JMTPxdC7Pb1MQ+3ncYpA2V/uWVBmkO7he5q1xW/Xqs2dIVwwlcmH4XXKI7BUYbDuWsB8uTcEnc
eo0SiQia0eLDNdtcCS4uqS7gmajwWb791MKPWnckOUynb645r77wNlKZsMAog7A2VWwkZXkrYD5o
uATwdTonezcb9lTne8uCpQg7vDRh+8WMXBWvElLtwDViNooMl45wCM5uP5OKa5MLCfGsnzzdrq8f
a0EaKOcEoE2yLooYLcH0zwm3K+OSoXLiy1w6AwPZFukVpVbge37JVEppOdevAmhMCiw5fy0P5MoB
pU2/HiU/8F8Sm+K18Yj+mxtN8K0pyveUt6NEJnHQ/RyyeIQa/IOEvwPWhru3B6x4nHzKSQwmYTuf
5qXndSWyS0zCW2+qocSvtLiOdNHxtyTnJt54oUwIH7RcnI73XuNiLmMBJlQr19Ci2lKF6NunHQVY
wr7RdB0vyctEXP+6nrZuxSMeP7EwKxSIAUlMCMUGOaQlQ4tYMteLO0Bqml0nBmLCieV+eOqMkoxJ
uUFUiJpHoBCK5bHuf/tNZv8Crx5LJc+FBa81A7CuFTdRdEyTJ1zPTm0RzPS76uvndN3wCq4xEYOd
W/9oOSzNQDYI4qFUMxmIwoyE3thnFGfVAO+47oZZ6cDDhth48nLI0MmJ3RLqirCuAg8Z34XzLbPO
tGnDlJRPvEblPv9Il5zYu4fAEkW2dUJEDOQqjg1c1FqoBm0pDrJ8d9mt78xxBBc/bAnxllfcMZkT
D83QYlWIHDwjfYt6vU281v6PLPEz8GuPaaqieI5dNHVvO+XDK+Aq248dyV5qV48yW8xW1qeU1Tyc
0mqHcAhfZkqxNfCMja5ifuDR3a2czWmmwAqrqE40h7iGsv5nbWV6kSn9y3IAXm2XblQaignDrnEi
mf0zWOF7ceOLjPupEaVXGjio13gPaSwpk+d2BBmrU2rScnY4OJlfY3PIXvPg/ukh0GJ+zjPYxTPU
KLOV9WeVjWLivxgkLDhaQBD7QJXzvtx2f7Q3bxjib8rlu14JLP+Th6peFI9aVuEqdBcfbE935/ZB
uJnPdOq5XXYf9OKwLQhAg1aJyNZnv+1+MenCPTFkpf8hjnWAegpqQ54VbhTMCxe6m0KvJdcUyblv
+yoaD5wv8HDtEiiuB82a0YeMXVNNELzDDjHY+P2CcducnwkQKzcaaYm3X3MgOw9GSVC+ztv02Evo
/2WATp/ksCIesNa8829iTXxG0S5qWIShXndH1SOy8HDga46Xqpd7B5388ndpxQw7V0JJA7qdRD2+
reqxty1KaSbIa54VXhEV12s8TMt9L2w6diC7W1MRCxiMUtAolwbp8q2FP9aoYdw6fmuuzVohFqkF
ZxRgfcdkep3Azc5WTa83mCe9CUg3p7dGvzAqrL2+xhZA/wnqmyKo9ISEUtytv2zcoOuFjL4V7Tw1
yMcYAnLyirjFAVGrYiF9UiCJg4buoZgO0S0+u15WqHCGen2deZiHYfCGBzJDi7Mipf7rbvWS841+
gT4LAUm3fwgmqOY4ZmRh10s5ndW35Hcn7JHXP+/J7/QZq2o2xWDardcWAOhgCCJoFV9YPClvSvnC
EfbpJ4ss059ZARiHQ2m3L2mDNdSz5Xny342mk3aDBnDeTfhedmFa39jxgHlqCYdMSHy8JlkXorCR
x069eNUKOZWQ9mvsgnmsh+kCHt36TzEz+Id48fPxcM2QWDiH3HRYgodPAo2KnrRQucAw+Zn/MN8h
tq8pI3pF8fe8HCkOakzP+yYctaH3uHHer9a6EfgdK4GnEpX0tAxnK/AW8mwCSfNb0EcTdofQ4vOL
oj+bO1fPyf932rM0fSb0JVSFl8hVXQrjWOVhhX1hZmniKNDyUcu+a2H45wKv5/6ml8kjgQXP8mrN
2TjzitsZFL7RlQn08DXrxBjiIupl9FDEUPkYTullR+JLFNq47D/ird4VZe5VmgBO6sf0NwfiXVDI
8Negd0SoK+lDNKcTghTYwu+LJ6THxhDM4bOANX9hQos1WLMU+ipNt61IsaY9QBzuDaykRaq6OMwI
oSdCn2VNsCW3744Lng6lpc0tlNxO/oOwkpZ2sF1MKq+xJtwmloFL6N7BSiuoWLkstzVZ/uT2+qIA
UwF4bLhCm11koHE7HdStdzJ8cE+S83Cv0PFSZLM4wchBiXdD/eXNDh3+IYVuWJKnRadmAYEhkG77
ZOFjmQv7lxg9mMYUPBTCDtc4LQGHeVw737vfJ+oj+AMEbxc0jCU5RCAuD+FU+ai032W/cKRGBB7p
QL+AWSgLHpcymCDmyfAbtD99KjphqWJGvMAxEjE5QjFTIppnocreHGoJbPAftBCbttqRQQVheHYj
iv19BuFRaSj791lKnOkvRTJ2BSLvn6ZBpR0PT9cXcBT8hu/E3vXr/1nJy3loC/facOr3X7RH7qOS
adjIcHbcyfZbegzdgWKuyZsdXa7QGAKoHjpYhnMII0Le8r5C7K507i/FvDUiW/sb1X+UUHY5q9Gg
seAdr82VcpTJOijZd/0KIZyl/zj61E2l0u6jGHdpwJmUduT6Q+l4A14NgsJFXL2YhRzi96twihJE
cbBkBjjY80to0+7Gq/Z9Ngd+rxfFm0D3SaIxlgPWq5X6mIJ1p+qzJpSyAsC6jcib4iEmTOUxDV4D
91zJI9Ao016nBmZ4ueLe+tNmX1XKDNI1s2EAIQcIlqJKYopwy5B1sE9bZB6YE/M2E2a+s1xZV8dB
6bLfgA7FxASyoAW9VwVRJb57e0jezv2qPWpZPeXwtcHXTfknajtzmm6K9wG6afS/Kg87kBRAOY6a
bRYc0db6mVtakOP5uDiG8cq1EdevQDraUc57WSaOqV31w6FpyELiMjAj3bfKFUWR7vuNKr/IuejH
rBApBFHB1iBtJWbGY+mtAKfHdcN8HIv+7dPZ78ghR+jQzrPnETTv/z8ztN22W9ByEthwDJJ+JLh6
bSfp29aFFF9qprtGxVhfChpIQ3DLXLFSaqKbRqGzYfTfqC4GvlkQsBZ9QCBGgGgRmsSQwc/YfJKZ
sehn7KwOptQkxRoRrsSEJLkMeNMnkcZk93jfOzb9UHAX5aH6eaiy/CAz5ZgBPRfGmx15QYB64jB/
t/5D0yjrV3tH6wb5bfkQWl++BzvD9KqKrkAvL5bM08Ntv9NgOFEhkaDkpNewjfqBMIWN34JGi/UY
o5LKIcNyUT+D51y+CI8cNPzs1dQ4cv94PCR8vHujHd4C4JrsChofwBUEKdh7NAZx98ZyhpZntpBj
TS1jjvh/gLtaHk5hM3kJH3A/U0AFIm5hCYj7Yr6oOthsZcVGigTWikdS5FDShQYWxC1KQjk0gm/z
EkcfId16v7jth4lVLwwvtspJggYd/yJhVDC1uL4/COL1z0T4gqHY50Pk77xr2QJ1Ukuqf5ZS5aO2
mFm0RdSCdxlk6g3GSG8HEvtA7n5TYjWmVcYZWyb4xyKd3Pj7BT5bOIaPJx58mJg+TV2VX1ExsiBs
5MPoCCtu9CHYjxe4BpaM7ge99fcvdHTiZIxSSo8CbJuQ3RAkx6VnLGEBJ2OMoYKXkBGgr2YOZTQ6
5HdDcOMZOh1TnF590C5H/4VP/ueOHZUl+R91l76ZNfNMRAqMRjwsD8i98ND5UuLcLyJrjg4YRdtf
pXHwTzYVK4QdkDGW8YHL2mv0MsiEP/JR2TQX0Dj7WgNLmuExBhU+p1RRcTzeXTQ4QcJC0txFC4+x
i+xL+ZF1USEr00fqwIMlaeuEKJoemgrs79pVZ7ELCNpj8iBRwwO3SLV6tsxBhmbhauMz+at4x8AA
dpG9325QuG0dJy+BeK9uiZBJYosQ9fWw4wWgC3u3Gq0mD62tMvJU+aJ4hOA5f0j+7vGcNb+pVmxe
cCSppvmFnWchLhCeEYEwgfxQ74ZZxeQhLfu5hrx3PbHtM4ATCCGv9Qb8avbPvNqTrWeu1vY6UzSH
wnKI84L7D5elbNbGJbPN36Ekfb1kciOyQppU2BV0F4SXA2v9XG60vjpnibcIazeUZHbpg1nP+TqV
VnCZvOnTjFPbpXoKg8u91uFJANcNIlPg+ms9OfOV68bOkOF88//YYH8PPvFOnvvxxuIGZyzQfjBB
y3NnYu+2ifoJA3gHBp9qBnyANCVd7U+TUvasqjSv7fcZ1YCpFvmcouOxFZsXEP0oGUrehv0aXXgc
1sfW0c+HHfyGp6fYlLcPrBwHBeQrOeD+q/XxGPEFaGfwZHL1Qd318+u8PX5IEX4EpAbLGBWW6gHM
8QD2scuMvWf56Qx6ew7VjWD/IDscniVPrr7NghvLMNXj0ySlMj6C+MtvEJmg/Tk0YMcTWKW5bgpD
3JEN6Wc52M1a5nL2PWgR3PfEPlxmxmTmd0aO6BTAcmTU1xV9WHY+gK+CSfujEgDCIFK6RDu/yx8v
J870NSJGtxDNa76RqEXi+DIlplPeILmq6+0ZYs8pd00UFQEch21e9L3Z+DVEUD4gi/f/qPC9jxAn
4wR3vZahcr+EKM3tF2R+FiPYyZKfHsedo/+J6yPvj48lO3eVsIIeqE3YgvGi3jP4cZzKzIJ1HTwV
7ljksubD5snYMIz0qh8pJxfw9VH1onuIoTTWpdvX8Ew5Zjgl8TEvnlVIqP5GihglJZBCcNonTVhH
ECPFRc/gjhSglAh34hnFLMUQXtknxdrjR2LT6BnyfAe9p+Aog4XkHMf9WTkvdxcGOUZ6R7MmXBIJ
wwEPD2fPFcNLu9P25P09pRUTNLUfzAliYnXNlrrsoz0o9ETjIF2M7v4+zyDPuQG5J0yuaTeITslr
AifQ1ZaORUKX4j46rFqNolDOy5f0epTVLqZsrURljwGFiBytIhL9E/z6ZaRyi2NQhetNNmFDvIjm
HiRpuTjhq6jwVE3MznkNm7dx30Sqs69kh8Lf4pE13mw367Ug8JrLpJQ3K9/BiwbeW/13FaLiWKGt
jBxZK4oykt2cy8m4SrlwVu0dRB66aLvJriB75bjuIi/cNPdPbffFO+rK7tFPx3f9ynBIwtNgYTh/
Zn05qSk5W5YCqd7JGP1xXS0S5IZ+LE0OTFomiqpRwWPaBBk/M7ucbmb5iXQiA2J5KIuJXBOOcaic
V2SfzT9yS4Aqcwxi7VEz9GFHOt0c/Cwr/gCX18DuQWd2r2Fon+Pj4EGKbJGlHhF52TC9UK9JtgjP
vcSuq/7sFe1cvqFiqeiGye4nzasK8s+DrD1HWl47pqhl79+WrL3ktWpNsjbAA0/sz3douKjTCJ3/
+mUvhaV04TUWJyxMpPS0HsBOILeGGC4bo6RpFplpdxsRtAI4PWLklV16OWqMgIyiydwPY2g0NuYX
G4Sdm772nQoPUR0zTM49vSroP0ahAcE9eI+UXDhn8RRXWZBbTUWZn4SR44OD/RfvUm+SJX4NGGXS
h/9CCkYn5kyB9TtuptAP8ojGIWBA3gbGHTvn22IB5meTqykQPzDDOHSBcnkbRmGlE3JhfSdPKdw1
aY+XbyBUc/iyElNdSGxK6lQavDy+PrtXhjScxaqKx64XuQFTSrwQSj34RsWIBWsMHA/xC2Fki7YL
jOzFJP1AZsSM4uxxBX7Ek/QMqv1XNLFe1UnrDL9H0z18x28FDJanWHTvc9/yZhvrM/uEVaT1/cHo
sz6BFP13S+DKiTB1OxdJiEAeHXvJftmt35HRxmT8EqdqpF62sUkxEL+b9h/lIgIaZP5ZzWXjWFWA
Y4Fur0cfH1h1FcIZ+kXA/XTV92j0kJgtBv5BOUqOnIQzuZgi9PtpTKionzEFbhRnuS57XLnYz712
DhpC3DcFcEKJgrl+UM/0Oi1F2ATsWkSwStskpvJGdnwPlQuLZ83ml4oy6jHStV89g6nzYL4iGu9M
7cQAfarkX4fU91bevpzEMEP+N/g99RjVA1ZKSejP1nfhAaqyo2+LVYkQDxr4wqF/23XYNku4XvGW
qZgBvANOjzpCCzWaw5Pri+bkg7uuSRLyyYhh91KJe62fu00VQIrm6lquAfhsuSRffdjSGpK09tTi
MKshvx9bU6msgjT/BBXSFJMnzpwEtdzRnR9R4Wlqoi691VCNFYUeAPL1eD/kpAyxfHmcNc5zDsEQ
aw1SwQUF0wy4WzPcz2jccL04UpI7/Y/jy4UUHuGyuIsl7cF1191FA5ytYIWB0/iYqxLispWwqT8r
jyFHYih6DXhV4LWtAsIrOpEBlG069/wSotdFC6mnq3Y7v92cMgv/RQejCqmFDZkpvvCYx+G8+2xA
t0e/fqaKIvYbLIg6YN4GnbayGfrHHD+YKLcFgFZU1/ZWglvrKPqFL/4G5oML4kS3vAz8iOC1rrUH
5Ht24AygK5dCm5ni+LNbdQ65UxBxYxGruFYI54bQzdhWe5PGmrMhJY9KdvvCHKOAnfsemwo26umY
ArO9oYWm40+i5iCQ2/ZCXQ6cquf0Ji3PcHOGKcWovxbX4zsSBMCzATPbt0o9dGR7qKC//LWFOOOf
F5zGcwBl9AvznL3Bg+NmLsHjfqeRDVr0pgETbC2a8hTY6LIAGbA9uryCN45k6/aDduZnrn5QV24T
r/s94TEOqNzXIixbRU5fNUC7nKw7Ds/UiZlkdAwOK/GthhfCF4XpDSq1GemDv6TBsF9rq5FZfPb5
AN+Drfa66vO5HwCebQPqJVUGXEjQEooPHtwm+joHi3nrLMxcv5Rfzkw9gQSjNDrD6jJvOXfOVcW4
KPg45RE18/WLpH/IVR3mvRVpjmJLcJEL0igOuRCYO6XQcRsnj0MCPfxuVJ1eB2z17IvS5C482b5o
rpx7jIxAiV994roklDnsJJ+iZhFa2lztUiQC8jlN6xeLBsgEwvOIzzTV9yUhl6vmNe+fWCZXXD1E
wPbYN3G2qIhNQ7wMnoQyXz7iIoyH7wzw9U7Z7jt5F9UJroRyVQ28Wl9r2tKs6oxE0/rOBKUyTaB2
1hW6ZhZMGPS4pb/+Gvc6s+HUzBe79kzcvKC5nW+rTbaSwTJ+bAM3vO14/y0roeO+aeFsBSMN64kY
i5E0sbwzSMzv5HQny4qqI/akuRmR3O/WIHCA/OKJ5cgVwFa+xdIWWBfOTXS2ynobZLPs+pCKtqrA
1U7JfDpwX0XAtVWMlpg460PaXPcLIFG6rKadbSymjxNr8hSAY6GcuE6M68fMKJll+mjHAFbu4dBx
4Ty+dQgUjPNjfLzgNx69q+tk+BCG4wiMFpi9z08QuJBXTiRyBuZTRjBy5RaxrxFVBlDNW2AQSs+x
lsyXWI7Pap41msRqoN0BsgR8XmOUMo9FHR4hhUTXknt5W335ZIFY7nbTcgP44Ah8aJWzASwspXIB
zreMVRKGAzNzAeNQnzDz6ZrwjoTXN8leNeBKU/vJ7+RT9ZoH2Y+Tf18Fy1Gd+ETxtIp7FPtUgznv
KKH4ie0L0h4xry6dK99UpkiPr3l63JZzS+SZLAKr+VLFsB4SdZzRa60VDhQkYXdjiEpJRQdKfB6X
PdsPTlzh8kaGCvVM4lC9wnYLDe2WtX3wdD58BN7/oX2i9wZ4JfYHU96n5HqBOZFnfaUNRoBNoNF2
Qz2/sWfoFtonWNarVU2rye2RZOqCGPauNrye9s6JsTowLyUgpsr08A8Df5wu2DBJvhnr2+6VECOK
JLgjVTQIuD1bKBkkxEf/SY9MqJKZRyWONtWQ3cGg9vRjmpDpIB3dte+UYAerZdNrOSXbMFHy8JxF
Na69YOfiXUJ3lDuSvzQjGHKM/EeHKUZoWs20Fd2hHfw39AoMh1vDPbCSgRJ+a+YUm3uUtLttKFo4
b8S0DHWB3kTTScdqz79QdmSCzontCQDJD2tm62wecQVEVgR491bK25tGW+zcKe/LK/A6GZLeke9m
OyhOFAetEi3bImMxUlu93ECjKD4QTbV20TuLQ28Xog1o8oF//ENl8xOJJF4GmVRZayCEuXsGy29w
FtwhdE3QkgRjrf6HjnCyPgNIw3WB/4YyMrEUpkU7J5l0c7ypbu5/vaF2FlxlVd0YL/KAA9C0Qt/f
C4fe5uYwpD5x96jrw7jN7avBGL8fQu+UY15age0HyfO2Hhu7OJt0wtjHvmRq1Xty3/8jWSUdvOOZ
Pf2pbDGgrPY3BhuA4QQFwg2bKNgNFQ1vaMSA2WsUNeOSkkopXqU6DCvU6VCDuDp4IGURWftsoEFq
KyfoeO8EKEEyJzRfcgxWKfUMwPjn/yuI3twb0Bt6DpaQfUXG+APVtnd2diCnChLgSMsqqt/kGEhd
we1prXb9hxEKqHU56bC+AoRfNr+Gpy/lonp1K3LVRe8x7HxrajJurOY9LFbmuZ16UTV5gaCIv0/H
s82YB4SycX+LbIgyGw4VoN76hdURBd7zuwTIlR6T//Z4iX2b3pvegF3HbXyo2rbeU3PMQNUYg58g
C/2eVubKxrLgbilEiuKACCHvY5oz38vWGWgTjgVBy86C0Gh9Ie5md4Bla9j9enVOGbi2m+ZoNvm7
FE53csqG61bmaY9CuJrqok2NmOM2IK56Uac8AfEpZWnFVrWVmoQC3zSqd3hvo4o0oHrO/ocijrY8
J7l68wOg8wL+1jYMuvSpgCCHcgYW/04W9wedtoYRFhgFeiYPL/LfAIQ2nledqEfEpHgQMHFve5pU
aX8nMtexIVmQ11TtkNP8HTVJylg29aJ7r4ZmKkrOnVfSOhVQAhISbckYPh6ceOoExcdlU/+okxIN
nB3XtFCEvHGHpJqk06cHUjjxQalopeokkW3QDvKkTrTwNGkDx6sIy8Wa/InK3IjN+5s8hdwmKv8z
blHaPyIDvgb7Zw+kfg2LCjbON8dR6bm6SupXvch4fixhafNmAegzZrEpfz6yr8wOHIsXC1z5Tv5V
CS9JxjUngmfJTX9BQwoMLw4NyJUXt40Cd98jsRcNBaAvx+jLkAvxC3MqUBDlX29h08tHCjRVYEsN
cMNjbsU6CkPOGPJmhcII9I1E0yeXxcDMWb+nBNrVNJ6a2SaagITM9S8noi/Mh11+b62UG6TH6UZ8
XYBz0rG58vxhshnyyYoswvOGWBeJkiN1mlEcdk6FWpJMNzIi5LQiVMA0j3FgdvYYJpD6nB4Wo9v8
FvKj20mmNCatNoy/3ruC2BzQydKjKOTK/2kRpaNvuvUdxiAfedNw5s7rfN0ojTDtY1fVO/A4ilZ4
85ax3lLH/1N4iPnXy9sai8b5+tfrHT3N/zCWscwaadWq+KvhMegJQKpp++cJ3ZLpz1iYi5L2uXQV
qLW+DT1WQC6OLoZIHuc5SkaUnZ0IP0gKaWz9KyOzYLNjMmGFV6qntGR7kMtzNOCnylE6og1kqFFE
MSycsXKHf0EsfQi9KxUkWS6lAOAUWhnlXVC4RmxiCe4bdlCDzcH5ONIPmhxhb2zh9mJ/HTZT3cCq
IeS/GI+2GygXy5vjmSS4L4MMRsXGJXzE91ALwJtpAHEIVKrzr3TinbZh0Y8JR9szEnSZSBnv+qej
HrbhKdZevHV/UFadfIZHZHUysV6Q0PPd1eJDJJhAAQ0cFktDgKmhIe4gDznwZHLfqYIyOf8smzZT
wk0yHZzZ2FdcWe+uS6T27P61tSeMoRGNnFKSvypgTsN7u4+58y4maajbPmjiz3BPQUXixpKUd59G
tafZeAlEq/M7HTudwtd8Y0CBRQpqxU9gffmosYf21xvX1xRsjyhPWTqCzjjidreLnaQe5JSRdkJD
0dVRM2owXLWlsJOVXDYh83tzi7BeAmFfG6OOdi+t0dO+Do3z6Lbb/jkicCbs+Jdv2nX5MvFM/UU3
kVyPNJWT1tCd4oSXJMuJQ1hZR5nXFZAcb5KYW/r76a8apKS7Wak1mERmlXKe6LkUhfowRHBTgNHa
BThBEdTJtJdd59mp3wWqCIK0Uw+PEDlZtEpbPoIE/bKHH9IgY5Vcn4I1ET/7xlVg4XPXOKTIfpCL
9lFwLYGDQBjwo1ncjlIZ6prlP+P2V279rKsGGvWaAvuT4SzeN1KbDxVzyL9DAK+Fb3jqoaWdk+HG
u5WCQ/IFvguHjzJm2dmrWZZaMQ/JYIqZkQFGhyX67nj1b2SNmYRAjqvMB24votMxxOVEJD1praXt
e8yZh7q/ywk5TBPPmWoioXmoZ5Dt9od0Z/7O2omHDbJeTZ1uPIBsOevhjt+eONmZaiITybIefsh9
ncGqiZCK8u3MXxtOmL7N8qEPNnTb5H4l3PwSHuhkCrSX6D+p2cFOGNVr9VDRCgqfWtT/D1bsZybU
eIGac2ftmeoaaFIBnlefYLc8c5aXQe6ytjKIAXfB/emT/cbjRtT6KFUSrBNZNDvWhRL1rJOT28Li
Sd1c8+/NvbiGR5MjbhbG39KNlluIimpUAXTNc4D7r4wTsCp4JuSiCaeH/e6Ck7ZFtIPMk5y36bVr
m6u0ujWzM2eeZ3ChA2w5bOm3dfegAsL4ZsNpbTKgWErLOu4yiq3PMsmTi8wGgGYSk2zRpY1JbhCU
vIUQmRQbZdcqznHach9kQJlDX6fU3DYMe3Bdms2lfzuxpQHuwAkm/Qlowo8Jn9fC6Xx/wAeKDxxu
22oyxg2uoOw9y+RCAeaIjMILs4nTmT6Uh60q9OqXFl8Zjhv/rBudpkBpmTyv7CYTSnyPXDjJdtKW
+PZCoILuSZUvV+8M2JAZCOsSOZjCz9z2UZEo7vfK5gjfkIUFbiUypCfhjIl3ENRYzU/lezwrZiaU
ZqoGNQAoVE2LSZajSYc5Q4Kd2JtOhEGuxLgSNshgD6BuwdkQkKDt5AbpWtJFnZmaR3PSzb2znIKo
p/UoxGilRA+0Znk06U/3R5Mxj8WeKciN0NkUBApga+1mZrhGK2fi9DAUht+X9q1cYlHfZgenkkL5
l2g+PrUt0PGP3sMU9RQ3AOewpFyqyPW+pKIyakv5kILYtyAt0GTUs6cvwCiQyBMC2FCwigSfn/JP
qYQRCbMTBSg6ja0s3qVaXUpqKKku42zCyrXN9llI/JkyFIv8aWZq7MboP8mLKjjwes5ToB3KnNBx
L7G5FrE1zBk+HxhH4dM/fKS4h+IeLJMSZ5IgnSbfmzLcdhqIxkzVzmIiObIih9Y+quR/kWduHsvl
g3WWL0DEY5yMQGw1RxTb9CM9tscBY7gc8zCSeXsiEOZH3SRrDFBrTQ9HggdZqr6yrO4znwddvAdf
1H6KP6uh1Ih1x2ebTddxD6GOlR2for7ThYB9i2rwHPeHKNGo5N3QjRbgjrtMKyyEjEHBNxvUZsOQ
pEXfF2GltpKgX/ARtjmk0X+QlfFVnFT64KrHWGDOnsO0VSKq3X7tfAYh1rKANlJgwfe6vLk9DXt5
jKG9dFGzFeEcFBuatXsXqb8WJRxtEHxwEtTsxMbH+62HZh2cClAW5fGfFWVspJaxToqqR7QCoR6c
WKLHSLJTECK6vM0JgICXsWpt0uCCH/ZXuPJ+zqBzmLOtwulbYzAVnrdOrFTQZaSvcjGh3eHEvEnA
STD4TFgHpJ0GZgZGafd3pkhQNvlvlMyvGjtAmKAR09oqVwwn91Dqivr4CI2r00a8mu8ZppJPzNVD
5kR3tuyrl5A6vyoOFFLhktQs7NP8uzvb9f3mz9DYJ0sGibd2kfmaAhBlV5VsVJd0DPoJiQ821WPi
xnrvT0utegmKu3TDckEQbqbhSjmg8ryB+1gGKvctbTANV+GE/JjRksECDyPysO2y+SQJGbg/Pkn2
9DP9lLdXyFv7ALA0+BgIAxmNek6bZ0uw/rpLv6mO5f0DacQhDj/SBYdYv3TH/0nf8RNiXGNnh4zH
HbLC5oj2WTUmHEGRy01q7gpJksAGaqQ+UvqmjYj8HxVGhtbGeunMzYa9h35QiHhFyCNaVWfhXdpk
uXfk1Na6pVmnkPe9w1mwmw/+yx677uomwe692D2TUL6DfcgXG6VwI3oDdERwG9gjrQLW82/pt1Cy
VzNxEK4i0CKZK/aXyLstjpR9uQTLS1odDcFMSjNeTHs7sV6LHt9xhjFQOGsJmw8iMh0VZDVMvKVD
xZJ8TWUPMrbanQvR4KXaTNfrU/7QT6Bfnza4XRmniA3uI1HzIkDhHV9Dacyj2rHebjNjYejEiNBv
O5JOB0yVMWBtYmULKPMqBVSVAZHQIOrCYj+HBM/L3LWjXEWOAqr+nB55AxNYqRtU/SjzkUFIHG5t
7h3otN7BKMLhqcbChglvRR5LbeKOiH284mPDzeO7Wn43b283LkgrD6VkKs6qGJtjvB7YHy63pg1b
FB3VGCI40PNLDtfDGbfTbcC/9LhEMDTFp5Rg8VLZhOKrgNyEINAztAkLnSD8SATMuQiKtFadqqk0
A0AfzbhUMC2M5AXDJHJ6ZcE5pu94eZhUBU448/6nY8qX21LTuplCGCobM1ZNnWvMawM0z0VGVzLT
g+i7C3H/JXU4iqC6a42G3vK5Tn86tKX4ebKVp8SrDrA4HmhmNI37Cv7HWqMTdA+GjhvolqdQbVWv
nfehnfa5Ge5SkIIvatvKc0XBnQ35dVy+gTZ+PZT8eIj6CQcgw6gDk5yyJzLVPsuH1C+Rj99kM1li
a5TmpSrjM5w8beeQLD1hbIi6T95Q9tvMXoYlPtSpoUpEGvVK5DnPA35IEL05PqSEEn6WOa/IENAF
MgM84taBlcncJIwFDoe+8IsdGTNLKJLYU9QbTyKX/le2J37DfU5544fX/AK4funq0AN3JxVTktzk
mCxnwE9bTL+n/IphFRVzTocy+uQLiw2QROHjDWbCPKcQW9gVEh1N2VNVbCYrFiZbknmXI46B544n
ULF/Au5mYWOTn6NbkYswp+Z9TyJ2BxfDHxdlTX1s6ljlqCdh1gERkJB4zLIlOgDpCHPquJsTeyq+
wCXDJz9ScAVf/g7XtpeuPAx/whYqrvHwUtSdBfL5tY4atg6drci5EcOZDwLejm47PwhqtkEIQSO+
uuIUpossHKwslx47alz4hJoid7aj9JvIAqMa0V+IIjeaBbXrb0jm/AHmwCGtsrrmnbZ6npzYaWeb
0YcUtPy/vTGBBN9y1kDzzhHRRwwhv3ceCpE5SLHCQcGvZ2o0IZ3GLh/ayIHsq/A13T6OEJ4k2Dh9
623J4LffOLTILeNIc56B2GLWi/emuuwBEkDoRwdLifPaIfnezx6Kipm+RpCHAWdnaBLDR3gKgjfL
1xDiLCIHFFV4VTzEqKbP2sTwnutIjux/kdBrscEonOHjuLJgOQWDIIK3Jf4kstwe6r1ydu0TtEvq
9yugT/dpI/jr9Vai/DQaiJlyf+m6i6m3LtdPtBDWiSs4IDW2XnzVown5dqqgEhtoya+iaBGt3WbV
RKZZugDE46OlNhnr4QZDd+5dDcHyg3G/b88gk19VA9UsD5f+5PYzcczWZJ5OKhyV7bMHVbBAylUD
c2rCPmhKhZN9dn/mDacMBOvnOHQyYNprbX/PwjipvflvtsApllI4WfBm7RUz4S2uAPXweFp8DdCm
6W6coWfVXSdOT0eVpdz+SX1mVeAqEecQig9j9lfGK13P0ctFUSZIUcjgJivag3/bP5lziMttWT3z
YvRqXzay/1ZycDq35I0gUamziYfLJ9NfZZi9XRY6RVUv26gh0T7BEkAbDteZEMITpb7q1O93Q5Q/
wx1GGXEvW287plMrTHOgo651YdgQ/NMxDnZ5ibWvthAN+/YaEhDH2hTMRprtg62nftr//SACi8Ts
E7+GM0ahayTDCt8lpRbNmLfFY9yhDmSOUVsOgpyHGtqAo/yFhDE0/kCNkVpxoz8Zb7lUDKSgkZi8
KJ3rl3oUD1BCzAIIn9Sqi5bgZiQ+IlYfowdAhjmWy1e0wOgZuSj4A540+I5vnGjTROq1XPBAHYE5
eJGnK9EWZ5tFlPYuVl3CHUhZSTZYUm5s0rRiJ4sd7XLBm6hYz9M4ma36RP8WJDGN/NoJJJZcx/Yj
bgObsTWHC7kVRTr4jbUw6i6Hv/hJx+v2fHaXiTOGLBB15m11m3EN5gBtvPBpuDXugXVvfJ2RY0HS
dCrDjfGFqK6jDwitFBli6p50OKBaoVV/Vl4MOtS0U7Cg4IK2ao7Q/BdVEPLz683ls7S3oqG9kW70
md+j3JMgNZyVjK9pVRg9wYBRNzsMQjIk/5dvP+B9LbJrRunqVeqF9m/IN8xFPKd2tXRFqoL1Gp+4
ndns+fcbA/zlWvL7Dy8s7lOCmA+buz8WmaQ3WG0XTm57GO/qOC2rU34jUdo3UbyP/Ts4ZIy2Ga8w
dcs+OoeRoaw0FLAm+7MlalqlbcZgpL7CPsk7vIcLWjMbmBsYTYjwynsFGyMExV060d++Y/n98nVM
fZ4p5WATo3PoW+JoD8dBPdFrfkwgDadZPct7ndegA+yd/kZYmI4fgqrLZsPNELTHDa30TYq+UqFU
fnSJGiECgZiK44t2YHg2kyVVOcmzt7DEjpf8Tgf7QocHlkOHPjs/IFRMjZjgAmCNgl4iiRA51g3k
jhaR18T49w9VtLyR42kKwX04ULooevIdMjqLmwS7fFWJXzMh6AW5ENhzsW8brr5WqQOgCzNJ/j3I
1qDcJa9PhElzZ0xr+REYOl5H6AC9M87+4A66h0Y5Furwn8m/Rhk4FURUr4WGM6wFDPV9ggcV09LZ
rTbMyCyPiaIDUG9KEEnoVju3L71G+i3aO/s3r9LpBfaNeg4XmRzsolOgR0csW2nQ+6nRjmc3EqQV
LksioSpFmzRn1VkAUOJGaVxq14jIvbovgVoO5ZpEHrXCzWaeOE4O6Wnmi2dKlPXH0qye94i///JI
Hg0S5+fmGcsctaAOgSOlWUSyh37EeUzgEbSIDY5obWsptkDU7lGzS+TJ2t8bSVYUgI/ihaamNevt
PZswKeEDJ1g2MTXW7eVRDUD0yXifZJdTZCB95F2ex/Ad8XeEUyJyHT3mxS4ssm9hGiTObzhhRG8w
l8/IkOUiQFguWQZ31WR+lOEOjYuCkJDdQB6AoNBh9vMIurkENGmYUfW8nxccLmcLMKTUpwfPiyjS
BkHdvTtjMn3AjlH9/wkGtL5EF+wor+9LREFK4FteR880mPGB2Ze6QjsUBJYQZ5tbUxtfRohkWxGs
cyguHE6ZjLOQ6OjX+mIzgHEiVPXaDw3C7+MxTRNCy+MfHiMu6dZ4klcd+NtS3GjXul7VJ95zUPN3
B3zTspaTpSIPhmog0pUObht68LvaGm8My6yOQkGstr/Cg/fBkzalmA269cLoqL4CMq35342WsBXb
/5hvyeuDVlwDSI6EvJrUZwYAbV/nhj6WQeqRqB05QuMVgWB1xk4lkP+Ac6T3DiRNXGOX8CN3gezF
JwubCNqKNZ7NVLDTmEGEl5A7k2SkVyb00n1jPPRiWBYM4Ql9IDGtgFgqLKtLyu3I9dYcFmSgPd0n
A0880Xufd5v+wuguo2aXWDAsI+CDjeC2CPlxBoPCXy+0hXgXLI940rRfp5fv0XKzQBqb20mPJD55
89kufFDdXH7yLpZDyGL6swBIMszKMWdf3KXZKIvTrDBDnifcTgsou7NRp68OpOq+UdQUoX5wpvo2
awww/fCwVIVpJe5Kc1kzk1QBdkX3yMIneu1LsbCB/0BKejNxulI0lhReif0Pf2R4dpXrJK2n2Zre
6ttHIkiO92HfFCErz3O1v9+HpkB7GKfOyA2Vph60WfZD/eQvIuEmrb+FMWUHLLTxV4lgio+diKGB
+M83cVmx1dajCF1B9tH5jCq8UsKbyFOxswCfAEQGjP1ph4B16DUAeykpnWalvmmRCi5vNr+/ds5n
p+T2OzLtbOW7DipDUDD4pKJVnBL/SAeOGELv2TH9/Z46jS4x4lvC/5jq0JzRhJqcqRlOwSOdWuLF
sGKbB74Kik8Y0O4F4dASuK3XiVJ9gkzih28YAWYHW02TPKmIyY0QdD13/vguIH6L3ZZDyQokN5d9
W5EjKLtJQk/vBUTg4RWnzErxKQ16UruUuph3AxWQ2hILOd8Yhj0l96lV7sqDO5HrdGyacfIL44Ks
w/MY3qVJucj6A3VSIwPy3GLS/ooB3/YWW4joCGE2VuBSJkc3uQrp4xdaf4Fc5SDAI8laHw0WwoFy
1JwYl15QDxPmHgWtlt6BNrdKRAmAXIpjIzakIQhiNVboMNjAJDycmCEM4ZsU19ALTRSu3ja3lMyA
9yrQwx7wF11sKSDA8B0x5CdFpTJNi3iVAEWBPBRp/Tw/Sw+4amO3rhMdQO2wG0FUo5jz7VG/N5mh
D74BteK5H1/VO85ZsSG96KRW6trj+71qh3UmEDdvtfVL+49WWw3nfgWsBLZnsHQC2KVCCo3wLJTy
rsnaVNySACDj/0v+k9QZ8tYYHfH1H2mi6iht0fisPHuyi3moaFNNFqc01m9CFsVmiNd/yweMj0Mv
6vT9UQWFioKM8PCA5KjftPN5kO7GHDqJcia/pszEceVCzGiSa43ycJFtzPIYXHP7mZw4rE3BDOOE
TAi3y82wSs4y3/3+NdlcF+ylmmeUBfqwXVLOVObaq2oJ48/RGWmY8s3uZ7rAYADJ/FxFszkkjIOo
M2cDqThuWoFk+53u0ZalxTwb5CIJi9XivAXdEeQ7IAall/0W3FSOxzUv3rU90LMJDKj3Nf+TSQL7
urS16Aa88xcsj+fITPMJClvRRCmGwZvi2fYib/9qH1sww1E8Yn8Mn9FMzo8uwGYqttk5hcCTFz8P
l+WueTR+LJJaQ5bviAdyNjmSJIKiBCNyNHgjg0gd2SZVeQHl/SwK7TghuP/B6WRk8Uxpa4UcaFhA
NDHy16BtvSTWSBmKGfetjd7hzS6mqxKFJ8DWUDW7SgA0zwkPuyIM68+MM1t5nEaU6XgC2paZ0jok
rAmE0FETnFmP5wU+oOSu3K3keUX38jm6FLBBqNisHdQxdm8Jia3Rh5cozjsw8N3cCFh/gKWO9iq9
S7Rp9fOanQqcXrf0eCIeCXT8YVZv/8/jM6W4w4GUHysqj+3mqwYdoa95pP29j4HzN09YdGEbO2iT
exCOXwF4RpXq5Wz82XbU2dO8qTETKX58+TuvERyZvkWiKoHJS1+QSn5kfcr70P9fEkixTF197a9j
rkADbe4eRz5aSuQUJsgijRJSzSevSiHdkej0yL8dijt2ZZy1LVrA6Y4tHioUw7SNv4sX/gtCB7r1
SpMgsnDMsM9fJrbRhluLYN7EoRAAezhO+dwujVY1a65SNSS9PD0uLDMNtDp3uXuy1lC7kdxwRvNE
6qqFovs56b8hH87G22CKbpoA4a9NEU/WDC/TEyWu00LucTOPbq56CJ2XQzYSO/jW12uuJv7gdttt
4N8H3RNUZSQksTZgtZ5l4Wtv5uSPu9NlQY+/fGZHz9D9Du/AEakYNk/ZW3dAB34qSGGe1YXRPLmw
WfPZKg/YuMf62UDqtJM4CplYZ2KxI1R6scXHf5w6JgGkSard1VIut5ANvea45NlieeABq/tgII+X
lhEvGEquBHuasieh6Sdwup9Xf3DksNAZMJAjNHLxnSI0kOBipcaTdCwl0vLyE6q8VYw4cIurEtUX
Jr81RE3DeKec0WZS6C6eFditrY1k77kyCKyiVxEWwv6KTKMLrMx0bJHah1fRm8DIgtjNU/i5c1w4
fIynq0S3U3STwOa6NilCTLZmMp4cmB2UigdEeFvM5r8m9YPNgFOve/pRxfU7/waPJbvsR6u5gc/N
CumLRvKkstfP/GBS2EmK5xN85GlwXKkBrxmD1lNaAQjc6LBY0FDYKGLuqiBTVQYSnDLLE4gYtbel
HOU+Z1NHox23vIeqNqRpYUx8TEjjJp5beUva5wf3/YSjWMJfC0cTPGZmz0PIsg62kgy/WFma4/IR
/nMyBzXpu13r/+bmfq3C/JT3J5XEoTNHb8chCT0PNTNIWymojj3YjC3vTO6irO8uNT2t6uyM4/UK
tjShTDiwyiWFyiZ0ZYV/aB1iifJ2Fm7YAVNym8YEmHzg1eeGDwP2G77IuXNoY1LX4ENvr+Imij7V
mWD5SeQMZ9gQvS4pNXzvFSoXzmHksn07eRzmq9s7IvMLjuP1yomqdUgzaR3FbO+1qniGZuw5Kds8
lUc8AObwTItdz9ul7HzvEkIydE8ArjTUAj68CpSDd8fhy3fHPiLb7RQS3kpuAQdm1Yr4nUDoL8te
nHDD+byE/rLkHcofrO5gv6+zAhI5gSn1EtghjQHaVLA0Vd+U92N/4tAAQ1Dod0P22xRw74AwCwdA
9iyaat983DqrpdJ1zerHmVbGk5oDriNg7KhuZ1kinNJ8EQE3x5UsEZtSBJoGSHaaSGrl69j54vC6
xXqjl37HNhNjyT8ExasWcEWq1e6+QQNqJQAUWTrnMEQ7vq8fHj2u7aWx1qXMJD6w9XMKXkbpqSxd
3+oIjPCONGa2vNv4iN/e0VdrFZwqjVKQGN6lUGfLars9Hgn4qbA0eSeNLNKMtSIYJKIeO++BBstI
GRzdMlLM3weEqgUc36Ktn0MqmXDkFYEH/EL3OgJwi30NVU/e9OyqJ5WRdm1t7djApKxefMjM82uL
EUXNcDwzeDyZPSYY8QkRWOJuxibJF554K0SRvBEfbdTUVAtWM0aP/ZLIGATx9KshHCOBm9e0Ltvn
ytBPQ3fPm8A01jxDWE7oYoTEfH/ntFH/OBnYe8cGzGxUQbmxsAVSAgN+ZPvfh0UcEDDaKqVmE6VZ
4kBlx/hlofTzy437AosOU8XhaGrImPbtU8r8zIfQs/vcW9ZGREf1WsL7EX7riXkbZsyXF/2JND5V
aTHRqujc1xsYCj3ag14YUzoam2ZK8NQ5NW9ut94hiNdHBVj4hmriG0B8mJJwBh09KWiqWM5bmZ5g
5eBPRqarT0mPcZ4//2LmPmR8W60gtAh2i1LUv1M0AcdQhKANY1Cn7dtrZK0UsWtjdxKePudyN2zb
ZGacLCfMvHH0LC98GuWSTV3GQvS3IJ/bSCf2UFYcr7SL+5Zi9Ws4hLk8ttyWK3X13MkDHKK9gsmp
v09DdFnYp/Xlibsh8K4uHJB468q/BXvU3seHtXK6I97IjtZsYo9mOQiZxdKlLWZ3SpXYa3HmAZ8K
MllalzU8FBzgy+8qUYvIMdmzJqPKSCyC7PDQRDL9+bWCvIjxh7w1EBOZO2favg/IlV1RblKRzNyZ
KwD6gSV9kPsxQQebScaZWLVlBs5SDWJTNz9bRxC4OniF0d+29qeHA93CwOeBVk9/lCmDmYAuj+3Y
6HhkFgCEx+5SPBfBXCz8oUl+BWfVcaIKdD7aGDh5O3XzJhXSlneNZB9xGqJoin4sobsH8jCdLSFN
dqpzC4gAnUQuheWpAljYFI9b7mQ9PosL70in4xx7DrhEmY9bMqvmztDApa12+rzKCjoN/a9/SCB7
gCuWDRVDxBUytCdBq8O84ltTuP2hM2Gj0tOHeed07CB5aVDtgUAkwa4YYweC4I3Ltx2DbDPxMKdK
zr8jx/IA+V6uPIIKRICV4Cx4o+El4ck+MioMWj2y75RMh4FoJX63r1q2DuczJuXpYiPtb13Fovp7
+3yVmDLo22+7D0B6w1gnEwzqMVD3QfdxzO2yLIaTGJFu7yusvjfpJWAJ0/bY3wyR5msiwk7Y6MKj
NVuJKwIHQ+L2sfO7waaFQXWIZ3c4YG4H37IP3IXa8t9B8kbuIbQhb8bnPDK3Wm4snJf69XypkvlV
sPHLOyAFTs6859UkjlwDNfGajC3vJtvVsCq5fYh/njATna02YkUHRVj7m2aCKfp0Y0K2HARvZRDW
OCIa6FnjjucnEQXP/Hzos6nB4wJHwbvdadVbZcurMDtPI6OoUXg58VToyPvtNsq387LkZ1ygLFVG
SlovFAm9kM2Z5A6m7XHvyG4o8j89NQjNvK0nMTdC8Z2v485BxHUXz2+ueQU3uRfTbrwoC/3ZdMPF
adWcsHEEZZwSJ6Sed4U/LKv4pzs//3Q5Rh3rrLDUtXt8yPM2ket4xsirz6zkyoHN1Ygk69/WWWWG
ZtF4mTEEUCg8iC2qKC9+Sr0+xrkmhUsOwZ+onJBq1iYTvgG9MPUYRinlPgU5aW/Sry8QDyShpk7A
UssJ0z5rvXuE4gRSxnJt2t/JUiHsFIcd9oJ59Y76HJfRghSNUDDOW/ynGKuy7PfFZh2rxfo5xbon
xvZx2BDCAZAYRAiZfTGPWJlgZUC1umw3DmFDDSZgFPNWVBUkM+bkJMo/eP2SJai6t8L8RHP9boRk
koOgs3foGS6Xoqvx/OqSSt+YDotAp4t96WLpuIpnDNLcvLzfg/SD7QlvFqe62KeCX66U+BG6Q/1m
VYgUtNGlfeXmmVmidQSccAcmVjwZrHAEVeDwufWwEvRGW5SEojoAoUDzKSHSs4IP1h8JagtHovH4
ccy0t55xS2NJVcJeGpRXfnA9AcSMB5Qq/mdyYwRwJ/2Px7IiLGZxhS7Kl1fxnSTnzwawLhnCeJ6a
kRC/D0QHejsQo1yt0GPpSTLHbpvRq/mLvWZOJD4u1+sMhX+p63RpZz8GW8VLy+/Lr9KWoA1Dj/H4
FmhmJGXB2x4HanNm8RPuUYZW8lQsMJf0g0xWzcJGjr+AmCK3KPkJ2sHIWf7ncKcT8+22rgHBUN5R
+taiTaLUUJykk4OATJUVfe4P/QQHmv9Q7FH79bltpBv6GgsE6LCHtwa/48A/tSiHRCRoZxCI2yLv
9JlfEN79mDee0f74KRBAr3HW8mhErGVNPfrDVHnfRoSQACSmjTkgabLWd3ELkjXupb7PSOCGsPSO
oVazxh4SwsnRZqhFnpAwDCUgUF57Q8bP9APuvMgy4/otHaOzBcl4AzuCUv44ARfjjfBT4HrblRGY
8r11qgUBw/IBfhgrMvzYRd4JoOVUspTNjfjOw+fjMkFDsJ+HaaEqaLcFnGkl8Z4wQwJh+wJQpxJ0
YfHBRRANxIbBiUgAXrtsHg1yFaQK9jXTcsvXMzesHYfLWr2GqburXySIswK6XRjoakct+LhEPwP6
lT1067sncucOIBJO36oFX+V0pYOR9dhLaBU6SJhI0ow80XYFxBAjQSpXwxivC2BYRwVPeSSorKGR
JG7pA7GkO7+zjHFnCdbHluWT3y5yBzL/24Kt1l91194TiHnuomrCsF3CVdfD5eqe0E8EMjj+Mlse
hYHFehT/9PGtTnT4xac0cjgJKXONH7YywF8cLj6zabv2LCII0wTRtYfs6qRYy9zWy50Z5nIby3oY
zzLRXHeTEGX37aJ4nWZ+O3Mbra0KSMKcW1jvhENeoEGu3uN/s1tcmU602hmvlQgVDbnIJpS2aatx
0+2RUBcozY72HN7/PTYHlJhQpZos/HPtfEg7rdiwRFqGuClFpgF5a5LcY/U2pYa411/1JzHKIX9M
q5synd4tdnxh4aTUzjW69cPO8EzpD1I/F+G1qzv97KRdYiuNvvqfQTGhDShLusbh7lv511MG/k9W
hJz5o1iXJb5l7jnMbaEsF/H5q/4E3lfvWhaf/UzI3NsMeOD1h1MFZZIWz0qhri0Ra4J080pVFJlm
mDZJ6GcpFcA59hfJ+gLyl2vqFDZmKvdjg5HZ+hPVmrCLvF0b06UMBH0dxoWMNzguHWMykIDTPK0H
XhI54Aws3gQtEWXBkKz7lUwx9Ak4S03alVl/PhXoSLdvqgK2lSIC9S5lJ/nVMExDpK9uCHr9GeC1
OQwsfdJWf0Gw2UYgIjg1D5l2ZipJcTT5eQK95fsRrntuM1KQ1z3EDSlM4lNh7AKg0Iz7OwjAJRDL
4qpNedCwuvtd/LGx9nEqipmRS5TgE89L1TTUmxJj0hkD2kkxR1V560f09iZ2wEFYOsZ//FpewmXl
CAey13hFTdUht+IAq2e3fXv9BBzgS85Z3Ov17heDajDggKe9lTDCTBDwb0N2r9nQHxfkGc5q/qwo
nR2415xgeRG2RXvXcFJfL4iDX4azwPkmDUbHU26Em/B4z0Rdt5UPKFX6pqlo/+I4tktOjwyb72g/
FYeBHTr5vxtH/6rhbUrM+XeS4xPWpprOyKh2lB/8RT9Hr5CmkROdDd+T8ja46nbbS3pPf5hM/IEl
4GzShM9mCEl3eSQTJmLPYyqJG6IPVCw+fCe64lTyBxvF62IL92/nrfv9ZsomyDevCt9NbtvwRm9j
pzmEgqSLDD2bQh4GxzCwQW7dFbbca+kQ0/585a3bzittnfdME8nTJvfWn5qzsAkXHdTEDi9uWn52
0x1WKusIZ8ElidnIXL+yhMsDeA+IwjAH3G7W0oWJvYM946SLW+wux+EuinvlhQErMRhUkkpM1pDU
3nCSdDHqaZ1UqM+jGZPLX755x6rrAtrOvxroKMAE492YQqzE9QRhL3kETQyNa+JQZtOB9hL9YjCN
qfacCKRAYCV8lsJSycXedBpqTZMUEaKtjyQO+Q82yA3rUMlt8CUu8qFDd0W5Gw/grAIwkRUp0E6z
9kMG6Nq7gZtOYWP/2cc0SzVySiD74O1a0qKwWDnI1H/gAKAz9PL3JPyAZZPVShj8juyk+vjiRT4m
yWeazfDQ1DR5HuwkSK9S+lHaCBAGor7lEHQySm4cDfOWakanGRgaRta6933rWpnSEfs8mzus25mt
T/ZBgzVIPnDVxX60BZtx5ie0KvjKJvJVnDQWvYGcEQWVXkuqoycZ/sFQFjzDCyGV4jBYH+dYXY7e
Q3ZVGFlHChjNJAaFw9nCGFaKgSs8UexCfvf1sSkrjW9+JsV52WXlmGlymdq2cHVhu+4dOStVEUpA
aK/sfkJh8CpbT9Od2N0fM+qJedbFKauxaccKGT1BsBGILFB2MAFXycJ4qcJ4CxIRxVJjPF2PkxAG
wtdo0mtrBlegJRp0lwgNoa/0YkBbmILpxYshOaUsHGFixV/rzlv1ZILAhRU9xXl3yt2KumK8wbPd
O8TNM/YS93T07xPmjbc8ICRHahkkfBP4D9D7v6iVW+I8NXT2yitASq+rTfdawn0GVRnWbTKXvXFy
guiibRekMMRaXxClzFUvaK7wbby+O4/dfCypSS62HQqyyO2i+Pu3cVi29228mjgCOzq9qZl5TMEy
LQ0nPkrQtqyoA9h2wfeoPE2Qn8rwwhDuAT1z5VOYroNWlXOTNnMoGsJflvtcpvDwCmIwvOoC8+Oz
QPslvNIta4mluVkqGoC1PpULRAiwFrjV24/BhSQLA7v9CGeEnG/ahnrk66upNR5YBQK3neGLyA2c
f88uMBj1avYvxIdNfPksfNCNilej7BqD17P0/lKEC3rNXKf+xBrYi1JaIaOy1mzsK/nSaiLXaWzN
CiD2HX7qq39+LprVoWb5jtCZ4CKpEjSDV6TDbFwJLfWGMpJQUhnImPMUHaX+93fXVwoefdwz8BRY
S6CgSz5PQWoRn0NL4iMtMGYI7SuUfrFYkL709PeWNC/KcHPSp5QT+BtNPGZRmHSzzWcCffo24/Lb
kyRfS6+AcgsRW/UjfGfgnq6NpwHL8xhzH137D2FsjxQNT5mC+4/IA7vOik2JhmpSfGs4qkH36WC7
Knibqyfs072SiG9V8VC+MH4MT7qwqNWmUHdz37EQrLKMBV8GgEHJyKBYGtsmUMo3cd/PDoTyGKyw
ZnvRddtmeXm/gbw5dyujwFtfWHuQm/5wMWhYFcIJWp4yIi3SmNmGFXcuyLM7FcccPwDd7TfFw7V1
QyjZBnayiEMZskMYF1yB+oUUDQG0UgwmJlHebt4wsO4naHMFoSAKzYNtTNuxeJaoFuayRmrosGo5
mhB3PsKHVgzsZnhw++rJ035AwIOBfdXFxest3+IRF67KptF+iYDFFoJAgzbvBj97hvK5uzHFFTqu
XlVzhhk/3wjW/pK7mMFEf8NRnnBykKCo1PKggGmUbNi0g55jUYURm36FWEN8oh3lZj/JZ4MlZNQv
q7VWTq0JtixbBj0GiK/dScVV6N8rqTtnWL1oQvcNUycAZbNglp4L8VhhLYrQgdN1CJLNqtfbkfgQ
mztKovekwX7ddSm5x9lpIZv+2yx5VYe1vi8ySZH8e3JO2OXA0LHOtYEMUYdXdw5Ln6PL6Qe82XrI
A7xwtJuChXIYe3U8JnA+nC6atwCeTU4O/0kIJxmpVP0Yhb4lrgvK6EVp/LpUvhfSc+lg/ybtsTol
aVRrHRj1NHC6A5jYjXcFEvKwMv4eHCMjfUxz59WuKsaee9xUds/Zt6yG0Wil7mRXAlYEhB55xcZY
77PCj2bPev7xFNwLVpVW5MNeAKvKbby8aRzp+7KhRaO3FNKDUyB/dcd20ytMSER4kH9r+ivyom7/
cDeCJCiLyUDBudN7ZWKj7jr35nLsfGQu3rddUSanYa5yn2VSP6PMYPUx5Jkizd92+4YhIX8TSF9J
hF+peNw3Wpo/g9HTOvOyrPZoYq+KwicJVr7/MmzuV5HTk+QnNIzAnqVIyKze9pM+oMjYVxmPedgA
V9278egY1u7drtobvPtpHUPEKm+qNws1imj1uFQucSTodlwiQElL4kmqiOkWbBWH5IMNZQx9diFt
NpJAE7Tvc6dtlvmLfqj7DGVe1ZyUmwMBp50uqgAfGchzUcCQRKXOA+Kt67MhbTaPxcXWacOwk4FK
ylC1m8vH2NfaAGzU6p0lYYI3GkkgRTigTsTTxmK3ELMniExp1LbOw8yasUnTIDmXeI9f9RJpH0rd
ot3pMk24tTN6FDoqZMPHjtjOxCz0mDHbikGHmlO/pFkBFY3xN62OCQ3C2fTtpnVj4Quu9IkZEZJr
kB9IikIDpJ9oMI04oTPDW3lKSHmp/2NA2lckp+/LclPOb9S5viC50fPaKsRKT2jfNafomiK1ykLZ
pB9CbzPiqIRysBu3bR0Ob8dqewCmFXbOXB2jD3RYoDWvvvrbJtThSNBn9QBc76NDOd+0tg7WOTgB
jVpPISZyV2TZravOU8Yo3Xy3WDuxd0wbL6iyKFOkcE9tI1nGt/70oJXOStFcGce+MLS6hNkHIU0E
EhW4JQLrIWN+LpAOGKtmMgDtw+RIb1emi7SfahRbSDNs3r3z/W1Ohy1lrEjRfX4HLDsXh0Da7rJi
kak5zXpSCfQTiuaqp/AVdL+m7qHKmw7hj2+sBLzn0hoo6vg4R6yclauxY2sP7a8f/irf2LUKebK/
TRtMcOIBbxH9fH/UeFxPF6rudwFO7yKYdXIoRbZv4ZLBE3LStVFv2C51wfNAYzqMfPCVgcP2LnXC
raYnFLTK7XEiVP44yeZQHsheleqsf4KvmQBFn2r3jufv+Q62DtCCVqgTMLwayomxh8lOFVW2x2+l
BZKw6Bv43OIpJyK0pCSI9IIMEZYNzYqgAORwn2Vp6nd8wjkJnn6x+91MM/xkp1lgrozEIKAVDj/o
k0AlMqBp4JZsOZf6WKpmwyHYWzjBrCk/y+Gj8Lytne3oclzNwn81CZSWMxJ+V4fUYW3p9Rv7QxS+
tbYQfnIC4aQqYFvpxyC1CM/L77IrR0349aLyTDnaypziAZLsDSXU5JlupiE1BbK9OhsvoIkgq4i9
YEP+C/2vC3ip7eFWa/JL5ap73vmHCkrg77AIGXtKzAP1Fbv58W6xMCYnFaFsN8IhNaBW+7WPsffb
Ntxg4gmeBC5xTWI+6JqtfTfrOGyhWCRUElZ1k5DPs+nCg4EBSthoWLJ8IInmdCb+Qn+3WM1hv/yF
8/KCjbcTfMTsMw7RPpCP2vS8YssShOBlOKwdyuPZeIdgn/2pR0b2W8PHlmImJ6ML+CYt6brSWdut
isKcLB3BWS8v6u04z2Do3F2x3IRS7/Yh3UEgfVl92tv34r+24WwNfpZYNskjwmmIM+sarG9vEmqY
a6Xvf1jeBaGSKey+Q0Y7IBVnYQtEjSkBA5JBopTLxUslMcEU0awdttfoS1E7x3wD+Azsle3USwQP
K2c0BcsP5FEdj731A1ttaD7IRHo1iioOEc7s2Wb3KXSuLy4p7OUIAD5GzeYAOvuqwN1o9zviH/cp
dlUfZbidIQ3xhNteQR6zvpTaZtQ9bPNHCngHxUxwaCLJMP29303TuNTwlvCPFJuXRQE0XXsR1SS4
Or/NchiOpXOvF3EX7HR5SBNOy/DBUGPyjs1H5G4kSuRg3egTRK7VJgA6a7uxDGsbEDlKu3isVzb5
mB/vAaKqHy5sBsJPhhegWW196VyjQw/7aKbB0nWaRsEljcDo63Lkym5U+QcHY0zDoyuHcWRQPeAy
GTxRxyAtdjGDX8wXi+q/Cvd2ULJ9ANiIImAbNZgbK4WGXBEW3tfStMQh/C5e8M06YpkUcdDGvM8O
6uWKJZixs1xLIAuL9C0xFbTX2sWNITsfZv8WlHOftJ/K8KeFMyHVViTNftmaywvHbcs8zmOYp5vh
7SlBrwZGIkFgIDeCjfISIRAA8CBUOWl7l30jN8iQhfl5yPZXaUkToWwZoXglN0XzqYto4oQwl7Qu
U+OssysDHBKKcaKwe2rsLcBX20+1Scz1tALXCWxx6G76WVHlgkBdVzHzyCayz86cEd59L9BcuZWc
ubQfeO5dCzC1Tsrwu3+UqMmgH/wZ+TU9TqDgVySzYWinIQi6Sr7MzUUoYiRXDN/x7bXJdzIddV1v
Ob5SqwENiFFsDXw6ZWiOn8LAjFFrsNnvKK5VjBFXkZLOskIdLfDUOiloq3LQsZYUWrB9dfjtNXpZ
6wErk+rzqx7IQ9JbrFTG8DjsWPFiNDe56u8Pqcukmgbnmg6xHnl0B6ior+SOFR6mxMQYzZWf99+Q
TIQKSKw6Xet9W4hpXlipDholqlhLHi2WF9Fc9C4Qsvg8fK6wcELiohfu+lPpYum76oiMV9NKrP5i
YTGS4dJl5aSe/8p/W+olqPX3UbPwJAlF99MsZY4Y5Cbho6fzlqqMnnJMVzw41XwZquqUgnJY/Rgq
ipwE72p3slEiGcaa2c+Dy5RmYSd4ivwEo19AW3Pds8s3ZXn9MO26eE95amhSVIStDGgE+g72zQ71
mqAHTEexyXj00NbH3DQz+8liPFY60zb8infyhSnSd/1nlQV/gqc9nmw4aftaQ2ET8NX1nvpU3Hxk
nnPCkt1TMTlgIRp9hlVaLq+cnq62S5X5HjnIMimR+IyESjJ/et3vwMH/Qu9KMIsgwsgBUQPDsvdT
G4zfNgUlJ6zmZOtgBjaOFGmgEeT011zfLYcR+wKOeQR4jL1eH7ii0grmsI/yUnkk1nCzab3+UopI
bQrUyRZClTrbtpMk9gEOUA9B365fBJKGsMa9cRzRpZsB4cho23dKWZv7rSpo3YsGGMfhYwy32z5h
6uYl8FMguBJDYD59ZbIai1TKdmJ9qU8Vin3gbaWzUt0TrHpyq9NL+hkqNV2kCz7aAB3/YtSsdqC2
lE0Uo2mPfN37Jlw6a9VzjFBDGgz1D43Vdu9CRCwQGAqlv9DIJDrapaCszltinjoTKCs8Ij+zXe8Y
nneifRoK6naQY9be7nyYVBrsSN2Icdt98ZR43Ckwj00im+zelGRBt5Px5OrnNHWki0Q6wEbkfLAK
2YGEcSmki1PvD7WNv0DgyV//JTSqUsXsiwi/iZAMOEka13K0NoEX6nDwICNxc1twWL2B9jJMjVyD
kM/MgD3KvdTbQdhkGNprR4lGQ88SOMOjey/178q2vLV8sfFQTf9IQ3sJNAfTYQv+fi+2VzfpB6uN
W+yqX0WHZHMK8fEBS0cgVyAjA3O+H+NxWUlmvYsS/J467gkJR6ciijFtEN6QYRznxwbtL/i/1mOX
f8EO0meHeYQi3ez0vFk/1a+lTB/abhg963iH/gYjBSoiLzzx4rgBZmZkXc+G1iiDLwT4PM8Z8LiY
DFPNsV0NhQdiayh/XRRXJCMfC0inodKnxTMqdsn4UZD9vcBnA90KQs1U10Gi3+q8YsQi64H8adoE
7bP6tNa2+a5hNbUAUzCMz1vgnRBlk1EtLFrq2NBYjGLK+cGXB1Mr24crpwqP8tdtMh0rCex0fMeh
jWDSzr1qMiRNAkhDCCXf6FR7Mar+7RJ+8haOSnHSS6pjZ3cvDIRzuG3eF7jHQWungv6ixjZXq56h
Zfn00L3zU2r493PmwVF/9E+eRo+1+sHSHYqgr1u3mRixHIfigcuFIu5qLMF6+3K60iNYXNpvUOq4
RzkQgdDUexvjiJfb/I3eGNoQnmTdM017URtwZzlBKlDAYbp7JaboIQDZStETca64oU5oZDanruVs
WflJumGTVSro7TgmlYfjvEdxZnbRfvVCI8LlFoYsR6mP/MHK2YTSg2Ydovk89RwyU5tjY7B9JYN5
z/dXtKbFdTYfL+RoSG3W00NivzWqlKh/hFKZ3E14L77wQtS+RL6fpk14xAvwVQ6zILK90DhcxVZu
Wm4E7IKwysLMGhMh/suA94B/c/GD59en8uayCFxLMsRcbTHGZtRi/NIOhfhKgnRf/sDgpZ1/Zddl
nfM6/GPJwGA1Gbk2aIQvHN8sPX25hdxHrVwz7RA6AzDcJI5O+yG0O9eFCxRUfOCvkd5tp2wH2HtC
4Ql0EKkgJN0tCOk5zPc1PesDuWJL5Xuu5w9ERzbviKD7FU3eWU6uM3JibQzLk65c0GNri5/9b5Qc
8mC+pGI31kEKKm/lFIr28XE1wGNLz00hEHz7ZlPDmkK8PWb+SietIenZxEIoBgzuie2eL3l+AEJs
NDZ23DwovPKTDgHvl6s+wdPUxLt/E7+3+Q13lFMtR4dr/c7iSRV/c4PAD3RVyL3IFtL9aJJ9fkIH
yoUeQ2fOTIDPsQH5weOgHRSHyl32aPSjqSQ9PDoB4w/wIAGNr71xJiyi9jZlMcRNgbSKV39DLliY
B4JLH4dmh/R/TY/e3ZbS4UXP8LO6UsERMqdqXc30s1Emt1Zn9IV6qbdcwWitpCEgHCl2aF4P2UiM
t481GVsGkH7tCXDfS6qwxyadTSyrut8hfl+MxMZN7Q7ug3afHz1Ls/hNzzVm/KOJI/2egpHuv85s
3bXGVm4CTRrc8pdLxD6CQzR4UfT/L8wZ71k28xTMTthiBygdnt0mkWVNruU1XrM2Rf1XG5ttq2Is
BsW6YJLlM32I3gtrvc04NnxyqhSAt255jZSP4rsht6EVsy01WtsjUKNFIxc8Gc5Uc0EjJ3dEQl33
TIdPCG1AvzsPB5Or0Wt7rvaSuWfzdgOLgEAGztScS2SbqkNOOe+LYRlcLco+YRc0bH7S/iu+C27t
Ovhz9XjRJtfQiCHeza0DAAFaQA6GofxCh2iAcnjTmPGtoUz50ZpMWKx3BPx0rgVoSbEqIkCB2Ab5
xQI1QqfjZ/jmA63Gh0EpYkKXyXybkFQrtnikOdisf0SJEc+9Uz0OPOkE/L1/pDEe7OtCkd7lGUbc
cK5SC37rj/IUjVsIPCJS3BIYH9rzcOgeqU5dLLWjzQOGwLA08RGfIsTH28LgBACAL472woUMe/dx
iOQjM6Tb8SOdxmxheWH6uruEoJReGXcKqW5qN6kqFwxpn+Z2ZnxoWxfB2eZJv/E4ceOoPp+Qbd0M
l/QpIvEutD868bVZqKl4iEHsIDE5RLgJfmb5oo5yjquu6SR7ovyHjZ9AEd1xH0IFl0guAfX3A8jD
XbyC9QaWFbETvdXY3eidlJsuUyoBFIgbriWFl7ywh4ITeWnft2s6aoWtUhX6Fa9xc8RolZFSqmsC
3wred8VVJwGn0tTFY30rO0uIFSNSgRqEcTLD7p2wIYCgYFL2jW5GV5hE7BbEexQmzSrjEl1NaBy5
wtfOa/Sch+PYE6Kk0C/arMWpLeHlKNDpJsHJLYVrzR+UZ6fMdBJxW9R9DQ9Na1TOPmufPgQffrc4
4BExz6rtMGcpDJh+UsmsuAnEB3ukyoxVd78nea96caYipmRvf9Zk4J06P0EWfxi1VqGk89qt4ydg
TJk0oZo95PL1Tksx2oei7Vi1jsvpR0dP2H/JmlvzflDsicXQmJaKKV6b2mCcKfe1xj99WlrIGocs
vpQJWqZ4r646Gnxl/PZiPIiVkpKzHl9sdb0j+mvQxwwVqqt7EbHVyaLL7iSH2QO0wzUSHMUyLvzB
RmAqB0GHyarbyeTEERJy8JGnmuJn9XNOpQ+juPozVxrl//Eb65DS2YdhqVQhA5ZPiBrH2eVwF6XJ
LF+FgC0mC1N/Qc2JYDbPLqkKFd0C/GuajWPbhi4aQcEJNmMIa468no4wsGMlnw+sP0eR+UYeeJXs
zrlFqDDKpcSioby6Ev1cREaF/TptF+nWJT279wev2A6gpdZ9GKvCSUUQGCazZ2MjrfWN4o19/3O+
vBFp+CQDGyv1xKHyJc8h3XwKTtS96lL6JpF96lA22LQVXyfa4+AAGtfFDLXbAV7JkGHIVW3qb2nn
4WVe0/JnjIpvUacZiiu8E7LQQaDnePJ+fz1pQpoE6JCFjgMx3bu8abOhk8VlOvvzjIUhbNqKqTqt
TVeX8vGnLmfpCTj9OStWcezwY4muHHS7bmExL1uq7FUz2hCbduOrelmweQ0N+iDQkmKVyxK0nIBe
VAViFc5e8/trQgw2FTVRRwI6VF8yK7vTIUG/QsL1QcGzMh+dEENGlWCnc9TcscHQqv6hyVydb76M
ejaEUNrPbOgM0vOZJvz3W2acrd+zSyoFAzquEClb7UYni5JGpPZsBZEUgShajdP4HxdPhU46+IGj
jU9Q6WmaWqvDLDdDeS55SeteVnS/nJQGucFSNgp1NpquiX0V676O9o7h/E9kJa8Pcaw5Pcd2LZIc
5jyyp1jXmFdb/tKzLPDPDmNuzGdPpDvYIwpIBGWsxxOYYKUTg5Cme8eP+10dyM/XKwHU458ZyzLI
IboBAxAduqSQuSQTL8ECfE2lTt4t193xFrpfjBXb/J2ZBOfb+vQXiP55vw3xSnQ4r0GbIrb3b6AM
rMEO2rGUQEys+pPo5d7X4D2NUUCYL7iMEpkfY5erF78bQxFn9cWA5eKblVEHihpaOKWyOPzpB5mh
yF2PqgP1gPBEMMGPj20wdUID/cWEjAIqs8ViTWhUqKNjdojnUrvYvDn3AZmxzj0g7FjfUPHjtzPx
vk/5nNSuib2N+1D7e7M4H/9nHjQzMxKO94opfP84M9LYKcilxxVwQoEK5E9/slQRNAFNkOFbM2KN
jhgnNhVdGWDVA9jWvT3xBNiy7zY0+1JQ56X6Lw24FkHupKg4v/hYJxM2/RKs07OomoDnjuYHzaIT
P4RlXwg8xJPst1J2vytPxP+T9DLVBhxfGRnaRyDX95YIEUmvn5uJzwOaQFPtIojZzWM/mdWa/9fv
lJWNCg/nAbZ+KuXaGM1R84DaVo1V981X4KI64jYevJMl18h8QbyqYEQCvRHnJqZRYxTCHlcInTzK
Lq2lbFK+HEuWadfr+Tr53fBLPqyDE3fC3Mf1DrmktmQIrgSFBPfuwE/V02WShDXTOJ1xz2V9NJ8M
uiNXIKhTVcvHJWeBOhEKfuQ8wFT3U45RaYKywWaP/dwJHLxeZneywZKxGMWQE9RUo2JjgM/BWCw2
LaOlzzhtn++LK9GodTJacBkMyI0vfeemcbLAqkqerfFIE2J1aHDnpipOGZngUQWif4GQbIuicjvC
gM0qOayOU0evPZ+5FFSP9tFVUS8PHgGWzNeJ0XrekOcG2INyvpGuQHylZdnnSde1GHmIkPl9gdnh
PgnVVq5totc6mgvA5iXfgqHL0insveSv5A2AihJoSnFX4OzfsUvP5yy/iC+uIk331/HRHIDro1nN
w+IfoCEuRUqu1109lmtdIXXaNJyS+SVFSw3XLJcqMUiamwraUKpmE+Yh2Js9YkKMHtVJ6o8wh6/p
2Y8CscHMiuVWN31g7xA7NQjmMtLqfDWvbU8u0J7Q4vS1aPI+Goi1QHcmnH/h68/0wmX1ZJaFE5bb
5cHi5hmnL+pUK8JZf4/2IfyxpIY4T1SJc3qNopm9HqypI2+pO+xFNY8csljCXuAj99PowpcAUzR4
qIetC55z4OiGZMbEyhvFdrRerRfet/MEjM73nX+k4qx919FvuB85gNHG8QsM1IXODajm9sgCYwFa
xfFuZAXyltHZjWEI0L4F7GpesgwZPCIBbzwEN42QsXCc7lqaMHHYg0v5hS9m8OB2Ng2ldt9n8SJG
pLHohdN+4KT4roRZcPUaMy/wT6cHiW5UHkg5wgw/pfXMxYafsTIReYJ61EIFyxroqkvDxMoXew7O
nNVVOQJas2Jd4g9JmBru6y/qv13hLXQOjd+NLLS+bGk82TegRZp8KFSx30UxO6KVQgC/6JsRoEKg
PkiNTCbdhMKXnL8ZBmN7OI7bPe5NykEDDVrdTig50ddNMYqU4YY4QA2r4Z3TRFiGfTHOTrW3KojU
1Fyr2+o+PvLwLPYtXN/lc5+l7IsmMZV5YOEOUSlwtmlYO8304KXFKj1IEylE1CD803jrjpxzWNru
caC72WPo4UeixW5GWO1WOvEkArN9oKXnOJ7y4TSkCVCahHXb9YqoupBJJ0MT7ZXASu/fWwpI5kSK
lNP14vYX6CnLwXaajO4HOW8iIEnH9sKgg5IMkXaOx49WKt/vPdblp4i2+/TfqzA9XI7aCipgPXQ5
/Dd4z4yQrbfnq6KGgAAJIi37sArSSAbbRmLCa0sskfuF2PrfcVZpcJ0RMt2EbQfOXn8Sxmwz8DVH
GoJcgFUOuUrN7oLpcVb8lAHsMVDFgsbBo9rVLzKllKdtHnjyAE3KLGos6YaOsmUNspIBOi1Z5EhC
3U5iVSgeOn1oovSMjGNUfj7GPcWwV9OD9BDZvDlpaIA6RzDuhu+LhEcA30IhmgoYhUvP6sGRQ8Mj
A0uZIT8DamB6up2vQDC/DTHP4wcZq3zhEwuxVBMI3mxsjrjZu9QbX4a0gXhprH9v+HF/bTt94IlI
fwtjSIl4vgaplUt3J1+N8C/36bYN/9SoOtGuREVXVA4hjSnkOTjWMOEk6WDs4xQSBiMzj5MrZjuL
hqCHH7GDnChw9K5i2xJr7Cjfwg3htllVKSnZVOj1zUGe2Rn9b7pjaAAqaSYIKQxr8YTrR9ViBbCt
vlgExK7OqxUOymp+932lBvSdHTV+KUcpX971hMyjstSAURqWchF95Fy1gZWeHQlaDTfgNAE+t+LQ
cUd2tFFzvnvnTZtL7oZT1WFmmFtAOtT7S5fUVssLuBPBiRDrQcE7uf7GvZ3W3R/ElVUAwbmBFx95
EleCCuHHFIR2Xlu00ypXusMGFXb/dddaQFN2T6L5FKLei1BYY/Sfe5TcbqC/cQlHGoBTdJc7SwsX
xS4v96RGsuMQalK7TGYV67pTQLxGhgP0aY1/WnNQ1IXTzQPXJrL2o/jk2GiLSxJooVjuFzNeSYRa
dPA6PS4LAjGSFluesvH9MZ864VO5oOYjhztX4xjGjxv3ks8DkJyQm+mqIhMOPXbMVh5MPCn+T9Rh
Gu+JDrGfTfEUo/yt13ZXhArucTN+Gb8iuaNgxB/frsnH4WNCTxBanLqEPRxDjfuDHb+WyCAY0Tb6
xD6/A+v3FOb/ZlSujUTv4j7gfgfzeaeWZp85wE+X2p6BkQu0W4o+vWQSOo2lBPyNfqjjf1MSv4D8
GqqAXGGQvec3fC07hbtMGxUSVOz3Tinc0+45vAc4opTMR+20dFVSaLZiO4wVUK8F++O6isMTlPPA
f0NiUkUyL4/Bte2GGTPh5vG2NBb4ZLU28AMIVXmcMcBybAmfmtRkLIKHmtvHLUbAjDWf3rB3STnx
kJajwZUQF0/cUr1P/EBDty6BfA6ovCkBvH/XfzZIFxuXhjvqZV5ETsigrpfLW5s3cXEqUV67jwKo
nU5BIxZYf4emUJi4WdZtKKMkMPVqoXyF6V039hLwqE52n50h0hcqXJOWZClXkbHS5dLcPFfkCy6f
/ir7ilHn/cRag9A6OBdojSsWDxei8m4mTwTMGuOj16yL6uWM5FDIgsWtc6t9uOK5FR5cNoKTleVJ
1YCzmuAEt3nFM8WEwiXn8zuQ9ZQe3Ozy0tCNhNmUyVcSOfrgZrvorA8MsTC1HwYxonoxKL3FrDUg
aOe/iF/s5Iam28GstCBcnYocKDivCnjl+DQSfa72mLj+cRIO+XnBFips1M2fh0qq5AbLBA3SlnZu
9+RlirmYJXGNKfCUpLQvKXRf+X0K0JOwrfYf06zP9BgSb3d34NhOwy6+/0KxbEyQSX0qdTGZfBDU
cooLYR3AoDyMMR4zWqYYGdzNakCK1HbP2OWQYszrFpK2nZ1A0jRtWSuTWgdzsq9zlSSJ75LOqGjs
tXnQN+yc5f/iqEY762bhqK6ESCYRu3M8KtCwB3rrhdpFykWw6qo9U24e8TdVTw7rhOvM3rUaOq3U
EcdpioIetvdYFuD6Wu7JiNdF2Zd70HQqg8FgrTnFehku6WEnj49NtLQ1vvIMFNQWWZJJvGSwZfrD
aaSc/g3B+8rMQpOBkTaupkS24OS2DT+hlP9zXhuqxNWAP8IHEHq5ROprEcM/WMRTMfyP9XwSMQvW
b28W/HSCP1uVVE34u9vn8M/EZV2KjTfMqSiOC4eHwrnug/wn51vw0ZayfCX4+ZaX+VSh60oHFdG1
31A+mdrf02xli4PiKquir6IsypKnqhismJGjDiXw4LiRj1beCOoYiDKNeetHqUJ8CoH/TSsZYFox
dBr4tMLKtdelLU9X7jJST+PXmtXCwI/8qSks8f9E3kOCsbfiPcC6gF1MB4dFcy5MJY1snWrcAG7h
O3Q3nokEVwCrfwo/Tg8t1TKFnfhf30w0TP0/Gaj7PF7X0iQ0y6xcDUBlwCHfpwLg2D3slNq+UOAg
ZlYCFbjNhOCUFiZ3ejg1eFYWFdWnsWvpbvzUoRx6vOCC7chIg402xZlCCEdG8/oXITqKv9TM+XkL
QXEqAXlBmK4LSYBvYt5cRSKkrwXRUrFAEnGkz1bpoMTkT4wVAfTgiPB07At2qz+xkbUGUIU63y2V
X8PkLizQr7/fyiiu2qy75sCMRtmwW56eatdedKjj1ukFbqFQHBxj5rzQU1rPN1cTUo49Elh07LC3
1Ushu0G2A7DgIUcgkSZONEbCpjwYY4l2ASxSLQHmLEu8Bv84oSgBVuJOryW6TUYD2EwirULebt6r
NrUNZbg1GiWePHEr96BqQ9JoFYnTGpjjguLHrEUZh0PHI0QnUidPC1skKuqHn0vFZgARrvsZXImL
ihaz5NNmAU9F2yTBkBExV/FThjsaoiT08hyJlUWMOXGDNwbsv78xdGCeLlbIvJ8lrCkFgnPjTdzp
U1STkPzgjvY9ML5gKC1je/UT71za8+NONhvmyj42z7nRn5uulvO73XFEYNmYgniigMABR9D3TYDp
pqGY+4w3rcUJEAo9xF1lWkrgStO7LRIxX6jS3OZYT63W+QGwEY7Kvl0Dt3wdAmPivWE0CllwUbY4
aE7pVa4U+acXl39CjThnhOHzBexInoGBXqZeI888yAw4SpvBo5fhlNoD/LotP9p5SkB9Dgr9OdBu
sYED8lXWcybrnd9Vnm3odY/VTtTlSEaOKjH7JTTAn20dMEeHTI+LYOcTxzYFWwQxofserVZC4wIa
nGWoiReDgVJ4pdsUwUmUxT7fGlIbe9IvzfFwtXxtQzpo6RCuHFf4lQovyuaBg0eOxXl7K0OkYwAr
aUk1tlaApKiAZm4JvYpXZLoks/ehWExEtCRH+ht1qGPgNFeB28KodTPR2a506ch4Mh1IxLM9PE25
+r0dcQfyZO8TFjzHkLPJEeDEH3gM4bFdfRqBpDfVSJ5KNeIxpLazwNWq9nyjAQ/oKOfr25cSZDti
XYz7YajuKHtPH0ledr+gfxEG44JoJZk/qCee8WDR20cw8N3IdheDtNPNFtZKvy6gE3KrVRYD11Uj
F6EDbGggQuGKLx7m5NLwIoMzHL+rJ6z0xcJqzWcrbTDhTUbv88PD6V3i4r4yUPZCuJfOutaOqldr
IlAEt1E3xhHh/nAqOhilu2djXFpAtNWRFXG9jFU4D3l1MiwvFtxmJnci2LvTJQeVd/oLlEyZRhx6
MnF2GC8ZQQ+X0hbNU/iro8VJTjw+M51OX3L3l7hPWbyKr+eDBMFK0FvbcJ35rHOTJJ7sRybxqxP7
0eSa1Gk+yj8P30obiDSh6I3qCqtxIhkfaUBoj/ppRUm3tNbc6Tn/bAQ6EqEtx1gRi2dvZtSEDLbc
OK/qx0ttu+9wl3WrWYppLKkBfmD0QiQVq516xGFxPxTphIp1v/2KYnhKrBdLyTRFqbXnmXM2ahuI
qZlp4p+7wVpwJhLNmWLJDc12l/N8ankM2S5SU11zIO07CUfeuZm518pwENIaN0RS9RURdpbKXTcf
Mf7+KZN9NuYwGRpv0wXeMu521KJ9lnNyFi72h91wMb4ti92/LRPrEUk7lkfN23rVIT0H2SbMHuRm
dmhplQGfmlmxFOf8MGHYZDkdqNx+MMOQ27S2fU8GzdHYfPA+6mSncPYgXVOFUptu2RxqKGPlD6jm
Ebp1TkiCvJbTZcUL18bi/xR/km3LIHWTr9VOdByQKzuEaxLmKJ6BkpDydOSqdSbNOXTjvYC6CXEG
G2MiPEfzhvlMR3B9ElOFvR0pufPjDYsmk34Lu2s/CqYQZnqRDO/lOI/sacanXGTMD4M32TL6HjvY
MkI/sueF/GFRRjruN31JZIGWh3FTr8L6mOgzy81RKyX7M+IwFpsCuxMBEXxDCSutHNdL5MVrhuuD
3Ea20MVeIVCZV4c1dvLs5uy6iA/MsgLD6Nx8mqwX4udhUBNBCQD2blLuPzaR5GxLptTu2AdnGju6
ClJNgxN4rQF4mplWDMejqen58crZeBFUMs/eHpXlQNH/1Tgo2frPl6jibWkyHG1OGDG13xsI65PM
DSUnsFYOfn6JQ4JM4IcTb7IBYTD0kaltrkkDGSAjZhajBkLS3cLbPa7eVYQFL9g9LAO4iVB85eZB
O+KzHl+hoaljVACBKHWEkvNAs79qbPxHN47+iDvq6Q7x1RHilUmvXpAOm4Fkh6gz15PRqonR2INk
dPIDMV67nBX7iPlvlwPw5YE4qvtuRGnYUHOPJFM2EzxcMQeLhnjyUztWZDMh/wJxgXQ5rVHg8F9J
1O4UCrwf+1NQTTzfm6U0JVmBaAWm8hZ1VDQH8wZdtU2byWy2aCulBGF+MjQNheRlmpOWarvrUxrZ
NtYDhEM/ITXSZW2r4wCqoTHQ8YfkOb086cyi8enWAr9F7ujve97hGykFkGAzWnw7lUJ20bmA29nq
2yeQmNlHZZho3decHF9aGlg25VKyqJtpjtu3D3jsxk1XpkFgNd2d2hchIwzj0f3YaARj8Nw6wOTn
sF8XkLkQ6VKrCZ4e8FudT3mbfQT7DU855O8sZ/agVyO98W29TxHQ3nhZKpIuaW2KingzlODeiMHB
xcY2w5Mk7d5eW7bc5SAtv87thtxviN+gJi8axMhMAyP6fOvsUTNreXn0/SfD/Z+don2J3rKjajtO
22V3jvcH01eGMQzbxTexXmrRR5nXBiGpVMjR1h5BlQBcfNnff+vjX7yien2TqZ+lFEKLVBQCfKz+
fOfNWCAcQc5lwTIv7P40aHupGKh4duofDttIn26Be94KeE6RWYWUjFsZNmO3XLCz4hfvJkSl7nfG
IyDFR8uLjbRrpJUaNcmoDDGL4ELh9tvbezQ/Y/Ys7QhFCDcz34skHjkXcRhlw+bmfYgEicv7zOnr
Qrs41Skkwq82ebj8foYY8iipNudjUw698olm7GywqI+ReZAzsJ2vLgfstWfQUMGTUnQCBvUlOR/N
wd1lZ2r18FFrTnUMkKknt2Ub8kQvsqCVeOL9a+BAtzTNKibN3o5/MXv8jAuKAIv15kaFazWcZ4bH
QcfYQBcbQpBEZjUvtgC7DGJUNreNmXoDB8sP6RmWz8lM8RS7zaTGOb+mh/6w4BiReY9GBZMBAIig
t2ev0HOGKAhkznBTy7hRPt7LC7SyDPl3pdBvHS2Jj1XQUUCnILCyGwpIjVH0kHYTv7MiEWtXsxl7
8he+lW4m9fnx3Atv16/R/X8UOz+spIHQB81qjiLv4rcrsrQOJf+23neupT4VRVZ59DkqyZTQxPQm
ilzGVLaokm5bcvvqG3LyuoamkEUJbMwJkjbYsjy/2FcthUWQbRPkLPSlNNc4BAMavyS1Szn7aCLI
6tteL8Na77u1NSp6SFmglORQFYeKJZv0reOC9vMmX3Gjc2Qa4lEvG2vpoXvs+pbR3Dku7kJuIX+j
o2o3YXh5rEpkkEzc5Izug0n+J6UZGaDF6NiS0ccCgXdkVW3w2ERjKT54EgHJL3Muq+R8VZ7rp3Xd
kfeC+1YQHdnbesYhXafwBM+/lu1m+WgvnIndtnFBjcesA2l/m1S19Iw/uANk7MIwLaulT8KeL1W8
JLq89jFL0ooCHQeX2m9lq2hTt28leT21+iKMfXuDjK09fmVZEBkgrf4dc43Zbh9jXUj8yaYZldaF
FSlM1C8Vw20vF0+jABgjpwwg/b2docE6TWvPVhnpzD2zBmessIApVZNT8ZWiCUG+qavMPkLvr7ya
ilapStGS7R46/Mt121ZdD1JINSVaZt1jBJ/Xd0M/n1f1H8/HmTNq3iBAY2CB8VgfThBdL6U3FkFS
/Bt1qvzeUnoTZtWyCSJwjCOmabPhep11C+GmimfgPObfbO7u/DSfw7Z5ngl+rydbePK56CTl/Ywa
Sk6xaEt1gDhLlcsVzCdn64nQqkXwvw+vnHFIO93HhGsQejG+qDGGkdy6Iib0rRifzn078AZVrVvQ
0E9/7crFD7uimRF/fucrSbuc0Oam/ujABdMBuZnF1sHaSsRlz4UegmutKOXZ8yoKpjT6MxXKbNis
8P+EJcLxis8K1+mwb5S4z0q/6Pm52TH3OG8lMI2o1H40iDUSc3awdBLFrMbIIYElSq6Wapgp7c5d
cXZcq0DiF7mjjACUpldba9kgkPec8MWP8x62zDqeMP7BTp0qee3YTQkuDfan08eL4aPrC8TnpFOM
l2G9nlT51uDZyd4sT0lKUZ+yFfjXHS7X1lKhZofaK2PckDFvtGiUh4Rxxi1jHdlx/+NBwmjEmWIi
jQoZI9VAVkvXaKGVh0DCatqtmwQQbo86+JkyQW7lDWUESYh2ITZopL+fsvLuo7jLvPq9CunsUHNL
I50Z31SziY7ZRx+UPo64S+k2CiaWYBaKCZ7spTjD6sbE5EgKf8mOm/t9T2SyiDUr2UySCZeb2g8W
KFDJ6V3uLOR/bzDlwQiNP0r/n6s2Qo94dJcK2msQzjd43YX0PhlVtKVqwrFDqf+bqj4Oa2xbR2Ru
EMLoRvusisuFYqE0anr8dSXsXwloash+s5oFwlFMaIDIFW5Gf38+2okF7tVMxT/QUIHN2Ulw/MXd
QBkRpkTv1KwWB7j3MzCYImP1tL0J+dSxQF25wgenzNOdck4mNvUjuYFkZEpaNWUhDAerVQ6ICe7b
VDkNuVKnAhtDFYVHR2l1+k5TOiOuTE4b7XPsUKSyUz1YvfXV1Mgo0F3T87t0d8IoM0r/MhLyr+TA
EZJtW7lDUaGu05/YXCSmgbQzv83X/haABRG1JerxvJ1uXb+r19i0Q86e/4QbirCWPPYYU7KmTBma
xCy9W0kbwPCoB/i2ntDB6blYhNOp+aWPAy/OZKYtCwB0SixXaYeb15oZNhIg9zz03Y3E4Fw8WRNA
8CgisZSNZ+tGXbYW+geB4fdaKNrPiPXzebfzy/heADms3PW6LTur6uzHCmFSmLpzWEXxUfDuDFHt
MnrCB7r0jYOXhRgALhpYb1xw7aFSaTYit2DLUnUC1JOJyNHfv+2fwi6U3bXFtbGbz7YCQUf1At8q
kmkKmoHduyvLUILLAJmnCuxcQnGlyHB833yIwbUh+f/0JsBN17InCKO/XXLd54v5wpyD/oZQhtqJ
v9Qc53Mm+FkdROjTS+kLYoRwNEy6RntK7JCmA32wV89Btq8R++F+DUyQIT9u5bHVX9i2/PeM4Dlr
mB6mDhxkyGZh7fdy0kC5B9feP2h/gC3d1PoP503MNqA/Il5zZY2y83w4JIw9vXslmq0B0XqGxknV
L4HGy8izwaC87W8s3G+Dw403z9+sYXHRBU/qfVeAC2LtR5lcCbxL+8259XCfp9zvuUBgJH0GbZk4
k0Y3HqZyGwbU8zN/kPu9aweFraWARno0GLurrVHCP0xug9REKw4R6wiaueFM+Iy3svPYmQZHKk8B
SegLX0YEQjYbUrBSfwSsERfZKH/zEtDjwIaOOCeFkHxzdjDVe5IrS5gO0jrzSr9Nwr4J1i+h/zAe
G6DbrIpWtWVsVSxRGtrUwbWWqU1rDpxpK6UHhHE6akWPKTg1ms8HAtxpjgBxBNJhNEkqO9IX5gS2
ho8qKuRGWDjncLI+CgOoojFBQnayfkt92N4EZoaYfaQ5MhJX+rfnSGT44dUn1SgHDuDA/iAgyCZu
fcece3kqE2V9/tL8bCA1mka0OcUwAVtrw3Nf8GCChk5XQZidOR4aJ+rKbWRZcAoU4SeH0VmPidfK
DRzmu3F0kAcy/H8nWHhfWucQHMKu/mP7sAK8KK3+np8ifyfT5OJgf/2oT2BIjHAGRv7xsb8Dlsut
Y+IvSdS6uJJ+/eSsCKR6/rj+/CNif7v0PBfmshzJPpzPi2r0mj/IaukonL9ArnsaAKR0FumC8yXA
nd3HP11qOZlza3hQ/S4Lzf+D5QqGwOeHIR6ibCgUUDeKxrJVZscOt+yFtXTax/OBuJuGC1RRFLps
Rfdy7eMm9OwJ2sERPihXQTTm+L34//BiNqNEzVeF50tB6APcb082RSSsrEqRpSRznoX35z4wrx+A
0HNG57x6l+EMjPA46nm112iQ4DEQbq3kGg+BtjmB/MAo1D4+ldE9ZAve1+HEVqSz9Pz63PM51opU
s0WFGns54oLWA1tDr1QunqryG++oApXfrU+KXrpl21Qk82ZH/EZTNCLdkZdXwrwQdvYmtW/1hHaP
l521efkO3Tkd9luA0t93Gip6dP4Nnp/BRh71faUWAiJPjLhIpzGHDkNrL1dRLFJ4d7tVbGY31tQ+
EU4tidAJPboR+fEHBu61gH25nEhtoQkv3d/+REtGPi6KBiJmOG616cMK5Qwy7gwim8WPBlpOfwhY
T1+f50dkSscFKssEeOBDefQHHihO6msxGtdZKTAPBOztY//U/mMLuH6YPFuopXWBmNWHRMZhMPfL
X9PPftjAcGJIm4O3MerSmY0OXG2rl2HkhKjc2S3ppVrsY3+GKcqp7kZ0CQfjnyyk1WFnBrNfoqNj
re0RDNEcFp55+amF/vKFDTOt1kE7W/OhHrCo4qi5rd9m4c8+NneczIwTU+RMJp27In1IMkpY2p9w
yMNjpmBovY69PnxClRNnmqIEdJEHzT74RiFCGtwaxkH9M/YhZyKlVfMBrYZ+c1cWeWm1tjl5oHQb
t0tpgZYZRGjegyLH/sgn+yuNh26vsdQ6M08xV4fg6T0SJL19PTxw2eKDH+sLKedezQyfBEXxZHlk
biIL6kbSvTy8H095RrFWKRs337XUbcCS2BHq4jBft40QEyUP6kxyXWH/aJ3cOaxi3ow2caRx0KaU
iJWsnyWNZEdWPlwBuST1YXtRAmaVQ4ZsUu32n6sLwKY6JnZH6A7pI5nfogm1OMF7nKfGoDdY3RTY
fnEamPumN6A/IGAakKVSoO3WzpDzCz2rHd/az22YjsFsDXuFOajW2ulkeVPrVHKQpafAMeJjs1bw
//y1MiC2U2/T6sugyWoLG4KHcX6WdkRGimlBCoksH/OoP8dnU32GB0WMcpFbip3i5QslnrX7DzbN
B+kcMU5NIWdCRgZr/7D8BWEdzOy5IO2Ce7jVuGBngSlId6ubVN1TVl9uAjVxGKjjlrYqgI/SQ/uA
Bi9P3haZQtSDxsysP6xxEVJx4ouxkvI8vTI4H+e8sDh7aghMDnVh0Lq6cJJiUXSxa+GcR3yKYGCa
CDnii7eQuHgPNzKtUVZfomLmGElG+EYy0KFMrrBw0zRz8c2E3vYSgZi+9aVAyj4v/Ij0iUERtLkp
LFetARKMz2e+JokpSYNHMhkZL5WjdFu2uwEgd5nhBUdgY1cia6P/ir2BCsFNVJaUA4f6MI6MTwek
G+IxfulrG7aKx5czQyKJfMbnWT6Nb8jZLm+6Vas4+NZC4UQqec87RSJDAwqJXEO4mWLy84I4G7X4
sgFO5VHaMXmRDR72TvDxuMzFPpWn0nSTcPnVnkDAIeMfJU9zrE+kd6o+XNcy4+q7B3rus/YfvH7N
5mCwHlKK187FcP1scJxj4q26DyJnpNInA/9zS+g9zZVyiNbqDVrhRPpc172qpsTFDz3WiVb1BAL6
tTYb9wtJCdVFA0SULSFT3+F+PyuBkA597fGnnQo+Ycums3HOLauv8qk4nudUpbbDrWUPjytlsNHP
3irHUKgicScFecog2qLHvsDJoMEd7S54k0/Ga+YbUfGYs2OwS+/0OG7ltfv4bKC3IX5jOUUCnXu/
vc9djHClMb49Z5+9d8tq3h6yt94S2JfrP0RyCXbPOBxQjkkMmqhEgC+pK3p+1K3lK+TSV78CCcSS
bsDpS878lZgOBS7M75XXL+ecGy2ZfByedz9YTCxgWtZl7W+356fJKDOXMX7FAfAIYoJ/gLAuXCBb
gkBWZt/Ume6qyHleunNXhcfsK/HMs3x4roTn40BHsIWFbw2NgUPRBUJx5oNVHUXoB6N6i9hYpq+f
bUcAbuIeT13SaEllNJv20VpRtKPgcmaPRUXweE9/MhJ6ybCsCHRjlhf+gZZW0g1V5WgLsgAOHt7F
lBAumb2LNn5r3FX0vx65weLQ3qWhHiyZmDqlXQ32vCzNng2H8rRzfYvnMvWNTJKyAMmRhPAQkBa2
yuFeerRjK9XIw34U6SyOfGAMumpgd3jWgUiHkzKIwKsKpI3zVMa3gw2NNnUmNOM2OoxVpEavvI9P
ClpQC+jmToTv5ZpPxK/LB+QvuxJliFKhknPYItpWtUG2OmquLnu3T6V/i+zqghNDKnB9qf1Q0zGP
+tEIie8+QXhxeeTTBspd+aEUMX1v9aHQNtn9h1dgMXesDwZRHlXIQYfD9wN9xRM3NhvUlSYAD7Yy
DUlIBSMqgfk4tZUtwJWWZPI88ReyyvLdp2hdpVRAqf/p/p3yDIeFbOPKeW8ekWRYo3w5M77zEs1p
eGmw8a/f/5xJ/jZPxTtc7Q/+C8y9w+Al1H2BiSQRvhCd1lMKcqsBF0aCiCFnGUgXne/htwJ2t0k0
F6q/Kj4dH5PeF9ocifnCXRHoTF/IsRwvJvVJoviiDyvT3oQx56M7BcgHwpglbb0DP0tvp9e0mnih
I+EWVpnaLXjGHO64V9aLcKOuUdWr9xAFB84fJ+MrjIZPHxjRxwlpEOLRhS7nlrRsJa4517tS8cJY
nHJ3fRyKDXbDkFtzKn+zPceI9Ga4JBhIxmASfUbebmowTXEqiRljyR26IkK4aCwPPvq7TbseUTki
s/lqHk724nkeTRhiHDz1Go/am+XWyCSiIVsgIB0zJM3u8Y8Qkp6+INdOqxFb5Xp0dH3vFGeN3tFt
t+MaG196uqYbrnrJ1BStjeRGRJ70Sn86lNMiqhvBA+paAjU47o25Rp8ONbyJNwyp498UCM4pjK+f
nHHfK0/8MoFMZ6QFYIKGaKq514he64LPqLcAYBxgv+XlwQHAq2HYmrCajUd3UZr8aOb1q0oT+NiF
EaEaUIKMazndbkHi99MHQIf9tQztqDbkQH1oSlqqHn6sWpNTxBqew5RHgUJRBtrGQ/FItke1S/+9
ViB2gDAO41aFETHCC4N/FFUFyVFHabOoMNDMPvOrplpe0G7sWKuPUGi6sVOgWWmfWXSR2A37eimh
XjPSsyyC/jWwoFPMNJ9tRMUy8hCxnAs0h/vGmtbHLjCTaZmSLN+PxyYLdIA0zcD6H4cbaeIgwdzv
6JKtqOtUKWMpp59JZEoiHg6Zei92XXXcSZh+BTPx5FrshEijb6MLYMThCkh2q5xtzpPgtlcfvdtX
7rT+4TGyR2f8y54oRUQbzCi6vIiS0g+Za64wiveXbe2lOu1P2GH66Pes2VRZk4MKMRbh7gbLdT4c
D2bglEnMReXZY6N/7iz7if0qfDfrRccJS63q+PkPl0m7hglQ2DTOC2GhLaqKcvm0kREKOAVTfS1U
fOdrbsxOnLDeZsGLuhYh75LCpqJ88w0sq/9UWJNp8A/S2qQ1eLyxYXFRgWxdFNhPcAbYsiLkWYfh
ogaTMTrlUl8SZCc3F8gVPI2K2cJBkdLx7oUH7OUkQB0uQ7WOqu9ouHf5TLFwEB0TGAS9zYkXtm5b
awwy74qP4Endns+Z+mrcpFrT/h9+U7WB99YGbAmAHXQShMP/kWxIXnrrP9V/DToQX/3LXgFmEF4F
RYK+2Ig08MGSEP1bdXAZKh45gZ00KNYpKvU/w3LsnFPpfgPwVezJvINXKy+b+JEOVyd1aPT+kVLP
3loUd1FpQUl5TlkTaFMD0qj9L1p5GKydOU7T7KyA3ZtE09PzSYRp6Xwz3OzT3ju9pwworhnWJZPK
8G8Om6LjaLPYYnrB+2pjUG1yFWhydoVEiIcJemKFkaKPFUy3QshnkyT3CyXwOA7Qt5WN/rFDCjir
px3bdJarBeyKxi/9l5nyYL8k2z+XgHn4OpxQadgyNocB1vP/QfugTCvFSXdflTTm/60z8u+gCHeF
w1AMDUNAk/clsIiTfdLYZYBEEv5fFJZU4Kmo8ljVSzjLlaowrEQbKld9w+lDaNOrtMz/m+dnfpn3
5YzGCTcGMrtrq8wNsfOdvz77xHmzqEnnltOoBv6zq/dxF8uoOqJtcfPOGbXLYMJIWItv0t0npBBV
9J+Y+gZ2UNhyljdez1yVXRIyXLesO6Tbyhr/WRdFeC1y/pJ6S7IHB0OXws6El2jeCrhbG8ma/jy4
Em9chu0aIvJgcZ3mDlZ/qnZYGKmaLAJIWHJ0vThav0hh0A92u2kG88mapwhDufzhgwtp+HtWTOI5
Ld4zuYAJP1w6DaA7vRP4D0vB3samwA56C5Fp+W+3CPNHUSH68/kTUuyMTwk/wGo3c9a4bBD9P9yt
YF6SyUGL6CIKXok/HKtQ/ZLb3UpPoEYv30LOYDBacs7pjYYZcVwJNMNBd4MNEk9++OOXe5mwSybZ
YX84WswNyy+zKJjc4+1gAD/ulkKCQMT6yKwEeEEStrgzUowy5cSfVR1g42sNaVyNMcjgKwUjHcn1
k3OMCMEBe6/0jny2WSCwJv49wRN7YkVcAYehdG8rZAr05yeERnJqo1fbRfUAcVlRZkueI+uVHFDF
egs6BKa2O4N8dMjsuMiyKCgT7ZLDn+PyJlkesbR9Gh9U2S779fo/I3raPwp/qtWY4EJB+xkmPWtW
KSzmsmlae8Ow3rXjboTiNFtyk1eohgQcncHb2y0ItcTL6k9OtttMN/fA+lyCfFqQfpSLIiRM7vY/
LAaUPVNYOHZ+O32Cyfty26wQgP+zuqDJF1IADpJ1c87ZR1L2glFX+7dXWWog9hIqnTViUJIv+PEM
wS+mAxWRWT12JjefBtQzWEvMa58hfHBQCT4Zfi2t/pfKor09USksVZKvynPyealvIGnHwiGhn1AQ
M/Aj5IjpgaHTAeg9hk/GUMoZ84yg1CQ+/7OSqun0CZ8Zp1almrKG22AfY+VNMjT9biByeVBLXiF7
e0DRn775i8v8lulEV6YZA+TKOl+5wys3Lf3D1eFzsCMwfDaougT9XjiBki1OjucgQ5EpS2gAHUSA
EGzfy6OXvCE+B/QBslprUvw9jEMhJSEsJxJT5REo9f4K7W70g+W4W4y/witzjpkFFv2csH8p3ZjC
mqjVYFu7nPjaXfb5BNjhmZOSNelM0X9XYXSVn9jrOSYV9FcApym5Bni6O2AOtjiRGUSfB18pFZuy
8qmeQOh9dMb3xgC2o0gNr4QHamC6GaxjjDlFdeM3giSuQEUFzN6MF9xWnaghIAMUq55P61VIcriy
3g9xHBuO4SyC9Qc2K2ROA1iH1ibVCNbbUXgyLOiCZBU8PlL+wh5ztrmN7OXeIfZZ5Dwp/KeLLXFS
vcQJqLVJiHmyOxKI+LaPLAhbPBiWUTzYqzgdqUIuSTwW7mx/9TZl9jVPIfqxWVzfRg4H9kMpRh00
eVAw8+STAyKfBURa0A1qa84XtmPI24bofyoHfmFetcVR6DRzZkiDNiCnr7uCXF0mMWWjnyfiGGg+
TG8aYh00SskH2Lwg9CZnLvTFL6JvdxSq7m+6Tcrcs0/qzbmbv3/PUyzru5oDP63hlAlDkobbS/sb
rNlmxLcZddJ8SlSRAz3cnoebuSSyJOfMXL8tc0h/udWUQU2xzji3wn2oHu1v9VOb27yAO1EiusCu
UhapF5yRg+nx5MBI8gEvEadMKJbXQtUe+81m5OfQoHP52LpBJ/VptCzFjwQ+pwuXCY9hPer3ArEU
T6m03KU8O5a1D2KRETtKUNZ57tkfX8/mxk2a/OWUUznu3jmjL2uGiKPy+9CrvJzQj7yyYk2RD40l
4raEBM1cYh/mv12IlH0NNk2AOTyBBvybMeAL3QztcVg81ealCmpImyrHvVWtfm18aErxSw8nRrDt
1joecMIT8oJQ8vD0KZn0g7r2CPqyM3rAiI8+23udA+y7vNIyUY36kNXvs7jfpwI5F+J8BIoZAQVe
gRosOpmk6/QWOlWhDnipYIcnQ/WrvZeLEQ2ej1gLSkrotBP6MP2thpgGy7/NguK+Ftfw4BEjRqn3
clrDPwZ7/OAVxMRk89GtJOtKlIolYxpsqettYx9zV0kqDWQyltqO1ZRDfPvR/qRFfnRZmEBCHGz+
mAyrjpUPgc34iZ1OUUit3eCeIoY+7vtJV/f85D9cn9h5iCAJUJScnpNfaekKPg0X+hoNFlQAHdjd
gjG27S1LZzsCZ9FygXu9URxt2DhmSR25kFU1hkLxU94urRis/sJXiVhdAXIP8Rh1mzQOoxBWmah+
5KSxiNdKEvkPzHJ+6r683TXFzkTQqnJYnSYQ3m1zq7GYQkjLvRV2QTmED80Sr1h0jkZQHDzLTLv8
jKqs+moU9VfocrYMZjcuGEcHoECJ1QWG8uhQeBC4KfJlWyTNzuMQHlum38/RMiSyCZ1EsX6QNxHz
hkexSOtUDcJ7dZfahj05RbjDgpKWsYeEnsMcvzidFo15EIb0/8Nyn/pVARbSMjOfRxiICMLsB6EN
xrlExTirTUjyi0pGZ7lEZW37zqNgsbDPAMW2oN7k/KLQ1sOdphzjP7vocvlUmwpigyw8A5+kzeR5
cmGzAsSyR8EORkKL0//IZ68J9rWc5ydYWUSNYjGyDqbHoVAXWx/MibO94BfK9Zsk+wAy9l9yPU3m
IETJ6CBXcVZJjOcBizKDJAGLiKeG6mxLbj5X/GyV390clCVtFjX3EEzc83a3/vcDtEnx6fyZQFe1
XsvQBcc+ePwJX6WYd8yXHo3Hy5/erlJSBlW0W0vLqltEc0szr+GyaCDIFrf6jiyxbGG+mAijpXTC
SMaWaSFHSt/I2mclUK0BQsmvKOADwzWOLVfFqZByL8dXzeKVWLGMp1I3EaJO2+nYxAha/YBizmlP
3KdYJNjW1WW4eOU2NsYvus/LE3m5Mkpt4GLZ98ixvTmHbgQVgNgyHSyR0VjKgi/k8JkhAWf+iToG
Tluz2ZX2dT6EuNn/02Z6UwZoXFJdx5p3wX7fvtbBK7AUK/BI38IBn76sYUB3DMhIV61NVfJwFb31
qIhck3OB7SDyQgbUB6I4U0epIBdYWS5EzchGOXg+YkQCEeBhoLu9WD8ENOVrLx5zWHjwgfmjIw/V
jLX68Il2IJu8tTxReJFLq4qONA+N9GWg2EfWxFsr7c4oIYq5ccNq4upqhluehSwxv/Gkod19UeBy
MpuYzBfFhcbkJtD/H4deNFbIxBVzTWQdWnJdnu8XW0vqWXPbpnjyIHcxNIOgU1UEzr2l6TGyG6O+
xEdMXLFYBCFiTi07gJoSoiu0TbdIaQrhWYTbApYRVjQfXnWvKdzwdH58FsEUEWskrswa6lf17+0d
UQdEetzdkbcP7T6LO8wg9zlqNp7J6uKyeF3yzyrrsjjD5f/oLCQlFlOUIjBlyKZzcm/DIKi4fqaO
QdnuOySnq0cza5OHVmGVLnx80eUmlkPxI/JxQhZszUANUSaEnyufgfY2olbkkezFirto5kTw4hX2
IRnaJrIcTwGF/ngjyPCX2t9YRtEpce+43rGc7rXPS6+tmcCV9FfGJZwmLrIkOv/J+veTJUeYwzXN
BonTdWFDrCcw+3MOPF27h3ozj+71zdr1H2YxG2O93Xtc+RydjPtKA2iuc6e86T3wc+Wpv1n10GjN
Jz9CinjrGWxMOJf6uVw1+i4ehlXIcaJBfs6pz40uCq5rqLG5smrrt6bYzVnibsfq73U/uWDKGk7d
ERd9nosEgAxlEvsNL6Ua5408QMBcpW+jICY/SHeumtPzc5DfZMehkGFon0y5xSXnLWMH1T1ltexA
bpXop5k6raoj3pN27CiB/q+9ufpftZqR/t8sN68G0izbyJJ4Us1PaXiQaMGbdbg8sd7C/0nChxbn
6PcPj/jZ3dkEJPMNG1YCH0/pRElNBamayGhn+omR4rY+TZmk1droQg22CA6qVRK0KB8dBH+bNXce
uZDld3s4gusPMZ9mwwhbepKkVKkd8gsXD2AUiAsOaaGdBUZtg1vagV5q8U8M6BIHhFqdXICk82Gy
wAhiy1bCSVNckZs7jMcFxtgqR3lFouHMcD9WxNdQk4DTO1SR7s9QOFCWh/+eAIYWjjVI8oe6uSnB
bwhCeoQamKFsf5N3R9I/yIGkWYp+Qfg9Zn2uWu0FfVAYEw/56IIgfFnwprEriBLmEPliAeg2gW+r
kpt28uJcqlZi9qPEY3mI1AVxiKMfBaHC4YNaqcaRvn36cA71QMnwy1mXetVBdjufLRjUhD6Lumqd
YkPTqs6IYjPGBpKSmTpWeo55myPXRaQiku1x2HCmEVM17YjuRCwDbvpUFbvJX5tWSvKxmebFYipy
Hue8CVQCD2jjckey9NmM7opZl+YtntopYX/9H6/4Q+dcnVQkkU9Fu8U8zzZgv3Cf1ciudMJm8fk2
lEatdVkP82upOy8iusH5/AjcgyBYym4mV9WbiWWGo6wA1PVZg0iBRSF063Ewtwmoo8aMq3trQCDm
VfwIUyrz6sQyJfXyZuM69Ma19BNGcTSL0N5sefpcPzZuzAd9Cuyl5wB35v7heoblHFiJK1iTGJKV
yiz96c6XsK9NgzIpZo2EpZeeImrZpCKLuv6RQ5SoDwgg4cHHamJp0JW2F0KniVTf9dm+t+z73rKo
Tz9K0zBhRWe84ekuASedY9FK6nys3Ol+mJxLenq2L4o5kv8ea1sCcox/SR+Q0ekubRsFtiH6mx2w
MNQr5bIAOJ5TF4zIvvbVKaec2OxbtqdHGnmr5nz0b1E294AuOnDzNsBYJhBLi8ownvN52+zyAR5J
sMA98RUUVUbq+YVaNXe9uporg0JdIg2Z//oJZBAlrPkbyonm1OZYCc56/+shn7QdgvqD3MWMkKuK
lfvjXUBYffrHLGgNY0IFJPA4dXMZ8NYzwmxnWIQUDL3DnCrwekxGtLNE/epj61/zWG9DSBCUPNJQ
jfsCAzKZYkLQmISKGTnCbpnU+dvY0BTRNQu+a4PwwvkSs+Nw7yPNkr6FMrm8MurEfkKpNPYkPOYR
OCZaxhY4cSF8WizdCsEM2TsLKS5dMaFIs24/rBDe7p7dp966B2yX9ktbam7YZOH6tPDcCcdDVeLd
z/Pt4OZF0wzGYmW6Cyi0PvQ8G0F7z5IEeUcWjPFGn+oiknBmzt5Ds705y/9bhKraPZhUTp1p8WKU
gzBIuALdgege65RGuO3Sfp10Ghx3JY7tEabJqgf6r5eDEtWgtfvGW2AYO2AveqJHYsEgJj5mBhCk
795lmpATKIGwiuu6RrBvaemLlqTL1m3Z0HeMz4mw+yruQtt4K/8a8Q5Ljsp0XIaJvGATIxwfkgCy
k+kKmApoZWCE28NKLhDdYDBLx/yJwjA5KVSTrusUEvppLPyw1ZOuT0Kh2VS0cGJK6kz1m5DXqE3r
J0CEu6wJbkDZ5DJyBviLR0MjCHPpIq6tzNVZCKCC+yJqY2D2h1e0zu7vlxnpwmtpcMbANcNgwwg/
JULHA6SuD21WhavnWDbTUmOFxmdd78sjJGrXNAk+N/i+uz7nEIaQMGTHEuSy+Eh85QgtDggFw+ee
oYrZxaKQCu4TrCntAyAbZRfxn5Fe4pUfvertB+QF6YmkS/hUxvCGKDJfR8MQDmtuqZICRB1/zA2p
3IT2dziXVX+g6wdHKtcfUeX0708yhZaiuahOcxuyGj2fp8MFOUvmoDFnnEIcISB4hv0cnFowarT9
5ymNOmN1XwzqKW/fcQeyugb4dQYvjPq/BQrFvpKNZVKzvaLUwTdmf4+LskH6tTtngIVSrcc2LCJ5
bJL3FDO0m1loVhzDsnnMmYHRndYCskTnAzJnb7SRwns1A7orPdjoU/O4LITWats3bbouLLnLbvHc
z1ohzTgX7Bfd5XBpjBZTV1NyXwHMJ+lWpvrFBZs+IhYTxfIe2pS0KzisDN4cB6H7Bjs2Ty+hag8J
GesZ7yseu/oktkdMOGmIzJMtqUWe2JEw5zT0IX54I8z/EVtN7G0KLhW/Gqt0cWuQ4CiCSttd0sv5
GP9QtDKd+AOV4dM5XsdXdS21ZkgX1zID2ZOoH+85kqByOP1UbOzqabWkpXpkA+fhBcavtCML1cBF
ij6S5FxrIwNaiu0eJ4cEUTzo9l4e3Ficir3/ID3/QpxzdkdGblcROsgDLoNtZ5dYoojAgYcaogkZ
1ZiPC9kCrQF2Cdia2XKj9kin7rJj01PYjpBZ3Bwt0EO+zSCt57gtz3jQteDY5axdqly5Z8DNHipa
OQmGwWX1lRArU9mxKC26lGYP4h052EdsUQ0GERqQxy1LLqxcv2/Ef1uQjoRM1OmpRJJ3zjCQ9q5F
DdvEgc9UdiyWWX3odhMeLud8ZinDVqZv2UqZ0Z52/I0AwEPmUwfKGqes7j9eflPDhIfL8meAtG8K
SgFOSHfJGBSFs2noqsCWPoJBttSFaVEusBWm3kjN5/UybKG5AShQI36DMfHOBua7myJOWSq02JdR
kbwwJGtQxjmbi8mby4kWJdnS4sLwooPFme8IESkaUzKJ+MRjJK8taXFWAGKaTEeSdecgn1iDo2ul
DT9TLnRCwkLPbg6J6aWp6dVhAeaccuelbcVDGBCrAWunDGwyJBIz4qFs4+vYKJ8dzrOSsNZKb4jj
uSYUgGpgKS7KwE1oTYrOQacuAciZuVHv/9rPIzJE2CbWO8FE6QtkAvdntMjHUvGEakbhQAyajG83
SKjEKdIjF2zwLV6JlJx7mGm0qcdEPaZZjcqSOiik2POmVHB3FYw9FRQ7om7z4gB+dLc+FsUIQDMY
lsYxuF0AoVOGE86g164xB+gpQJIcCXvM0BBdr1FykG4MeXk6QAVTt5zkke63fpb3SOfJgpe9YU5o
pB0FuzHTvt37tIu5KMHFn77e7T5k4WeG/6vzfUWjup9oICjbLoCVebHgqellHJT5cTFZrkN46xpR
XKs6FoxDPdfHxrIA+/vFNpxgGi5EPe+WoWVOk7oz736z9L8vlPgeCxfzJExkC+sc5DksMY20il2E
NFXxLkMV8ysCjniShaBWlq8sMRdqHBgjY+7VDe6a8t+wo9Y1/r5ExrYE7vYN6ugyD2kT5haufyA/
ISsbXi+oQAYkIsBulqK6HSJF9nji8W56gpUOLY66NsOkvfd/YWQFkPVvhFndYZP6D4YrYj0cGiae
+exCck2cOxlsdr9euqjCtCaa0msMaZJJUrrKif8b86eu0bygwzJOktdKxTOeaIWyz1PANT/dM4k8
ZhzWsffS7rPJ2QwCaf3AXUVTEuZY0TsOFpYt0ZakwMsehlbRzTUSw2Ldux2BIagPVCVluKRbmVnX
rJt+x7LWdoQbbUx34LRJOERBq5ST9ga6VAVlhhxitfRuMKGudnTJljdrwFdapQTMu1RtCRzDb70R
Cpl8hIRJF4nFKlU9BYvlFUO4Bm8e35FDeTai/o7oK5w21IgxAojl06rkP0dqS2fFm/tCtGayyBa6
M5tCYuDijpusF12pauffi/X8Tqh37YHbwNOHwsm9PydvAEgDEGkRIEYe1sTT/98IS7EaXwBTOa9O
l46VUzDyVIN2saUck/4W5LfASnJFAPJ6OED6yVjqLDzOFybeObLCqVIujg2r3bUOYqcmP+7PzneV
m6RfKSkhZmmO99lPPxpz+FfkQurb2BidpB2gNUO5U9zDU1jD7QWzacD7HtztxLptOCCSNORp2i6V
mehgOajxOKOm0tRqnWEJ5PVD1tXNAJxA3misIRgl1PvGBcJrCErQh4HQ1AQKZKwI7Bcc/hvGcdG+
OYVsxA8IypBihgCgsEK5pzgeC/IKjU2rfCZY1EaZe7OZzwKsb8pHOYyRa8U+bVObUooCMM04V+JE
mdymX+BxV4UE8l0XkFV21S8Fw0ybAQfYUvVYiHpInZwaTG5xXX+o0rFxRBVefzwBHe8eL8Kv/rxv
D7imdLowSQuxyck53YT8Go2Dq1q7B9cInx62D8jGnt6kMFAw72bmHnZrdvKM/SMABgsZpcCf1I8H
SZnGclxgJ6HSsEowQlMz8DyA5eAKNBgDmf7zkzlW4Pn9MNAzALwqsZ1TcnnI6WVe8GX4o4WIoemc
OrPd4aW2/Cps0fQM99aWPTmCjwqYtvSOkjy3W6tmSGr6CRQPB5Ua+JNBxYGr9HZUd1hruTxxcuIH
REqP/iQS9bQOon9EgOD+0Yzo3EMCsDE9hUR6vAR7ezskX3TEsXwvQHICaLTfBGA2Agi8UgoX9bXQ
MRU//wlNpYaH1O4dhtyZooOI6PxIf1kjw49ekNaPBSrlx/Gl+cfY5h0LRJcHJ3Q7eMF8jkjdxLMJ
gcpjgYzWWe8WFhRbvuWoDY7ZT0zBw1e4p3J40Np/E+LkAl6Q6Wq/97BBtlr+O4UUZBU8GVVpHDIN
wHqeOqN59ZQjktl9k58jNLlPyhuQROxvCrXNX0IXx6qKF5MjRJfo7ogtvqY6ynxxzWVqZajeJRwv
/5Pc+nq6+7qgUGTR2whKDbb5EFR21a2FcLQYoOUcPiW1Nkq6PIrz8z3RaIrkdF8bV0B7LxBfmPLR
pT6ahM8OsqV/LCs07ivVuhqYR7G1vX9On51SSNG4jSsgVpwnQzWltoQZzxpT5GgPLfEXruoSMFKq
ci0MS+6LBncsaI7XZ7xyMv4JW7evvdlFnxsGnwZosoE0ufMtFFD0V19UQ3eIuJNBpqdklgVPX7/5
ZxZysjYr3x/HFZ5tNyrmqA9HSK7E+PhuGXHOmP3se39oxEFdDnfWrm5DZOvM1lejUR0vEm0wz+dk
WFbXG3fEpI2b/poPH4d7SWhs1zJPdudk86ZmJIijDr8F/Nl3Vc+dfbvEGtIyx4xCNINpjHcfHHPX
N50j+mBnzyHhfvhzbV8y2beRIY/OBXU9piSqA9UuUn0sfTONvQjgZqA9DYTgU3FuBth+8lHWnAmf
FLKAnF+Tvq4lVAtRVrMMMJm7nS4JZvf6slPQauNw1rLcrddi2yaEiel4vhZmd8qFzFdrwSWBl8Di
cTlNK//wJgEtaNxjLC5u95P51ENs7/7F5U1R7WuVvavXD8FTUcCc/F3s357jHr7xf47NPyyvq5oR
bXLnscgbxtrH4BBL+O5D00Lu88Lkd4U5P9RqSzxF47HvXwynnmOunPw7mjHq0uKsDLD5ydvhK7OC
5vwMZW2fx51glaHw7MvLVPDm23sQGhyC6oEqVa6cb+Pa4lrUd48qJTQCbsQ3VJwlCe0gB1i4MHGj
6NAppnAUbFLsBEs070FJzHSOY15rOpQIYvCZwgot808BfLIue2+THtTIYmslM1Qb1GKgod9w3QU3
VYBAulhmc39dd4mBhCkF+JvMvp7+dmf7ZWQ/AxJbCCcK0DWcsZA4nyteo5NVSjrrt2HJfDFwm1Bw
FrqckQdXZNA7u3VAZS0DdpqRtzN0wgR6nNdLaf4nhqA43fzrlQSC39QUUSr+vdacB//PoEQt+H0y
cVpoz1OkYm8PlknfA/TRkO8Lsy6dww8MUzk2KpREHVVOsdr5JRako9h1QJewjX6ax52aAYLbArIM
AR3glv+spFXVomUB4CfH8ZMw+16lXX0tKu0EdIDYLPy/hR3zZgGtCcMlgsYWqkMI75qNZy7cZb6P
jvDnOBk+BrCnAFQlTUG7YUmgvucQYS3Mq7mIUwV6nN4ikunsLnfJVzKleaRxA15vjcDB+oEoJq6n
WP04I59zKKvt9gnVBlx4Hg1ycSesQSC03JnTr0b36BcEdBIk48PO9V3b4bXgCVDLqBlVEYE4rU63
02aozeZXg3KemmtVmmNtbTYvHGQAFWoaCWAF3KaFORGSOumxjvvkBlti2bsZf39vsUxx6/ct1Fqa
IvOhBNSG0ASkiPa6SVFeFv6EhG3TctcG57vletIVamIpgoBal+UqEhHZ852ownOrI71Qoek7ngX7
IbPTvSVCnPTBChtG7q09N6/pbQ6gEJ23oJYv38qJL3/UeZm6BjttaBP5+OC5z8hNGv74U6+wbYNK
Ttpjpc9net8rKWr9zzBx/bj3WTgootbCKDYQzUZiYf9jzoCAyAXEmDH1DW7uNDYTPKpK+rlkmi4q
gImr0Uriim8ZWb7nBjRFRPDnGqtkhgvVIqacCuOTI7QvPbh7xxYv/DWOuEDHYU3UotGKhcfpmkaO
nBe1D6tAy7KWYx01LzPvTjg9bsRuGrN18o73Xpk+cZgKeiQEymIMSp4YcLC1v69m9jNilfOU5OPO
DluMVIxGHtKj1i7+OR2KOAiQ2L0Mwpa/tH6/8ubVg5T3eqICRn85TZXO7vMxjtFb5yOOenWanrkg
rVRyIJSLBkupOvjvzONeXrS+2NFVARIJB9k1x9d5ip1RRUd7HXyYlThw23cQza57WqcL6JyJQxh4
KS8bgxM7MC3L/sHktkRk9rjPhSaA4saA17VZb3ozx/tOX2t7X81NCh5oJqWdxmPtUts8yGZt3XxU
FpelxLoqIG3lBCbGXI3o0pAvGsb2f34GDBhhaQNHy8je7Ks5Q+Eu0sfT4sKhcPEEWDGrcEtlCps4
T1vk6aEjS98bjP6/cih5lWYA/oUbpOUrX6n468Zgyv4nMeCyvQx7lX3AxH4qHumRlvhFBWEB7Yq5
tzgjTTDDD/Vq74k6puov3YXvSseK2jHhJkewub46FOlvWwX7YHHBkX7mAjw+vlEwHigQdkE9cxnb
p+iIa0oHH6xr6QG24VK+Iuvkx/tVXCt+AEkJt+SzOdv7UoYuXvKceLHAPtTeMpydi3ikBWEK24eE
Fsa1q0Ca/KAZCc6ThU0PoTVMNL+H63p8ALgOwfimZEK4k5AtQokwzk7QqsuFZRYl8UfwhQwx2V1i
fNqPIA3LO8mjt44OadOw68Y/02b1Q7T5KGa5pnTTdyVPGDgI8yf7hT14Lb3ihfWDSqOVifmNXIPU
FNX1IoK6u/Fx3uz2z74Mdu2iN2ZFk0R6xkemy4yv74nwYdI9WxSMbc1Bdt2/UwP3pPV+5M4YPyUj
97Lo+ShzVSjCfJGyMa5l0UaQDilEW7SvtU5OOIxqtE5dAkswF4PUWxsPUaeuBBhTa/gp0urR8Kda
J39MrDLpjyWjh3CGqk6Znns/VrnP004exaF3eqhZsMk5blX+JV5XHQvQaYZAJh0/dCnRDJoJqGAU
075jjYrFuXJs1mqAkp8blMI2s373J64NT3/zqNOLOLeeetuQT+qpgiARb6QiSzp2ZKgOx/x7pFM9
94i4f+Tg5968XnYyy2IQ1RTFWXEcPjzAKntq1Gr7TLpw3dYaEBmlrFdnWIwvNdE8Y+c7QXltIMDk
aLHmurvDpD/rhUOjtTEW0K66Q7XFhhjg2hggRBkt8eB6wroKzV5fzWE1dx+sce4IMOFr4VGOPOq6
espNtvJntB1dtwPT7y1Y9//zCzgeOMroHayRFSfFNW+Vu7V9iYD4Y33ZDLi2iXV+yI4+P3wdkoiR
EBTEIAPawYEO6rgQzMCu8wyWZB02Zgx036lqhDkZ/WQyGcNYYgcSFH0KTneIFDHlG5L3HCLYy+b7
LA4QePg9DArwLKM86+zsTzLAc4hHRPg4h7T+A2UoF1H7hTnIhr8jvnZSEnoo1WYbEFyuEGq5ldPN
qIl2eR5uLijVVnLbPnDlX3kJMoAy+YqvxAvgaRnwvmfPa1EMmk7lSI/ivj9+OLyebyQse27A1zrZ
IQmTbffPDSi7Yxkm72aQui5hAO8X3gacWwaHqB5sChY1ZVPbOg7/AKniSNnYYpK1uOMQqOwdFaxR
05gRGDbxWBEoboz3V+L07l+nUrCYDzx+Iw5lkVt03cpmLWGrchdY+bLbGlWvMYH3r+i4KelbItqA
5IQRsU8GpxzaBlCO77nsxud8huo63/fc5yWbPQFCIu/8OcsJGoKnNchLwmZ3hN3C6pPC9k5Hk60z
BiS1X8VAE0jv32EefFvqqnicISFixroxHMjpMlUjibx1k9JeaVGqcg8adUVJLTxCLKNjr2M0SUy2
FZmF+GNaKLf17uo84TIpGDOpBR9fRQHK/JiK5eItlwFxNjzf8KIkNgD4aZFz9J+44cfqgBRo6lnE
DPL4QAfsZyVEcg0E+bMeMV4U4atrDvjaj0fMQrbqRNHsr9WcFxsojse7pfCIeYfyS4I8kcwE83NC
EoC2Tf8uWEw2sR7mSmw3VELgyrGzYByJE/Kg3A/IvypFPkLhnMvc/CXpyzmsP6NrDu6MttrJv2M6
gongTXY0ludNw7SD/5fsdl5eKKs0eLidiTJV4NbTGoC3BC5osyRDuR2VTrTX2l0ITZZtODPY/kNB
QHJeCl/2yBc26CF0HbygYU3c7XxzZuo88zP8f3u4bc5z4tSG12cjjkPKE4OF58/zBcLkNprPtd6D
TBJOiVCan6+wxKFvnnxbR2vSFeRluFvo0of690BLmkO1/SCyU4bK1XEcgk4LFepW1PEZdrgg+tRu
qoDtsbpHcWtrxmh9WtFk07JuWmfskMWfmCpAZA2FycFI5garMhKjqJoCJaiudTgrJPxoOliyC8HK
PFzB1LjLMFNFMA47UGrfVayrTg2UE9Q62cO02mqNRFKiMQxaTSZbjV6s5O6+F/FKrIe7eY75IMYP
eim3zQAwN4C9oLtEMtuUhqwnM1XesYdF0pCX91HMYSL4jG0Kv/pOsvb/1yGRBjSjsvHqf9pOZe+z
nDJTzBzXcZ6dRzs3cmdkFuaVsvum6OtwzvB2zoSNtb21+Ra0o4kR6AiEB0rDppeVcGlf69U83X4s
JWhXg4+3PDry97u49EwxKy1IpBofVMMPvVOVm5W+bDkZMGBUvMScWSJv0SWNUHBHH0I8U3VRa02Q
XAibuY59x6/uPD77MZDHK6tofaydi5JJXLczHFJVpTABj+cAZbDfTZmPZyphRoNczwL/+9eaMwg2
tBqA/gw//QD+eGwwYbrYEcrfOwyeO/Wpd71OZKbn8HJQGeobZ/qXJWN8YabGgLERiKILPjsiL5PR
jVgAL2VsSTUdr8v6n5wZT4F58wO5zhUrLDiPbOl2HQtoxr6TPbyi5INn81b9MF9GUBDXiAU0PQYD
mfoCT8U6sh+Io7YSpa7sywEcMcQV3NA88FyPMWEtTi6mQX6dD95rAj4bnb6J7kFS8e6hRbGyih/c
otGkMSa8lQCQl2cIqI+xyAH2Xp10RCIewZAuihFqy9uusiIUM49sqwHgaZZVYJdtwR6bN9s27yyu
Tbjf0O4UlBjBDtxX+90/k57SM7rILlrS+lY/nftRAtk0SHK/tUgI8DD/BrATrBz/N/NNQ4n8laQX
k4dY33bQGCruZbuWKtlG4oDeJqm94iwsgjKaNfj/thJ8jjOP8wDLFfP/q6TpAxTgEIpGCMUctt05
/RsXC7TFNLUYc6bJl2EY6bv1Zu80mQx2nEmw4/8OvGIpMgNLOlA2NKjTygBAib804iNJ861JE6oC
r+aJO9OCTaW/VEK3rF541yUUxQWrHztccLLO4VWVRqXaXYZj9EhAptmQH1LzB0K4fAI3Scsx8TKc
iuMRtesV/2o2/wEBj4AYjjWt3o/ksy+tsWf/WXITU9cn5wSHTMko5WXMVTBY1ouv8Hi1keVX7nKx
2U7JLPeaLzcMS2SshZaZ3yHSBBiEXUFi71Zgh0JbUWSGX8unDWzBQIc8rEgTTabYZRMTsuqFJG+E
nBl7OeKoLDadeCa/y1drkPM7Qfnc9HHWfzoYYOT59K+KnPUnNhW1+J/pAMQkCLIQbV+i+xtqeGmA
aEK9mFqQGdaATihgh3l6fIAUI3ZFNVn352P+wUXeanO9HWAgahCxCjgbzbNY18qHX9FkrAfwYpSw
+AaN6wLak+Y7Tcl/xZXxyhhPGO+dYlEJtxQfYVnMT4SbU2BmSzZSfzGBwA6MiFYSwzgjfHeVMO+V
WOZH4iVOvh4UjV3Z3tHt1m9eY9UBKcXPZW8PgltorohhWoU/lO91BaiKTJSjXdxXiepOl1q83QJe
3NDrJiEAGnm61PTzcSOv8kiYo8o2DDHcB2dFGPRmJ7+j6p1tx02RFPcllvVu5ZszHcJdQxOIvczH
96RpD1h2UpA2j/ewXOo8ajMdFu4p1/FkL68N1EJvjSh2uIxWQHBry1txmLm+olJ4ZdX3TA0EmlE2
unmAnyzGmYRgp9Oni3c+7WbnC0Owm4LOvZGvuDkWN/9P6OAUzYArE4JS4xSIBBMn+w6CEhHRn+5B
TzbGOoBD59906O4LEl0tQ+i5Hr+chzHkVOpUieQjsjZkGwmd6pY1exAGjxaHEhj0Z3/nMeQiHyWG
84az/CpzF6H4/duTIHcQqecsXbWTuSy9G02JtMGDzEfR9wEJPVIiQTwiY+Hap6thSiM69RqjHxRY
c3GeVQMVHxJ3czaV/1FvAO4FDcBAF/UmlUlAPpVgWNk7TW4Mba1gPvTGBbYzFdL/HtSfisWXzkGQ
iAA7nU9xV5v6psk5X3fPzC3cZsiU3bb+EGbTySWKCLf9RrhTauMKlYw5SFYe7CPmwkjgyzrKJPAC
LDcR+vhCYAJ/HxiH6aEMdLBLnk9AVWmqZHB0K8p1S/aWJMZ/JLi6le9Fj7rrQGIg+32Q+s0Gfg+i
fsKBS3BurUJln7L16Wr7IxtzAdgqeve/rhY6V/Bs37jIUgLZ7igsHJ0M5Q/BIcwUQ4v1nPetmx36
IRt1CvOofICeVRY52tame7n4xI7I6z35rNL7iF0fpIIrQty8M6P8YKmMA3kkOuCfRImDl8yqLVBu
A/kXbBRsMJeek7NtfULRbXAkQJNYzKRxrOJ7IvAnrXm8F4jsv1CjlDuAN8xycRN7cjnBROdKvDN0
dIBNc3gA1tNvND5suq4Hrzmruo0fq6Q8BDlZtlXkR8KdiGmMbUaKq0FYvZ7GFD0EhBYVFi9tCgQf
wIEI8kPGotRahC0MDCgazz/TOMcy/Zfh5DWkpCPNu4Q49seQnmhWLB5ZJKUZNBYMw4CUJehKQ3Fn
szuRLsiTLUlk/MHcfauh2cj9aMWlvrwW/SRcKDc3dzko+3VWeIMX4bE6XdKxuJDAq+ltZ7bVzB6l
4bthPhe+yGI4L4c3INoqFFeL1QvgXs1/4LghlUxe7RYnZsYYsUvtiooE3c3WvWn+dX5k/acY3xVy
CMecJusYlwIHSw==
`protect end_protected

