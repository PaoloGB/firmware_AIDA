--=============================================================================
--! @file arrivalTimeLUT_rtl.vhd
--=============================================================================
--
-------------------------------------------------------------------------------
-- --
-- University of Bristol, High Energy Physics Group.
-- --
------------------------------------------------------------------------------- --
-- VHDL Architecture work.ArivalTimeLUT.rtl
--
--------------------------------------------------------------------------------
-- 
-- Created using using Mentor Graphics HDL Designer(TM) 2010.3 (Build 21)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

--! @brief Uses a look-up-table to convert the eight bits from the two 1:4 deserializers\n
--! into a 5-bit time ( 3 bits from the position in 8-bit deserialized data \n
--! plus two bits from position w.r.t. the strobe_4x_logic_i signal ( one pulse
--! every 4 cycles of clk_4x_logic_i 
--
--! @author David Cussans , David.Cussans@bristol.ac.uk
--
--! @date 12:46:34 11/21/12
--
--! @version v0.1
--
--! @details
--! Rising and falling edge times encoded as a LUT. Contents:
--! MRFrrrfff
--! \li M = multiple edges present ( more than one rising or falling edge)
--! \li R = at least one rising edge present
--! \li F = at least one falling edge present.
--! \li rrr = time of first rising edge
--! \li fff = time of first falling edge
ENTITY arrivalTimeLUT IS
   GENERIC( 
      g_NUM_FINE_BITS   : positive := 3;
      g_NUM_COARSE_BITS : positive := 2
   );
   PORT( 
      clk_4x_logic_i           : IN     std_logic;                                                        --! Rising edge active
      strobe_4x_logic_i        : IN     std_logic;                                                        --! Pulses high once every 4 cycles of clk_4x_logic
      deserialized_data_i      : IN     std_logic_vector (8 DOWNTO 0);                                    --! Output from the two 4-bit deserializers, concatenated with most recent bit of previous clock cycle. Clocked by clk_4x_logic_i . bit-8 is the most recent data
      first_rising_edge_time_o : OUT    std_logic_vector (g_NUM_FINE_BITS+g_NUM_COARSE_BITS-1 DOWNTO 0);  --! Position of rising edge w.r.t. 40MHz strobe. Clocked by clk_4x_logic_i
      last_falling_edge_time_o : OUT    std_logic_vector (g_NUM_FINE_BITS+g_NUM_COARSE_BITS-1 DOWNTO 0);  --! Position of rising edge w.r.t. 40MHz strobe. Clocked by clk_4x_logic_i
      rising_edge_o            : OUT    std_logic;                                                        --! goes high if there is a rising edge in the data. Clocked by clk_4x_logic_i
      falling_edge_o           : OUT    std_logic;                                                        --! goes high if there is a falling edge in the data.Clocked by clk_4x_logic_i
      multiple_edges_o         : OUT    std_logic                                                         --! there is more than one rising or falling edge transition.
   );

-- Declarations

END ENTITY arrivalTimeLUT ;

--
ARCHITECTURE rtl OF arrivalTimeLUT IS

  constant c_FALLING_EDGE_BIT : positive := 2*g_NUM_FINE_BITS;  --! Bit position of bit set when falling edge detected
  constant c_RISING_EDGE_BIT : positive :=  2*g_NUM_FINE_BITS+1;  --! Bit position of bit set when rising edge detected
  constant c_MULTI_EDGE_BIT : positive :=  2*g_NUM_FINE_BITS+2;  --! Bit position of bit set when rising edge detected


  signal s_coarse_bits : std_logic_vector(g_NUM_COARSE_BITS-1 downto 0) := "00";  --! phase w.r.t. strobe

  signal s_LUT_ENTRY : std_logic_vector(g_NUM_FINE_BITS*2 +3-1 downto 0);  -- stores intermediate LUT value.
  
  type t_LUT is array (natural range <>) of std_logic_vector(g_NUM_FINE_BITS*2 + 3 -1 downto 0);
  --! Lookup table for arrival time and rising/falling edge detection (3bits
  --! for position in 9-bit deserialized data plus two bits for rising/falling 
  constant c_LUT : t_LUT(0 to 511) := (
    "000000000", "001000000", "011000001", "001000001", "011001010", "011001010", "011000010", "001000010", --0 [0, 7]
    "011010011", "011010011", "111000011", "011010011", "011001011", "011001011", "011000011", "001000011", --1 [8, 15]
    "011011100", "011011100", "111000100", "011011100", "111001100", "111001100", "111000100", "011011100", --2 [16, 23]
    "011010100", "011010100", "111000100", "011010100", "011001100", "011001100", "011000100", "001000100", --3 [24, 31]
    "011100101", "011100101", "111000101", "011100101", "111001101", "111001101", "111000101", "011100101", --4 [32, 39]
    "111010101", "111010101", "111000101", "111010101", "111001101", "111001101", "111000101", "011100101", --5 [40, 47]
    "011011101", "011011101", "111000101", "011011101", "111001101", "111001101", "111000101", "011011101", --6 [48, 55]
    "011010101", "011010101", "111000101", "011010101", "011001101", "011001101", "011000101", "001000101", --7 [56, 63]
    "011101110", "011101110", "111000110", "011101110", "111001110", "111001110", "111000110", "011101110", --8 [64, 71]
    "111010110", "111010110", "111000110", "111010110", "111001110", "111001110", "111000110", "011101110", --9 [72, 79]
    "111011110", "111011110", "111000110", "111011110", "111001110", "111001110", "111000110", "111011110", --10 [80, 87]
    "111010110", "111010110", "111000110", "111010110", "111001110", "111001110", "111000110", "011101110", --11 [88, 95]
    "011100110", "011100110", "111000110", "011100110", "111001110", "111001110", "111000110", "011100110", --12 [96, 103]
    "111010110", "111010110", "111000110", "111010110", "111001110", "111001110", "111000110", "011100110", --13 [104, 111]
    "011011110", "011011110", "111000110", "011011110", "111001110", "111001110", "111000110", "011011110", --14 [112, 119]
    "011010110", "011010110", "111000110", "011010110", "011001110", "011001110", "011000110", "001000110", --15 [120, 127]
    "011110111", "011110111", "111000111", "011110111", "111001111", "111001111", "111000111", "011110111", --16 [128, 135]
    "111010111", "111010111", "111000111", "111010111", "111001111", "111001111", "111000111", "011110111", --17 [136, 143]
    "111011111", "111011111", "111000111", "111011111", "111001111", "111001111", "111000111", "111011111", --18 [144, 152]
    "111010111", "111010111", "111000111", "111010111", "111001111", "111001111", "111000111", "011110111", --19 [152, 159]
    "111100111", "111100111", "111000111", "111100111", "111001111", "111001111", "111000111", "111100111", --20 [160, 167]
    "111010111", "111010111", "111000111", "111010111", "111001111", "111001111", "111000111", "111100111", --21 [168, 175]
    "111011111", "111011111", "111000111", "111011111", "111001111", "111001111", "111000111", "111011111", --22 [176, 183]
    "111010111", "111010111", "111000111", "111010111", "111001111", "111001111", "111000111", "011110111", --23 [184, 191]
    "011101111", "011101111", "111000111", "011101111", "111001111", "111001111", "111000111", "011101111", --24 [192, 199]
    "111010111", "111010111", "111000111", "111010111", "111001111", "111001111", "111000111", "011101111", --25 [200, 207]
    "111011111", "111011111", "111000111", "111011111", "111001111", "111001111", "111000111", "111011111", --26 [208, 215]
    "111010111", "111010111", "111000111", "111010111", "111001111", "111001111", "111000111", "011101111", --27 [216, 223]
    "011100111", "011100111", "111000111", "011100111", "111001111", "111001111", "111000111", "011100111", --28 [224, 231]
    "111010111", "111010111", "111000111", "111010111", "111001111", "111001111", "111000111", "011100111", --29 [232, 239]
    "011011111", "011011111", "111000111", "011011111", "111001111", "111001111", "111000111", "011011111", --30 [240, 247]
    "011010111", "011010111", "111000111", "011010111", "011001111", "011001111", "011000111", "001000111", --31 [248, 255]
    "010111000", "011111000", "111000001", "011111001", "111001010", "111001010", "111000010", "011111010", --32 [256, 263]
    "111010011", "111010011", "111000011", "111010011", "111001011", "111001011", "111000011", "011111011", --33 [264, 271]
    "111011100", "111011100", "111000100", "111011100", "111001100", "111001100", "111000100", "111011100", --34 [272, 279]
    "111010100", "111010100", "111000100", "111010100", "111001100", "111001100", "111000100", "011111100", --35 [280, 287]
    "111100101", "111100101", "111000101", "111100101", "111001101", "111001101", "111000101", "111100101", --36 [288, 295]
    "111010101", "111010101", "111000101", "111010101", "111001101", "111001101", "111000101", "111100101", --37 [296, 303]
    "111011101", "111011101", "111000101", "111011101", "111001101", "111001101", "111000101", "111011101", --38 [304, 311]
    "111010101", "111010101", "111000101", "111010101", "111001101", "111001101", "111000101", "011111101", --39 [312, 319]
    "111101110", "111101110", "111000110", "111101110", "111001110", "111001110", "111000110", "111101110", --40 [320, 327]
    "111010110", "111010110", "111000110", "111010110", "111001110", "111001110", "111000110", "111101110", --41 [328, 333]
    "111011110", "111011110", "111000110", "111011110", "111001110", "111001110", "111000110", "111011110", --42 [336, 343]
    "111010110", "111010110", "111000110", "111010110", "111001110", "111001110", "111000110", "111101110", --43 [344, 351]
    "111100110", "111100110", "111000110", "111100110", "111001110", "111001110", "111000110", "111100110", --44 [352, 359]
    "111010110", "111010110", "111000110", "111010110", "111001110", "111001110", "111000110", "111100110", --45 [360, 367]
    "111011110", "111011110", "111000110", "111011110", "111001110", "111001110", "111000110", "111011110", --46 [368, 375]
    "111010110", "111010110", "111000110", "111010110", "111001110", "111001110", "111000110", "011111110", --47 [376, 383]
    "010110000", "011110000", "111000001", "011110001", "111001010", "111001010", "111000010", "011110010", --48 [384, 391]
    "111010011", "111010011", "111000011", "111010011", "111001011", "111001011", "111000011", "011110011", --49 [392, 399]
    "111011100", "111011100", "111000100", "111011100", "111001100", "111001100", "111000100", "111011100", --50 [400, 407]
    "111010100", "111010100", "111000100", "111010100", "111001100", "111001100", "111000100", "011110100", --51 [408, 415]
    "111100101", "111100101", "111000101", "111100101", "111001101", "111001101", "111000101", "111100101", --52 [416, 423]
    "111010101", "111010101", "111000101", "111010101", "111001101", "111001101", "111000101", "111100101", --53 [424, 431]
    "111011101", "111011101", "111000101", "111011101", "111001101", "111001101", "111000101", "111011101", --54 [432, 439]
    "111010101", "111010101", "111000101", "111010101", "111001101", "111001101", "111000101", "011110101", --55 [440, 447]
    "010101000", "011101000", "111000001", "011101001", "111001010", "111001010", "111000010", "011101010", --56 [448, 455]
    "111010011", "111010011", "111000011", "111010011", "111001011", "111001011", "111000011", "011101011", --57 [456, 463]
    "111011100", "111011100", "111000100", "111011100", "111001100", "111001100", "111000100", "111011100", --58 [464, 471]
    "111010100", "111010100", "111000100", "111010100", "111001100", "111001100", "111000100", "011101100", --59 [472, 479]
    "010100000", "011100000", "111000001", "011100001", "111001010", "111001010", "111000010", "011100010", --60 [480, 487]
    "111010011", "111010011", "111000011", "111010011", "111001011", "111001011", "111000011", "011100011", --61 [488, 495]
    "010011000", "011011000", "111000001", "011011001", "111001010", "111001010", "111000010", "011011010", --62 [496, 503]
    "010010000", "011010000", "111000001", "011010001", "010001000", "011001000", "010000000", "000000000" -- 63 [504, 511]
    );  
  
BEGIN

  -- purpose: uses the deserialized data as a index into
  --          a lookup table holding the position of the first rising edge (if any)
  --          and if there is a rising or falling edge
  -- type   : combinational
  -- inputs : clk_4x_logic_i
  -- outputs: arrival_time_o , rising_edge_o , falling_edge_o
  examine_lut: process (clk_4x_logic_i) -- , deserialized_data_i)
--    variable v_LUT_entry : std_logic_vector(g_NUM_FINE_BITS+2-1 downto 0);  --! Entry in LUT pointed to by deserialized data
  begin  -- process examine_lut
    
--    v_LUT_entry := c_LUT(to_integer(unsigned(deserialized_data_i)));

    if rising_edge(clk_4x_logic_i) then
      s_LUT_ENTRY <= c_LUT(to_integer(unsigned(deserialized_data_i)));
      first_rising_edge_time_o <= s_coarse_bits & s_LUT_ENTRY(g_NUM_FINE_BITS*2-1 downto g_NUM_FINE_BITS);
      last_falling_edge_time_o <= s_coarse_bits & s_LUT_ENTRY(g_NUM_FINE_BITS-1 downto 0);
      rising_edge_o  <= s_LUT_ENTRY(c_RISING_EDGE_BIT);
      falling_edge_o <= s_LUT_ENTRY(c_FALLING_EDGE_BIT);
      multiple_edges_o <= s_LUT_ENTRY(c_MULTI_EDGE_BIT); 
    end if;

  end process examine_lut;
  
  --! Coarse time stamp. Phase w.r.t. strobe
--	c_coarse_ts : entity work.CounterUp
--   PORT MAP (
--     clk   => clk_4x_logic_i,
--     ce    => '1',
--     sinit => strobe_4x_logic_i, --'0',
--	  q(31 downto 2) => open,
--     q(1 downto 0)  => s_coarse_bits
--	);
--  
  	c_coarse_ts : entity work.CounterWithReset
  	GENERIC MAP (
  	  g_COUNTER_WIDTH => 2 )
   PORT MAP (
     clock_i   => clk_4x_logic_i,
     enable_i   => '1',
     reset_i => strobe_4x_logic_i,        -- Synchronous reset, so the counter will present result_o="11" when reset_i='1'
     result_o => s_coarse_bits
	);
	
END ARCHITECTURE rtl;

